magic
tech sky130A
magscale 1 2
timestamp 1615910487
<< nwell >>
rect -1550 -800 1550 800
<< pmos >>
rect -1456 -700 -1316 700
rect -1258 -700 -1118 700
rect -1060 -700 -920 700
rect -862 -700 -722 700
rect -664 -700 -524 700
rect -466 -700 -326 700
rect -268 -700 -128 700
rect -70 -700 70 700
rect 128 -700 268 700
rect 326 -700 466 700
rect 524 -700 664 700
rect 722 -700 862 700
rect 920 -700 1060 700
rect 1118 -700 1258 700
rect 1316 -700 1456 700
<< pdiff >>
rect -1514 688 -1456 700
rect -1514 -688 -1502 688
rect -1468 -688 -1456 688
rect -1514 -700 -1456 -688
rect -1316 688 -1258 700
rect -1316 -688 -1304 688
rect -1270 -688 -1258 688
rect -1316 -700 -1258 -688
rect -1118 688 -1060 700
rect -1118 -688 -1106 688
rect -1072 -688 -1060 688
rect -1118 -700 -1060 -688
rect -920 688 -862 700
rect -920 -688 -908 688
rect -874 -688 -862 688
rect -920 -700 -862 -688
rect -722 688 -664 700
rect -722 -688 -710 688
rect -676 -688 -664 688
rect -722 -700 -664 -688
rect -524 688 -466 700
rect -524 -688 -512 688
rect -478 -688 -466 688
rect -524 -700 -466 -688
rect -326 688 -268 700
rect -326 -688 -314 688
rect -280 -688 -268 688
rect -326 -700 -268 -688
rect -128 688 -70 700
rect -128 -688 -116 688
rect -82 -688 -70 688
rect -128 -700 -70 -688
rect 70 688 128 700
rect 70 -688 82 688
rect 116 -688 128 688
rect 70 -700 128 -688
rect 268 688 326 700
rect 268 -688 280 688
rect 314 -688 326 688
rect 268 -700 326 -688
rect 466 688 524 700
rect 466 -688 478 688
rect 512 -688 524 688
rect 466 -700 524 -688
rect 664 688 722 700
rect 664 -688 676 688
rect 710 -688 722 688
rect 664 -700 722 -688
rect 862 688 920 700
rect 862 -688 874 688
rect 908 -688 920 688
rect 862 -700 920 -688
rect 1060 688 1118 700
rect 1060 -688 1072 688
rect 1106 -688 1118 688
rect 1060 -700 1118 -688
rect 1258 688 1316 700
rect 1258 -688 1270 688
rect 1304 -688 1316 688
rect 1258 -700 1316 -688
rect 1456 688 1514 700
rect 1456 -688 1468 688
rect 1502 -688 1514 688
rect 1456 -700 1514 -688
<< pdiffc >>
rect -1502 -688 -1468 688
rect -1304 -688 -1270 688
rect -1106 -688 -1072 688
rect -908 -688 -874 688
rect -710 -688 -676 688
rect -512 -688 -478 688
rect -314 -688 -280 688
rect -116 -688 -82 688
rect 82 -688 116 688
rect 280 -688 314 688
rect 478 -688 512 688
rect 676 -688 710 688
rect 874 -688 908 688
rect 1072 -688 1106 688
rect 1270 -688 1304 688
rect 1468 -688 1502 688
<< poly >>
rect -1456 781 -1316 797
rect -1456 747 -1440 781
rect -1332 747 -1316 781
rect -1456 700 -1316 747
rect -1258 781 -1118 797
rect -1258 747 -1242 781
rect -1134 747 -1118 781
rect -1258 700 -1118 747
rect -1060 781 -920 797
rect -1060 747 -1044 781
rect -936 747 -920 781
rect -1060 700 -920 747
rect -862 781 -722 797
rect -862 747 -846 781
rect -738 747 -722 781
rect -862 700 -722 747
rect -664 781 -524 797
rect -664 747 -648 781
rect -540 747 -524 781
rect -664 700 -524 747
rect -466 781 -326 797
rect -466 747 -450 781
rect -342 747 -326 781
rect -466 700 -326 747
rect -268 781 -128 797
rect -268 747 -252 781
rect -144 747 -128 781
rect -268 700 -128 747
rect -70 781 70 797
rect -70 747 -54 781
rect 54 747 70 781
rect -70 700 70 747
rect 128 781 268 797
rect 128 747 144 781
rect 252 747 268 781
rect 128 700 268 747
rect 326 781 466 797
rect 326 747 342 781
rect 450 747 466 781
rect 326 700 466 747
rect 524 781 664 797
rect 524 747 540 781
rect 648 747 664 781
rect 524 700 664 747
rect 722 781 862 797
rect 722 747 738 781
rect 846 747 862 781
rect 722 700 862 747
rect 920 781 1060 797
rect 920 747 936 781
rect 1044 747 1060 781
rect 920 700 1060 747
rect 1118 781 1258 797
rect 1118 747 1134 781
rect 1242 747 1258 781
rect 1118 700 1258 747
rect 1316 781 1456 797
rect 1316 747 1332 781
rect 1440 747 1456 781
rect 1316 700 1456 747
rect -1456 -747 -1316 -700
rect -1456 -781 -1440 -747
rect -1332 -781 -1316 -747
rect -1456 -797 -1316 -781
rect -1258 -747 -1118 -700
rect -1258 -781 -1242 -747
rect -1134 -781 -1118 -747
rect -1258 -797 -1118 -781
rect -1060 -747 -920 -700
rect -1060 -781 -1044 -747
rect -936 -781 -920 -747
rect -1060 -797 -920 -781
rect -862 -747 -722 -700
rect -862 -781 -846 -747
rect -738 -781 -722 -747
rect -862 -797 -722 -781
rect -664 -747 -524 -700
rect -664 -781 -648 -747
rect -540 -781 -524 -747
rect -664 -797 -524 -781
rect -466 -747 -326 -700
rect -466 -781 -450 -747
rect -342 -781 -326 -747
rect -466 -797 -326 -781
rect -268 -747 -128 -700
rect -268 -781 -252 -747
rect -144 -781 -128 -747
rect -268 -797 -128 -781
rect -70 -747 70 -700
rect -70 -781 -54 -747
rect 54 -781 70 -747
rect -70 -797 70 -781
rect 128 -747 268 -700
rect 128 -781 144 -747
rect 252 -781 268 -747
rect 128 -797 268 -781
rect 326 -747 466 -700
rect 326 -781 342 -747
rect 450 -781 466 -747
rect 326 -797 466 -781
rect 524 -747 664 -700
rect 524 -781 540 -747
rect 648 -781 664 -747
rect 524 -797 664 -781
rect 722 -747 862 -700
rect 722 -781 738 -747
rect 846 -781 862 -747
rect 722 -797 862 -781
rect 920 -747 1060 -700
rect 920 -781 936 -747
rect 1044 -781 1060 -747
rect 920 -797 1060 -781
rect 1118 -747 1258 -700
rect 1118 -781 1134 -747
rect 1242 -781 1258 -747
rect 1118 -797 1258 -781
rect 1316 -747 1456 -700
rect 1316 -781 1332 -747
rect 1440 -781 1456 -747
rect 1316 -797 1456 -781
<< polycont >>
rect -1440 747 -1332 781
rect -1242 747 -1134 781
rect -1044 747 -936 781
rect -846 747 -738 781
rect -648 747 -540 781
rect -450 747 -342 781
rect -252 747 -144 781
rect -54 747 54 781
rect 144 747 252 781
rect 342 747 450 781
rect 540 747 648 781
rect 738 747 846 781
rect 936 747 1044 781
rect 1134 747 1242 781
rect 1332 747 1440 781
rect -1440 -781 -1332 -747
rect -1242 -781 -1134 -747
rect -1044 -781 -936 -747
rect -846 -781 -738 -747
rect -648 -781 -540 -747
rect -450 -781 -342 -747
rect -252 -781 -144 -747
rect -54 -781 54 -747
rect 144 -781 252 -747
rect 342 -781 450 -747
rect 540 -781 648 -747
rect 738 -781 846 -747
rect 936 -781 1044 -747
rect 1134 -781 1242 -747
rect 1332 -781 1440 -747
<< locali >>
rect -1456 747 -1440 781
rect -1332 747 -1316 781
rect -1258 747 -1242 781
rect -1134 747 -1118 781
rect -1060 747 -1044 781
rect -936 747 -920 781
rect -862 747 -846 781
rect -738 747 -722 781
rect -664 747 -648 781
rect -540 747 -524 781
rect -466 747 -450 781
rect -342 747 -326 781
rect -268 747 -252 781
rect -144 747 -128 781
rect -70 747 -54 781
rect 54 747 70 781
rect 128 747 144 781
rect 252 747 268 781
rect 326 747 342 781
rect 450 747 466 781
rect 524 747 540 781
rect 648 747 664 781
rect 722 747 738 781
rect 846 747 862 781
rect 920 747 936 781
rect 1044 747 1060 781
rect 1118 747 1134 781
rect 1242 747 1258 781
rect 1316 747 1332 781
rect 1440 747 1456 781
rect -1502 688 -1468 704
rect -1502 -704 -1468 -688
rect -1304 688 -1270 704
rect -1304 -704 -1270 -688
rect -1106 688 -1072 704
rect -1106 -704 -1072 -688
rect -908 688 -874 704
rect -908 -704 -874 -688
rect -710 688 -676 704
rect -710 -704 -676 -688
rect -512 688 -478 704
rect -512 -704 -478 -688
rect -314 688 -280 704
rect -314 -704 -280 -688
rect -116 688 -82 704
rect -116 -704 -82 -688
rect 82 688 116 704
rect 82 -704 116 -688
rect 280 688 314 704
rect 280 -704 314 -688
rect 478 688 512 704
rect 478 -704 512 -688
rect 676 688 710 704
rect 676 -704 710 -688
rect 874 688 908 704
rect 874 -704 908 -688
rect 1072 688 1106 704
rect 1072 -704 1106 -688
rect 1270 688 1304 704
rect 1270 -704 1304 -688
rect 1468 688 1502 704
rect 1468 -704 1502 -688
rect -1456 -781 -1440 -747
rect -1332 -781 -1316 -747
rect -1258 -781 -1242 -747
rect -1134 -781 -1118 -747
rect -1060 -781 -1044 -747
rect -936 -781 -920 -747
rect -862 -781 -846 -747
rect -738 -781 -722 -747
rect -664 -781 -648 -747
rect -540 -781 -524 -747
rect -466 -781 -450 -747
rect -342 -781 -326 -747
rect -268 -781 -252 -747
rect -144 -781 -128 -747
rect -70 -781 -54 -747
rect 54 -781 70 -747
rect 128 -781 144 -747
rect 252 -781 268 -747
rect 326 -781 342 -747
rect 450 -781 466 -747
rect 524 -781 540 -747
rect 648 -781 664 -747
rect 722 -781 738 -747
rect 846 -781 862 -747
rect 920 -781 936 -747
rect 1044 -781 1060 -747
rect 1118 -781 1134 -747
rect 1242 -781 1258 -747
rect 1316 -781 1332 -747
rect 1440 -781 1456 -747
<< viali >>
rect -1440 747 -1332 781
rect -1242 747 -1134 781
rect -1044 747 -936 781
rect -846 747 -738 781
rect -648 747 -540 781
rect -450 747 -342 781
rect -252 747 -144 781
rect -54 747 54 781
rect 144 747 252 781
rect 342 747 450 781
rect 540 747 648 781
rect 738 747 846 781
rect 936 747 1044 781
rect 1134 747 1242 781
rect 1332 747 1440 781
rect -1502 -688 -1468 688
rect -1304 -688 -1270 688
rect -1106 -688 -1072 688
rect -908 -688 -874 688
rect -710 -688 -676 688
rect -512 -688 -478 688
rect -314 -688 -280 688
rect -116 -688 -82 688
rect 82 -688 116 688
rect 280 -688 314 688
rect 478 -688 512 688
rect 676 -688 710 688
rect 874 -688 908 688
rect 1072 -688 1106 688
rect 1270 -688 1304 688
rect 1468 -688 1502 688
rect -1440 -781 -1332 -747
rect -1242 -781 -1134 -747
rect -1044 -781 -936 -747
rect -846 -781 -738 -747
rect -648 -781 -540 -747
rect -450 -781 -342 -747
rect -252 -781 -144 -747
rect -54 -781 54 -747
rect 144 -781 252 -747
rect 342 -781 450 -747
rect 540 -781 648 -747
rect 738 -781 846 -747
rect 936 -781 1044 -747
rect 1134 -781 1242 -747
rect 1332 -781 1440 -747
<< metal1 >>
rect -1452 781 -1320 787
rect -1452 747 -1440 781
rect -1332 747 -1320 781
rect -1452 741 -1320 747
rect -1254 781 -1122 787
rect -1254 747 -1242 781
rect -1134 747 -1122 781
rect -1254 741 -1122 747
rect -1056 781 -924 787
rect -1056 747 -1044 781
rect -936 747 -924 781
rect -1056 741 -924 747
rect -858 781 -726 787
rect -858 747 -846 781
rect -738 747 -726 781
rect -858 741 -726 747
rect -660 781 -528 787
rect -660 747 -648 781
rect -540 747 -528 781
rect -660 741 -528 747
rect -462 781 -330 787
rect -462 747 -450 781
rect -342 747 -330 781
rect -462 741 -330 747
rect -264 781 -132 787
rect -264 747 -252 781
rect -144 747 -132 781
rect -264 741 -132 747
rect -66 781 66 787
rect -66 747 -54 781
rect 54 747 66 781
rect -66 741 66 747
rect 132 781 264 787
rect 132 747 144 781
rect 252 747 264 781
rect 132 741 264 747
rect 330 781 462 787
rect 330 747 342 781
rect 450 747 462 781
rect 330 741 462 747
rect 528 781 660 787
rect 528 747 540 781
rect 648 747 660 781
rect 528 741 660 747
rect 726 781 858 787
rect 726 747 738 781
rect 846 747 858 781
rect 726 741 858 747
rect 924 781 1056 787
rect 924 747 936 781
rect 1044 747 1056 781
rect 924 741 1056 747
rect 1122 781 1254 787
rect 1122 747 1134 781
rect 1242 747 1254 781
rect 1122 741 1254 747
rect 1320 781 1452 787
rect 1320 747 1332 781
rect 1440 747 1452 781
rect 1320 741 1452 747
rect -1508 688 -1462 700
rect -1508 -688 -1502 688
rect -1468 -688 -1462 688
rect -1508 -700 -1462 -688
rect -1310 688 -1264 700
rect -1310 -688 -1304 688
rect -1270 -688 -1264 688
rect -1310 -700 -1264 -688
rect -1112 688 -1066 700
rect -1112 -688 -1106 688
rect -1072 -688 -1066 688
rect -1112 -700 -1066 -688
rect -914 688 -868 700
rect -914 -688 -908 688
rect -874 -688 -868 688
rect -914 -700 -868 -688
rect -716 688 -670 700
rect -716 -688 -710 688
rect -676 -688 -670 688
rect -716 -700 -670 -688
rect -518 688 -472 700
rect -518 -688 -512 688
rect -478 -688 -472 688
rect -518 -700 -472 -688
rect -320 688 -274 700
rect -320 -688 -314 688
rect -280 -688 -274 688
rect -320 -700 -274 -688
rect -122 688 -76 700
rect -122 -688 -116 688
rect -82 -688 -76 688
rect -122 -700 -76 -688
rect 76 688 122 700
rect 76 -688 82 688
rect 116 -688 122 688
rect 76 -700 122 -688
rect 274 688 320 700
rect 274 -688 280 688
rect 314 -688 320 688
rect 274 -700 320 -688
rect 472 688 518 700
rect 472 -688 478 688
rect 512 -688 518 688
rect 472 -700 518 -688
rect 670 688 716 700
rect 670 -688 676 688
rect 710 -688 716 688
rect 670 -700 716 -688
rect 868 688 914 700
rect 868 -688 874 688
rect 908 -688 914 688
rect 868 -700 914 -688
rect 1066 688 1112 700
rect 1066 -688 1072 688
rect 1106 -688 1112 688
rect 1066 -700 1112 -688
rect 1264 688 1310 700
rect 1264 -688 1270 688
rect 1304 -688 1310 688
rect 1264 -700 1310 -688
rect 1462 688 1508 700
rect 1462 -688 1468 688
rect 1502 -688 1508 688
rect 1462 -700 1508 -688
rect -1452 -747 -1320 -741
rect -1452 -781 -1440 -747
rect -1332 -781 -1320 -747
rect -1452 -787 -1320 -781
rect -1254 -747 -1122 -741
rect -1254 -781 -1242 -747
rect -1134 -781 -1122 -747
rect -1254 -787 -1122 -781
rect -1056 -747 -924 -741
rect -1056 -781 -1044 -747
rect -936 -781 -924 -747
rect -1056 -787 -924 -781
rect -858 -747 -726 -741
rect -858 -781 -846 -747
rect -738 -781 -726 -747
rect -858 -787 -726 -781
rect -660 -747 -528 -741
rect -660 -781 -648 -747
rect -540 -781 -528 -747
rect -660 -787 -528 -781
rect -462 -747 -330 -741
rect -462 -781 -450 -747
rect -342 -781 -330 -747
rect -462 -787 -330 -781
rect -264 -747 -132 -741
rect -264 -781 -252 -747
rect -144 -781 -132 -747
rect -264 -787 -132 -781
rect -66 -747 66 -741
rect -66 -781 -54 -747
rect 54 -781 66 -747
rect -66 -787 66 -781
rect 132 -747 264 -741
rect 132 -781 144 -747
rect 252 -781 264 -747
rect 132 -787 264 -781
rect 330 -747 462 -741
rect 330 -781 342 -747
rect 450 -781 462 -747
rect 330 -787 462 -781
rect 528 -747 660 -741
rect 528 -781 540 -747
rect 648 -781 660 -747
rect 528 -787 660 -781
rect 726 -747 858 -741
rect 726 -781 738 -747
rect 846 -781 858 -747
rect 726 -787 858 -781
rect 924 -747 1056 -741
rect 924 -781 936 -747
rect 1044 -781 1056 -747
rect 924 -787 1056 -781
rect 1122 -747 1254 -741
rect 1122 -781 1134 -747
rect 1242 -781 1254 -747
rect 1122 -787 1254 -781
rect 1320 -747 1452 -741
rect 1320 -781 1332 -747
rect 1440 -781 1452 -747
rect 1320 -787 1452 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
