magic
tech sky130A
timestamp 1615910487
<< nwell >>
rect -775 -1128 775 1128
<< pmos >>
rect -728 397 -658 1097
rect -629 397 -559 1097
rect -530 397 -460 1097
rect -431 397 -361 1097
rect -332 397 -262 1097
rect -233 397 -163 1097
rect -134 397 -64 1097
rect -35 397 35 1097
rect 64 397 134 1097
rect 163 397 233 1097
rect 262 397 332 1097
rect 361 397 431 1097
rect 460 397 530 1097
rect 559 397 629 1097
rect 658 397 728 1097
rect -728 -350 -658 350
rect -629 -350 -559 350
rect -530 -350 -460 350
rect -431 -350 -361 350
rect -332 -350 -262 350
rect -233 -350 -163 350
rect -134 -350 -64 350
rect -35 -350 35 350
rect 64 -350 134 350
rect 163 -350 233 350
rect 262 -350 332 350
rect 361 -350 431 350
rect 460 -350 530 350
rect 559 -350 629 350
rect 658 -350 728 350
rect -728 -1097 -658 -397
rect -629 -1097 -559 -397
rect -530 -1097 -460 -397
rect -431 -1097 -361 -397
rect -332 -1097 -262 -397
rect -233 -1097 -163 -397
rect -134 -1097 -64 -397
rect -35 -1097 35 -397
rect 64 -1097 134 -397
rect 163 -1097 233 -397
rect 262 -1097 332 -397
rect 361 -1097 431 -397
rect 460 -1097 530 -397
rect 559 -1097 629 -397
rect 658 -1097 728 -397
<< pdiff >>
rect -757 1091 -728 1097
rect -757 403 -751 1091
rect -734 403 -728 1091
rect -757 397 -728 403
rect -658 1091 -629 1097
rect -658 403 -652 1091
rect -635 403 -629 1091
rect -658 397 -629 403
rect -559 1091 -530 1097
rect -559 403 -553 1091
rect -536 403 -530 1091
rect -559 397 -530 403
rect -460 1091 -431 1097
rect -460 403 -454 1091
rect -437 403 -431 1091
rect -460 397 -431 403
rect -361 1091 -332 1097
rect -361 403 -355 1091
rect -338 403 -332 1091
rect -361 397 -332 403
rect -262 1091 -233 1097
rect -262 403 -256 1091
rect -239 403 -233 1091
rect -262 397 -233 403
rect -163 1091 -134 1097
rect -163 403 -157 1091
rect -140 403 -134 1091
rect -163 397 -134 403
rect -64 1091 -35 1097
rect -64 403 -58 1091
rect -41 403 -35 1091
rect -64 397 -35 403
rect 35 1091 64 1097
rect 35 403 41 1091
rect 58 403 64 1091
rect 35 397 64 403
rect 134 1091 163 1097
rect 134 403 140 1091
rect 157 403 163 1091
rect 134 397 163 403
rect 233 1091 262 1097
rect 233 403 239 1091
rect 256 403 262 1091
rect 233 397 262 403
rect 332 1091 361 1097
rect 332 403 338 1091
rect 355 403 361 1091
rect 332 397 361 403
rect 431 1091 460 1097
rect 431 403 437 1091
rect 454 403 460 1091
rect 431 397 460 403
rect 530 1091 559 1097
rect 530 403 536 1091
rect 553 403 559 1091
rect 530 397 559 403
rect 629 1091 658 1097
rect 629 403 635 1091
rect 652 403 658 1091
rect 629 397 658 403
rect 728 1091 757 1097
rect 728 403 734 1091
rect 751 403 757 1091
rect 728 397 757 403
rect -757 344 -728 350
rect -757 -344 -751 344
rect -734 -344 -728 344
rect -757 -350 -728 -344
rect -658 344 -629 350
rect -658 -344 -652 344
rect -635 -344 -629 344
rect -658 -350 -629 -344
rect -559 344 -530 350
rect -559 -344 -553 344
rect -536 -344 -530 344
rect -559 -350 -530 -344
rect -460 344 -431 350
rect -460 -344 -454 344
rect -437 -344 -431 344
rect -460 -350 -431 -344
rect -361 344 -332 350
rect -361 -344 -355 344
rect -338 -344 -332 344
rect -361 -350 -332 -344
rect -262 344 -233 350
rect -262 -344 -256 344
rect -239 -344 -233 344
rect -262 -350 -233 -344
rect -163 344 -134 350
rect -163 -344 -157 344
rect -140 -344 -134 344
rect -163 -350 -134 -344
rect -64 344 -35 350
rect -64 -344 -58 344
rect -41 -344 -35 344
rect -64 -350 -35 -344
rect 35 344 64 350
rect 35 -344 41 344
rect 58 -344 64 344
rect 35 -350 64 -344
rect 134 344 163 350
rect 134 -344 140 344
rect 157 -344 163 344
rect 134 -350 163 -344
rect 233 344 262 350
rect 233 -344 239 344
rect 256 -344 262 344
rect 233 -350 262 -344
rect 332 344 361 350
rect 332 -344 338 344
rect 355 -344 361 344
rect 332 -350 361 -344
rect 431 344 460 350
rect 431 -344 437 344
rect 454 -344 460 344
rect 431 -350 460 -344
rect 530 344 559 350
rect 530 -344 536 344
rect 553 -344 559 344
rect 530 -350 559 -344
rect 629 344 658 350
rect 629 -344 635 344
rect 652 -344 658 344
rect 629 -350 658 -344
rect 728 344 757 350
rect 728 -344 734 344
rect 751 -344 757 344
rect 728 -350 757 -344
rect -757 -403 -728 -397
rect -757 -1091 -751 -403
rect -734 -1091 -728 -403
rect -757 -1097 -728 -1091
rect -658 -403 -629 -397
rect -658 -1091 -652 -403
rect -635 -1091 -629 -403
rect -658 -1097 -629 -1091
rect -559 -403 -530 -397
rect -559 -1091 -553 -403
rect -536 -1091 -530 -403
rect -559 -1097 -530 -1091
rect -460 -403 -431 -397
rect -460 -1091 -454 -403
rect -437 -1091 -431 -403
rect -460 -1097 -431 -1091
rect -361 -403 -332 -397
rect -361 -1091 -355 -403
rect -338 -1091 -332 -403
rect -361 -1097 -332 -1091
rect -262 -403 -233 -397
rect -262 -1091 -256 -403
rect -239 -1091 -233 -403
rect -262 -1097 -233 -1091
rect -163 -403 -134 -397
rect -163 -1091 -157 -403
rect -140 -1091 -134 -403
rect -163 -1097 -134 -1091
rect -64 -403 -35 -397
rect -64 -1091 -58 -403
rect -41 -1091 -35 -403
rect -64 -1097 -35 -1091
rect 35 -403 64 -397
rect 35 -1091 41 -403
rect 58 -1091 64 -403
rect 35 -1097 64 -1091
rect 134 -403 163 -397
rect 134 -1091 140 -403
rect 157 -1091 163 -403
rect 134 -1097 163 -1091
rect 233 -403 262 -397
rect 233 -1091 239 -403
rect 256 -1091 262 -403
rect 233 -1097 262 -1091
rect 332 -403 361 -397
rect 332 -1091 338 -403
rect 355 -1091 361 -403
rect 332 -1097 361 -1091
rect 431 -403 460 -397
rect 431 -1091 437 -403
rect 454 -1091 460 -403
rect 431 -1097 460 -1091
rect 530 -403 559 -397
rect 530 -1091 536 -403
rect 553 -1091 559 -403
rect 530 -1097 559 -1091
rect 629 -403 658 -397
rect 629 -1091 635 -403
rect 652 -1091 658 -403
rect 629 -1097 658 -1091
rect 728 -403 757 -397
rect 728 -1091 734 -403
rect 751 -1091 757 -403
rect 728 -1097 757 -1091
<< pdiffc >>
rect -751 403 -734 1091
rect -652 403 -635 1091
rect -553 403 -536 1091
rect -454 403 -437 1091
rect -355 403 -338 1091
rect -256 403 -239 1091
rect -157 403 -140 1091
rect -58 403 -41 1091
rect 41 403 58 1091
rect 140 403 157 1091
rect 239 403 256 1091
rect 338 403 355 1091
rect 437 403 454 1091
rect 536 403 553 1091
rect 635 403 652 1091
rect 734 403 751 1091
rect -751 -344 -734 344
rect -652 -344 -635 344
rect -553 -344 -536 344
rect -454 -344 -437 344
rect -355 -344 -338 344
rect -256 -344 -239 344
rect -157 -344 -140 344
rect -58 -344 -41 344
rect 41 -344 58 344
rect 140 -344 157 344
rect 239 -344 256 344
rect 338 -344 355 344
rect 437 -344 454 344
rect 536 -344 553 344
rect 635 -344 652 344
rect 734 -344 751 344
rect -751 -1091 -734 -403
rect -652 -1091 -635 -403
rect -553 -1091 -536 -403
rect -454 -1091 -437 -403
rect -355 -1091 -338 -403
rect -256 -1091 -239 -403
rect -157 -1091 -140 -403
rect -58 -1091 -41 -403
rect 41 -1091 58 -403
rect 140 -1091 157 -403
rect 239 -1091 256 -403
rect 338 -1091 355 -403
rect 437 -1091 454 -403
rect 536 -1091 553 -403
rect 635 -1091 652 -403
rect 734 -1091 751 -403
<< poly >>
rect -728 1097 -658 1110
rect -629 1097 -559 1110
rect -530 1097 -460 1110
rect -431 1097 -361 1110
rect -332 1097 -262 1110
rect -233 1097 -163 1110
rect -134 1097 -64 1110
rect -35 1097 35 1110
rect 64 1097 134 1110
rect 163 1097 233 1110
rect 262 1097 332 1110
rect 361 1097 431 1110
rect 460 1097 530 1110
rect 559 1097 629 1110
rect 658 1097 728 1110
rect -728 384 -658 397
rect -629 384 -559 397
rect -530 384 -460 397
rect -431 384 -361 397
rect -332 384 -262 397
rect -233 384 -163 397
rect -134 384 -64 397
rect -35 384 35 397
rect 64 384 134 397
rect 163 384 233 397
rect 262 384 332 397
rect 361 384 431 397
rect 460 384 530 397
rect 559 384 629 397
rect 658 384 728 397
rect -728 350 -658 363
rect -629 350 -559 363
rect -530 350 -460 363
rect -431 350 -361 363
rect -332 350 -262 363
rect -233 350 -163 363
rect -134 350 -64 363
rect -35 350 35 363
rect 64 350 134 363
rect 163 350 233 363
rect 262 350 332 363
rect 361 350 431 363
rect 460 350 530 363
rect 559 350 629 363
rect 658 350 728 363
rect -728 -363 -658 -350
rect -629 -363 -559 -350
rect -530 -363 -460 -350
rect -431 -363 -361 -350
rect -332 -363 -262 -350
rect -233 -363 -163 -350
rect -134 -363 -64 -350
rect -35 -363 35 -350
rect 64 -363 134 -350
rect 163 -363 233 -350
rect 262 -363 332 -350
rect 361 -363 431 -350
rect 460 -363 530 -350
rect 559 -363 629 -350
rect 658 -363 728 -350
rect -728 -397 -658 -384
rect -629 -397 -559 -384
rect -530 -397 -460 -384
rect -431 -397 -361 -384
rect -332 -397 -262 -384
rect -233 -397 -163 -384
rect -134 -397 -64 -384
rect -35 -397 35 -384
rect 64 -397 134 -384
rect 163 -397 233 -384
rect 262 -397 332 -384
rect 361 -397 431 -384
rect 460 -397 530 -384
rect 559 -397 629 -384
rect 658 -397 728 -384
rect -728 -1110 -658 -1097
rect -629 -1110 -559 -1097
rect -530 -1110 -460 -1097
rect -431 -1110 -361 -1097
rect -332 -1110 -262 -1097
rect -233 -1110 -163 -1097
rect -134 -1110 -64 -1097
rect -35 -1110 35 -1097
rect 64 -1110 134 -1097
rect 163 -1110 233 -1097
rect 262 -1110 332 -1097
rect 361 -1110 431 -1097
rect 460 -1110 530 -1097
rect 559 -1110 629 -1097
rect 658 -1110 728 -1097
<< locali >>
rect -751 1091 -734 1099
rect -751 395 -734 403
rect -652 1091 -635 1099
rect -652 395 -635 403
rect -553 1091 -536 1099
rect -553 395 -536 403
rect -454 1091 -437 1099
rect -454 395 -437 403
rect -355 1091 -338 1099
rect -355 395 -338 403
rect -256 1091 -239 1099
rect -256 395 -239 403
rect -157 1091 -140 1099
rect -157 395 -140 403
rect -58 1091 -41 1099
rect -58 395 -41 403
rect 41 1091 58 1099
rect 41 395 58 403
rect 140 1091 157 1099
rect 140 395 157 403
rect 239 1091 256 1099
rect 239 395 256 403
rect 338 1091 355 1099
rect 338 395 355 403
rect 437 1091 454 1099
rect 437 395 454 403
rect 536 1091 553 1099
rect 536 395 553 403
rect 635 1091 652 1099
rect 635 395 652 403
rect 734 1091 751 1099
rect 734 395 751 403
rect -751 344 -734 352
rect -751 -352 -734 -344
rect -652 344 -635 352
rect -652 -352 -635 -344
rect -553 344 -536 352
rect -553 -352 -536 -344
rect -454 344 -437 352
rect -454 -352 -437 -344
rect -355 344 -338 352
rect -355 -352 -338 -344
rect -256 344 -239 352
rect -256 -352 -239 -344
rect -157 344 -140 352
rect -157 -352 -140 -344
rect -58 344 -41 352
rect -58 -352 -41 -344
rect 41 344 58 352
rect 41 -352 58 -344
rect 140 344 157 352
rect 140 -352 157 -344
rect 239 344 256 352
rect 239 -352 256 -344
rect 338 344 355 352
rect 338 -352 355 -344
rect 437 344 454 352
rect 437 -352 454 -344
rect 536 344 553 352
rect 536 -352 553 -344
rect 635 344 652 352
rect 635 -352 652 -344
rect 734 344 751 352
rect 734 -352 751 -344
rect -751 -403 -734 -395
rect -751 -1099 -734 -1091
rect -652 -403 -635 -395
rect -652 -1099 -635 -1091
rect -553 -403 -536 -395
rect -553 -1099 -536 -1091
rect -454 -403 -437 -395
rect -454 -1099 -437 -1091
rect -355 -403 -338 -395
rect -355 -1099 -338 -1091
rect -256 -403 -239 -395
rect -256 -1099 -239 -1091
rect -157 -403 -140 -395
rect -157 -1099 -140 -1091
rect -58 -403 -41 -395
rect -58 -1099 -41 -1091
rect 41 -403 58 -395
rect 41 -1099 58 -1091
rect 140 -403 157 -395
rect 140 -1099 157 -1091
rect 239 -403 256 -395
rect 239 -1099 256 -1091
rect 338 -403 355 -395
rect 338 -1099 355 -1091
rect 437 -403 454 -395
rect 437 -1099 454 -1091
rect 536 -403 553 -395
rect 536 -1099 553 -1091
rect 635 -403 652 -395
rect 635 -1099 652 -1091
rect 734 -403 751 -395
rect 734 -1099 751 -1091
<< viali >>
rect -751 403 -734 1091
rect -652 403 -635 1091
rect -553 403 -536 1091
rect -454 403 -437 1091
rect -355 403 -338 1091
rect -256 403 -239 1091
rect -157 403 -140 1091
rect -58 403 -41 1091
rect 41 403 58 1091
rect 140 403 157 1091
rect 239 403 256 1091
rect 338 403 355 1091
rect 437 403 454 1091
rect 536 403 553 1091
rect 635 403 652 1091
rect 734 403 751 1091
rect -751 -344 -734 344
rect -652 -344 -635 344
rect -553 -344 -536 344
rect -454 -344 -437 344
rect -355 -344 -338 344
rect -256 -344 -239 344
rect -157 -344 -140 344
rect -58 -344 -41 344
rect 41 -344 58 344
rect 140 -344 157 344
rect 239 -344 256 344
rect 338 -344 355 344
rect 437 -344 454 344
rect 536 -344 553 344
rect 635 -344 652 344
rect 734 -344 751 344
rect -751 -1091 -734 -403
rect -652 -1091 -635 -403
rect -553 -1091 -536 -403
rect -454 -1091 -437 -403
rect -355 -1091 -338 -403
rect -256 -1091 -239 -403
rect -157 -1091 -140 -403
rect -58 -1091 -41 -403
rect 41 -1091 58 -403
rect 140 -1091 157 -403
rect 239 -1091 256 -403
rect 338 -1091 355 -403
rect 437 -1091 454 -403
rect 536 -1091 553 -403
rect 635 -1091 652 -403
rect 734 -1091 751 -403
<< metal1 >>
rect -754 1091 -731 1097
rect -754 403 -751 1091
rect -734 403 -731 1091
rect -754 397 -731 403
rect -655 1091 -632 1097
rect -655 403 -652 1091
rect -635 403 -632 1091
rect -655 397 -632 403
rect -556 1091 -533 1097
rect -556 403 -553 1091
rect -536 403 -533 1091
rect -556 397 -533 403
rect -457 1091 -434 1097
rect -457 403 -454 1091
rect -437 403 -434 1091
rect -457 397 -434 403
rect -358 1091 -335 1097
rect -358 403 -355 1091
rect -338 403 -335 1091
rect -358 397 -335 403
rect -259 1091 -236 1097
rect -259 403 -256 1091
rect -239 403 -236 1091
rect -259 397 -236 403
rect -160 1091 -137 1097
rect -160 403 -157 1091
rect -140 403 -137 1091
rect -160 397 -137 403
rect -61 1091 -38 1097
rect -61 403 -58 1091
rect -41 403 -38 1091
rect -61 397 -38 403
rect 38 1091 61 1097
rect 38 403 41 1091
rect 58 403 61 1091
rect 38 397 61 403
rect 137 1091 160 1097
rect 137 403 140 1091
rect 157 403 160 1091
rect 137 397 160 403
rect 236 1091 259 1097
rect 236 403 239 1091
rect 256 403 259 1091
rect 236 397 259 403
rect 335 1091 358 1097
rect 335 403 338 1091
rect 355 403 358 1091
rect 335 397 358 403
rect 434 1091 457 1097
rect 434 403 437 1091
rect 454 403 457 1091
rect 434 397 457 403
rect 533 1091 556 1097
rect 533 403 536 1091
rect 553 403 556 1091
rect 533 397 556 403
rect 632 1091 655 1097
rect 632 403 635 1091
rect 652 403 655 1091
rect 632 397 655 403
rect 731 1091 754 1097
rect 731 403 734 1091
rect 751 403 754 1091
rect 731 397 754 403
rect -754 344 -731 350
rect -754 -344 -751 344
rect -734 -344 -731 344
rect -754 -350 -731 -344
rect -655 344 -632 350
rect -655 -344 -652 344
rect -635 -344 -632 344
rect -655 -350 -632 -344
rect -556 344 -533 350
rect -556 -344 -553 344
rect -536 -344 -533 344
rect -556 -350 -533 -344
rect -457 344 -434 350
rect -457 -344 -454 344
rect -437 -344 -434 344
rect -457 -350 -434 -344
rect -358 344 -335 350
rect -358 -344 -355 344
rect -338 -344 -335 344
rect -358 -350 -335 -344
rect -259 344 -236 350
rect -259 -344 -256 344
rect -239 -344 -236 344
rect -259 -350 -236 -344
rect -160 344 -137 350
rect -160 -344 -157 344
rect -140 -344 -137 344
rect -160 -350 -137 -344
rect -61 344 -38 350
rect -61 -344 -58 344
rect -41 -344 -38 344
rect -61 -350 -38 -344
rect 38 344 61 350
rect 38 -344 41 344
rect 58 -344 61 344
rect 38 -350 61 -344
rect 137 344 160 350
rect 137 -344 140 344
rect 157 -344 160 344
rect 137 -350 160 -344
rect 236 344 259 350
rect 236 -344 239 344
rect 256 -344 259 344
rect 236 -350 259 -344
rect 335 344 358 350
rect 335 -344 338 344
rect 355 -344 358 344
rect 335 -350 358 -344
rect 434 344 457 350
rect 434 -344 437 344
rect 454 -344 457 344
rect 434 -350 457 -344
rect 533 344 556 350
rect 533 -344 536 344
rect 553 -344 556 344
rect 533 -350 556 -344
rect 632 344 655 350
rect 632 -344 635 344
rect 652 -344 655 344
rect 632 -350 655 -344
rect 731 344 754 350
rect 731 -344 734 344
rect 751 -344 754 344
rect 731 -350 754 -344
rect -754 -403 -731 -397
rect -754 -1091 -751 -403
rect -734 -1091 -731 -403
rect -754 -1097 -731 -1091
rect -655 -403 -632 -397
rect -655 -1091 -652 -403
rect -635 -1091 -632 -403
rect -655 -1097 -632 -1091
rect -556 -403 -533 -397
rect -556 -1091 -553 -403
rect -536 -1091 -533 -403
rect -556 -1097 -533 -1091
rect -457 -403 -434 -397
rect -457 -1091 -454 -403
rect -437 -1091 -434 -403
rect -457 -1097 -434 -1091
rect -358 -403 -335 -397
rect -358 -1091 -355 -403
rect -338 -1091 -335 -403
rect -358 -1097 -335 -1091
rect -259 -403 -236 -397
rect -259 -1091 -256 -403
rect -239 -1091 -236 -403
rect -259 -1097 -236 -1091
rect -160 -403 -137 -397
rect -160 -1091 -157 -403
rect -140 -1091 -137 -403
rect -160 -1097 -137 -1091
rect -61 -403 -38 -397
rect -61 -1091 -58 -403
rect -41 -1091 -38 -403
rect -61 -1097 -38 -1091
rect 38 -403 61 -397
rect 38 -1091 41 -403
rect 58 -1091 61 -403
rect 38 -1097 61 -1091
rect 137 -403 160 -397
rect 137 -1091 140 -403
rect 157 -1091 160 -403
rect 137 -1097 160 -1091
rect 236 -403 259 -397
rect 236 -1091 239 -403
rect 256 -1091 259 -403
rect 236 -1097 259 -1091
rect 335 -403 358 -397
rect 335 -1091 338 -403
rect 355 -1091 358 -403
rect 335 -1097 358 -1091
rect 434 -403 457 -397
rect 434 -1091 437 -403
rect 454 -1091 457 -403
rect 434 -1097 457 -1091
rect 533 -403 556 -397
rect 533 -1091 536 -403
rect 553 -1091 556 -403
rect 533 -1097 556 -1091
rect 632 -403 655 -397
rect 632 -1091 635 -403
rect 652 -1091 655 -403
rect 632 -1097 655 -1091
rect 731 -403 754 -397
rect 731 -1091 734 -403
rect 751 -1091 754 -403
rect 731 -1097 754 -1091
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 3 nf 15 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
