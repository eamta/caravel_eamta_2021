magic
tech sky130A
magscale 1 2
timestamp 1616176710
<< pwell >>
rect -2576 -1229 2576 1229
<< nmos >>
rect -2380 -1081 -2000 1019
rect -1942 -1081 -1562 1019
rect -1504 -1081 -1124 1019
rect -1066 -1081 -686 1019
rect -628 -1081 -248 1019
rect -190 -1081 190 1019
rect 248 -1081 628 1019
rect 686 -1081 1066 1019
rect 1124 -1081 1504 1019
rect 1562 -1081 1942 1019
rect 2000 -1081 2380 1019
<< ndiff >>
rect -2438 1007 -2380 1019
rect -2438 -1069 -2426 1007
rect -2392 -1069 -2380 1007
rect -2438 -1081 -2380 -1069
rect -2000 1007 -1942 1019
rect -2000 -1069 -1988 1007
rect -1954 -1069 -1942 1007
rect -2000 -1081 -1942 -1069
rect -1562 1007 -1504 1019
rect -1562 -1069 -1550 1007
rect -1516 -1069 -1504 1007
rect -1562 -1081 -1504 -1069
rect -1124 1007 -1066 1019
rect -1124 -1069 -1112 1007
rect -1078 -1069 -1066 1007
rect -1124 -1081 -1066 -1069
rect -686 1007 -628 1019
rect -686 -1069 -674 1007
rect -640 -1069 -628 1007
rect -686 -1081 -628 -1069
rect -248 1007 -190 1019
rect -248 -1069 -236 1007
rect -202 -1069 -190 1007
rect -248 -1081 -190 -1069
rect 190 1007 248 1019
rect 190 -1069 202 1007
rect 236 -1069 248 1007
rect 190 -1081 248 -1069
rect 628 1007 686 1019
rect 628 -1069 640 1007
rect 674 -1069 686 1007
rect 628 -1081 686 -1069
rect 1066 1007 1124 1019
rect 1066 -1069 1078 1007
rect 1112 -1069 1124 1007
rect 1066 -1081 1124 -1069
rect 1504 1007 1562 1019
rect 1504 -1069 1516 1007
rect 1550 -1069 1562 1007
rect 1504 -1081 1562 -1069
rect 1942 1007 2000 1019
rect 1942 -1069 1954 1007
rect 1988 -1069 2000 1007
rect 1942 -1081 2000 -1069
rect 2380 1007 2438 1019
rect 2380 -1069 2392 1007
rect 2426 -1069 2438 1007
rect 2380 -1081 2438 -1069
<< ndiffc >>
rect -2426 -1069 -2392 1007
rect -1988 -1069 -1954 1007
rect -1550 -1069 -1516 1007
rect -1112 -1069 -1078 1007
rect -674 -1069 -640 1007
rect -236 -1069 -202 1007
rect 202 -1069 236 1007
rect 640 -1069 674 1007
rect 1078 -1069 1112 1007
rect 1516 -1069 1550 1007
rect 1954 -1069 1988 1007
rect 2392 -1069 2426 1007
<< psubdiff >>
rect -2540 1159 -2444 1193
rect 2444 1159 2540 1193
rect -2540 1097 -2506 1159
rect 2506 1097 2540 1159
rect -2540 -1159 -2506 -1097
rect 2506 -1159 2540 -1097
rect -2540 -1193 -2444 -1159
rect 2444 -1193 2540 -1159
<< psubdiffcont >>
rect -2444 1159 2444 1193
rect -2540 -1097 -2506 1097
rect 2506 -1097 2540 1097
rect -2444 -1193 2444 -1159
<< poly >>
rect -2380 1091 -2000 1107
rect -2380 1057 -2364 1091
rect -2016 1057 -2000 1091
rect -2380 1019 -2000 1057
rect -1942 1091 -1562 1107
rect -1942 1057 -1926 1091
rect -1578 1057 -1562 1091
rect -1942 1019 -1562 1057
rect -1504 1091 -1124 1107
rect -1504 1057 -1488 1091
rect -1140 1057 -1124 1091
rect -1504 1019 -1124 1057
rect -1066 1091 -686 1107
rect -1066 1057 -1050 1091
rect -702 1057 -686 1091
rect -1066 1019 -686 1057
rect -628 1091 -248 1107
rect -628 1057 -612 1091
rect -264 1057 -248 1091
rect -628 1019 -248 1057
rect -190 1091 190 1107
rect -190 1057 -174 1091
rect 174 1057 190 1091
rect -190 1019 190 1057
rect 248 1091 628 1107
rect 248 1057 264 1091
rect 612 1057 628 1091
rect 248 1019 628 1057
rect 686 1091 1066 1107
rect 686 1057 702 1091
rect 1050 1057 1066 1091
rect 686 1019 1066 1057
rect 1124 1091 1504 1107
rect 1124 1057 1140 1091
rect 1488 1057 1504 1091
rect 1124 1019 1504 1057
rect 1562 1091 1942 1107
rect 1562 1057 1578 1091
rect 1926 1057 1942 1091
rect 1562 1019 1942 1057
rect 2000 1091 2380 1107
rect 2000 1057 2016 1091
rect 2364 1057 2380 1091
rect 2000 1019 2380 1057
rect -2380 -1107 -2000 -1081
rect -1942 -1107 -1562 -1081
rect -1504 -1107 -1124 -1081
rect -1066 -1107 -686 -1081
rect -628 -1107 -248 -1081
rect -190 -1107 190 -1081
rect 248 -1107 628 -1081
rect 686 -1107 1066 -1081
rect 1124 -1107 1504 -1081
rect 1562 -1107 1942 -1081
rect 2000 -1107 2380 -1081
<< polycont >>
rect -2364 1057 -2016 1091
rect -1926 1057 -1578 1091
rect -1488 1057 -1140 1091
rect -1050 1057 -702 1091
rect -612 1057 -264 1091
rect -174 1057 174 1091
rect 264 1057 612 1091
rect 702 1057 1050 1091
rect 1140 1057 1488 1091
rect 1578 1057 1926 1091
rect 2016 1057 2364 1091
<< locali >>
rect -2540 1159 -2444 1193
rect 2444 1159 2540 1193
rect -2540 1097 -2506 1159
rect 2506 1097 2540 1159
rect -2380 1057 -2364 1091
rect -2016 1057 -2000 1091
rect -1942 1057 -1926 1091
rect -1578 1057 -1562 1091
rect -1504 1057 -1488 1091
rect -1140 1057 -1124 1091
rect -1066 1057 -1050 1091
rect -702 1057 -686 1091
rect -628 1057 -612 1091
rect -264 1057 -248 1091
rect -190 1057 -174 1091
rect 174 1057 190 1091
rect 248 1057 264 1091
rect 612 1057 628 1091
rect 686 1057 702 1091
rect 1050 1057 1066 1091
rect 1124 1057 1140 1091
rect 1488 1057 1504 1091
rect 1562 1057 1578 1091
rect 1926 1057 1942 1091
rect 2000 1057 2016 1091
rect 2364 1057 2380 1091
rect -2426 1007 -2392 1023
rect -2426 -1085 -2392 -1069
rect -1988 1007 -1954 1023
rect -1988 -1085 -1954 -1069
rect -1550 1007 -1516 1023
rect -1550 -1085 -1516 -1069
rect -1112 1007 -1078 1023
rect -1112 -1085 -1078 -1069
rect -674 1007 -640 1023
rect -674 -1085 -640 -1069
rect -236 1007 -202 1023
rect -236 -1085 -202 -1069
rect 202 1007 236 1023
rect 202 -1085 236 -1069
rect 640 1007 674 1023
rect 640 -1085 674 -1069
rect 1078 1007 1112 1023
rect 1078 -1085 1112 -1069
rect 1516 1007 1550 1023
rect 1516 -1085 1550 -1069
rect 1954 1007 1988 1023
rect 1954 -1085 1988 -1069
rect 2392 1007 2426 1023
rect 2392 -1085 2426 -1069
rect -2540 -1159 -2506 -1097
rect 2506 -1159 2540 -1097
rect -2540 -1193 -2444 -1159
rect 2444 -1193 2540 -1159
<< viali >>
rect -2364 1057 -2016 1091
rect -1926 1057 -1578 1091
rect -1488 1057 -1140 1091
rect -1050 1057 -702 1091
rect -612 1057 -264 1091
rect -174 1057 174 1091
rect 264 1057 612 1091
rect 702 1057 1050 1091
rect 1140 1057 1488 1091
rect 1578 1057 1926 1091
rect 2016 1057 2364 1091
rect -2426 -1069 -2392 1007
rect -1988 -1069 -1954 1007
rect -1550 -1069 -1516 1007
rect -1112 -1069 -1078 1007
rect -674 -1069 -640 1007
rect -236 -1069 -202 1007
rect 202 -1069 236 1007
rect 640 -1069 674 1007
rect 1078 -1069 1112 1007
rect 1516 -1069 1550 1007
rect 1954 -1069 1988 1007
rect 2392 -1069 2426 1007
<< metal1 >>
rect -2376 1091 -2004 1097
rect -2376 1057 -2364 1091
rect -2016 1057 -2004 1091
rect -2376 1051 -2004 1057
rect -1938 1091 -1566 1097
rect -1938 1057 -1926 1091
rect -1578 1057 -1566 1091
rect -1938 1051 -1566 1057
rect -1500 1091 -1128 1097
rect -1500 1057 -1488 1091
rect -1140 1057 -1128 1091
rect -1500 1051 -1128 1057
rect -1062 1091 -690 1097
rect -1062 1057 -1050 1091
rect -702 1057 -690 1091
rect -1062 1051 -690 1057
rect -624 1091 -252 1097
rect -624 1057 -612 1091
rect -264 1057 -252 1091
rect -624 1051 -252 1057
rect -186 1091 186 1097
rect -186 1057 -174 1091
rect 174 1057 186 1091
rect -186 1051 186 1057
rect 252 1091 624 1097
rect 252 1057 264 1091
rect 612 1057 624 1091
rect 252 1051 624 1057
rect 690 1091 1062 1097
rect 690 1057 702 1091
rect 1050 1057 1062 1091
rect 690 1051 1062 1057
rect 1128 1091 1500 1097
rect 1128 1057 1140 1091
rect 1488 1057 1500 1091
rect 1128 1051 1500 1057
rect 1566 1091 1938 1097
rect 1566 1057 1578 1091
rect 1926 1057 1938 1091
rect 1566 1051 1938 1057
rect 2004 1091 2376 1097
rect 2004 1057 2016 1091
rect 2364 1057 2376 1091
rect 2004 1051 2376 1057
rect -2432 1007 -2386 1019
rect -2432 -1069 -2426 1007
rect -2392 -1069 -2386 1007
rect -2432 -1081 -2386 -1069
rect -1994 1007 -1948 1019
rect -1994 -1069 -1988 1007
rect -1954 -1069 -1948 1007
rect -1994 -1081 -1948 -1069
rect -1556 1007 -1510 1019
rect -1556 -1069 -1550 1007
rect -1516 -1069 -1510 1007
rect -1556 -1081 -1510 -1069
rect -1118 1007 -1072 1019
rect -1118 -1069 -1112 1007
rect -1078 -1069 -1072 1007
rect -1118 -1081 -1072 -1069
rect -680 1007 -634 1019
rect -680 -1069 -674 1007
rect -640 -1069 -634 1007
rect -680 -1081 -634 -1069
rect -242 1007 -196 1019
rect -242 -1069 -236 1007
rect -202 -1069 -196 1007
rect -242 -1081 -196 -1069
rect 196 1007 242 1019
rect 196 -1069 202 1007
rect 236 -1069 242 1007
rect 196 -1081 242 -1069
rect 634 1007 680 1019
rect 634 -1069 640 1007
rect 674 -1069 680 1007
rect 634 -1081 680 -1069
rect 1072 1007 1118 1019
rect 1072 -1069 1078 1007
rect 1112 -1069 1118 1007
rect 1072 -1081 1118 -1069
rect 1510 1007 1556 1019
rect 1510 -1069 1516 1007
rect 1550 -1069 1556 1007
rect 1510 -1081 1556 -1069
rect 1948 1007 1994 1019
rect 1948 -1069 1954 1007
rect 1988 -1069 1994 1007
rect 1948 -1081 1994 -1069
rect 2386 1007 2432 1019
rect 2386 -1069 2392 1007
rect 2426 -1069 2432 1007
rect 2386 -1081 2432 -1069
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2523 -1176 2523 1176
string parameters w 10.5 l 1.9 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
