magic
tech sky130A
magscale 1 2
timestamp 1615920820
<< nwell >>
rect -4223 -764 4223 798
<< pmos >>
rect -4129 -664 -3989 736
rect -3931 -664 -3791 736
rect -3733 -664 -3593 736
rect -3535 -664 -3395 736
rect -3337 -664 -3197 736
rect -3139 -664 -2999 736
rect -2941 -664 -2801 736
rect -2743 -664 -2603 736
rect -2545 -664 -2405 736
rect -2347 -664 -2207 736
rect -2149 -664 -2009 736
rect -1951 -664 -1811 736
rect -1753 -664 -1613 736
rect -1555 -664 -1415 736
rect -1357 -664 -1217 736
rect -1159 -664 -1019 736
rect -961 -664 -821 736
rect -763 -664 -623 736
rect -565 -664 -425 736
rect -367 -664 -227 736
rect -169 -664 -29 736
rect 29 -664 169 736
rect 227 -664 367 736
rect 425 -664 565 736
rect 623 -664 763 736
rect 821 -664 961 736
rect 1019 -664 1159 736
rect 1217 -664 1357 736
rect 1415 -664 1555 736
rect 1613 -664 1753 736
rect 1811 -664 1951 736
rect 2009 -664 2149 736
rect 2207 -664 2347 736
rect 2405 -664 2545 736
rect 2603 -664 2743 736
rect 2801 -664 2941 736
rect 2999 -664 3139 736
rect 3197 -664 3337 736
rect 3395 -664 3535 736
rect 3593 -664 3733 736
rect 3791 -664 3931 736
rect 3989 -664 4129 736
<< pdiff >>
rect -4187 724 -4129 736
rect -4187 -652 -4175 724
rect -4141 -652 -4129 724
rect -4187 -664 -4129 -652
rect -3989 724 -3931 736
rect -3989 -652 -3977 724
rect -3943 -652 -3931 724
rect -3989 -664 -3931 -652
rect -3791 724 -3733 736
rect -3791 -652 -3779 724
rect -3745 -652 -3733 724
rect -3791 -664 -3733 -652
rect -3593 724 -3535 736
rect -3593 -652 -3581 724
rect -3547 -652 -3535 724
rect -3593 -664 -3535 -652
rect -3395 724 -3337 736
rect -3395 -652 -3383 724
rect -3349 -652 -3337 724
rect -3395 -664 -3337 -652
rect -3197 724 -3139 736
rect -3197 -652 -3185 724
rect -3151 -652 -3139 724
rect -3197 -664 -3139 -652
rect -2999 724 -2941 736
rect -2999 -652 -2987 724
rect -2953 -652 -2941 724
rect -2999 -664 -2941 -652
rect -2801 724 -2743 736
rect -2801 -652 -2789 724
rect -2755 -652 -2743 724
rect -2801 -664 -2743 -652
rect -2603 724 -2545 736
rect -2603 -652 -2591 724
rect -2557 -652 -2545 724
rect -2603 -664 -2545 -652
rect -2405 724 -2347 736
rect -2405 -652 -2393 724
rect -2359 -652 -2347 724
rect -2405 -664 -2347 -652
rect -2207 724 -2149 736
rect -2207 -652 -2195 724
rect -2161 -652 -2149 724
rect -2207 -664 -2149 -652
rect -2009 724 -1951 736
rect -2009 -652 -1997 724
rect -1963 -652 -1951 724
rect -2009 -664 -1951 -652
rect -1811 724 -1753 736
rect -1811 -652 -1799 724
rect -1765 -652 -1753 724
rect -1811 -664 -1753 -652
rect -1613 724 -1555 736
rect -1613 -652 -1601 724
rect -1567 -652 -1555 724
rect -1613 -664 -1555 -652
rect -1415 724 -1357 736
rect -1415 -652 -1403 724
rect -1369 -652 -1357 724
rect -1415 -664 -1357 -652
rect -1217 724 -1159 736
rect -1217 -652 -1205 724
rect -1171 -652 -1159 724
rect -1217 -664 -1159 -652
rect -1019 724 -961 736
rect -1019 -652 -1007 724
rect -973 -652 -961 724
rect -1019 -664 -961 -652
rect -821 724 -763 736
rect -821 -652 -809 724
rect -775 -652 -763 724
rect -821 -664 -763 -652
rect -623 724 -565 736
rect -623 -652 -611 724
rect -577 -652 -565 724
rect -623 -664 -565 -652
rect -425 724 -367 736
rect -425 -652 -413 724
rect -379 -652 -367 724
rect -425 -664 -367 -652
rect -227 724 -169 736
rect -227 -652 -215 724
rect -181 -652 -169 724
rect -227 -664 -169 -652
rect -29 724 29 736
rect -29 -652 -17 724
rect 17 -652 29 724
rect -29 -664 29 -652
rect 169 724 227 736
rect 169 -652 181 724
rect 215 -652 227 724
rect 169 -664 227 -652
rect 367 724 425 736
rect 367 -652 379 724
rect 413 -652 425 724
rect 367 -664 425 -652
rect 565 724 623 736
rect 565 -652 577 724
rect 611 -652 623 724
rect 565 -664 623 -652
rect 763 724 821 736
rect 763 -652 775 724
rect 809 -652 821 724
rect 763 -664 821 -652
rect 961 724 1019 736
rect 961 -652 973 724
rect 1007 -652 1019 724
rect 961 -664 1019 -652
rect 1159 724 1217 736
rect 1159 -652 1171 724
rect 1205 -652 1217 724
rect 1159 -664 1217 -652
rect 1357 724 1415 736
rect 1357 -652 1369 724
rect 1403 -652 1415 724
rect 1357 -664 1415 -652
rect 1555 724 1613 736
rect 1555 -652 1567 724
rect 1601 -652 1613 724
rect 1555 -664 1613 -652
rect 1753 724 1811 736
rect 1753 -652 1765 724
rect 1799 -652 1811 724
rect 1753 -664 1811 -652
rect 1951 724 2009 736
rect 1951 -652 1963 724
rect 1997 -652 2009 724
rect 1951 -664 2009 -652
rect 2149 724 2207 736
rect 2149 -652 2161 724
rect 2195 -652 2207 724
rect 2149 -664 2207 -652
rect 2347 724 2405 736
rect 2347 -652 2359 724
rect 2393 -652 2405 724
rect 2347 -664 2405 -652
rect 2545 724 2603 736
rect 2545 -652 2557 724
rect 2591 -652 2603 724
rect 2545 -664 2603 -652
rect 2743 724 2801 736
rect 2743 -652 2755 724
rect 2789 -652 2801 724
rect 2743 -664 2801 -652
rect 2941 724 2999 736
rect 2941 -652 2953 724
rect 2987 -652 2999 724
rect 2941 -664 2999 -652
rect 3139 724 3197 736
rect 3139 -652 3151 724
rect 3185 -652 3197 724
rect 3139 -664 3197 -652
rect 3337 724 3395 736
rect 3337 -652 3349 724
rect 3383 -652 3395 724
rect 3337 -664 3395 -652
rect 3535 724 3593 736
rect 3535 -652 3547 724
rect 3581 -652 3593 724
rect 3535 -664 3593 -652
rect 3733 724 3791 736
rect 3733 -652 3745 724
rect 3779 -652 3791 724
rect 3733 -664 3791 -652
rect 3931 724 3989 736
rect 3931 -652 3943 724
rect 3977 -652 3989 724
rect 3931 -664 3989 -652
rect 4129 724 4187 736
rect 4129 -652 4141 724
rect 4175 -652 4187 724
rect 4129 -664 4187 -652
<< pdiffc >>
rect -4175 -652 -4141 724
rect -3977 -652 -3943 724
rect -3779 -652 -3745 724
rect -3581 -652 -3547 724
rect -3383 -652 -3349 724
rect -3185 -652 -3151 724
rect -2987 -652 -2953 724
rect -2789 -652 -2755 724
rect -2591 -652 -2557 724
rect -2393 -652 -2359 724
rect -2195 -652 -2161 724
rect -1997 -652 -1963 724
rect -1799 -652 -1765 724
rect -1601 -652 -1567 724
rect -1403 -652 -1369 724
rect -1205 -652 -1171 724
rect -1007 -652 -973 724
rect -809 -652 -775 724
rect -611 -652 -577 724
rect -413 -652 -379 724
rect -215 -652 -181 724
rect -17 -652 17 724
rect 181 -652 215 724
rect 379 -652 413 724
rect 577 -652 611 724
rect 775 -652 809 724
rect 973 -652 1007 724
rect 1171 -652 1205 724
rect 1369 -652 1403 724
rect 1567 -652 1601 724
rect 1765 -652 1799 724
rect 1963 -652 1997 724
rect 2161 -652 2195 724
rect 2359 -652 2393 724
rect 2557 -652 2591 724
rect 2755 -652 2789 724
rect 2953 -652 2987 724
rect 3151 -652 3185 724
rect 3349 -652 3383 724
rect 3547 -652 3581 724
rect 3745 -652 3779 724
rect 3943 -652 3977 724
rect 4141 -652 4175 724
<< poly >>
rect -4129 736 -3989 762
rect -3931 736 -3791 762
rect -3733 736 -3593 762
rect -3535 736 -3395 762
rect -3337 736 -3197 762
rect -3139 736 -2999 762
rect -2941 736 -2801 762
rect -2743 736 -2603 762
rect -2545 736 -2405 762
rect -2347 736 -2207 762
rect -2149 736 -2009 762
rect -1951 736 -1811 762
rect -1753 736 -1613 762
rect -1555 736 -1415 762
rect -1357 736 -1217 762
rect -1159 736 -1019 762
rect -961 736 -821 762
rect -763 736 -623 762
rect -565 736 -425 762
rect -367 736 -227 762
rect -169 736 -29 762
rect 29 736 169 762
rect 227 736 367 762
rect 425 736 565 762
rect 623 736 763 762
rect 821 736 961 762
rect 1019 736 1159 762
rect 1217 736 1357 762
rect 1415 736 1555 762
rect 1613 736 1753 762
rect 1811 736 1951 762
rect 2009 736 2149 762
rect 2207 736 2347 762
rect 2405 736 2545 762
rect 2603 736 2743 762
rect 2801 736 2941 762
rect 2999 736 3139 762
rect 3197 736 3337 762
rect 3395 736 3535 762
rect 3593 736 3733 762
rect 3791 736 3931 762
rect 3989 736 4129 762
rect -4129 -711 -3989 -664
rect -4129 -745 -4113 -711
rect -4005 -745 -3989 -711
rect -4129 -761 -3989 -745
rect -3931 -711 -3791 -664
rect -3931 -745 -3915 -711
rect -3807 -745 -3791 -711
rect -3931 -761 -3791 -745
rect -3733 -711 -3593 -664
rect -3733 -745 -3717 -711
rect -3609 -745 -3593 -711
rect -3733 -761 -3593 -745
rect -3535 -711 -3395 -664
rect -3535 -745 -3519 -711
rect -3411 -745 -3395 -711
rect -3535 -761 -3395 -745
rect -3337 -711 -3197 -664
rect -3337 -745 -3321 -711
rect -3213 -745 -3197 -711
rect -3337 -761 -3197 -745
rect -3139 -711 -2999 -664
rect -3139 -745 -3123 -711
rect -3015 -745 -2999 -711
rect -3139 -761 -2999 -745
rect -2941 -711 -2801 -664
rect -2941 -745 -2925 -711
rect -2817 -745 -2801 -711
rect -2941 -761 -2801 -745
rect -2743 -711 -2603 -664
rect -2743 -745 -2727 -711
rect -2619 -745 -2603 -711
rect -2743 -761 -2603 -745
rect -2545 -711 -2405 -664
rect -2545 -745 -2529 -711
rect -2421 -745 -2405 -711
rect -2545 -761 -2405 -745
rect -2347 -711 -2207 -664
rect -2347 -745 -2331 -711
rect -2223 -745 -2207 -711
rect -2347 -761 -2207 -745
rect -2149 -711 -2009 -664
rect -2149 -745 -2133 -711
rect -2025 -745 -2009 -711
rect -2149 -761 -2009 -745
rect -1951 -711 -1811 -664
rect -1951 -745 -1935 -711
rect -1827 -745 -1811 -711
rect -1951 -761 -1811 -745
rect -1753 -711 -1613 -664
rect -1753 -745 -1737 -711
rect -1629 -745 -1613 -711
rect -1753 -761 -1613 -745
rect -1555 -711 -1415 -664
rect -1555 -745 -1539 -711
rect -1431 -745 -1415 -711
rect -1555 -761 -1415 -745
rect -1357 -711 -1217 -664
rect -1357 -745 -1341 -711
rect -1233 -745 -1217 -711
rect -1357 -761 -1217 -745
rect -1159 -711 -1019 -664
rect -1159 -745 -1143 -711
rect -1035 -745 -1019 -711
rect -1159 -761 -1019 -745
rect -961 -711 -821 -664
rect -961 -745 -945 -711
rect -837 -745 -821 -711
rect -961 -761 -821 -745
rect -763 -711 -623 -664
rect -763 -745 -747 -711
rect -639 -745 -623 -711
rect -763 -761 -623 -745
rect -565 -711 -425 -664
rect -565 -745 -549 -711
rect -441 -745 -425 -711
rect -565 -761 -425 -745
rect -367 -711 -227 -664
rect -367 -745 -351 -711
rect -243 -745 -227 -711
rect -367 -761 -227 -745
rect -169 -711 -29 -664
rect -169 -745 -153 -711
rect -45 -745 -29 -711
rect -169 -761 -29 -745
rect 29 -711 169 -664
rect 29 -745 45 -711
rect 153 -745 169 -711
rect 29 -761 169 -745
rect 227 -711 367 -664
rect 227 -745 243 -711
rect 351 -745 367 -711
rect 227 -761 367 -745
rect 425 -711 565 -664
rect 425 -745 441 -711
rect 549 -745 565 -711
rect 425 -761 565 -745
rect 623 -711 763 -664
rect 623 -745 639 -711
rect 747 -745 763 -711
rect 623 -761 763 -745
rect 821 -711 961 -664
rect 821 -745 837 -711
rect 945 -745 961 -711
rect 821 -761 961 -745
rect 1019 -711 1159 -664
rect 1019 -745 1035 -711
rect 1143 -745 1159 -711
rect 1019 -761 1159 -745
rect 1217 -711 1357 -664
rect 1217 -745 1233 -711
rect 1341 -745 1357 -711
rect 1217 -761 1357 -745
rect 1415 -711 1555 -664
rect 1415 -745 1431 -711
rect 1539 -745 1555 -711
rect 1415 -761 1555 -745
rect 1613 -711 1753 -664
rect 1613 -745 1629 -711
rect 1737 -745 1753 -711
rect 1613 -761 1753 -745
rect 1811 -711 1951 -664
rect 1811 -745 1827 -711
rect 1935 -745 1951 -711
rect 1811 -761 1951 -745
rect 2009 -711 2149 -664
rect 2009 -745 2025 -711
rect 2133 -745 2149 -711
rect 2009 -761 2149 -745
rect 2207 -711 2347 -664
rect 2207 -745 2223 -711
rect 2331 -745 2347 -711
rect 2207 -761 2347 -745
rect 2405 -711 2545 -664
rect 2405 -745 2421 -711
rect 2529 -745 2545 -711
rect 2405 -761 2545 -745
rect 2603 -711 2743 -664
rect 2603 -745 2619 -711
rect 2727 -745 2743 -711
rect 2603 -761 2743 -745
rect 2801 -711 2941 -664
rect 2801 -745 2817 -711
rect 2925 -745 2941 -711
rect 2801 -761 2941 -745
rect 2999 -711 3139 -664
rect 2999 -745 3015 -711
rect 3123 -745 3139 -711
rect 2999 -761 3139 -745
rect 3197 -711 3337 -664
rect 3197 -745 3213 -711
rect 3321 -745 3337 -711
rect 3197 -761 3337 -745
rect 3395 -711 3535 -664
rect 3395 -745 3411 -711
rect 3519 -745 3535 -711
rect 3395 -761 3535 -745
rect 3593 -711 3733 -664
rect 3593 -745 3609 -711
rect 3717 -745 3733 -711
rect 3593 -761 3733 -745
rect 3791 -711 3931 -664
rect 3791 -745 3807 -711
rect 3915 -745 3931 -711
rect 3791 -761 3931 -745
rect 3989 -711 4129 -664
rect 3989 -745 4005 -711
rect 4113 -745 4129 -711
rect 3989 -761 4129 -745
<< polycont >>
rect -4113 -745 -4005 -711
rect -3915 -745 -3807 -711
rect -3717 -745 -3609 -711
rect -3519 -745 -3411 -711
rect -3321 -745 -3213 -711
rect -3123 -745 -3015 -711
rect -2925 -745 -2817 -711
rect -2727 -745 -2619 -711
rect -2529 -745 -2421 -711
rect -2331 -745 -2223 -711
rect -2133 -745 -2025 -711
rect -1935 -745 -1827 -711
rect -1737 -745 -1629 -711
rect -1539 -745 -1431 -711
rect -1341 -745 -1233 -711
rect -1143 -745 -1035 -711
rect -945 -745 -837 -711
rect -747 -745 -639 -711
rect -549 -745 -441 -711
rect -351 -745 -243 -711
rect -153 -745 -45 -711
rect 45 -745 153 -711
rect 243 -745 351 -711
rect 441 -745 549 -711
rect 639 -745 747 -711
rect 837 -745 945 -711
rect 1035 -745 1143 -711
rect 1233 -745 1341 -711
rect 1431 -745 1539 -711
rect 1629 -745 1737 -711
rect 1827 -745 1935 -711
rect 2025 -745 2133 -711
rect 2223 -745 2331 -711
rect 2421 -745 2529 -711
rect 2619 -745 2727 -711
rect 2817 -745 2925 -711
rect 3015 -745 3123 -711
rect 3213 -745 3321 -711
rect 3411 -745 3519 -711
rect 3609 -745 3717 -711
rect 3807 -745 3915 -711
rect 4005 -745 4113 -711
<< locali >>
rect -4175 724 -4141 740
rect -4175 -668 -4141 -652
rect -3977 724 -3943 740
rect -3977 -668 -3943 -652
rect -3779 724 -3745 740
rect -3779 -668 -3745 -652
rect -3581 724 -3547 740
rect -3581 -668 -3547 -652
rect -3383 724 -3349 740
rect -3383 -668 -3349 -652
rect -3185 724 -3151 740
rect -3185 -668 -3151 -652
rect -2987 724 -2953 740
rect -2987 -668 -2953 -652
rect -2789 724 -2755 740
rect -2789 -668 -2755 -652
rect -2591 724 -2557 740
rect -2591 -668 -2557 -652
rect -2393 724 -2359 740
rect -2393 -668 -2359 -652
rect -2195 724 -2161 740
rect -2195 -668 -2161 -652
rect -1997 724 -1963 740
rect -1997 -668 -1963 -652
rect -1799 724 -1765 740
rect -1799 -668 -1765 -652
rect -1601 724 -1567 740
rect -1601 -668 -1567 -652
rect -1403 724 -1369 740
rect -1403 -668 -1369 -652
rect -1205 724 -1171 740
rect -1205 -668 -1171 -652
rect -1007 724 -973 740
rect -1007 -668 -973 -652
rect -809 724 -775 740
rect -809 -668 -775 -652
rect -611 724 -577 740
rect -611 -668 -577 -652
rect -413 724 -379 740
rect -413 -668 -379 -652
rect -215 724 -181 740
rect -215 -668 -181 -652
rect -17 724 17 740
rect -17 -668 17 -652
rect 181 724 215 740
rect 181 -668 215 -652
rect 379 724 413 740
rect 379 -668 413 -652
rect 577 724 611 740
rect 577 -668 611 -652
rect 775 724 809 740
rect 775 -668 809 -652
rect 973 724 1007 740
rect 973 -668 1007 -652
rect 1171 724 1205 740
rect 1171 -668 1205 -652
rect 1369 724 1403 740
rect 1369 -668 1403 -652
rect 1567 724 1601 740
rect 1567 -668 1601 -652
rect 1765 724 1799 740
rect 1765 -668 1799 -652
rect 1963 724 1997 740
rect 1963 -668 1997 -652
rect 2161 724 2195 740
rect 2161 -668 2195 -652
rect 2359 724 2393 740
rect 2359 -668 2393 -652
rect 2557 724 2591 740
rect 2557 -668 2591 -652
rect 2755 724 2789 740
rect 2755 -668 2789 -652
rect 2953 724 2987 740
rect 2953 -668 2987 -652
rect 3151 724 3185 740
rect 3151 -668 3185 -652
rect 3349 724 3383 740
rect 3349 -668 3383 -652
rect 3547 724 3581 740
rect 3547 -668 3581 -652
rect 3745 724 3779 740
rect 3745 -668 3779 -652
rect 3943 724 3977 740
rect 3943 -668 3977 -652
rect 4141 724 4175 740
rect 4141 -668 4175 -652
rect -4129 -745 -4113 -711
rect -4005 -745 -3989 -711
rect -3931 -745 -3915 -711
rect -3807 -745 -3791 -711
rect -3733 -745 -3717 -711
rect -3609 -745 -3593 -711
rect -3535 -745 -3519 -711
rect -3411 -745 -3395 -711
rect -3337 -745 -3321 -711
rect -3213 -745 -3197 -711
rect -3139 -745 -3123 -711
rect -3015 -745 -2999 -711
rect -2941 -745 -2925 -711
rect -2817 -745 -2801 -711
rect -2743 -745 -2727 -711
rect -2619 -745 -2603 -711
rect -2545 -745 -2529 -711
rect -2421 -745 -2405 -711
rect -2347 -745 -2331 -711
rect -2223 -745 -2207 -711
rect -2149 -745 -2133 -711
rect -2025 -745 -2009 -711
rect -1951 -745 -1935 -711
rect -1827 -745 -1811 -711
rect -1753 -745 -1737 -711
rect -1629 -745 -1613 -711
rect -1555 -745 -1539 -711
rect -1431 -745 -1415 -711
rect -1357 -745 -1341 -711
rect -1233 -745 -1217 -711
rect -1159 -745 -1143 -711
rect -1035 -745 -1019 -711
rect -961 -745 -945 -711
rect -837 -745 -821 -711
rect -763 -745 -747 -711
rect -639 -745 -623 -711
rect -565 -745 -549 -711
rect -441 -745 -425 -711
rect -367 -745 -351 -711
rect -243 -745 -227 -711
rect -169 -745 -153 -711
rect -45 -745 -29 -711
rect 29 -745 45 -711
rect 153 -745 169 -711
rect 227 -745 243 -711
rect 351 -745 367 -711
rect 425 -745 441 -711
rect 549 -745 565 -711
rect 623 -745 639 -711
rect 747 -745 763 -711
rect 821 -745 837 -711
rect 945 -745 961 -711
rect 1019 -745 1035 -711
rect 1143 -745 1159 -711
rect 1217 -745 1233 -711
rect 1341 -745 1357 -711
rect 1415 -745 1431 -711
rect 1539 -745 1555 -711
rect 1613 -745 1629 -711
rect 1737 -745 1753 -711
rect 1811 -745 1827 -711
rect 1935 -745 1951 -711
rect 2009 -745 2025 -711
rect 2133 -745 2149 -711
rect 2207 -745 2223 -711
rect 2331 -745 2347 -711
rect 2405 -745 2421 -711
rect 2529 -745 2545 -711
rect 2603 -745 2619 -711
rect 2727 -745 2743 -711
rect 2801 -745 2817 -711
rect 2925 -745 2941 -711
rect 2999 -745 3015 -711
rect 3123 -745 3139 -711
rect 3197 -745 3213 -711
rect 3321 -745 3337 -711
rect 3395 -745 3411 -711
rect 3519 -745 3535 -711
rect 3593 -745 3609 -711
rect 3717 -745 3733 -711
rect 3791 -745 3807 -711
rect 3915 -745 3931 -711
rect 3989 -745 4005 -711
rect 4113 -745 4129 -711
<< viali >>
rect -4175 -652 -4141 724
rect -3977 -652 -3943 724
rect -3779 -652 -3745 724
rect -3581 -652 -3547 724
rect -3383 -652 -3349 724
rect -3185 -652 -3151 724
rect -2987 -652 -2953 724
rect -2789 -652 -2755 724
rect -2591 -652 -2557 724
rect -2393 -652 -2359 724
rect -2195 -652 -2161 724
rect -1997 -652 -1963 724
rect -1799 -652 -1765 724
rect -1601 -652 -1567 724
rect -1403 -652 -1369 724
rect -1205 -652 -1171 724
rect -1007 -652 -973 724
rect -809 -652 -775 724
rect -611 -652 -577 724
rect -413 -652 -379 724
rect -215 -652 -181 724
rect -17 -652 17 724
rect 181 -652 215 724
rect 379 -652 413 724
rect 577 -652 611 724
rect 775 -652 809 724
rect 973 -652 1007 724
rect 1171 -652 1205 724
rect 1369 -652 1403 724
rect 1567 -652 1601 724
rect 1765 -652 1799 724
rect 1963 -652 1997 724
rect 2161 -652 2195 724
rect 2359 -652 2393 724
rect 2557 -652 2591 724
rect 2755 -652 2789 724
rect 2953 -652 2987 724
rect 3151 -652 3185 724
rect 3349 -652 3383 724
rect 3547 -652 3581 724
rect 3745 -652 3779 724
rect 3943 -652 3977 724
rect 4141 -652 4175 724
rect -4113 -745 -4005 -711
rect -3915 -745 -3807 -711
rect -3717 -745 -3609 -711
rect -3519 -745 -3411 -711
rect -3321 -745 -3213 -711
rect -3123 -745 -3015 -711
rect -2925 -745 -2817 -711
rect -2727 -745 -2619 -711
rect -2529 -745 -2421 -711
rect -2331 -745 -2223 -711
rect -2133 -745 -2025 -711
rect -1935 -745 -1827 -711
rect -1737 -745 -1629 -711
rect -1539 -745 -1431 -711
rect -1341 -745 -1233 -711
rect -1143 -745 -1035 -711
rect -945 -745 -837 -711
rect -747 -745 -639 -711
rect -549 -745 -441 -711
rect -351 -745 -243 -711
rect -153 -745 -45 -711
rect 45 -745 153 -711
rect 243 -745 351 -711
rect 441 -745 549 -711
rect 639 -745 747 -711
rect 837 -745 945 -711
rect 1035 -745 1143 -711
rect 1233 -745 1341 -711
rect 1431 -745 1539 -711
rect 1629 -745 1737 -711
rect 1827 -745 1935 -711
rect 2025 -745 2133 -711
rect 2223 -745 2331 -711
rect 2421 -745 2529 -711
rect 2619 -745 2727 -711
rect 2817 -745 2925 -711
rect 3015 -745 3123 -711
rect 3213 -745 3321 -711
rect 3411 -745 3519 -711
rect 3609 -745 3717 -711
rect 3807 -745 3915 -711
rect 4005 -745 4113 -711
<< metal1 >>
rect -4181 724 -4135 736
rect -4181 -652 -4175 724
rect -4141 -652 -4135 724
rect -4181 -664 -4135 -652
rect -3983 724 -3937 736
rect -3983 -652 -3977 724
rect -3943 -652 -3937 724
rect -3983 -664 -3937 -652
rect -3785 724 -3739 736
rect -3785 -652 -3779 724
rect -3745 -652 -3739 724
rect -3785 -664 -3739 -652
rect -3587 724 -3541 736
rect -3587 -652 -3581 724
rect -3547 -652 -3541 724
rect -3587 -664 -3541 -652
rect -3389 724 -3343 736
rect -3389 -652 -3383 724
rect -3349 -652 -3343 724
rect -3389 -664 -3343 -652
rect -3191 724 -3145 736
rect -3191 -652 -3185 724
rect -3151 -652 -3145 724
rect -3191 -664 -3145 -652
rect -2993 724 -2947 736
rect -2993 -652 -2987 724
rect -2953 -652 -2947 724
rect -2993 -664 -2947 -652
rect -2795 724 -2749 736
rect -2795 -652 -2789 724
rect -2755 -652 -2749 724
rect -2795 -664 -2749 -652
rect -2597 724 -2551 736
rect -2597 -652 -2591 724
rect -2557 -652 -2551 724
rect -2597 -664 -2551 -652
rect -2399 724 -2353 736
rect -2399 -652 -2393 724
rect -2359 -652 -2353 724
rect -2399 -664 -2353 -652
rect -2201 724 -2155 736
rect -2201 -652 -2195 724
rect -2161 -652 -2155 724
rect -2201 -664 -2155 -652
rect -2003 724 -1957 736
rect -2003 -652 -1997 724
rect -1963 -652 -1957 724
rect -2003 -664 -1957 -652
rect -1805 724 -1759 736
rect -1805 -652 -1799 724
rect -1765 -652 -1759 724
rect -1805 -664 -1759 -652
rect -1607 724 -1561 736
rect -1607 -652 -1601 724
rect -1567 -652 -1561 724
rect -1607 -664 -1561 -652
rect -1409 724 -1363 736
rect -1409 -652 -1403 724
rect -1369 -652 -1363 724
rect -1409 -664 -1363 -652
rect -1211 724 -1165 736
rect -1211 -652 -1205 724
rect -1171 -652 -1165 724
rect -1211 -664 -1165 -652
rect -1013 724 -967 736
rect -1013 -652 -1007 724
rect -973 -652 -967 724
rect -1013 -664 -967 -652
rect -815 724 -769 736
rect -815 -652 -809 724
rect -775 -652 -769 724
rect -815 -664 -769 -652
rect -617 724 -571 736
rect -617 -652 -611 724
rect -577 -652 -571 724
rect -617 -664 -571 -652
rect -419 724 -373 736
rect -419 -652 -413 724
rect -379 -652 -373 724
rect -419 -664 -373 -652
rect -221 724 -175 736
rect -221 -652 -215 724
rect -181 -652 -175 724
rect -221 -664 -175 -652
rect -23 724 23 736
rect -23 -652 -17 724
rect 17 -652 23 724
rect -23 -664 23 -652
rect 175 724 221 736
rect 175 -652 181 724
rect 215 -652 221 724
rect 175 -664 221 -652
rect 373 724 419 736
rect 373 -652 379 724
rect 413 -652 419 724
rect 373 -664 419 -652
rect 571 724 617 736
rect 571 -652 577 724
rect 611 -652 617 724
rect 571 -664 617 -652
rect 769 724 815 736
rect 769 -652 775 724
rect 809 -652 815 724
rect 769 -664 815 -652
rect 967 724 1013 736
rect 967 -652 973 724
rect 1007 -652 1013 724
rect 967 -664 1013 -652
rect 1165 724 1211 736
rect 1165 -652 1171 724
rect 1205 -652 1211 724
rect 1165 -664 1211 -652
rect 1363 724 1409 736
rect 1363 -652 1369 724
rect 1403 -652 1409 724
rect 1363 -664 1409 -652
rect 1561 724 1607 736
rect 1561 -652 1567 724
rect 1601 -652 1607 724
rect 1561 -664 1607 -652
rect 1759 724 1805 736
rect 1759 -652 1765 724
rect 1799 -652 1805 724
rect 1759 -664 1805 -652
rect 1957 724 2003 736
rect 1957 -652 1963 724
rect 1997 -652 2003 724
rect 1957 -664 2003 -652
rect 2155 724 2201 736
rect 2155 -652 2161 724
rect 2195 -652 2201 724
rect 2155 -664 2201 -652
rect 2353 724 2399 736
rect 2353 -652 2359 724
rect 2393 -652 2399 724
rect 2353 -664 2399 -652
rect 2551 724 2597 736
rect 2551 -652 2557 724
rect 2591 -652 2597 724
rect 2551 -664 2597 -652
rect 2749 724 2795 736
rect 2749 -652 2755 724
rect 2789 -652 2795 724
rect 2749 -664 2795 -652
rect 2947 724 2993 736
rect 2947 -652 2953 724
rect 2987 -652 2993 724
rect 2947 -664 2993 -652
rect 3145 724 3191 736
rect 3145 -652 3151 724
rect 3185 -652 3191 724
rect 3145 -664 3191 -652
rect 3343 724 3389 736
rect 3343 -652 3349 724
rect 3383 -652 3389 724
rect 3343 -664 3389 -652
rect 3541 724 3587 736
rect 3541 -652 3547 724
rect 3581 -652 3587 724
rect 3541 -664 3587 -652
rect 3739 724 3785 736
rect 3739 -652 3745 724
rect 3779 -652 3785 724
rect 3739 -664 3785 -652
rect 3937 724 3983 736
rect 3937 -652 3943 724
rect 3977 -652 3983 724
rect 3937 -664 3983 -652
rect 4135 724 4181 736
rect 4135 -652 4141 724
rect 4175 -652 4181 724
rect 4135 -664 4181 -652
rect -4125 -711 -3993 -705
rect -4125 -745 -4113 -711
rect -4005 -745 -3993 -711
rect -4125 -751 -3993 -745
rect -3927 -711 -3795 -705
rect -3927 -745 -3915 -711
rect -3807 -745 -3795 -711
rect -3927 -751 -3795 -745
rect -3729 -711 -3597 -705
rect -3729 -745 -3717 -711
rect -3609 -745 -3597 -711
rect -3729 -751 -3597 -745
rect -3531 -711 -3399 -705
rect -3531 -745 -3519 -711
rect -3411 -745 -3399 -711
rect -3531 -751 -3399 -745
rect -3333 -711 -3201 -705
rect -3333 -745 -3321 -711
rect -3213 -745 -3201 -711
rect -3333 -751 -3201 -745
rect -3135 -711 -3003 -705
rect -3135 -745 -3123 -711
rect -3015 -745 -3003 -711
rect -3135 -751 -3003 -745
rect -2937 -711 -2805 -705
rect -2937 -745 -2925 -711
rect -2817 -745 -2805 -711
rect -2937 -751 -2805 -745
rect -2739 -711 -2607 -705
rect -2739 -745 -2727 -711
rect -2619 -745 -2607 -711
rect -2739 -751 -2607 -745
rect -2541 -711 -2409 -705
rect -2541 -745 -2529 -711
rect -2421 -745 -2409 -711
rect -2541 -751 -2409 -745
rect -2343 -711 -2211 -705
rect -2343 -745 -2331 -711
rect -2223 -745 -2211 -711
rect -2343 -751 -2211 -745
rect -2145 -711 -2013 -705
rect -2145 -745 -2133 -711
rect -2025 -745 -2013 -711
rect -2145 -751 -2013 -745
rect -1947 -711 -1815 -705
rect -1947 -745 -1935 -711
rect -1827 -745 -1815 -711
rect -1947 -751 -1815 -745
rect -1749 -711 -1617 -705
rect -1749 -745 -1737 -711
rect -1629 -745 -1617 -711
rect -1749 -751 -1617 -745
rect -1551 -711 -1419 -705
rect -1551 -745 -1539 -711
rect -1431 -745 -1419 -711
rect -1551 -751 -1419 -745
rect -1353 -711 -1221 -705
rect -1353 -745 -1341 -711
rect -1233 -745 -1221 -711
rect -1353 -751 -1221 -745
rect -1155 -711 -1023 -705
rect -1155 -745 -1143 -711
rect -1035 -745 -1023 -711
rect -1155 -751 -1023 -745
rect -957 -711 -825 -705
rect -957 -745 -945 -711
rect -837 -745 -825 -711
rect -957 -751 -825 -745
rect -759 -711 -627 -705
rect -759 -745 -747 -711
rect -639 -745 -627 -711
rect -759 -751 -627 -745
rect -561 -711 -429 -705
rect -561 -745 -549 -711
rect -441 -745 -429 -711
rect -561 -751 -429 -745
rect -363 -711 -231 -705
rect -363 -745 -351 -711
rect -243 -745 -231 -711
rect -363 -751 -231 -745
rect -165 -711 -33 -705
rect -165 -745 -153 -711
rect -45 -745 -33 -711
rect -165 -751 -33 -745
rect 33 -711 165 -705
rect 33 -745 45 -711
rect 153 -745 165 -711
rect 33 -751 165 -745
rect 231 -711 363 -705
rect 231 -745 243 -711
rect 351 -745 363 -711
rect 231 -751 363 -745
rect 429 -711 561 -705
rect 429 -745 441 -711
rect 549 -745 561 -711
rect 429 -751 561 -745
rect 627 -711 759 -705
rect 627 -745 639 -711
rect 747 -745 759 -711
rect 627 -751 759 -745
rect 825 -711 957 -705
rect 825 -745 837 -711
rect 945 -745 957 -711
rect 825 -751 957 -745
rect 1023 -711 1155 -705
rect 1023 -745 1035 -711
rect 1143 -745 1155 -711
rect 1023 -751 1155 -745
rect 1221 -711 1353 -705
rect 1221 -745 1233 -711
rect 1341 -745 1353 -711
rect 1221 -751 1353 -745
rect 1419 -711 1551 -705
rect 1419 -745 1431 -711
rect 1539 -745 1551 -711
rect 1419 -751 1551 -745
rect 1617 -711 1749 -705
rect 1617 -745 1629 -711
rect 1737 -745 1749 -711
rect 1617 -751 1749 -745
rect 1815 -711 1947 -705
rect 1815 -745 1827 -711
rect 1935 -745 1947 -711
rect 1815 -751 1947 -745
rect 2013 -711 2145 -705
rect 2013 -745 2025 -711
rect 2133 -745 2145 -711
rect 2013 -751 2145 -745
rect 2211 -711 2343 -705
rect 2211 -745 2223 -711
rect 2331 -745 2343 -711
rect 2211 -751 2343 -745
rect 2409 -711 2541 -705
rect 2409 -745 2421 -711
rect 2529 -745 2541 -711
rect 2409 -751 2541 -745
rect 2607 -711 2739 -705
rect 2607 -745 2619 -711
rect 2727 -745 2739 -711
rect 2607 -751 2739 -745
rect 2805 -711 2937 -705
rect 2805 -745 2817 -711
rect 2925 -745 2937 -711
rect 2805 -751 2937 -745
rect 3003 -711 3135 -705
rect 3003 -745 3015 -711
rect 3123 -745 3135 -711
rect 3003 -751 3135 -745
rect 3201 -711 3333 -705
rect 3201 -745 3213 -711
rect 3321 -745 3333 -711
rect 3201 -751 3333 -745
rect 3399 -711 3531 -705
rect 3399 -745 3411 -711
rect 3519 -745 3531 -711
rect 3399 -751 3531 -745
rect 3597 -711 3729 -705
rect 3597 -745 3609 -711
rect 3717 -745 3729 -711
rect 3597 -751 3729 -745
rect 3795 -711 3927 -705
rect 3795 -745 3807 -711
rect 3915 -745 3927 -711
rect 3795 -751 3927 -745
rect 3993 -711 4125 -705
rect 3993 -745 4005 -711
rect 4113 -745 4125 -711
rect 3993 -751 4125 -745
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 1 nf 42 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
