magic
tech sky130A
magscale 1 2
timestamp 1619109957
<< nwell >>
rect -1647 -759 1647 759
<< pmos >>
rect -1451 -540 -1361 540
rect -1303 -540 -1213 540
rect -1155 -540 -1065 540
rect -1007 -540 -917 540
rect -859 -540 -769 540
rect -711 -540 -621 540
rect -563 -540 -473 540
rect -415 -540 -325 540
rect -267 -540 -177 540
rect -119 -540 -29 540
rect 29 -540 119 540
rect 177 -540 267 540
rect 325 -540 415 540
rect 473 -540 563 540
rect 621 -540 711 540
rect 769 -540 859 540
rect 917 -540 1007 540
rect 1065 -540 1155 540
rect 1213 -540 1303 540
rect 1361 -540 1451 540
<< pdiff >>
rect -1509 528 -1451 540
rect -1509 -528 -1497 528
rect -1463 -528 -1451 528
rect -1509 -540 -1451 -528
rect -1361 528 -1303 540
rect -1361 -528 -1349 528
rect -1315 -528 -1303 528
rect -1361 -540 -1303 -528
rect -1213 528 -1155 540
rect -1213 -528 -1201 528
rect -1167 -528 -1155 528
rect -1213 -540 -1155 -528
rect -1065 528 -1007 540
rect -1065 -528 -1053 528
rect -1019 -528 -1007 528
rect -1065 -540 -1007 -528
rect -917 528 -859 540
rect -917 -528 -905 528
rect -871 -528 -859 528
rect -917 -540 -859 -528
rect -769 528 -711 540
rect -769 -528 -757 528
rect -723 -528 -711 528
rect -769 -540 -711 -528
rect -621 528 -563 540
rect -621 -528 -609 528
rect -575 -528 -563 528
rect -621 -540 -563 -528
rect -473 528 -415 540
rect -473 -528 -461 528
rect -427 -528 -415 528
rect -473 -540 -415 -528
rect -325 528 -267 540
rect -325 -528 -313 528
rect -279 -528 -267 528
rect -325 -540 -267 -528
rect -177 528 -119 540
rect -177 -528 -165 528
rect -131 -528 -119 528
rect -177 -540 -119 -528
rect -29 528 29 540
rect -29 -528 -17 528
rect 17 -528 29 528
rect -29 -540 29 -528
rect 119 528 177 540
rect 119 -528 131 528
rect 165 -528 177 528
rect 119 -540 177 -528
rect 267 528 325 540
rect 267 -528 279 528
rect 313 -528 325 528
rect 267 -540 325 -528
rect 415 528 473 540
rect 415 -528 427 528
rect 461 -528 473 528
rect 415 -540 473 -528
rect 563 528 621 540
rect 563 -528 575 528
rect 609 -528 621 528
rect 563 -540 621 -528
rect 711 528 769 540
rect 711 -528 723 528
rect 757 -528 769 528
rect 711 -540 769 -528
rect 859 528 917 540
rect 859 -528 871 528
rect 905 -528 917 528
rect 859 -540 917 -528
rect 1007 528 1065 540
rect 1007 -528 1019 528
rect 1053 -528 1065 528
rect 1007 -540 1065 -528
rect 1155 528 1213 540
rect 1155 -528 1167 528
rect 1201 -528 1213 528
rect 1155 -540 1213 -528
rect 1303 528 1361 540
rect 1303 -528 1315 528
rect 1349 -528 1361 528
rect 1303 -540 1361 -528
rect 1451 528 1509 540
rect 1451 -528 1463 528
rect 1497 -528 1509 528
rect 1451 -540 1509 -528
<< pdiffc >>
rect -1497 -528 -1463 528
rect -1349 -528 -1315 528
rect -1201 -528 -1167 528
rect -1053 -528 -1019 528
rect -905 -528 -871 528
rect -757 -528 -723 528
rect -609 -528 -575 528
rect -461 -528 -427 528
rect -313 -528 -279 528
rect -165 -528 -131 528
rect -17 -528 17 528
rect 131 -528 165 528
rect 279 -528 313 528
rect 427 -528 461 528
rect 575 -528 609 528
rect 723 -528 757 528
rect 871 -528 905 528
rect 1019 -528 1053 528
rect 1167 -528 1201 528
rect 1315 -528 1349 528
rect 1463 -528 1497 528
<< nsubdiff >>
rect -1611 689 -1515 723
rect 1515 689 1611 723
rect -1611 627 -1577 689
rect 1577 627 1611 689
rect -1611 -689 -1577 -627
rect 1577 -689 1611 -627
rect -1611 -723 -1515 -689
rect 1515 -723 1611 -689
<< nsubdiffcont >>
rect -1515 689 1515 723
rect -1611 -627 -1577 627
rect 1577 -627 1611 627
rect -1515 -723 1515 -689
<< poly >>
rect -1451 621 -1361 637
rect -1451 587 -1435 621
rect -1377 587 -1361 621
rect -1451 540 -1361 587
rect -1303 621 -1213 637
rect -1303 587 -1287 621
rect -1229 587 -1213 621
rect -1303 540 -1213 587
rect -1155 621 -1065 637
rect -1155 587 -1139 621
rect -1081 587 -1065 621
rect -1155 540 -1065 587
rect -1007 621 -917 637
rect -1007 587 -991 621
rect -933 587 -917 621
rect -1007 540 -917 587
rect -859 621 -769 637
rect -859 587 -843 621
rect -785 587 -769 621
rect -859 540 -769 587
rect -711 621 -621 637
rect -711 587 -695 621
rect -637 587 -621 621
rect -711 540 -621 587
rect -563 621 -473 637
rect -563 587 -547 621
rect -489 587 -473 621
rect -563 540 -473 587
rect -415 621 -325 637
rect -415 587 -399 621
rect -341 587 -325 621
rect -415 540 -325 587
rect -267 621 -177 637
rect -267 587 -251 621
rect -193 587 -177 621
rect -267 540 -177 587
rect -119 621 -29 637
rect -119 587 -103 621
rect -45 587 -29 621
rect -119 540 -29 587
rect 29 621 119 637
rect 29 587 45 621
rect 103 587 119 621
rect 29 540 119 587
rect 177 621 267 637
rect 177 587 193 621
rect 251 587 267 621
rect 177 540 267 587
rect 325 621 415 637
rect 325 587 341 621
rect 399 587 415 621
rect 325 540 415 587
rect 473 621 563 637
rect 473 587 489 621
rect 547 587 563 621
rect 473 540 563 587
rect 621 621 711 637
rect 621 587 637 621
rect 695 587 711 621
rect 621 540 711 587
rect 769 621 859 637
rect 769 587 785 621
rect 843 587 859 621
rect 769 540 859 587
rect 917 621 1007 637
rect 917 587 933 621
rect 991 587 1007 621
rect 917 540 1007 587
rect 1065 621 1155 637
rect 1065 587 1081 621
rect 1139 587 1155 621
rect 1065 540 1155 587
rect 1213 621 1303 637
rect 1213 587 1229 621
rect 1287 587 1303 621
rect 1213 540 1303 587
rect 1361 621 1451 637
rect 1361 587 1377 621
rect 1435 587 1451 621
rect 1361 540 1451 587
rect -1451 -587 -1361 -540
rect -1451 -621 -1435 -587
rect -1377 -621 -1361 -587
rect -1451 -637 -1361 -621
rect -1303 -587 -1213 -540
rect -1303 -621 -1287 -587
rect -1229 -621 -1213 -587
rect -1303 -637 -1213 -621
rect -1155 -587 -1065 -540
rect -1155 -621 -1139 -587
rect -1081 -621 -1065 -587
rect -1155 -637 -1065 -621
rect -1007 -587 -917 -540
rect -1007 -621 -991 -587
rect -933 -621 -917 -587
rect -1007 -637 -917 -621
rect -859 -587 -769 -540
rect -859 -621 -843 -587
rect -785 -621 -769 -587
rect -859 -637 -769 -621
rect -711 -587 -621 -540
rect -711 -621 -695 -587
rect -637 -621 -621 -587
rect -711 -637 -621 -621
rect -563 -587 -473 -540
rect -563 -621 -547 -587
rect -489 -621 -473 -587
rect -563 -637 -473 -621
rect -415 -587 -325 -540
rect -415 -621 -399 -587
rect -341 -621 -325 -587
rect -415 -637 -325 -621
rect -267 -587 -177 -540
rect -267 -621 -251 -587
rect -193 -621 -177 -587
rect -267 -637 -177 -621
rect -119 -587 -29 -540
rect -119 -621 -103 -587
rect -45 -621 -29 -587
rect -119 -637 -29 -621
rect 29 -587 119 -540
rect 29 -621 45 -587
rect 103 -621 119 -587
rect 29 -637 119 -621
rect 177 -587 267 -540
rect 177 -621 193 -587
rect 251 -621 267 -587
rect 177 -637 267 -621
rect 325 -587 415 -540
rect 325 -621 341 -587
rect 399 -621 415 -587
rect 325 -637 415 -621
rect 473 -587 563 -540
rect 473 -621 489 -587
rect 547 -621 563 -587
rect 473 -637 563 -621
rect 621 -587 711 -540
rect 621 -621 637 -587
rect 695 -621 711 -587
rect 621 -637 711 -621
rect 769 -587 859 -540
rect 769 -621 785 -587
rect 843 -621 859 -587
rect 769 -637 859 -621
rect 917 -587 1007 -540
rect 917 -621 933 -587
rect 991 -621 1007 -587
rect 917 -637 1007 -621
rect 1065 -587 1155 -540
rect 1065 -621 1081 -587
rect 1139 -621 1155 -587
rect 1065 -637 1155 -621
rect 1213 -587 1303 -540
rect 1213 -621 1229 -587
rect 1287 -621 1303 -587
rect 1213 -637 1303 -621
rect 1361 -587 1451 -540
rect 1361 -621 1377 -587
rect 1435 -621 1451 -587
rect 1361 -637 1451 -621
<< polycont >>
rect -1435 587 -1377 621
rect -1287 587 -1229 621
rect -1139 587 -1081 621
rect -991 587 -933 621
rect -843 587 -785 621
rect -695 587 -637 621
rect -547 587 -489 621
rect -399 587 -341 621
rect -251 587 -193 621
rect -103 587 -45 621
rect 45 587 103 621
rect 193 587 251 621
rect 341 587 399 621
rect 489 587 547 621
rect 637 587 695 621
rect 785 587 843 621
rect 933 587 991 621
rect 1081 587 1139 621
rect 1229 587 1287 621
rect 1377 587 1435 621
rect -1435 -621 -1377 -587
rect -1287 -621 -1229 -587
rect -1139 -621 -1081 -587
rect -991 -621 -933 -587
rect -843 -621 -785 -587
rect -695 -621 -637 -587
rect -547 -621 -489 -587
rect -399 -621 -341 -587
rect -251 -621 -193 -587
rect -103 -621 -45 -587
rect 45 -621 103 -587
rect 193 -621 251 -587
rect 341 -621 399 -587
rect 489 -621 547 -587
rect 637 -621 695 -587
rect 785 -621 843 -587
rect 933 -621 991 -587
rect 1081 -621 1139 -587
rect 1229 -621 1287 -587
rect 1377 -621 1435 -587
<< locali >>
rect -1611 689 -1515 723
rect 1515 689 1611 723
rect -1611 627 -1577 689
rect 1577 627 1611 689
rect -1451 587 -1435 621
rect -1377 587 -1361 621
rect -1303 587 -1287 621
rect -1229 587 -1213 621
rect -1155 587 -1139 621
rect -1081 587 -1065 621
rect -1007 587 -991 621
rect -933 587 -917 621
rect -859 587 -843 621
rect -785 587 -769 621
rect -711 587 -695 621
rect -637 587 -621 621
rect -563 587 -547 621
rect -489 587 -473 621
rect -415 587 -399 621
rect -341 587 -325 621
rect -267 587 -251 621
rect -193 587 -177 621
rect -119 587 -103 621
rect -45 587 -29 621
rect 29 587 45 621
rect 103 587 119 621
rect 177 587 193 621
rect 251 587 267 621
rect 325 587 341 621
rect 399 587 415 621
rect 473 587 489 621
rect 547 587 563 621
rect 621 587 637 621
rect 695 587 711 621
rect 769 587 785 621
rect 843 587 859 621
rect 917 587 933 621
rect 991 587 1007 621
rect 1065 587 1081 621
rect 1139 587 1155 621
rect 1213 587 1229 621
rect 1287 587 1303 621
rect 1361 587 1377 621
rect 1435 587 1451 621
rect -1497 528 -1463 544
rect -1497 -544 -1463 -528
rect -1349 528 -1315 544
rect -1349 -544 -1315 -528
rect -1201 528 -1167 544
rect -1201 -544 -1167 -528
rect -1053 528 -1019 544
rect -1053 -544 -1019 -528
rect -905 528 -871 544
rect -905 -544 -871 -528
rect -757 528 -723 544
rect -757 -544 -723 -528
rect -609 528 -575 544
rect -609 -544 -575 -528
rect -461 528 -427 544
rect -461 -544 -427 -528
rect -313 528 -279 544
rect -313 -544 -279 -528
rect -165 528 -131 544
rect -165 -544 -131 -528
rect -17 528 17 544
rect -17 -544 17 -528
rect 131 528 165 544
rect 131 -544 165 -528
rect 279 528 313 544
rect 279 -544 313 -528
rect 427 528 461 544
rect 427 -544 461 -528
rect 575 528 609 544
rect 575 -544 609 -528
rect 723 528 757 544
rect 723 -544 757 -528
rect 871 528 905 544
rect 871 -544 905 -528
rect 1019 528 1053 544
rect 1019 -544 1053 -528
rect 1167 528 1201 544
rect 1167 -544 1201 -528
rect 1315 528 1349 544
rect 1315 -544 1349 -528
rect 1463 528 1497 544
rect 1463 -544 1497 -528
rect -1451 -621 -1435 -587
rect -1377 -621 -1361 -587
rect -1303 -621 -1287 -587
rect -1229 -621 -1213 -587
rect -1155 -621 -1139 -587
rect -1081 -621 -1065 -587
rect -1007 -621 -991 -587
rect -933 -621 -917 -587
rect -859 -621 -843 -587
rect -785 -621 -769 -587
rect -711 -621 -695 -587
rect -637 -621 -621 -587
rect -563 -621 -547 -587
rect -489 -621 -473 -587
rect -415 -621 -399 -587
rect -341 -621 -325 -587
rect -267 -621 -251 -587
rect -193 -621 -177 -587
rect -119 -621 -103 -587
rect -45 -621 -29 -587
rect 29 -621 45 -587
rect 103 -621 119 -587
rect 177 -621 193 -587
rect 251 -621 267 -587
rect 325 -621 341 -587
rect 399 -621 415 -587
rect 473 -621 489 -587
rect 547 -621 563 -587
rect 621 -621 637 -587
rect 695 -621 711 -587
rect 769 -621 785 -587
rect 843 -621 859 -587
rect 917 -621 933 -587
rect 991 -621 1007 -587
rect 1065 -621 1081 -587
rect 1139 -621 1155 -587
rect 1213 -621 1229 -587
rect 1287 -621 1303 -587
rect 1361 -621 1377 -587
rect 1435 -621 1451 -587
rect -1611 -689 -1577 -627
rect 1577 -689 1611 -627
rect -1611 -723 -1515 -689
rect 1515 -723 1611 -689
<< viali >>
rect -1435 587 -1377 621
rect -1287 587 -1229 621
rect -1139 587 -1081 621
rect -991 587 -933 621
rect -843 587 -785 621
rect -695 587 -637 621
rect -547 587 -489 621
rect -399 587 -341 621
rect -251 587 -193 621
rect -103 587 -45 621
rect 45 587 103 621
rect 193 587 251 621
rect 341 587 399 621
rect 489 587 547 621
rect 637 587 695 621
rect 785 587 843 621
rect 933 587 991 621
rect 1081 587 1139 621
rect 1229 587 1287 621
rect 1377 587 1435 621
rect -1497 -528 -1463 528
rect -1349 -528 -1315 528
rect -1201 -528 -1167 528
rect -1053 -528 -1019 528
rect -905 -528 -871 528
rect -757 -528 -723 528
rect -609 -528 -575 528
rect -461 -528 -427 528
rect -313 -528 -279 528
rect -165 -528 -131 528
rect -17 -528 17 528
rect 131 -528 165 528
rect 279 -528 313 528
rect 427 -528 461 528
rect 575 -528 609 528
rect 723 -528 757 528
rect 871 -528 905 528
rect 1019 -528 1053 528
rect 1167 -528 1201 528
rect 1315 -528 1349 528
rect 1463 -528 1497 528
rect -1435 -621 -1377 -587
rect -1287 -621 -1229 -587
rect -1139 -621 -1081 -587
rect -991 -621 -933 -587
rect -843 -621 -785 -587
rect -695 -621 -637 -587
rect -547 -621 -489 -587
rect -399 -621 -341 -587
rect -251 -621 -193 -587
rect -103 -621 -45 -587
rect 45 -621 103 -587
rect 193 -621 251 -587
rect 341 -621 399 -587
rect 489 -621 547 -587
rect 637 -621 695 -587
rect 785 -621 843 -587
rect 933 -621 991 -587
rect 1081 -621 1139 -587
rect 1229 -621 1287 -587
rect 1377 -621 1435 -587
<< metal1 >>
rect -1447 621 -1365 627
rect -1447 587 -1435 621
rect -1377 587 -1365 621
rect -1447 581 -1365 587
rect -1299 621 -1217 627
rect -1299 587 -1287 621
rect -1229 587 -1217 621
rect -1299 581 -1217 587
rect -1151 621 -1069 627
rect -1151 587 -1139 621
rect -1081 587 -1069 621
rect -1151 581 -1069 587
rect -1003 621 -921 627
rect -1003 587 -991 621
rect -933 587 -921 621
rect -1003 581 -921 587
rect -855 621 -773 627
rect -855 587 -843 621
rect -785 587 -773 621
rect -855 581 -773 587
rect -707 621 -625 627
rect -707 587 -695 621
rect -637 587 -625 621
rect -707 581 -625 587
rect -559 621 -477 627
rect -559 587 -547 621
rect -489 587 -477 621
rect -559 581 -477 587
rect -411 621 -329 627
rect -411 587 -399 621
rect -341 587 -329 621
rect -411 581 -329 587
rect -263 621 -181 627
rect -263 587 -251 621
rect -193 587 -181 621
rect -263 581 -181 587
rect -115 621 -33 627
rect -115 587 -103 621
rect -45 587 -33 621
rect -115 581 -33 587
rect 33 621 115 627
rect 33 587 45 621
rect 103 587 115 621
rect 33 581 115 587
rect 181 621 263 627
rect 181 587 193 621
rect 251 587 263 621
rect 181 581 263 587
rect 329 621 411 627
rect 329 587 341 621
rect 399 587 411 621
rect 329 581 411 587
rect 477 621 559 627
rect 477 587 489 621
rect 547 587 559 621
rect 477 581 559 587
rect 625 621 707 627
rect 625 587 637 621
rect 695 587 707 621
rect 625 581 707 587
rect 773 621 855 627
rect 773 587 785 621
rect 843 587 855 621
rect 773 581 855 587
rect 921 621 1003 627
rect 921 587 933 621
rect 991 587 1003 621
rect 921 581 1003 587
rect 1069 621 1151 627
rect 1069 587 1081 621
rect 1139 587 1151 621
rect 1069 581 1151 587
rect 1217 621 1299 627
rect 1217 587 1229 621
rect 1287 587 1299 621
rect 1217 581 1299 587
rect 1365 621 1447 627
rect 1365 587 1377 621
rect 1435 587 1447 621
rect 1365 581 1447 587
rect -1503 528 -1457 540
rect -1503 -528 -1497 528
rect -1463 -528 -1457 528
rect -1503 -540 -1457 -528
rect -1355 528 -1309 540
rect -1355 -528 -1349 528
rect -1315 -528 -1309 528
rect -1355 -540 -1309 -528
rect -1207 528 -1161 540
rect -1207 -528 -1201 528
rect -1167 -528 -1161 528
rect -1207 -540 -1161 -528
rect -1059 528 -1013 540
rect -1059 -528 -1053 528
rect -1019 -528 -1013 528
rect -1059 -540 -1013 -528
rect -911 528 -865 540
rect -911 -528 -905 528
rect -871 -528 -865 528
rect -911 -540 -865 -528
rect -763 528 -717 540
rect -763 -528 -757 528
rect -723 -528 -717 528
rect -763 -540 -717 -528
rect -615 528 -569 540
rect -615 -528 -609 528
rect -575 -528 -569 528
rect -615 -540 -569 -528
rect -467 528 -421 540
rect -467 -528 -461 528
rect -427 -528 -421 528
rect -467 -540 -421 -528
rect -319 528 -273 540
rect -319 -528 -313 528
rect -279 -528 -273 528
rect -319 -540 -273 -528
rect -171 528 -125 540
rect -171 -528 -165 528
rect -131 -528 -125 528
rect -171 -540 -125 -528
rect -23 528 23 540
rect -23 -528 -17 528
rect 17 -528 23 528
rect -23 -540 23 -528
rect 125 528 171 540
rect 125 -528 131 528
rect 165 -528 171 528
rect 125 -540 171 -528
rect 273 528 319 540
rect 273 -528 279 528
rect 313 -528 319 528
rect 273 -540 319 -528
rect 421 528 467 540
rect 421 -528 427 528
rect 461 -528 467 528
rect 421 -540 467 -528
rect 569 528 615 540
rect 569 -528 575 528
rect 609 -528 615 528
rect 569 -540 615 -528
rect 717 528 763 540
rect 717 -528 723 528
rect 757 -528 763 528
rect 717 -540 763 -528
rect 865 528 911 540
rect 865 -528 871 528
rect 905 -528 911 528
rect 865 -540 911 -528
rect 1013 528 1059 540
rect 1013 -528 1019 528
rect 1053 -528 1059 528
rect 1013 -540 1059 -528
rect 1161 528 1207 540
rect 1161 -528 1167 528
rect 1201 -528 1207 528
rect 1161 -540 1207 -528
rect 1309 528 1355 540
rect 1309 -528 1315 528
rect 1349 -528 1355 528
rect 1309 -540 1355 -528
rect 1457 528 1503 540
rect 1457 -528 1463 528
rect 1497 -528 1503 528
rect 1457 -540 1503 -528
rect -1447 -587 -1365 -581
rect -1447 -621 -1435 -587
rect -1377 -621 -1365 -587
rect -1447 -627 -1365 -621
rect -1299 -587 -1217 -581
rect -1299 -621 -1287 -587
rect -1229 -621 -1217 -587
rect -1299 -627 -1217 -621
rect -1151 -587 -1069 -581
rect -1151 -621 -1139 -587
rect -1081 -621 -1069 -587
rect -1151 -627 -1069 -621
rect -1003 -587 -921 -581
rect -1003 -621 -991 -587
rect -933 -621 -921 -587
rect -1003 -627 -921 -621
rect -855 -587 -773 -581
rect -855 -621 -843 -587
rect -785 -621 -773 -587
rect -855 -627 -773 -621
rect -707 -587 -625 -581
rect -707 -621 -695 -587
rect -637 -621 -625 -587
rect -707 -627 -625 -621
rect -559 -587 -477 -581
rect -559 -621 -547 -587
rect -489 -621 -477 -587
rect -559 -627 -477 -621
rect -411 -587 -329 -581
rect -411 -621 -399 -587
rect -341 -621 -329 -587
rect -411 -627 -329 -621
rect -263 -587 -181 -581
rect -263 -621 -251 -587
rect -193 -621 -181 -587
rect -263 -627 -181 -621
rect -115 -587 -33 -581
rect -115 -621 -103 -587
rect -45 -621 -33 -587
rect -115 -627 -33 -621
rect 33 -587 115 -581
rect 33 -621 45 -587
rect 103 -621 115 -587
rect 33 -627 115 -621
rect 181 -587 263 -581
rect 181 -621 193 -587
rect 251 -621 263 -587
rect 181 -627 263 -621
rect 329 -587 411 -581
rect 329 -621 341 -587
rect 399 -621 411 -587
rect 329 -627 411 -621
rect 477 -587 559 -581
rect 477 -621 489 -587
rect 547 -621 559 -587
rect 477 -627 559 -621
rect 625 -587 707 -581
rect 625 -621 637 -587
rect 695 -621 707 -587
rect 625 -627 707 -621
rect 773 -587 855 -581
rect 773 -621 785 -587
rect 843 -621 855 -587
rect 773 -627 855 -621
rect 921 -587 1003 -581
rect 921 -621 933 -587
rect 991 -621 1003 -587
rect 921 -627 1003 -621
rect 1069 -587 1151 -581
rect 1069 -621 1081 -587
rect 1139 -621 1151 -587
rect 1069 -627 1151 -621
rect 1217 -587 1299 -581
rect 1217 -621 1229 -587
rect 1287 -621 1299 -587
rect 1217 -627 1299 -621
rect 1365 -587 1447 -581
rect 1365 -621 1377 -587
rect 1435 -621 1447 -587
rect 1365 -627 1447 -621
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1594 -706 1594 706
string parameters w 5.4 l 0.45 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
