magic
tech sky130A
magscale 1 2
timestamp 1615600491
<< error_s >>
rect 65 1497 468 1498
rect 46 1341 468 1497
rect 214 1330 487 1341
rect 1166 1340 1398 1341
rect 214 1329 233 1330
rect 300 1262 487 1330
rect 75 852 113 1072
rect 226 852 260 1072
rect 75 818 480 852
rect 831 747 871 979
rect 846 730 1085 747
rect 871 725 1085 730
<< pwell >>
rect -1083 329 6 356
rect -469 6 6 329
<< metal1 >>
rect -517 1612 -220 1658
rect -32 1612 23 1659
rect 1462 1393 1471 1427
rect 99 1278 100 1349
rect -1059 1197 -1049 1249
rect -997 1197 -987 1249
rect -1084 811 -170 858
rect -98 852 1467 858
rect -98 818 322 852
rect 561 818 906 852
rect 1370 818 1467 852
rect -98 811 1467 818
rect -762 454 -752 506
rect -700 454 -690 506
rect -37 391 -27 443
rect 25 425 35 443
rect 25 392 64 425
rect 25 391 63 392
rect -1029 337 -1019 389
rect -967 337 -957 389
rect -551 356 -477 387
rect -469 13 5 58
rect 1103 52 1496 58
rect 1103 18 1115 52
rect 1484 18 1496 52
rect 1103 12 1496 18
<< via1 >>
rect -1049 1197 -997 1249
rect -752 454 -700 506
rect -27 391 25 443
rect -1019 337 -967 389
<< metal2 >>
rect -1040 1553 1423 1587
rect -1040 1259 -1006 1553
rect -1049 1249 -997 1259
rect -1049 1187 -997 1197
rect -1040 399 -1006 1187
rect -768 506 -700 516
rect -768 464 -752 506
rect -255 498 -221 968
rect -700 464 -221 498
rect -752 444 -700 454
rect -17 453 17 1314
rect 1389 1295 1423 1553
rect -27 443 25 453
rect -1040 389 -967 399
rect -1040 345 -1019 389
rect -27 381 25 391
rect -1019 327 -967 337
rect 31 182 32 216
use and  and_0
timestamp 1615600491
transform 1 0 -1017 0 1 494
box -67 -481 548 400
use xor  xor_0
timestamp 1615600491
transform 1 0 -864 0 -1 1689
box -220 31 881 917
use ffd  ffd_0
timestamp 1615600491
transform 1 0 -1403 0 1 -1111
box 1310 1103 2980 2788
<< labels >>
rlabel metal2 1389 1295 1423 1587 1 Dn
rlabel space 1246 1393 1466 1427 1 Dnb
rlabel metal2 -700 464 -221 498 1 CE
rlabel metal1 -480 356 -477 387 1 Sout
rlabel metal1 1470 1393 1471 1427 1 Dnb
rlabel metal2 31 182 32 216 1 CLR
rlabel metal1 99 1278 100 1349 1 CLK
<< end >>
