magic
tech sky130A
magscale 1 2
timestamp 1622937437
<< error_p >>
rect -927 921 -865 927
rect -799 921 -737 927
rect -671 921 -609 927
rect -543 921 -481 927
rect -415 921 -353 927
rect -287 921 -225 927
rect -159 921 -97 927
rect -31 921 31 927
rect 97 921 159 927
rect 225 921 287 927
rect 353 921 415 927
rect 481 921 543 927
rect 609 921 671 927
rect 737 921 799 927
rect 865 921 927 927
rect -927 887 -915 921
rect -799 887 -787 921
rect -671 887 -659 921
rect -543 887 -531 921
rect -415 887 -403 921
rect -287 887 -275 921
rect -159 887 -147 921
rect -31 887 -19 921
rect 97 887 109 921
rect 225 887 237 921
rect 353 887 365 921
rect 481 887 493 921
rect 609 887 621 921
rect 737 887 749 921
rect 865 887 877 921
rect -927 881 -865 887
rect -799 881 -737 887
rect -671 881 -609 887
rect -543 881 -481 887
rect -415 881 -353 887
rect -287 881 -225 887
rect -159 881 -97 887
rect -31 881 31 887
rect 97 881 159 887
rect 225 881 287 887
rect 353 881 415 887
rect 481 881 543 887
rect 609 881 671 887
rect 737 881 799 887
rect 865 881 927 887
rect -927 -887 -865 -881
rect -799 -887 -737 -881
rect -671 -887 -609 -881
rect -543 -887 -481 -881
rect -415 -887 -353 -881
rect -287 -887 -225 -881
rect -159 -887 -97 -881
rect -31 -887 31 -881
rect 97 -887 159 -881
rect 225 -887 287 -881
rect 353 -887 415 -881
rect 481 -887 543 -881
rect 609 -887 671 -881
rect 737 -887 799 -881
rect 865 -887 927 -881
rect -927 -921 -915 -887
rect -799 -921 -787 -887
rect -671 -921 -659 -887
rect -543 -921 -531 -887
rect -415 -921 -403 -887
rect -287 -921 -275 -887
rect -159 -921 -147 -887
rect -31 -921 -19 -887
rect 97 -921 109 -887
rect 225 -921 237 -887
rect 353 -921 365 -887
rect 481 -921 493 -887
rect 609 -921 621 -887
rect 737 -921 749 -887
rect 865 -921 877 -887
rect -927 -927 -865 -921
rect -799 -927 -737 -921
rect -671 -927 -609 -921
rect -543 -927 -481 -921
rect -415 -927 -353 -921
rect -287 -927 -225 -921
rect -159 -927 -97 -921
rect -31 -927 31 -921
rect 97 -927 159 -921
rect 225 -927 287 -921
rect 353 -927 415 -921
rect 481 -927 543 -921
rect 609 -927 671 -921
rect 737 -927 799 -921
rect 865 -927 927 -921
<< nwell >>
rect -1127 -1059 1127 1059
<< pmos >>
rect -931 -840 -861 840
rect -803 -840 -733 840
rect -675 -840 -605 840
rect -547 -840 -477 840
rect -419 -840 -349 840
rect -291 -840 -221 840
rect -163 -840 -93 840
rect -35 -840 35 840
rect 93 -840 163 840
rect 221 -840 291 840
rect 349 -840 419 840
rect 477 -840 547 840
rect 605 -840 675 840
rect 733 -840 803 840
rect 861 -840 931 840
<< pdiff >>
rect -989 828 -931 840
rect -989 -828 -977 828
rect -943 -828 -931 828
rect -989 -840 -931 -828
rect -861 828 -803 840
rect -861 -828 -849 828
rect -815 -828 -803 828
rect -861 -840 -803 -828
rect -733 828 -675 840
rect -733 -828 -721 828
rect -687 -828 -675 828
rect -733 -840 -675 -828
rect -605 828 -547 840
rect -605 -828 -593 828
rect -559 -828 -547 828
rect -605 -840 -547 -828
rect -477 828 -419 840
rect -477 -828 -465 828
rect -431 -828 -419 828
rect -477 -840 -419 -828
rect -349 828 -291 840
rect -349 -828 -337 828
rect -303 -828 -291 828
rect -349 -840 -291 -828
rect -221 828 -163 840
rect -221 -828 -209 828
rect -175 -828 -163 828
rect -221 -840 -163 -828
rect -93 828 -35 840
rect -93 -828 -81 828
rect -47 -828 -35 828
rect -93 -840 -35 -828
rect 35 828 93 840
rect 35 -828 47 828
rect 81 -828 93 828
rect 35 -840 93 -828
rect 163 828 221 840
rect 163 -828 175 828
rect 209 -828 221 828
rect 163 -840 221 -828
rect 291 828 349 840
rect 291 -828 303 828
rect 337 -828 349 828
rect 291 -840 349 -828
rect 419 828 477 840
rect 419 -828 431 828
rect 465 -828 477 828
rect 419 -840 477 -828
rect 547 828 605 840
rect 547 -828 559 828
rect 593 -828 605 828
rect 547 -840 605 -828
rect 675 828 733 840
rect 675 -828 687 828
rect 721 -828 733 828
rect 675 -840 733 -828
rect 803 828 861 840
rect 803 -828 815 828
rect 849 -828 861 828
rect 803 -840 861 -828
rect 931 828 989 840
rect 931 -828 943 828
rect 977 -828 989 828
rect 931 -840 989 -828
<< pdiffc >>
rect -977 -828 -943 828
rect -849 -828 -815 828
rect -721 -828 -687 828
rect -593 -828 -559 828
rect -465 -828 -431 828
rect -337 -828 -303 828
rect -209 -828 -175 828
rect -81 -828 -47 828
rect 47 -828 81 828
rect 175 -828 209 828
rect 303 -828 337 828
rect 431 -828 465 828
rect 559 -828 593 828
rect 687 -828 721 828
rect 815 -828 849 828
rect 943 -828 977 828
<< nsubdiff >>
rect -1091 989 -995 1023
rect 995 989 1091 1023
rect -1091 927 -1057 989
rect 1057 927 1091 989
rect -1091 -989 -1057 -927
rect 1057 -989 1091 -927
rect -1091 -1023 -995 -989
rect 995 -1023 1091 -989
<< nsubdiffcont >>
rect -995 989 995 1023
rect -1091 -927 -1057 927
rect 1057 -927 1091 927
rect -995 -1023 995 -989
<< poly >>
rect -931 921 -861 937
rect -931 887 -915 921
rect -877 887 -861 921
rect -931 840 -861 887
rect -803 921 -733 937
rect -803 887 -787 921
rect -749 887 -733 921
rect -803 840 -733 887
rect -675 921 -605 937
rect -675 887 -659 921
rect -621 887 -605 921
rect -675 840 -605 887
rect -547 921 -477 937
rect -547 887 -531 921
rect -493 887 -477 921
rect -547 840 -477 887
rect -419 921 -349 937
rect -419 887 -403 921
rect -365 887 -349 921
rect -419 840 -349 887
rect -291 921 -221 937
rect -291 887 -275 921
rect -237 887 -221 921
rect -291 840 -221 887
rect -163 921 -93 937
rect -163 887 -147 921
rect -109 887 -93 921
rect -163 840 -93 887
rect -35 921 35 937
rect -35 887 -19 921
rect 19 887 35 921
rect -35 840 35 887
rect 93 921 163 937
rect 93 887 109 921
rect 147 887 163 921
rect 93 840 163 887
rect 221 921 291 937
rect 221 887 237 921
rect 275 887 291 921
rect 221 840 291 887
rect 349 921 419 937
rect 349 887 365 921
rect 403 887 419 921
rect 349 840 419 887
rect 477 921 547 937
rect 477 887 493 921
rect 531 887 547 921
rect 477 840 547 887
rect 605 921 675 937
rect 605 887 621 921
rect 659 887 675 921
rect 605 840 675 887
rect 733 921 803 937
rect 733 887 749 921
rect 787 887 803 921
rect 733 840 803 887
rect 861 921 931 937
rect 861 887 877 921
rect 915 887 931 921
rect 861 840 931 887
rect -931 -887 -861 -840
rect -931 -921 -915 -887
rect -877 -921 -861 -887
rect -931 -937 -861 -921
rect -803 -887 -733 -840
rect -803 -921 -787 -887
rect -749 -921 -733 -887
rect -803 -937 -733 -921
rect -675 -887 -605 -840
rect -675 -921 -659 -887
rect -621 -921 -605 -887
rect -675 -937 -605 -921
rect -547 -887 -477 -840
rect -547 -921 -531 -887
rect -493 -921 -477 -887
rect -547 -937 -477 -921
rect -419 -887 -349 -840
rect -419 -921 -403 -887
rect -365 -921 -349 -887
rect -419 -937 -349 -921
rect -291 -887 -221 -840
rect -291 -921 -275 -887
rect -237 -921 -221 -887
rect -291 -937 -221 -921
rect -163 -887 -93 -840
rect -163 -921 -147 -887
rect -109 -921 -93 -887
rect -163 -937 -93 -921
rect -35 -887 35 -840
rect -35 -921 -19 -887
rect 19 -921 35 -887
rect -35 -937 35 -921
rect 93 -887 163 -840
rect 93 -921 109 -887
rect 147 -921 163 -887
rect 93 -937 163 -921
rect 221 -887 291 -840
rect 221 -921 237 -887
rect 275 -921 291 -887
rect 221 -937 291 -921
rect 349 -887 419 -840
rect 349 -921 365 -887
rect 403 -921 419 -887
rect 349 -937 419 -921
rect 477 -887 547 -840
rect 477 -921 493 -887
rect 531 -921 547 -887
rect 477 -937 547 -921
rect 605 -887 675 -840
rect 605 -921 621 -887
rect 659 -921 675 -887
rect 605 -937 675 -921
rect 733 -887 803 -840
rect 733 -921 749 -887
rect 787 -921 803 -887
rect 733 -937 803 -921
rect 861 -887 931 -840
rect 861 -921 877 -887
rect 915 -921 931 -887
rect 861 -937 931 -921
<< polycont >>
rect -915 887 -877 921
rect -787 887 -749 921
rect -659 887 -621 921
rect -531 887 -493 921
rect -403 887 -365 921
rect -275 887 -237 921
rect -147 887 -109 921
rect -19 887 19 921
rect 109 887 147 921
rect 237 887 275 921
rect 365 887 403 921
rect 493 887 531 921
rect 621 887 659 921
rect 749 887 787 921
rect 877 887 915 921
rect -915 -921 -877 -887
rect -787 -921 -749 -887
rect -659 -921 -621 -887
rect -531 -921 -493 -887
rect -403 -921 -365 -887
rect -275 -921 -237 -887
rect -147 -921 -109 -887
rect -19 -921 19 -887
rect 109 -921 147 -887
rect 237 -921 275 -887
rect 365 -921 403 -887
rect 493 -921 531 -887
rect 621 -921 659 -887
rect 749 -921 787 -887
rect 877 -921 915 -887
<< locali >>
rect -1091 989 -995 1023
rect 995 989 1091 1023
rect -1091 927 -1057 989
rect 1057 927 1091 989
rect -931 887 -915 921
rect -877 887 -861 921
rect -803 887 -787 921
rect -749 887 -733 921
rect -675 887 -659 921
rect -621 887 -605 921
rect -547 887 -531 921
rect -493 887 -477 921
rect -419 887 -403 921
rect -365 887 -349 921
rect -291 887 -275 921
rect -237 887 -221 921
rect -163 887 -147 921
rect -109 887 -93 921
rect -35 887 -19 921
rect 19 887 35 921
rect 93 887 109 921
rect 147 887 163 921
rect 221 887 237 921
rect 275 887 291 921
rect 349 887 365 921
rect 403 887 419 921
rect 477 887 493 921
rect 531 887 547 921
rect 605 887 621 921
rect 659 887 675 921
rect 733 887 749 921
rect 787 887 803 921
rect 861 887 877 921
rect 915 887 931 921
rect -977 828 -943 844
rect -977 -844 -943 -828
rect -849 828 -815 844
rect -849 -844 -815 -828
rect -721 828 -687 844
rect -721 -844 -687 -828
rect -593 828 -559 844
rect -593 -844 -559 -828
rect -465 828 -431 844
rect -465 -844 -431 -828
rect -337 828 -303 844
rect -337 -844 -303 -828
rect -209 828 -175 844
rect -209 -844 -175 -828
rect -81 828 -47 844
rect -81 -844 -47 -828
rect 47 828 81 844
rect 47 -844 81 -828
rect 175 828 209 844
rect 175 -844 209 -828
rect 303 828 337 844
rect 303 -844 337 -828
rect 431 828 465 844
rect 431 -844 465 -828
rect 559 828 593 844
rect 559 -844 593 -828
rect 687 828 721 844
rect 687 -844 721 -828
rect 815 828 849 844
rect 815 -844 849 -828
rect 943 828 977 844
rect 943 -844 977 -828
rect -931 -921 -915 -887
rect -877 -921 -861 -887
rect -803 -921 -787 -887
rect -749 -921 -733 -887
rect -675 -921 -659 -887
rect -621 -921 -605 -887
rect -547 -921 -531 -887
rect -493 -921 -477 -887
rect -419 -921 -403 -887
rect -365 -921 -349 -887
rect -291 -921 -275 -887
rect -237 -921 -221 -887
rect -163 -921 -147 -887
rect -109 -921 -93 -887
rect -35 -921 -19 -887
rect 19 -921 35 -887
rect 93 -921 109 -887
rect 147 -921 163 -887
rect 221 -921 237 -887
rect 275 -921 291 -887
rect 349 -921 365 -887
rect 403 -921 419 -887
rect 477 -921 493 -887
rect 531 -921 547 -887
rect 605 -921 621 -887
rect 659 -921 675 -887
rect 733 -921 749 -887
rect 787 -921 803 -887
rect 861 -921 877 -887
rect 915 -921 931 -887
rect -1091 -989 -1057 -927
rect 1057 -989 1091 -927
rect -1091 -1023 -995 -989
rect 995 -1023 1091 -989
<< viali >>
rect -915 887 -877 921
rect -787 887 -749 921
rect -659 887 -621 921
rect -531 887 -493 921
rect -403 887 -365 921
rect -275 887 -237 921
rect -147 887 -109 921
rect -19 887 19 921
rect 109 887 147 921
rect 237 887 275 921
rect 365 887 403 921
rect 493 887 531 921
rect 621 887 659 921
rect 749 887 787 921
rect 877 887 915 921
rect -977 -828 -943 828
rect -849 -828 -815 828
rect -721 -828 -687 828
rect -593 -828 -559 828
rect -465 -828 -431 828
rect -337 -828 -303 828
rect -209 -828 -175 828
rect -81 -828 -47 828
rect 47 -828 81 828
rect 175 -828 209 828
rect 303 -828 337 828
rect 431 -828 465 828
rect 559 -828 593 828
rect 687 -828 721 828
rect 815 -828 849 828
rect 943 -828 977 828
rect -915 -921 -877 -887
rect -787 -921 -749 -887
rect -659 -921 -621 -887
rect -531 -921 -493 -887
rect -403 -921 -365 -887
rect -275 -921 -237 -887
rect -147 -921 -109 -887
rect -19 -921 19 -887
rect 109 -921 147 -887
rect 237 -921 275 -887
rect 365 -921 403 -887
rect 493 -921 531 -887
rect 621 -921 659 -887
rect 749 -921 787 -887
rect 877 -921 915 -887
<< metal1 >>
rect -927 921 -865 927
rect -927 887 -915 921
rect -877 887 -865 921
rect -927 881 -865 887
rect -799 921 -737 927
rect -799 887 -787 921
rect -749 887 -737 921
rect -799 881 -737 887
rect -671 921 -609 927
rect -671 887 -659 921
rect -621 887 -609 921
rect -671 881 -609 887
rect -543 921 -481 927
rect -543 887 -531 921
rect -493 887 -481 921
rect -543 881 -481 887
rect -415 921 -353 927
rect -415 887 -403 921
rect -365 887 -353 921
rect -415 881 -353 887
rect -287 921 -225 927
rect -287 887 -275 921
rect -237 887 -225 921
rect -287 881 -225 887
rect -159 921 -97 927
rect -159 887 -147 921
rect -109 887 -97 921
rect -159 881 -97 887
rect -31 921 31 927
rect -31 887 -19 921
rect 19 887 31 921
rect -31 881 31 887
rect 97 921 159 927
rect 97 887 109 921
rect 147 887 159 921
rect 97 881 159 887
rect 225 921 287 927
rect 225 887 237 921
rect 275 887 287 921
rect 225 881 287 887
rect 353 921 415 927
rect 353 887 365 921
rect 403 887 415 921
rect 353 881 415 887
rect 481 921 543 927
rect 481 887 493 921
rect 531 887 543 921
rect 481 881 543 887
rect 609 921 671 927
rect 609 887 621 921
rect 659 887 671 921
rect 609 881 671 887
rect 737 921 799 927
rect 737 887 749 921
rect 787 887 799 921
rect 737 881 799 887
rect 865 921 927 927
rect 865 887 877 921
rect 915 887 927 921
rect 865 881 927 887
rect -983 828 -937 840
rect -983 -828 -977 828
rect -943 -828 -937 828
rect -983 -840 -937 -828
rect -855 828 -809 840
rect -855 -828 -849 828
rect -815 -828 -809 828
rect -855 -840 -809 -828
rect -727 828 -681 840
rect -727 -828 -721 828
rect -687 -828 -681 828
rect -727 -840 -681 -828
rect -599 828 -553 840
rect -599 -828 -593 828
rect -559 -828 -553 828
rect -599 -840 -553 -828
rect -471 828 -425 840
rect -471 -828 -465 828
rect -431 -828 -425 828
rect -471 -840 -425 -828
rect -343 828 -297 840
rect -343 -828 -337 828
rect -303 -828 -297 828
rect -343 -840 -297 -828
rect -215 828 -169 840
rect -215 -828 -209 828
rect -175 -828 -169 828
rect -215 -840 -169 -828
rect -87 828 -41 840
rect -87 -828 -81 828
rect -47 -828 -41 828
rect -87 -840 -41 -828
rect 41 828 87 840
rect 41 -828 47 828
rect 81 -828 87 828
rect 41 -840 87 -828
rect 169 828 215 840
rect 169 -828 175 828
rect 209 -828 215 828
rect 169 -840 215 -828
rect 297 828 343 840
rect 297 -828 303 828
rect 337 -828 343 828
rect 297 -840 343 -828
rect 425 828 471 840
rect 425 -828 431 828
rect 465 -828 471 828
rect 425 -840 471 -828
rect 553 828 599 840
rect 553 -828 559 828
rect 593 -828 599 828
rect 553 -840 599 -828
rect 681 828 727 840
rect 681 -828 687 828
rect 721 -828 727 828
rect 681 -840 727 -828
rect 809 828 855 840
rect 809 -828 815 828
rect 849 -828 855 828
rect 809 -840 855 -828
rect 937 828 983 840
rect 937 -828 943 828
rect 977 -828 983 828
rect 937 -840 983 -828
rect -927 -887 -865 -881
rect -927 -921 -915 -887
rect -877 -921 -865 -887
rect -927 -927 -865 -921
rect -799 -887 -737 -881
rect -799 -921 -787 -887
rect -749 -921 -737 -887
rect -799 -927 -737 -921
rect -671 -887 -609 -881
rect -671 -921 -659 -887
rect -621 -921 -609 -887
rect -671 -927 -609 -921
rect -543 -887 -481 -881
rect -543 -921 -531 -887
rect -493 -921 -481 -887
rect -543 -927 -481 -921
rect -415 -887 -353 -881
rect -415 -921 -403 -887
rect -365 -921 -353 -887
rect -415 -927 -353 -921
rect -287 -887 -225 -881
rect -287 -921 -275 -887
rect -237 -921 -225 -887
rect -287 -927 -225 -921
rect -159 -887 -97 -881
rect -159 -921 -147 -887
rect -109 -921 -97 -887
rect -159 -927 -97 -921
rect -31 -887 31 -881
rect -31 -921 -19 -887
rect 19 -921 31 -887
rect -31 -927 31 -921
rect 97 -887 159 -881
rect 97 -921 109 -887
rect 147 -921 159 -887
rect 97 -927 159 -921
rect 225 -887 287 -881
rect 225 -921 237 -887
rect 275 -921 287 -887
rect 225 -927 287 -921
rect 353 -887 415 -881
rect 353 -921 365 -887
rect 403 -921 415 -887
rect 353 -927 415 -921
rect 481 -887 543 -881
rect 481 -921 493 -887
rect 531 -921 543 -887
rect 481 -927 543 -921
rect 609 -887 671 -881
rect 609 -921 621 -887
rect 659 -921 671 -887
rect 609 -927 671 -921
rect 737 -887 799 -881
rect 737 -921 749 -887
rect 787 -921 799 -887
rect 737 -927 799 -921
rect 865 -887 927 -881
rect 865 -921 877 -887
rect 915 -921 927 -887
rect 865 -927 927 -921
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1074 -1006 1074 1006
string parameters w 8.4 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
