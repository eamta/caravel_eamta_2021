magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect 667 1042 702 1076
rect 129 919 187 925
rect 129 885 141 919
rect 129 879 187 885
rect 316 804 386 1042
rect 668 1023 702 1042
rect 687 980 702 1023
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect -53 766 386 804
rect 466 766 500 800
rect 554 766 588 800
rect 668 766 702 980
rect 721 989 756 1023
rect 721 766 755 989
rect 2512 957 2547 991
rect 2513 938 2547 957
rect 867 921 925 927
rect 867 887 879 921
rect 1037 898 1071 927
rect 867 881 925 887
rect 1037 862 1107 898
rect 1037 828 1125 862
rect 1405 828 1440 862
rect 1828 845 1863 863
rect 1037 804 1124 828
rect 1406 809 1440 828
rect 1792 830 1863 845
rect 1425 804 1440 809
rect 1459 804 1775 809
rect 1792 804 1862 830
rect 835 766 869 800
rect 923 766 957 800
rect 1037 766 1862 804
rect 1952 766 2054 796
rect 2163 766 2178 864
rect -53 762 2106 766
rect -53 735 2058 762
rect -53 732 2106 735
rect 2163 732 2182 766
rect -53 660 386 732
rect 454 713 494 732
rect 532 713 600 732
rect 470 694 584 700
rect 510 678 554 684
rect 479 666 591 678
rect 398 660 414 666
rect 479 663 594 666
rect -53 650 424 660
rect -53 640 430 650
rect -53 634 386 640
rect -53 626 378 634
rect -53 547 369 626
rect 380 564 386 634
rect 404 634 430 640
rect 404 616 424 634
rect 494 632 594 663
rect 599 650 620 678
rect 668 660 702 732
rect 721 678 755 732
rect 860 704 869 732
rect 806 684 835 690
rect 852 684 881 704
rect 806 678 881 684
rect 636 650 702 660
rect 630 640 702 650
rect 630 634 667 640
rect 494 626 556 632
rect 494 616 532 626
rect 574 600 594 632
rect 646 616 667 634
rect 668 634 702 640
rect 668 626 680 634
rect 681 626 702 634
rect 668 616 702 626
rect 668 564 680 616
rect 380 553 425 564
rect 352 530 356 547
rect 380 541 414 553
rect 369 530 425 541
rect 474 530 620 564
rect 635 553 680 564
rect 646 541 680 553
rect 681 541 702 616
rect 635 530 702 541
rect 706 530 756 678
rect 806 672 869 678
rect 806 666 835 672
rect 860 656 869 672
rect 894 661 903 732
rect 944 684 969 732
rect 923 678 969 684
rect 1037 678 1862 732
rect 2018 712 2036 732
rect 1908 694 2098 709
rect 2030 681 2040 685
rect 923 672 957 678
rect 883 660 911 661
rect 998 660 1023 678
rect 829 600 840 647
rect 882 619 940 660
rect 867 613 940 619
rect 863 579 940 613
rect 1037 650 1874 678
rect 1930 660 1983 681
rect 2018 678 2070 681
rect 2019 669 2070 678
rect 2024 666 2070 669
rect 2144 678 2182 732
rect 1996 661 2006 666
rect 1892 650 1983 660
rect 1988 650 2006 661
rect 867 573 929 579
rect 882 563 929 573
rect 219 498 347 519
rect 474 498 532 519
rect 721 511 755 530
rect 1037 511 1862 650
rect 1886 640 2006 650
rect 1886 634 1921 640
rect 1902 616 1921 634
rect 1930 616 2006 640
rect 721 506 940 511
rect 998 506 1862 511
rect 721 498 1862 506
rect 1930 516 1936 616
rect 1942 516 1976 616
rect 1996 600 2006 616
rect 2030 650 2064 666
rect 2030 616 2094 650
rect 1930 513 1976 516
rect 2030 513 2064 616
rect 1930 501 1951 513
rect 298 482 300 488
rect 472 482 488 488
rect 256 472 268 482
rect 298 472 310 482
rect 446 472 457 482
rect 472 473 498 482
rect 721 477 1845 498
rect 487 472 498 473
rect 1054 472 1845 477
rect 250 462 278 472
rect 288 462 316 472
rect 250 456 276 462
rect 266 448 276 456
rect 290 456 316 462
rect 440 463 504 472
rect 440 462 467 463
rect 477 462 504 463
rect 440 456 466 462
rect 290 448 310 456
rect 266 438 310 448
rect 456 448 466 456
rect 478 456 504 462
rect 478 448 498 456
rect 456 438 467 448
rect 477 438 498 448
rect 687 443 1845 472
rect 1988 470 2018 501
rect 284 428 310 438
rect 487 428 498 438
rect 284 422 300 428
rect 487 422 488 428
rect 90 404 106 410
rect 282 404 298 410
rect 562 404 564 410
rect 72 394 116 404
rect 256 394 308 404
rect 520 394 532 404
rect 562 394 574 404
rect 1054 394 1845 443
rect 1970 460 2018 470
rect 2020 460 2067 501
rect 1970 420 2067 460
rect 1970 414 2032 420
rect 1851 394 1862 405
rect 1970 404 2018 414
rect 72 384 122 394
rect 96 378 122 384
rect 250 384 314 394
rect 250 378 276 384
rect 96 370 116 378
rect 72 360 116 370
rect 266 370 276 378
rect 288 378 314 384
rect 514 384 542 394
rect 552 384 580 394
rect 1054 388 1862 394
rect 514 378 540 384
rect 266 360 278 370
rect 288 360 308 378
rect 530 370 540 378
rect 554 378 580 384
rect 554 370 574 378
rect 530 360 574 370
rect 1322 370 1332 388
rect 1342 384 1370 388
rect 1344 378 1370 384
rect 1344 370 1364 378
rect 1322 360 1364 370
rect 90 350 116 360
rect 548 350 574 360
rect 1338 350 1364 360
rect 1423 352 1862 388
rect 2144 352 2194 678
rect 90 344 106 350
rect 548 344 564 350
rect 715 318 843 349
rect 1338 344 1354 350
rect 1423 341 1947 352
rect 1423 336 1936 341
rect 1960 336 2194 352
rect 1423 335 2194 336
rect 1828 318 2194 335
rect 2197 318 2231 918
rect 2343 889 2401 895
rect 2343 855 2355 889
rect 2343 849 2401 855
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 794 312 796 318
rect 752 302 764 312
rect 794 302 806 312
rect 2136 310 2138 316
rect 2094 302 2106 310
rect 2136 302 2148 310
rect 746 292 774 302
rect 784 292 812 302
rect 746 286 772 292
rect 762 278 772 286
rect 786 286 812 292
rect 786 278 806 286
rect 1794 284 2154 302
rect 2197 284 2212 318
rect 150 236 160 270
rect 174 236 194 270
rect 762 268 774 278
rect 784 268 806 278
rect 2104 278 2114 284
rect 2128 278 2148 284
rect 2104 268 2116 278
rect 2126 268 2148 278
rect 794 258 806 268
rect 2136 258 2148 268
rect 2532 265 2547 938
rect 2566 904 2601 938
rect 2566 265 2600 904
rect 2712 836 2770 842
rect 2712 802 2724 836
rect 2712 796 2770 802
rect 2882 633 2916 651
rect 4726 639 4761 673
rect 2882 597 2952 633
rect 4727 620 4761 639
rect 2899 563 2970 597
rect 3250 563 3285 597
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 794 252 796 258
rect 2136 252 2138 258
rect 1086 244 1088 250
rect 2048 244 2052 250
rect 1044 234 1056 244
rect 1086 234 1098 244
rect 2048 234 2062 244
rect 138 224 196 228
rect 380 200 390 234
rect 404 200 424 234
rect 1038 224 1066 234
rect 1076 224 1104 234
rect 1038 218 1064 224
rect 1054 210 1064 218
rect 1078 218 1104 224
rect 1078 210 1098 218
rect 1054 200 1066 210
rect 1076 200 1098 210
rect 1436 200 1446 234
rect 1460 200 1480 234
rect 2018 200 2028 234
rect 2038 224 2068 234
rect 2566 231 2581 265
rect 2042 218 2068 224
rect 2042 210 2062 218
rect 2038 200 2062 210
rect 110 196 200 200
rect 1086 190 1098 200
rect 2048 190 2062 200
rect 2899 212 2969 563
rect 3251 544 3285 563
rect 3081 495 3139 501
rect 3081 461 3093 495
rect 3081 455 3139 461
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 1086 184 1088 190
rect 2048 184 2052 190
rect 998 176 1014 182
rect 2899 176 2952 212
rect 980 166 1024 176
rect 980 156 1030 166
rect 1004 150 1030 156
rect 1004 148 1024 150
rect 980 132 1024 148
rect 1170 148 1180 166
rect 1170 132 1182 148
rect 1194 132 1214 166
rect 3270 159 3285 544
rect 3304 510 3339 544
rect 3619 510 3654 544
rect 4042 527 4077 545
rect 3304 159 3338 510
rect 3620 491 3654 510
rect 4006 512 4077 527
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 998 122 1024 132
rect 3304 125 3319 159
rect 998 116 1014 122
rect 112 82 116 110
rect 150 58 160 82
rect 174 58 194 82
rect 150 48 194 58
rect 210 48 222 110
rect 342 82 356 110
rect 608 82 620 110
rect 380 58 394 82
rect 404 58 424 82
rect 380 48 424 58
rect 646 58 658 82
rect 670 58 690 82
rect 646 48 690 58
rect 706 48 718 110
rect 1132 82 1144 110
rect 1398 82 1410 110
rect 1170 58 1182 82
rect 1194 58 1214 82
rect 1170 48 1214 58
rect 1436 58 1448 82
rect 1460 58 1480 82
rect 1436 48 1480 58
rect 1496 48 1508 110
rect 1628 82 1642 110
rect 1666 58 1680 82
rect 1690 58 1710 82
rect 1666 48 1710 58
rect 1728 48 1738 110
rect 1864 82 1874 110
rect 1902 58 1912 82
rect 1926 58 1946 82
rect 1902 48 1946 58
rect 1960 48 1974 110
rect 3639 106 3654 491
rect 3673 457 3708 491
rect 3673 106 3707 457
rect 3819 389 3877 395
rect 3819 355 3831 389
rect 3819 349 3877 355
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4006 53 4076 512
rect 4188 444 4246 450
rect 4188 410 4200 444
rect 4188 404 4246 410
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 168 38 194 48
rect 398 38 424 48
rect 664 38 690 48
rect 1188 38 1214 48
rect 1454 38 1480 48
rect 1684 38 1710 48
rect 1920 38 1946 48
rect 168 32 184 38
rect 398 32 414 38
rect 664 32 680 38
rect 1188 32 1204 38
rect 1454 32 1470 38
rect 1684 32 1700 38
rect 1920 32 1936 38
rect 4006 17 4059 53
rect 4377 0 4392 546
rect 4411 0 4445 600
rect 4557 571 4615 577
rect 4557 537 4569 571
rect 4557 531 4615 537
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 620
rect 4780 586 4815 620
rect 4780 -53 4814 586
rect 4926 518 4984 524
rect 4926 484 4938 518
rect 4926 478 4984 484
rect 5096 315 5130 333
rect 5096 279 5166 315
rect 5113 245 5184 279
rect 5464 245 5499 279
rect 5887 262 5922 280
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5113 -106 5183 245
rect 5465 226 5499 245
rect 5851 247 5922 262
rect 5295 177 5353 183
rect 5295 143 5307 177
rect 5295 137 5353 143
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5113 -142 5166 -106
rect 5484 -159 5499 226
rect 5518 192 5553 226
rect 5518 -159 5552 192
rect 5664 124 5722 130
rect 5664 90 5676 124
rect 5664 84 5722 90
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5518 -193 5533 -159
rect 5851 -212 5921 247
rect 6033 179 6091 185
rect 6033 145 6045 179
rect 6203 156 6237 174
rect 6033 139 6091 145
rect 6203 120 6273 156
rect 6220 86 6291 120
rect 6571 86 6606 120
rect 6994 103 7029 121
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5851 -248 5904 -212
rect 6220 -265 6290 86
rect 6572 67 6606 86
rect 6958 88 7029 103
rect 7309 88 7344 122
rect 6402 18 6460 24
rect 6402 -16 6414 18
rect 6402 -22 6460 -16
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6220 -301 6273 -265
rect 6591 -318 6606 67
rect 6625 33 6660 67
rect 6625 -318 6659 33
rect 6771 -35 6829 -29
rect 6771 -69 6783 -35
rect 6771 -75 6829 -69
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6625 -352 6640 -318
rect 6958 -371 7028 88
rect 7310 69 7344 88
rect 7140 20 7198 26
rect 7140 -14 7152 20
rect 7140 -20 7198 -14
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6958 -407 7011 -371
rect 7329 -424 7344 69
rect 7363 35 7398 69
rect 7363 -424 7397 35
rect 7509 -33 7567 -27
rect 7509 -67 7521 -33
rect 7679 -56 7713 -38
rect 7509 -73 7567 -67
rect 7679 -92 7749 -56
rect 7696 -126 7767 -92
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7363 -458 7378 -424
rect 7696 -477 7766 -126
rect 7878 -194 7936 -188
rect 7878 -228 7890 -194
rect 7878 -234 7936 -228
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7696 -513 7749 -477
<< nwell >>
rect -66 280 2230 804
<< nmos >>
rect 28 20 58 110
rect 268 20 298 110
rect 532 20 562 110
rect 764 20 794 110
rect 852 20 882 110
rect 1056 20 1086 110
rect 1322 20 1352 110
rect 1554 20 1584 110
rect 1786 20 1816 110
rect 2018 20 2048 110
rect 2106 20 2136 110
<< pmos >>
rect 28 498 58 678
rect 268 498 298 678
rect 532 498 562 678
rect 764 318 794 678
rect 852 318 882 678
rect 1056 498 1086 678
rect 1322 498 1352 678
rect 1554 498 1584 678
rect 1786 498 1816 678
rect 2018 318 2048 678
rect 2106 318 2136 678
<< ndiff >>
rect -30 82 28 110
rect -30 48 -18 82
rect 16 48 28 82
rect -30 20 28 48
rect 58 82 116 110
rect 58 48 70 82
rect 104 48 116 82
rect 210 82 268 110
rect 210 48 222 82
rect 256 48 268 82
rect 58 20 116 48
rect 210 20 268 48
rect 298 82 356 110
rect 298 48 310 82
rect 344 48 356 82
rect 474 82 532 110
rect 474 48 486 82
rect 520 48 532 82
rect 298 20 356 48
rect 474 20 532 48
rect 562 82 620 110
rect 562 48 574 82
rect 608 48 620 82
rect 706 82 764 110
rect 706 48 718 82
rect 752 48 764 82
rect 562 20 620 48
rect 706 20 764 48
rect 794 82 852 110
rect 794 48 806 82
rect 840 48 852 82
rect 794 20 852 48
rect 882 82 940 110
rect 882 48 894 82
rect 928 48 940 82
rect 882 20 940 48
rect 998 82 1056 110
rect 998 48 1010 82
rect 1044 48 1056 82
rect 998 20 1056 48
rect 1086 82 1144 110
rect 1086 48 1098 82
rect 1132 48 1144 82
rect 1264 82 1322 110
rect 1264 48 1276 82
rect 1310 48 1322 82
rect 1086 20 1144 48
rect 1264 20 1322 48
rect 1352 82 1410 110
rect 1352 48 1364 82
rect 1398 48 1410 82
rect 1496 82 1554 110
rect 1496 48 1508 82
rect 1542 48 1554 82
rect 1352 20 1410 48
rect 1496 20 1554 48
rect 1584 82 1642 110
rect 1584 48 1596 82
rect 1630 48 1642 82
rect 1728 82 1786 110
rect 1728 48 1740 82
rect 1774 48 1786 82
rect 1584 20 1642 48
rect 1728 20 1786 48
rect 1816 82 1874 110
rect 1816 48 1828 82
rect 1862 48 1874 82
rect 1960 82 2018 110
rect 1960 48 1972 82
rect 2006 48 2018 82
rect 1816 20 1874 48
rect 1960 20 2018 48
rect 2048 82 2106 110
rect 2048 48 2060 82
rect 2094 48 2106 82
rect 2048 20 2106 48
rect 2136 82 2194 110
rect 2136 48 2148 82
rect 2182 48 2194 82
rect 2136 20 2194 48
<< pdiff >>
rect -30 650 28 678
rect -30 616 -18 650
rect 16 616 28 650
rect -30 498 28 616
rect 58 650 116 678
rect 210 650 268 678
rect 58 616 70 650
rect 104 616 116 650
rect 58 498 116 616
rect 210 616 222 650
rect 256 616 268 650
rect 210 498 268 616
rect 298 650 356 678
rect 474 650 532 678
rect 298 616 310 650
rect 344 616 356 650
rect 298 498 356 616
rect 474 616 486 650
rect 520 616 532 650
rect 474 498 532 616
rect 562 650 620 678
rect 706 650 764 678
rect 562 616 574 650
rect 608 616 620 650
rect 562 498 620 616
rect 706 616 718 650
rect 752 616 764 650
rect 706 318 764 616
rect 794 650 852 678
rect 794 616 806 650
rect 840 616 852 650
rect 794 318 852 616
rect 882 650 940 678
rect 882 616 894 650
rect 928 616 940 650
rect 882 318 940 616
rect 998 650 1056 678
rect 998 616 1010 650
rect 1044 616 1056 650
rect 998 498 1056 616
rect 1086 650 1144 678
rect 1264 650 1322 678
rect 1086 616 1098 650
rect 1132 616 1144 650
rect 1086 498 1144 616
rect 1264 616 1276 650
rect 1310 616 1322 650
rect 1264 498 1322 616
rect 1352 650 1410 678
rect 1496 650 1554 678
rect 1352 616 1364 650
rect 1398 616 1410 650
rect 1352 498 1410 616
rect 1496 616 1508 650
rect 1542 616 1554 650
rect 1496 498 1554 616
rect 1584 650 1642 678
rect 1728 650 1786 678
rect 1584 616 1596 650
rect 1630 616 1642 650
rect 1584 498 1642 616
rect 1728 616 1740 650
rect 1774 616 1786 650
rect 1728 498 1786 616
rect 1816 650 1874 678
rect 1960 650 2018 678
rect 1816 616 1828 650
rect 1862 616 1874 650
rect 1816 498 1874 616
rect 1960 616 1972 650
rect 2006 616 2018 650
rect 1960 318 2018 616
rect 2048 650 2106 678
rect 2048 616 2060 650
rect 2094 616 2106 650
rect 2048 318 2106 616
rect 2136 650 2194 678
rect 2136 616 2148 650
rect 2182 616 2194 650
rect 2136 318 2194 616
<< ndiffc >>
rect -18 48 16 82
rect 70 48 104 82
rect 222 48 256 82
rect 310 48 344 82
rect 486 48 520 82
rect 574 48 608 82
rect 718 48 752 82
rect 806 48 840 82
rect 894 48 928 82
rect 1010 48 1044 82
rect 1098 48 1132 82
rect 1276 48 1310 82
rect 1364 48 1398 82
rect 1508 48 1542 82
rect 1596 48 1630 82
rect 1740 48 1774 82
rect 1828 48 1862 82
rect 1972 48 2006 82
rect 2060 48 2094 82
rect 2148 48 2182 82
<< pdiffc >>
rect -18 616 16 650
rect 70 616 104 650
rect 222 616 256 650
rect 310 616 344 650
rect 486 616 520 650
rect 574 616 608 650
rect 718 616 752 650
rect 806 616 840 650
rect 894 616 928 650
rect 1010 616 1044 650
rect 1098 616 1132 650
rect 1276 616 1310 650
rect 1364 616 1398 650
rect 1508 616 1542 650
rect 1596 616 1630 650
rect 1740 616 1774 650
rect 1828 616 1862 650
rect 1972 616 2006 650
rect 2060 616 2094 650
rect 2148 616 2182 650
<< psubdiff >>
rect 14 -68 58 -34
rect 2106 -68 2154 -34
<< nsubdiff >>
rect 4 732 58 766
rect 2106 732 2154 766
<< psubdiffcont >>
rect 58 -68 2106 -34
<< nsubdiffcont >>
rect 58 732 2106 766
<< poly >>
rect 28 678 58 704
rect 268 678 298 704
rect 532 678 562 704
rect 764 678 794 704
rect 852 678 882 704
rect 1056 678 1086 704
rect 1322 678 1352 704
rect 1554 678 1584 704
rect 1786 678 1816 704
rect 2018 678 2048 704
rect 2106 678 2136 704
rect 28 394 58 498
rect 28 360 72 394
rect 28 110 58 360
rect 150 270 184 616
rect 268 472 298 498
rect 150 82 184 236
rect 268 110 298 360
rect 380 234 414 616
rect 457 472 487 473
rect 457 312 487 438
rect 532 394 562 498
rect 457 282 562 312
rect 380 82 414 200
rect 532 110 562 282
rect 646 82 680 616
rect 764 302 794 318
rect 764 110 794 268
rect 852 166 882 318
rect 1056 234 1086 498
rect 852 132 980 166
rect 852 110 882 132
rect 1056 110 1086 200
rect 1170 166 1204 616
rect 1246 314 1280 438
rect 1322 394 1352 498
rect 1246 280 1352 314
rect 1170 82 1204 132
rect 1322 110 1352 280
rect 1436 234 1470 616
rect 1554 472 1584 498
rect 1554 394 1584 396
rect 1436 82 1470 200
rect 1554 110 1584 360
rect 1666 82 1700 616
rect 1786 394 1816 498
rect 1902 394 1936 616
rect 1786 360 1936 394
rect 1786 110 1816 360
rect 1902 82 1936 360
rect 2018 234 2048 318
rect 2106 300 2136 318
rect 2018 110 2048 200
rect 2106 110 2136 268
rect 28 -6 58 20
rect 268 -6 298 20
rect 532 -6 562 20
rect 764 -6 794 20
rect 852 -6 882 20
rect 1056 -6 1086 20
rect 1322 -6 1352 20
rect 1554 -6 1584 20
rect 1786 -6 1816 20
rect 2018 -6 2048 20
rect 2106 -6 2136 20
<< polycont >>
rect 150 616 184 650
rect 72 360 106 394
rect 380 616 414 650
rect 266 438 300 472
rect 266 360 298 394
rect 150 236 184 270
rect 646 616 680 650
rect 456 438 488 472
rect 530 360 564 394
rect 380 200 414 234
rect 150 48 184 82
rect 380 48 414 82
rect 1170 616 1204 650
rect 762 268 796 302
rect 1054 200 1088 234
rect 980 132 1014 166
rect 1436 616 1470 650
rect 1246 438 1280 472
rect 1322 360 1354 394
rect 1170 132 1204 166
rect 646 48 680 82
rect 1666 616 1700 650
rect 1552 438 1586 472
rect 1552 360 1586 394
rect 1436 200 1470 234
rect 1170 48 1204 82
rect 1436 48 1470 82
rect 1902 616 1936 650
rect 1666 48 1700 82
rect 2104 268 2138 300
rect 2018 200 2052 234
rect 1902 48 1936 82
<< locali >>
rect 14 732 58 766
rect 2106 732 2182 766
rect -18 650 16 666
rect -18 472 16 616
rect 70 650 104 732
rect 70 600 104 616
rect 150 650 256 666
rect 184 616 222 650
rect 150 600 256 616
rect 310 650 520 666
rect 344 616 380 650
rect 414 616 486 650
rect 310 600 520 616
rect 574 650 752 666
rect 608 616 646 650
rect 680 616 718 650
rect 574 600 752 616
rect 806 650 840 666
rect 806 600 840 616
rect 894 650 928 732
rect 894 600 928 616
rect 1010 650 1044 732
rect 1010 600 1044 616
rect 1098 650 1310 666
rect 1132 616 1170 650
rect 1204 616 1276 650
rect 1098 600 1310 616
rect 1364 650 1542 666
rect 1398 616 1436 650
rect 1470 616 1508 650
rect 1364 600 1542 616
rect 1596 650 1774 666
rect 1630 616 1666 650
rect 1700 616 1740 650
rect 1596 600 1774 616
rect 1828 650 1862 732
rect 1828 600 1862 616
rect 1902 650 2006 666
rect 1936 616 1972 650
rect 1902 600 2006 616
rect 2060 650 2094 666
rect 2060 600 2094 616
rect 2148 650 2182 732
rect 2148 600 2182 616
rect -18 438 266 472
rect 300 438 456 472
rect 488 438 1246 472
rect 1280 438 1552 472
rect 1586 438 1602 472
rect -18 82 16 438
rect 56 360 72 394
rect 106 360 266 394
rect 298 360 530 394
rect 564 360 1322 394
rect 1354 360 1552 394
rect 1586 360 1602 394
rect 150 270 184 286
rect 746 268 762 302
rect 796 300 2154 302
rect 796 268 2104 300
rect 2138 268 2154 300
rect 150 220 184 236
rect 364 200 380 234
rect 414 200 1054 234
rect 1088 200 1104 234
rect 1420 200 1436 234
rect 1470 200 2018 234
rect 2052 200 2068 234
rect 718 132 928 166
rect 964 132 980 166
rect 1014 132 1170 166
rect 1204 132 1220 166
rect 1972 132 2182 166
rect 718 98 752 132
rect -18 32 16 48
rect 70 82 104 98
rect 70 -34 104 48
rect 150 82 256 98
rect 184 48 222 82
rect 150 32 256 48
rect 310 82 520 98
rect 344 48 380 82
rect 414 48 486 82
rect 310 32 520 48
rect 574 82 752 98
rect 608 48 646 82
rect 680 48 718 82
rect 574 32 752 48
rect 806 82 840 98
rect 806 -34 840 48
rect 894 82 928 132
rect 1972 98 2006 132
rect 894 32 928 48
rect 1010 82 1044 98
rect 1010 -34 1044 48
rect 1098 82 1310 98
rect 1132 48 1170 82
rect 1204 48 1276 82
rect 1098 32 1310 48
rect 1364 82 1542 98
rect 1398 48 1436 82
rect 1470 48 1508 82
rect 1364 32 1542 48
rect 1596 82 1774 98
rect 1630 48 1666 82
rect 1700 48 1740 82
rect 1596 32 1774 48
rect 1828 82 1862 98
rect 1828 -34 1862 48
rect 1902 82 2006 98
rect 1936 48 1972 82
rect 1902 32 2006 48
rect 2060 82 2094 98
rect 2060 -34 2094 48
rect 2148 82 2182 132
rect 2148 32 2182 48
rect 14 -68 58 -34
rect 2106 -68 2138 -34
<< viali >>
rect 58 732 2106 766
rect 72 360 106 394
rect 150 236 184 270
rect 762 268 796 302
rect 1666 48 1700 82
rect 1902 48 1936 82
rect 58 -68 2106 -34
<< metal1 >>
rect -66 766 2230 804
rect -66 732 58 766
rect 2106 732 2230 766
rect -66 694 2230 732
rect 60 394 118 406
rect 60 360 72 394
rect 106 360 118 394
rect 60 348 118 360
rect 750 302 808 314
rect 138 270 196 282
rect 138 236 150 270
rect 184 236 196 270
rect 750 268 762 302
rect 796 268 808 302
rect 750 256 808 268
rect 138 224 196 236
rect 0 4 200 200
rect 1654 82 1714 94
rect 1654 48 1666 82
rect 1700 48 1714 82
rect 1654 36 1714 48
rect 1890 82 1948 94
rect 1890 48 1902 82
rect 1936 48 1948 82
rect 1890 36 1948 48
rect -66 -34 2230 4
rect -66 -68 58 -34
rect 2106 -68 2230 -34
rect -66 -106 2230 -68
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use sky130_fd_pr__pfet_01v8_XYCVAL  XM6
timestamp 1624053917
transform 1 0 2372 0 1 628
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM7
timestamp 1624053917
transform 1 0 2741 0 1 575
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM8
timestamp 1624053917
transform 1 0 3110 0 1 378
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM10
timestamp 1624053917
transform 1 0 3848 0 1 272
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM14
timestamp 1624053917
transform 1 0 5324 0 1 60
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM13
timestamp 1624053917
transform 1 0 4955 0 1 257
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM12
timestamp 1624053917
transform 1 0 4586 0 1 310
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XSLFBL  XM11
timestamp 1624053917
transform 1 0 4217 0 1 273
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM18
timestamp 1624053917
transform 1 0 6800 0 1 -152
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM17
timestamp 1624053917
transform 1 0 6431 0 1 -99
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM16
timestamp 1624053917
transform 1 0 6062 0 1 8
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM15
timestamp 1624053917
transform 1 0 5693 0 1 7
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM21
timestamp 1624053917
transform 1 0 7907 0 1 -311
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM20
timestamp 1624053917
transform 1 0 7538 0 1 -204
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM19
timestamp 1624053917
transform 1 0 7169 0 1 -151
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM0
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM3
timestamp 1624053917
transform 1 0 1265 0 1 643
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1624053917
transform 1 0 1634 0 1 590
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
<< labels >>
rlabel metal1 1072 -106 1072 -106 5 VSS
rlabel metal1 1070 804 1070 804 1 VDD
rlabel metal1 88 348 88 348 5 CLK
rlabel metal1 138 252 138 252 7 D
rlabel metal1 780 256 780 256 5 CLR
rlabel metal1 1684 36 1684 36 5 Qb
rlabel metal1 1920 36 1920 36 5 Q
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Q
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 D
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLK
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLR
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Qb
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 VDD
port 9 nsew
<< end >>
