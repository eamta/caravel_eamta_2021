magic
tech sky130A
magscale 1 2
timestamp 1619545672
<< nwell >>
rect -67 913 22681 1152
rect -67 895 14887 913
rect -67 890 11553 895
rect -67 685 8569 890
rect 14241 845 14887 895
rect 14241 821 14480 845
rect 14485 821 14887 845
rect -67 9 8251 685
rect -67 -12 519 9
rect 796 -12 8251 9
rect 14241 176 14887 821
rect 14241 139 14781 176
rect 14818 139 14887 176
rect 796 -3837 832 -308
rect 14241 -990 14887 139
rect 20846 -990 22681 913
rect 796 -7373 819 -3837
<< pwell >>
rect 11043 -10013 22905 -7071
rect 793 -10164 22905 -10013
<< pdiff >>
rect 7133 -2308 7167 -2296
rect 7669 -2308 7703 -2296
rect 7133 -3696 7167 -3684
rect 7669 -3696 7703 -3684
rect 1237 -3997 1271 -3985
rect 1773 -3997 1807 -3985
rect 2309 -3997 2343 -3985
rect 2845 -3997 2879 -3985
rect 3381 -3997 3415 -3985
rect 4453 -3997 4487 -3985
rect 4989 -3997 5023 -3985
rect 5525 -3997 5559 -3985
rect 6061 -3997 6095 -3985
rect 6597 -3997 6631 -3985
rect 7133 -3997 7167 -3985
rect 7669 -3997 7703 -3985
rect 1237 -5385 1271 -5373
rect 1773 -5385 1807 -5373
rect 2309 -5385 2343 -5373
rect 2845 -5385 2879 -5373
rect 3381 -5385 3415 -5373
rect 4453 -5385 4487 -5373
rect 4989 -5385 5023 -5373
rect 5525 -5385 5559 -5373
rect 6061 -5385 6095 -5373
rect 6597 -5385 6631 -5373
rect 7133 -5385 7167 -5373
rect 7669 -5385 7703 -5373
rect 1237 -5837 1271 -5825
rect 1773 -5837 1807 -5825
rect 2309 -5837 2343 -5825
rect 2845 -5837 2879 -5825
rect 3381 -5837 3415 -5825
rect 3917 -5837 3951 -5825
rect 4453 -5837 4487 -5825
rect 4989 -5837 5023 -5825
rect 5525 -5837 5559 -5825
rect 6061 -5837 6095 -5825
rect 6597 -5837 6631 -5825
rect 7133 -5837 7167 -5825
rect 7669 -5837 7703 -5825
rect 1237 -7225 1271 -7213
rect 1773 -7225 1807 -7213
rect 2309 -7225 2343 -7213
rect 2845 -7225 2879 -7213
rect 3381 -7225 3415 -7213
rect 3917 -7225 3951 -7213
rect 4453 -7225 4487 -7213
rect 4989 -7225 5023 -7213
rect 5525 -7225 5559 -7213
rect 6061 -7225 6095 -7213
rect 6597 -7225 6631 -7213
rect 7133 -7225 7167 -7213
rect 7669 -7225 7703 -7213
<< psubdiff >>
rect 11119 -8354 12657 -8330
rect 11119 -9919 12657 -9895
rect 812 -10122 836 -10066
rect 10951 -10122 10975 -10066
rect 12666 -10122 12690 -9975
rect 22854 -10122 22878 -9975
<< nsubdiff >>
rect 31 1089 8226 1091
rect 31 973 66 1089
rect 8178 973 8226 1089
rect 31 970 8226 973
rect 8280 1085 20805 1086
rect 8280 970 8316 1085
rect 20769 970 20805 1085
rect 8280 969 20805 970
rect 20889 1002 22604 1060
rect 20889 -790 20945 1002
rect 22549 -790 22604 1002
rect 20889 -842 22604 -790
<< psubdiffcont >>
rect 11119 -9895 12657 -8354
rect 836 -10122 10951 -10066
rect 12690 -10122 22854 -9975
<< nsubdiffcont >>
rect 66 973 8178 1089
rect 8316 970 20769 1085
rect 951 -378 7721 -344
rect 7783 -1943 7817 -441
rect 20945 -790 22549 1002
rect 7783 -3711 7817 -2209
<< locali >>
rect 42 973 66 1089
rect 8178 973 8216 1089
rect 8290 970 8316 1085
rect 20769 970 20796 1085
rect 20909 1002 22587 1042
rect 20909 -790 20945 1002
rect 22549 -790 22587 1002
rect 20909 -823 22587 -790
rect 7133 -2308 7167 -2292
rect 7669 -2308 7703 -2292
rect 7133 -3700 7167 -3684
rect 7669 -3700 7703 -3684
rect 1237 -3997 1271 -3981
rect 1773 -3997 1807 -3981
rect 2309 -3997 2343 -3981
rect 2845 -3997 2879 -3981
rect 3381 -3997 3415 -3981
rect 3917 -3997 3951 -3981
rect 4453 -3997 4487 -3981
rect 4989 -3997 5023 -3981
rect 5525 -3997 5559 -3981
rect 6061 -3997 6095 -3981
rect 6597 -3997 6631 -3981
rect 7133 -3997 7167 -3981
rect 7669 -3997 7703 -3981
rect 1237 -5389 1271 -5373
rect 1773 -5389 1807 -5373
rect 2309 -5389 2343 -5373
rect 2845 -5389 2879 -5373
rect 3381 -5389 3415 -5373
rect 3917 -5389 3951 -5373
rect 4453 -5389 4487 -5373
rect 4989 -5389 5023 -5373
rect 5525 -5389 5559 -5373
rect 6061 -5389 6095 -5373
rect 6597 -5389 6631 -5373
rect 7133 -5389 7167 -5373
rect 7669 -5389 7703 -5373
rect 1237 -5837 1271 -5821
rect 1773 -5837 1807 -5821
rect 2309 -5837 2343 -5821
rect 2845 -5837 2879 -5821
rect 3381 -5837 3415 -5821
rect 3917 -5837 3951 -5821
rect 4453 -5837 4487 -5821
rect 4989 -5837 5023 -5821
rect 5525 -5837 5559 -5821
rect 6061 -5837 6095 -5821
rect 6597 -5837 6631 -5821
rect 7133 -5837 7167 -5821
rect 7669 -5837 7703 -5821
rect 1237 -7229 1271 -7213
rect 1773 -7229 1807 -7213
rect 2309 -7229 2343 -7213
rect 2845 -7229 2879 -7213
rect 3381 -7229 3415 -7213
rect 3917 -7229 3951 -7213
rect 4453 -7229 4487 -7213
rect 4989 -7229 5023 -7213
rect 5525 -7229 5559 -7213
rect 6061 -7229 6095 -7213
rect 6597 -7229 6631 -7213
rect 7133 -7229 7167 -7213
rect 7669 -7229 7703 -7213
rect 11119 -8354 12657 -8338
rect 11119 -9911 12657 -9895
rect 820 -10122 836 -10066
rect 10951 -10122 10967 -10066
rect 12674 -10122 12690 -9975
rect 22854 -10122 22870 -9975
<< viali >>
rect 66 973 8178 1089
rect 8316 970 20769 1085
rect 8384 858 14354 892
rect 14766 858 20736 892
rect 2160 708 8130 742
rect 65 557 1905 591
rect -31 145 3 494
rect 1967 183 2001 494
rect 2064 183 2098 645
rect 8192 178 8226 645
rect 8288 179 8322 795
rect 20798 93 20832 795
rect 951 -378 7721 -344
rect 855 -1860 889 -441
rect 7783 -1943 7817 -441
rect 8288 -857 8322 -155
rect 20798 -857 20832 -155
rect 20945 -790 22549 1002
rect 8384 -954 14354 -920
rect 14766 -954 20736 -920
rect 855 -3711 889 -2292
rect 7783 -3711 7817 -2209
rect 855 -5389 889 -3970
rect 7783 -5472 7817 -3970
rect 855 -7240 889 -5821
rect 7783 -7240 7817 -5738
rect 951 -7337 7721 -7303
rect 22835 -7660 22869 -7204
rect 830 -9896 864 -7702
rect 5876 -9896 5910 -7800
rect 5964 -9896 5998 -7800
rect 11010 -9896 11044 -7702
rect 11119 -9895 12657 -8354
rect 22835 -8380 22869 -7924
rect 22835 -9100 22869 -8644
rect 22835 -9820 22869 -9364
rect 836 -10122 10951 -10066
rect 12690 -10122 22854 -9975
<< metal1 >>
rect 35 1091 22578 1095
rect -31 1089 22578 1091
rect -31 973 66 1089
rect 8178 1085 22578 1089
rect 8178 973 8316 1085
rect -31 970 8316 973
rect 20769 1002 22578 1085
rect 20769 970 20945 1002
rect -31 892 20945 970
rect -31 858 8384 892
rect 14354 858 14766 892
rect 20736 858 20945 892
rect -31 847 20945 858
rect -31 807 8323 847
rect 8467 846 20945 847
rect -31 795 8328 807
rect -31 742 8288 795
rect -31 708 2160 742
rect 8130 708 8288 742
rect -31 698 8288 708
rect -31 645 2104 698
rect -31 591 2064 645
rect -31 557 65 591
rect 1905 557 2064 591
rect -31 543 2064 557
rect -31 506 9 543
rect -37 494 9 506
rect -37 145 -31 494
rect 3 145 9 494
rect 83 472 117 543
rect 319 477 353 543
rect 555 477 589 543
rect 791 478 825 543
rect 1027 478 1061 543
rect 1263 477 1297 543
rect 1499 477 1533 543
rect 1735 479 1769 543
rect 1961 494 2064 543
rect -37 133 9 145
rect 201 138 235 196
rect 437 138 471 200
rect 673 138 707 200
rect 909 138 943 198
rect 1145 138 1179 202
rect 1381 138 1415 199
rect 1617 138 1651 203
rect 1853 138 1887 202
rect 1961 183 1967 494
rect 2001 183 2064 494
rect 2098 183 2104 645
rect 1961 171 2104 183
rect 2157 176 2167 634
rect 2223 176 2233 634
rect 2296 625 2330 698
rect 2393 176 2403 634
rect 2459 176 2469 634
rect 2532 630 2566 698
rect 2629 176 2639 634
rect 2695 176 2705 634
rect 2768 630 2802 698
rect 2865 176 2875 634
rect 2931 176 2941 634
rect 3004 630 3038 698
rect 3101 176 3111 634
rect 3167 176 3177 634
rect 3240 630 3274 698
rect 3337 176 3347 634
rect 3403 176 3413 634
rect 3476 630 3510 698
rect 3573 176 3583 634
rect 3639 176 3649 634
rect 3712 630 3746 698
rect 3809 176 3819 634
rect 3875 176 3885 634
rect 3948 630 3982 698
rect 4045 176 4055 634
rect 4111 176 4121 634
rect 4184 621 4218 698
rect 4281 176 4291 634
rect 4347 176 4357 634
rect 4420 621 4454 698
rect 4517 176 4527 634
rect 4583 176 4593 634
rect 4656 621 4690 698
rect 4753 176 4763 634
rect 4819 176 4829 634
rect 4892 621 4926 698
rect 4989 176 4999 634
rect 5055 176 5065 634
rect 5128 621 5162 698
rect 5225 176 5235 634
rect 5291 176 5301 634
rect 5364 621 5398 698
rect 5461 176 5471 634
rect 5527 176 5537 634
rect 5600 621 5634 698
rect 5697 176 5707 634
rect 5763 176 5773 634
rect 5836 621 5870 698
rect 5933 176 5943 634
rect 5999 176 6009 634
rect 6072 621 6106 698
rect 6169 176 6179 634
rect 6235 176 6245 634
rect 6308 621 6342 698
rect 6405 176 6415 634
rect 6471 176 6481 634
rect 6544 621 6578 698
rect 6641 176 6651 634
rect 6707 176 6717 634
rect 6780 627 6814 698
rect 6877 176 6887 634
rect 6943 176 6953 634
rect 7016 627 7050 698
rect 7113 176 7123 634
rect 7179 176 7189 634
rect 7252 626 7286 698
rect 7349 176 7359 634
rect 7415 176 7425 634
rect 7488 626 7522 698
rect 7585 176 7595 634
rect 7651 176 7661 634
rect 7724 626 7758 698
rect 7821 176 7831 634
rect 7887 176 7897 634
rect 7960 626 7994 698
rect 8191 657 8288 698
rect 8186 645 8288 657
rect 8057 176 8067 634
rect 8123 176 8133 634
rect 8186 178 8192 645
rect 8226 179 8288 645
rect 8322 179 8328 795
rect 8226 178 8328 179
rect 8186 167 8328 178
rect 8381 176 8391 784
rect 8447 176 8457 784
rect 8499 176 8509 784
rect 8565 176 8575 784
rect 8617 176 8627 784
rect 8683 176 8693 784
rect 8735 176 8745 784
rect 8801 176 8811 784
rect 8853 176 8863 784
rect 8919 176 8929 784
rect 8971 176 8981 784
rect 9037 176 9047 784
rect 9089 176 9099 784
rect 9155 176 9165 784
rect 9207 176 9217 784
rect 9273 176 9283 784
rect 9325 176 9335 784
rect 9391 176 9401 784
rect 9443 176 9453 784
rect 9509 176 9519 784
rect 9561 176 9571 784
rect 9627 176 9637 784
rect 9679 176 9689 784
rect 9745 176 9755 784
rect 9797 176 9807 784
rect 9863 176 9873 784
rect 9915 176 9925 784
rect 9981 176 9991 784
rect 10033 176 10043 784
rect 10099 176 10109 784
rect 10151 176 10161 784
rect 10217 176 10227 784
rect 10269 176 10279 784
rect 10335 176 10345 784
rect 10387 176 10397 784
rect 10453 176 10463 784
rect 10505 176 10515 784
rect 10571 176 10581 784
rect 10623 176 10633 784
rect 10689 176 10699 784
rect 10741 176 10751 784
rect 10807 176 10817 784
rect 10859 176 10869 784
rect 10925 176 10935 784
rect 10977 176 10987 784
rect 11043 176 11053 784
rect 11095 176 11105 784
rect 11161 176 11171 784
rect 11213 176 11223 784
rect 11279 176 11289 784
rect 11331 176 11341 784
rect 11397 176 11407 784
rect 11449 176 11459 784
rect 11515 176 11525 784
rect 11567 176 11577 784
rect 11633 176 11643 784
rect 11685 176 11695 784
rect 11751 176 11761 784
rect 11803 176 11813 784
rect 11869 176 11879 784
rect 11921 176 11931 784
rect 11987 176 11997 784
rect 12039 176 12049 784
rect 12105 176 12115 784
rect 12157 176 12167 784
rect 12223 176 12233 784
rect 12275 176 12285 784
rect 12341 176 12351 784
rect 12393 176 12403 784
rect 12459 176 12469 784
rect 12511 176 12521 784
rect 12577 176 12587 784
rect 12629 176 12639 784
rect 12695 176 12705 784
rect 12747 176 12757 784
rect 12813 176 12823 784
rect 12865 176 12875 784
rect 12931 176 12941 784
rect 12983 176 12993 784
rect 13049 176 13059 784
rect 13101 176 13111 784
rect 13167 176 13177 784
rect 13219 176 13229 784
rect 13285 176 13295 784
rect 13337 176 13347 784
rect 13403 176 13413 784
rect 13455 176 13465 784
rect 13521 176 13531 784
rect 13573 176 13583 784
rect 13639 176 13649 784
rect 13691 176 13701 784
rect 13757 176 13767 784
rect 13809 176 13819 784
rect 13875 176 13885 784
rect 13927 176 13937 784
rect 13993 176 14003 784
rect 14045 176 14055 784
rect 14111 176 14121 784
rect 14163 176 14173 784
rect 14229 176 14239 784
rect 14281 176 14291 784
rect 14347 176 14357 784
rect 14416 590 14704 846
rect 20792 795 20945 846
rect 14416 377 14706 590
rect 14406 318 14416 377
rect 14704 318 14714 377
rect 14763 176 14773 784
rect 14829 176 14839 784
rect 14881 176 14891 784
rect 14947 176 14957 784
rect 14999 176 15009 784
rect 15065 176 15075 784
rect 15117 176 15127 784
rect 15183 176 15193 784
rect 15235 176 15245 784
rect 15301 176 15311 784
rect 15353 176 15363 784
rect 15419 176 15429 784
rect 15471 176 15481 784
rect 15537 176 15547 784
rect 15589 176 15599 784
rect 15655 176 15665 784
rect 15707 176 15717 784
rect 15773 176 15783 784
rect 15825 176 15835 784
rect 15891 176 15901 784
rect 15943 176 15953 784
rect 16009 176 16019 784
rect 16061 176 16071 784
rect 16127 176 16137 784
rect 16179 176 16189 784
rect 16245 176 16255 784
rect 16297 176 16307 784
rect 16363 176 16373 784
rect 16415 176 16425 784
rect 16481 176 16491 784
rect 16533 176 16543 784
rect 16599 176 16609 784
rect 16651 176 16661 784
rect 16717 176 16727 784
rect 16769 176 16779 784
rect 16835 176 16845 784
rect 16887 176 16897 784
rect 16953 176 16963 784
rect 17005 176 17015 784
rect 17071 176 17081 784
rect 17123 176 17133 784
rect 17189 176 17199 784
rect 17241 176 17251 784
rect 17307 176 17317 784
rect 17359 176 17369 784
rect 17425 176 17435 784
rect 17477 176 17487 784
rect 17543 176 17553 784
rect 17595 176 17605 784
rect 17661 176 17671 784
rect 17713 176 17723 784
rect 17779 176 17789 784
rect 17831 176 17841 784
rect 17897 176 17907 784
rect 17949 176 17959 784
rect 18015 176 18025 784
rect 18067 176 18077 784
rect 18133 176 18143 784
rect 18185 176 18195 784
rect 18251 176 18261 784
rect 18303 176 18313 784
rect 18369 176 18379 784
rect 18421 176 18431 784
rect 18487 176 18497 784
rect 18539 176 18549 784
rect 18605 176 18615 784
rect 18657 176 18667 784
rect 18723 176 18733 784
rect 18775 176 18785 784
rect 18841 176 18851 784
rect 18893 176 18903 784
rect 18959 176 18969 784
rect 19011 176 19021 784
rect 19077 176 19087 784
rect 19129 176 19139 784
rect 19195 176 19205 784
rect 19247 176 19257 784
rect 19313 176 19323 784
rect 19365 176 19375 784
rect 19431 176 19441 784
rect 19483 176 19493 784
rect 19549 176 19559 784
rect 19601 176 19611 784
rect 19667 176 19677 784
rect 19719 176 19729 784
rect 19785 176 19795 784
rect 19837 176 19847 784
rect 19903 176 19913 784
rect 19955 176 19965 784
rect 20021 176 20031 784
rect 20073 176 20083 784
rect 20139 176 20149 784
rect 20191 176 20201 784
rect 20257 176 20267 784
rect 20309 176 20319 784
rect 20375 176 20385 784
rect 20427 176 20437 784
rect 20493 176 20503 784
rect 20545 176 20555 784
rect 20611 176 20621 784
rect 20663 176 20673 784
rect 20729 176 20736 784
rect 8186 166 8232 167
rect 8360 138 20675 139
rect 63 92 20675 138
rect 63 -425 471 92
rect 796 -97 2167 -5
rect 8123 -97 8133 -5
rect 796 -344 8133 -97
rect 796 -378 951 -344
rect 7721 -378 8133 -344
rect 796 -420 8133 -378
rect 796 -441 1003 -420
rect 796 -1860 855 -441
rect 889 -1537 1003 -441
rect 889 -1856 992 -1537
rect 889 -1860 1003 -1856
rect 1216 -1860 1226 -452
rect 1282 -1860 1292 -452
rect 1505 -458 1539 -420
rect 1752 -1860 1762 -452
rect 1818 -1860 1828 -452
rect 2041 -458 2075 -420
rect 2288 -1860 2298 -452
rect 2354 -1860 2364 -452
rect 2577 -458 2611 -420
rect 2824 -1860 2834 -452
rect 2890 -1860 2900 -452
rect 3113 -458 3147 -420
rect 3360 -1860 3370 -452
rect 3426 -1860 3436 -452
rect 3649 -459 3683 -420
rect 3896 -1860 3906 -452
rect 3962 -1860 3972 -452
rect 4185 -457 4219 -420
rect 4432 -1860 4442 -452
rect 4498 -1860 4508 -452
rect 4721 -458 4755 -420
rect 796 -1872 1003 -1860
rect 4968 -1861 4978 -453
rect 5034 -1861 5044 -453
rect 5257 -459 5291 -420
rect 5504 -1860 5514 -452
rect 5570 -1860 5580 -452
rect 5793 -458 5827 -420
rect 6040 -1860 6050 -452
rect 6106 -1860 6116 -452
rect 6329 -457 6363 -420
rect 6576 -1860 6586 -452
rect 6642 -1860 6652 -452
rect 6865 -458 6899 -420
rect 7112 -1860 7122 -452
rect 7178 -1860 7188 -452
rect 7401 -459 7435 -420
rect 7755 -441 8133 -420
rect 7649 -1861 7659 -453
rect 7715 -1861 7725 -453
rect 64 -2249 7657 -1903
rect 7755 -1943 7783 -441
rect 7817 -1943 8133 -441
rect 8282 -155 8328 -143
rect 8282 -857 8288 -155
rect 8322 -857 8328 -155
rect 8360 -201 20675 92
rect 20792 93 20798 795
rect 20832 93 20945 795
rect 20792 -155 20945 93
rect 8381 -846 8391 -238
rect 8447 -846 8457 -238
rect 8499 -846 8509 -238
rect 8565 -846 8575 -238
rect 8617 -846 8627 -238
rect 8683 -846 8693 -238
rect 8735 -846 8745 -238
rect 8801 -846 8811 -238
rect 8853 -846 8863 -238
rect 8919 -846 8929 -238
rect 8971 -846 8981 -238
rect 9037 -846 9047 -238
rect 9089 -846 9099 -238
rect 9155 -846 9165 -238
rect 9207 -846 9217 -238
rect 9273 -846 9283 -238
rect 9325 -846 9335 -238
rect 9391 -846 9401 -238
rect 9443 -846 9453 -238
rect 9509 -846 9519 -238
rect 9561 -846 9571 -238
rect 9627 -846 9637 -238
rect 9679 -846 9689 -238
rect 9745 -846 9755 -238
rect 9797 -846 9807 -238
rect 9863 -846 9873 -238
rect 9915 -846 9925 -238
rect 9981 -846 9991 -238
rect 10033 -846 10043 -238
rect 10099 -846 10109 -238
rect 10151 -846 10161 -238
rect 10217 -846 10227 -238
rect 10269 -846 10279 -238
rect 10335 -846 10345 -238
rect 10387 -846 10397 -238
rect 10453 -846 10463 -238
rect 10505 -846 10515 -238
rect 10571 -846 10581 -238
rect 10623 -846 10633 -238
rect 10689 -846 10699 -238
rect 10741 -846 10751 -238
rect 10807 -846 10817 -238
rect 10859 -846 10869 -238
rect 10925 -846 10935 -238
rect 10977 -846 10987 -238
rect 11043 -846 11053 -238
rect 11095 -846 11105 -238
rect 11161 -846 11171 -238
rect 11213 -846 11223 -238
rect 11279 -846 11289 -238
rect 11331 -846 11341 -238
rect 11397 -846 11407 -238
rect 11449 -846 11459 -238
rect 11515 -846 11525 -238
rect 11567 -846 11577 -238
rect 11633 -846 11643 -238
rect 11685 -846 11695 -238
rect 11751 -846 11761 -238
rect 11803 -846 11813 -238
rect 11869 -846 11879 -238
rect 11921 -846 11931 -238
rect 11987 -846 11997 -238
rect 12039 -846 12049 -238
rect 12105 -846 12115 -238
rect 12157 -846 12167 -238
rect 12223 -846 12233 -238
rect 12275 -846 12285 -238
rect 12341 -846 12351 -238
rect 12393 -846 12403 -238
rect 12459 -846 12469 -238
rect 12511 -846 12521 -238
rect 12577 -846 12587 -238
rect 12629 -846 12639 -238
rect 12695 -846 12705 -238
rect 12747 -846 12757 -238
rect 12813 -846 12823 -238
rect 12865 -846 12875 -238
rect 12931 -846 12941 -238
rect 12983 -846 12993 -238
rect 13049 -846 13059 -238
rect 13101 -846 13111 -238
rect 13167 -846 13177 -238
rect 13219 -846 13229 -238
rect 13285 -846 13295 -238
rect 13337 -846 13347 -238
rect 13403 -846 13413 -238
rect 13455 -846 13465 -238
rect 13521 -846 13531 -238
rect 13573 -846 13583 -238
rect 13639 -846 13649 -238
rect 13691 -846 13701 -238
rect 13757 -846 13767 -238
rect 13809 -846 13819 -238
rect 13875 -846 13885 -238
rect 13927 -846 13937 -238
rect 13993 -846 14003 -238
rect 14045 -846 14055 -238
rect 14111 -846 14121 -238
rect 14163 -846 14173 -238
rect 14229 -846 14239 -238
rect 14281 -846 14291 -238
rect 14347 -846 14357 -238
rect 14414 -381 14704 -376
rect 14406 -435 14416 -381
rect 14704 -435 14714 -381
rect 14414 -648 14704 -435
rect 8282 -914 8328 -857
rect 14416 -914 14704 -648
rect 14763 -846 14773 -238
rect 14829 -846 14839 -238
rect 14881 -846 14891 -238
rect 14947 -846 14957 -238
rect 14999 -846 15009 -238
rect 15065 -846 15075 -238
rect 15117 -846 15127 -238
rect 15183 -846 15193 -238
rect 15235 -846 15245 -238
rect 15301 -846 15311 -238
rect 15353 -846 15363 -238
rect 15419 -846 15429 -238
rect 15471 -846 15481 -238
rect 15537 -846 15547 -238
rect 15589 -846 15599 -238
rect 15655 -846 15665 -238
rect 15707 -846 15717 -238
rect 15773 -846 15783 -238
rect 15825 -846 15835 -238
rect 15891 -846 15901 -238
rect 15943 -846 15953 -238
rect 16009 -846 16019 -238
rect 16061 -846 16071 -238
rect 16127 -846 16137 -238
rect 16179 -846 16189 -238
rect 16245 -846 16255 -238
rect 16297 -846 16307 -238
rect 16363 -846 16373 -238
rect 16415 -846 16425 -238
rect 16481 -846 16491 -238
rect 16533 -846 16543 -238
rect 16599 -846 16609 -238
rect 16651 -846 16661 -238
rect 16717 -846 16727 -238
rect 16769 -846 16779 -238
rect 16835 -846 16845 -238
rect 16887 -846 16897 -238
rect 16953 -846 16963 -238
rect 17005 -846 17015 -238
rect 17071 -846 17081 -238
rect 17123 -846 17133 -238
rect 17189 -846 17199 -238
rect 17241 -846 17251 -238
rect 17307 -846 17317 -238
rect 17359 -846 17369 -238
rect 17425 -846 17435 -238
rect 17477 -846 17487 -238
rect 17543 -846 17553 -238
rect 17595 -846 17605 -238
rect 17661 -846 17671 -238
rect 17713 -846 17723 -238
rect 17779 -846 17789 -238
rect 17831 -846 17841 -238
rect 17897 -846 17907 -238
rect 17949 -846 17959 -238
rect 18015 -846 18025 -238
rect 18067 -846 18077 -238
rect 18133 -846 18143 -238
rect 18185 -846 18195 -238
rect 18251 -846 18261 -238
rect 18303 -846 18313 -238
rect 18369 -846 18379 -238
rect 18421 -846 18431 -238
rect 18487 -846 18497 -238
rect 18539 -846 18549 -238
rect 18605 -846 18615 -238
rect 18657 -846 18667 -238
rect 18723 -846 18733 -238
rect 18775 -846 18785 -238
rect 18841 -846 18851 -238
rect 18893 -846 18903 -238
rect 18959 -846 18969 -238
rect 19011 -846 19021 -238
rect 19077 -846 19087 -238
rect 19129 -846 19139 -238
rect 19195 -846 19205 -238
rect 19247 -846 19257 -238
rect 19313 -846 19323 -238
rect 19365 -846 19375 -238
rect 19431 -846 19441 -238
rect 19483 -846 19493 -238
rect 19549 -846 19559 -238
rect 19601 -846 19611 -238
rect 19667 -846 19677 -238
rect 19719 -846 19729 -238
rect 19785 -846 19795 -238
rect 19837 -846 19847 -238
rect 19903 -846 19913 -238
rect 19955 -846 19965 -238
rect 20021 -846 20031 -238
rect 20073 -846 20083 -238
rect 20139 -846 20149 -238
rect 20191 -846 20201 -238
rect 20257 -846 20267 -238
rect 20309 -846 20319 -238
rect 20375 -846 20385 -238
rect 20427 -846 20437 -238
rect 20493 -846 20503 -238
rect 20545 -846 20555 -238
rect 20611 -846 20621 -238
rect 20663 -846 20673 -238
rect 20729 -846 20736 -238
rect 20792 -857 20798 -155
rect 20832 -790 20945 -155
rect 22549 -790 22578 1002
rect 20832 -853 22578 -790
rect 20832 -857 20838 -853
rect 20792 -914 20838 -857
rect 8282 -920 20838 -914
rect 8282 -954 8384 -920
rect 14354 -954 14766 -920
rect 20736 -954 20838 -920
rect 8282 -960 20838 -954
rect 7755 -2209 8133 -1943
rect 849 -2292 895 -2280
rect 796 -3711 855 -2292
rect 889 -3711 1003 -2292
rect 1216 -3700 1226 -2292
rect 1282 -3700 1292 -2292
rect 796 -3729 1003 -3711
rect 1505 -3729 1539 -3691
rect 1752 -3700 1762 -2292
rect 1818 -3700 1828 -2292
rect 2041 -3729 2075 -3694
rect 2288 -3700 2298 -2292
rect 2354 -3700 2364 -2292
rect 2577 -3729 2611 -3694
rect 2824 -3700 2834 -2292
rect 2890 -3700 2900 -2292
rect 3113 -3729 3147 -3693
rect 3360 -3701 3370 -2283
rect 3426 -3701 3436 -2283
rect 3649 -3729 3683 -3695
rect 3896 -3701 3906 -2283
rect 3962 -3701 3972 -2283
rect 4185 -3729 4219 -3693
rect 4432 -3701 4442 -2283
rect 4498 -3701 4508 -2283
rect 4721 -3729 4755 -3692
rect 4968 -3701 4978 -2283
rect 5034 -3701 5044 -2283
rect 5257 -3729 5291 -3693
rect 5504 -3701 5514 -2283
rect 5570 -3701 5580 -2283
rect 5793 -3729 5827 -3693
rect 6040 -3701 6050 -2283
rect 6106 -3701 6116 -2283
rect 6329 -3729 6363 -3693
rect 6576 -3701 6586 -2283
rect 6642 -3701 6652 -2283
rect 6865 -3729 6899 -3692
rect 7113 -3701 7123 -2283
rect 7179 -3701 7189 -2283
rect 7401 -3729 7435 -3693
rect 7649 -3701 7659 -2284
rect 7715 -3701 7725 -2284
rect 7755 -3711 7783 -2209
rect 7817 -3711 8133 -2209
rect 7755 -3719 8133 -3711
rect 7754 -3729 8133 -3719
rect 796 -3952 8133 -3729
rect 796 -3970 1003 -3952
rect 796 -5389 855 -3970
rect 889 -5389 1003 -3970
rect 1216 -5389 1226 -3981
rect 1282 -5389 1292 -3981
rect 1505 -3988 1539 -3952
rect 1752 -5389 1762 -3981
rect 1818 -5389 1828 -3981
rect 2041 -3988 2075 -3952
rect 2288 -5389 2298 -3981
rect 2354 -5389 2364 -3981
rect 2577 -3988 2611 -3952
rect 2824 -5389 2834 -3981
rect 2890 -5389 2900 -3981
rect 3113 -3987 3147 -3952
rect 3360 -5389 3370 -3981
rect 3426 -5389 3436 -3981
rect 3649 -3988 3683 -3952
rect 3896 -5389 3906 -3981
rect 3962 -5389 3972 -3981
rect 4185 -3988 4219 -3952
rect 4432 -5389 4442 -3981
rect 4498 -5389 4508 -3981
rect 4721 -3987 4755 -3952
rect 849 -5401 895 -5389
rect 4968 -5390 4978 -3982
rect 5034 -5390 5044 -3982
rect 5257 -3987 5291 -3952
rect 5504 -5389 5514 -3981
rect 5570 -5389 5580 -3981
rect 5793 -3987 5827 -3952
rect 6040 -5389 6050 -3981
rect 6106 -5389 6116 -3981
rect 6329 -3987 6363 -3952
rect 6576 -5389 6586 -3981
rect 6642 -5389 6652 -3981
rect 6865 -3987 6899 -3952
rect 7112 -5389 7122 -3981
rect 7178 -5389 7188 -3981
rect 7401 -3987 7435 -3952
rect 7754 -3970 8133 -3952
rect 7649 -5390 7659 -3982
rect 7715 -5390 7725 -3982
rect 514 -5778 7725 -5432
rect 7754 -5472 7783 -3970
rect 7817 -5472 8133 -3970
rect 7754 -5738 8133 -5472
rect 796 -5821 1003 -5809
rect 796 -7240 855 -5821
rect 889 -7240 1003 -5821
rect 1216 -7229 1226 -5821
rect 1282 -7229 1292 -5821
rect 796 -7258 1003 -7240
rect 1505 -7258 1539 -7216
rect 1752 -7229 1762 -5821
rect 1818 -7229 1828 -5821
rect 2041 -7258 2075 -7217
rect 2288 -7229 2298 -5821
rect 2354 -7229 2364 -5821
rect 2577 -7258 2611 -7217
rect 2824 -7229 2834 -5821
rect 2890 -7229 2900 -5821
rect 3113 -7258 3147 -7218
rect 3360 -7230 3370 -5812
rect 3426 -7230 3436 -5812
rect 3649 -7258 3683 -7219
rect 3896 -7230 3906 -5812
rect 3962 -7230 3972 -5812
rect 4185 -7258 4219 -7219
rect 4432 -7230 4442 -5812
rect 4498 -7230 4508 -5812
rect 4721 -7258 4755 -7219
rect 4968 -7230 4978 -5812
rect 5034 -7230 5044 -5812
rect 5257 -7258 5291 -7222
rect 5504 -7230 5514 -5812
rect 5570 -7230 5580 -5812
rect 5793 -7258 5827 -7220
rect 6040 -7230 6050 -5812
rect 6106 -7230 6116 -5812
rect 6329 -7258 6363 -7220
rect 6576 -7230 6586 -5812
rect 6642 -7230 6652 -5812
rect 6865 -7258 6899 -7221
rect 7113 -7230 7123 -5812
rect 7179 -7230 7189 -5812
rect 7401 -7258 7435 -7222
rect 7649 -7230 7659 -5813
rect 7715 -7230 7725 -5813
rect 7754 -7240 7783 -5738
rect 7817 -7240 8133 -5738
rect 7754 -7258 8133 -7240
rect 795 -7303 8133 -7258
rect 795 -7337 951 -7303
rect 7721 -7337 8133 -7303
rect 795 -7431 8133 -7337
rect 8162 -2146 8172 -2006
rect 8292 -2146 8302 -2006
rect 8162 -7641 8302 -2146
rect 824 -7699 870 -7690
rect 820 -7702 870 -7699
rect 820 -9896 830 -7702
rect 864 -9896 870 -7702
rect 944 -7748 10884 -7641
rect 11004 -7702 11050 -7690
rect 944 -7788 978 -7748
rect 1361 -9884 1371 -7776
rect 1427 -9884 1437 -7776
rect 1820 -7783 1854 -7748
rect 2237 -9884 2247 -7776
rect 2303 -9884 2313 -7776
rect 2696 -7783 2730 -7748
rect 3113 -9884 3123 -7776
rect 3179 -9884 3189 -7776
rect 3572 -7782 3606 -7748
rect 3989 -9884 3999 -7776
rect 4055 -9884 4065 -7776
rect 4448 -7782 4482 -7748
rect 4865 -9884 4875 -7776
rect 4931 -9884 4941 -7776
rect 5324 -7782 5358 -7748
rect 5741 -9884 5751 -7776
rect 5807 -9884 5817 -7776
rect 5870 -7800 6004 -7788
rect 820 -9930 870 -9896
rect 5870 -9896 5876 -7800
rect 5910 -9896 5964 -7800
rect 5998 -9896 6004 -7800
rect 6057 -9884 6067 -7776
rect 6123 -9884 6133 -7776
rect 6495 -9884 6505 -7776
rect 6561 -9884 6571 -7776
rect 6933 -9884 6943 -7776
rect 6999 -9884 7009 -7776
rect 7371 -9884 7381 -7776
rect 7437 -9884 7447 -7776
rect 7809 -9884 7819 -7776
rect 7875 -9884 7885 -7776
rect 8247 -9884 8257 -7776
rect 8313 -9884 8323 -7776
rect 8685 -9884 8695 -7776
rect 8751 -9884 8761 -7776
rect 9123 -9884 9133 -7776
rect 9189 -9884 9199 -7776
rect 9561 -9884 9571 -7776
rect 9627 -9884 9637 -7776
rect 9999 -9884 10009 -7776
rect 10065 -9884 10075 -7776
rect 10437 -9884 10447 -7776
rect 10503 -9884 10513 -7776
rect 10875 -9884 10885 -7776
rect 10941 -9884 10948 -7776
rect 5870 -9930 6004 -9896
rect 11004 -9896 11010 -7702
rect 11044 -8333 11050 -7702
rect 11716 -7722 12074 -960
rect 12726 -7204 22688 -7189
rect 11209 -8084 11219 -7776
rect 11279 -8084 11289 -7776
rect 11320 -8141 11366 -8050
rect 11397 -8084 11407 -7776
rect 11471 -8084 11481 -7776
rect 11518 -8141 11552 -8076
rect 11589 -8084 11599 -7776
rect 11663 -8084 11673 -7776
rect 11710 -8141 11744 -8077
rect 11781 -8084 11791 -7776
rect 11855 -8084 11865 -7776
rect 11902 -8141 11936 -8071
rect 11973 -8084 11983 -7776
rect 12047 -8084 12057 -7776
rect 12094 -8141 12128 -8074
rect 12165 -8084 12175 -7776
rect 12239 -8084 12249 -7776
rect 12286 -8141 12320 -8071
rect 12357 -8084 12367 -7776
rect 12431 -8084 12441 -7776
rect 12478 -8141 12512 -8071
rect 12549 -8084 12559 -7776
rect 12623 -8084 12633 -7776
rect 11310 -8195 11320 -8141
rect 12512 -8195 12522 -8141
rect 11044 -8354 12663 -8333
rect 11044 -9895 11119 -8354
rect 12657 -9793 12663 -8354
rect 12719 -9409 12726 -7204
rect 12923 -7248 22688 -7204
rect 22808 -7204 22905 -7192
rect 12923 -7910 12954 -7248
rect 22808 -7633 22835 -7204
rect 22778 -7660 22835 -7633
rect 22869 -7660 22905 -7204
rect 22778 -7762 22905 -7660
rect 12923 -7969 22688 -7910
rect 22808 -7924 22905 -7762
rect 12923 -8630 12954 -7969
rect 22808 -8353 22835 -7924
rect 22785 -8380 22835 -8353
rect 22869 -8380 22905 -7924
rect 22785 -8482 22905 -8380
rect 12923 -8689 22688 -8630
rect 22808 -8644 22905 -8482
rect 12923 -9350 12954 -8689
rect 22808 -9073 22835 -8644
rect 22785 -9100 22835 -9073
rect 22869 -9100 22905 -8644
rect 22785 -9202 22905 -9100
rect 12923 -9409 22688 -9350
rect 22808 -9364 22905 -9202
rect 22808 -9793 22835 -9364
rect 12657 -9820 22835 -9793
rect 22869 -9820 22905 -9364
rect 12657 -9895 22905 -9820
rect 11044 -9896 22905 -9895
rect 11004 -9930 22905 -9896
rect 820 -9975 22905 -9930
rect 820 -10066 12690 -9975
rect 820 -10122 836 -10066
rect 10951 -10122 12690 -10066
rect 22854 -10122 22905 -9975
rect 820 -10133 22905 -10122
<< via1 >>
rect 8316 970 20769 1085
rect 2167 176 2223 634
rect 2403 176 2459 634
rect 2639 176 2695 634
rect 2875 176 2931 634
rect 3111 176 3167 634
rect 3347 176 3403 634
rect 3583 176 3639 634
rect 3819 176 3875 634
rect 4055 176 4111 634
rect 4291 176 4347 634
rect 4527 176 4583 634
rect 4763 176 4819 634
rect 4999 176 5055 634
rect 5235 176 5291 634
rect 5471 176 5527 634
rect 5707 176 5763 634
rect 5943 176 5999 634
rect 6179 176 6235 634
rect 6415 176 6471 634
rect 6651 176 6707 634
rect 6887 176 6943 634
rect 7123 176 7179 634
rect 7359 176 7415 634
rect 7595 176 7651 634
rect 7831 176 7887 634
rect 8067 176 8123 634
rect 8391 176 8447 784
rect 8509 176 8565 784
rect 8627 176 8683 784
rect 8745 176 8801 784
rect 8863 176 8919 784
rect 8981 176 9037 784
rect 9099 176 9155 784
rect 9217 176 9273 784
rect 9335 176 9391 784
rect 9453 176 9509 784
rect 9571 176 9627 784
rect 9689 176 9745 784
rect 9807 176 9863 784
rect 9925 176 9981 784
rect 10043 176 10099 784
rect 10161 176 10217 784
rect 10279 176 10335 784
rect 10397 176 10453 784
rect 10515 176 10571 784
rect 10633 176 10689 784
rect 10751 176 10807 784
rect 10869 176 10925 784
rect 10987 176 11043 784
rect 11105 176 11161 784
rect 11223 176 11279 784
rect 11341 176 11397 784
rect 11459 176 11515 784
rect 11577 176 11633 784
rect 11695 176 11751 784
rect 11813 176 11869 784
rect 11931 176 11987 784
rect 12049 176 12105 784
rect 12167 176 12223 784
rect 12285 176 12341 784
rect 12403 176 12459 784
rect 12521 176 12577 784
rect 12639 176 12695 784
rect 12757 176 12813 784
rect 12875 176 12931 784
rect 12993 176 13049 784
rect 13111 176 13167 784
rect 13229 176 13285 784
rect 13347 176 13403 784
rect 13465 176 13521 784
rect 13583 176 13639 784
rect 13701 176 13757 784
rect 13819 176 13875 784
rect 13937 176 13993 784
rect 14055 176 14111 784
rect 14173 176 14229 784
rect 14291 176 14347 784
rect 14416 318 14704 377
rect 14773 176 14829 784
rect 14891 176 14947 784
rect 15009 176 15065 784
rect 15127 176 15183 784
rect 15245 176 15301 784
rect 15363 176 15419 784
rect 15481 176 15537 784
rect 15599 176 15655 784
rect 15717 176 15773 784
rect 15835 176 15891 784
rect 15953 176 16009 784
rect 16071 176 16127 784
rect 16189 176 16245 784
rect 16307 176 16363 784
rect 16425 176 16481 784
rect 16543 176 16599 784
rect 16661 176 16717 784
rect 16779 176 16835 784
rect 16897 176 16953 784
rect 17015 176 17071 784
rect 17133 176 17189 784
rect 17251 176 17307 784
rect 17369 176 17425 784
rect 17487 176 17543 784
rect 17605 176 17661 784
rect 17723 176 17779 784
rect 17841 176 17897 784
rect 17959 176 18015 784
rect 18077 176 18133 784
rect 18195 176 18251 784
rect 18313 176 18369 784
rect 18431 176 18487 784
rect 18549 176 18605 784
rect 18667 176 18723 784
rect 18785 176 18841 784
rect 18903 176 18959 784
rect 19021 176 19077 784
rect 19139 176 19195 784
rect 19257 176 19313 784
rect 19375 176 19431 784
rect 19493 176 19549 784
rect 19611 176 19667 784
rect 19729 176 19785 784
rect 19847 176 19903 784
rect 19965 176 20021 784
rect 20083 176 20139 784
rect 20201 176 20257 784
rect 20319 176 20375 784
rect 20437 176 20493 784
rect 20555 176 20611 784
rect 20673 176 20729 784
rect 2167 -97 8123 -5
rect 1226 -1860 1282 -452
rect 1762 -1860 1818 -452
rect 2298 -1860 2354 -452
rect 2834 -1860 2890 -452
rect 3370 -1860 3426 -452
rect 3906 -1860 3962 -452
rect 4442 -1860 4498 -452
rect 4978 -1861 5034 -453
rect 5514 -1860 5570 -452
rect 6050 -1860 6106 -452
rect 6586 -1860 6642 -452
rect 7122 -1860 7178 -452
rect 7659 -1861 7715 -453
rect 8391 -846 8447 -238
rect 8509 -846 8565 -238
rect 8627 -846 8683 -238
rect 8745 -846 8801 -238
rect 8863 -846 8919 -238
rect 8981 -846 9037 -238
rect 9099 -846 9155 -238
rect 9217 -846 9273 -238
rect 9335 -846 9391 -238
rect 9453 -846 9509 -238
rect 9571 -846 9627 -238
rect 9689 -846 9745 -238
rect 9807 -846 9863 -238
rect 9925 -846 9981 -238
rect 10043 -846 10099 -238
rect 10161 -846 10217 -238
rect 10279 -846 10335 -238
rect 10397 -846 10453 -238
rect 10515 -846 10571 -238
rect 10633 -846 10689 -238
rect 10751 -846 10807 -238
rect 10869 -846 10925 -238
rect 10987 -846 11043 -238
rect 11105 -846 11161 -238
rect 11223 -846 11279 -238
rect 11341 -846 11397 -238
rect 11459 -846 11515 -238
rect 11577 -846 11633 -238
rect 11695 -846 11751 -238
rect 11813 -846 11869 -238
rect 11931 -846 11987 -238
rect 12049 -846 12105 -238
rect 12167 -846 12223 -238
rect 12285 -846 12341 -238
rect 12403 -846 12459 -238
rect 12521 -846 12577 -238
rect 12639 -846 12695 -238
rect 12757 -846 12813 -238
rect 12875 -846 12931 -238
rect 12993 -846 13049 -238
rect 13111 -846 13167 -238
rect 13229 -846 13285 -238
rect 13347 -846 13403 -238
rect 13465 -846 13521 -238
rect 13583 -846 13639 -238
rect 13701 -846 13757 -238
rect 13819 -846 13875 -238
rect 13937 -846 13993 -238
rect 14055 -846 14111 -238
rect 14173 -846 14229 -238
rect 14291 -846 14347 -238
rect 14416 -435 14704 -381
rect 14773 -846 14829 -238
rect 14891 -846 14947 -238
rect 15009 -846 15065 -238
rect 15127 -846 15183 -238
rect 15245 -846 15301 -238
rect 15363 -846 15419 -238
rect 15481 -846 15537 -238
rect 15599 -846 15655 -238
rect 15717 -846 15773 -238
rect 15835 -846 15891 -238
rect 15953 -846 16009 -238
rect 16071 -846 16127 -238
rect 16189 -846 16245 -238
rect 16307 -846 16363 -238
rect 16425 -846 16481 -238
rect 16543 -846 16599 -238
rect 16661 -846 16717 -238
rect 16779 -846 16835 -238
rect 16897 -846 16953 -238
rect 17015 -846 17071 -238
rect 17133 -846 17189 -238
rect 17251 -846 17307 -238
rect 17369 -846 17425 -238
rect 17487 -846 17543 -238
rect 17605 -846 17661 -238
rect 17723 -846 17779 -238
rect 17841 -846 17897 -238
rect 17959 -846 18015 -238
rect 18077 -846 18133 -238
rect 18195 -846 18251 -238
rect 18313 -846 18369 -238
rect 18431 -846 18487 -238
rect 18549 -846 18605 -238
rect 18667 -846 18723 -238
rect 18785 -846 18841 -238
rect 18903 -846 18959 -238
rect 19021 -846 19077 -238
rect 19139 -846 19195 -238
rect 19257 -846 19313 -238
rect 19375 -846 19431 -238
rect 19493 -846 19549 -238
rect 19611 -846 19667 -238
rect 19729 -846 19785 -238
rect 19847 -846 19903 -238
rect 19965 -846 20021 -238
rect 20083 -846 20139 -238
rect 20201 -846 20257 -238
rect 20319 -846 20375 -238
rect 20437 -846 20493 -238
rect 20555 -846 20611 -238
rect 20673 -846 20729 -238
rect 1226 -3700 1282 -2292
rect 1762 -3700 1818 -2292
rect 2298 -3700 2354 -2292
rect 2834 -3700 2890 -2292
rect 3370 -3701 3426 -2283
rect 3906 -3701 3962 -2283
rect 4442 -3701 4498 -2283
rect 4978 -3701 5034 -2283
rect 5514 -3701 5570 -2283
rect 6050 -3701 6106 -2283
rect 6586 -3701 6642 -2283
rect 7123 -3701 7179 -2283
rect 7659 -3701 7715 -2284
rect 1226 -5389 1282 -3981
rect 1762 -5389 1818 -3981
rect 2298 -5389 2354 -3981
rect 2834 -5389 2890 -3981
rect 3370 -5389 3426 -3981
rect 3906 -5389 3962 -3981
rect 4442 -5389 4498 -3981
rect 4978 -5390 5034 -3982
rect 5514 -5389 5570 -3981
rect 6050 -5389 6106 -3981
rect 6586 -5389 6642 -3981
rect 7122 -5389 7178 -3981
rect 7659 -5390 7715 -3982
rect 1226 -7229 1282 -5821
rect 1762 -7229 1818 -5821
rect 2298 -7229 2354 -5821
rect 2834 -7229 2890 -5821
rect 3370 -7230 3426 -5812
rect 3906 -7230 3962 -5812
rect 4442 -7230 4498 -5812
rect 4978 -7230 5034 -5812
rect 5514 -7230 5570 -5812
rect 6050 -7230 6106 -5812
rect 6586 -7230 6642 -5812
rect 7123 -7230 7179 -5812
rect 7659 -7230 7715 -5813
rect 8172 -2146 8292 -2006
rect 1371 -9884 1427 -7776
rect 2247 -9884 2303 -7776
rect 3123 -9884 3179 -7776
rect 3999 -9884 4055 -7776
rect 4875 -9884 4931 -7776
rect 5751 -9884 5807 -7776
rect 6067 -9884 6123 -7776
rect 6505 -9884 6561 -7776
rect 6943 -9884 6999 -7776
rect 7381 -9884 7437 -7776
rect 7819 -9884 7875 -7776
rect 8257 -9884 8313 -7776
rect 8695 -9884 8751 -7776
rect 9133 -9884 9189 -7776
rect 9571 -9884 9627 -7776
rect 10009 -9884 10065 -7776
rect 10447 -9884 10503 -7776
rect 10885 -9884 10941 -7776
rect 11219 -8084 11279 -7776
rect 11407 -8084 11471 -7776
rect 11599 -8084 11663 -7776
rect 11791 -8084 11855 -7776
rect 11983 -8084 12047 -7776
rect 12175 -8084 12239 -7776
rect 12367 -8084 12431 -7776
rect 12559 -8084 12623 -7776
rect 11320 -8195 12512 -8141
rect 12726 -9409 12923 -7204
rect 836 -10122 10951 -10066
<< metal2 >>
rect 8289 1085 20914 1179
rect 8289 970 8316 1085
rect 20769 970 20914 1085
rect 8289 908 14375 970
rect 8334 822 14375 908
rect 14745 908 20914 970
rect 14745 905 20913 908
rect 14745 822 20862 905
rect 8391 784 8447 822
rect 2167 634 2223 644
rect 2167 5 2223 176
rect 2403 634 2459 644
rect 2403 5 2459 176
rect 2639 634 2695 644
rect 2639 5 2695 176
rect 2875 634 2931 644
rect 2875 5 2931 176
rect 3111 634 3167 644
rect 3111 5 3167 176
rect 3347 634 3403 644
rect 3347 5 3403 176
rect 3583 634 3639 644
rect 3583 5 3639 176
rect 3819 634 3875 644
rect 3819 5 3875 176
rect 4055 634 4111 644
rect 4055 5 4111 176
rect 4291 634 4347 644
rect 4291 5 4347 176
rect 4527 634 4583 644
rect 4527 5 4583 176
rect 4763 634 4819 644
rect 4763 5 4819 176
rect 4999 634 5055 644
rect 4999 5 5055 176
rect 5235 634 5291 644
rect 5235 5 5291 176
rect 5471 634 5527 644
rect 5471 5 5527 176
rect 5707 634 5763 644
rect 5707 5 5763 176
rect 5943 634 5999 644
rect 5943 5 5999 176
rect 6179 634 6235 644
rect 6179 5 6235 176
rect 6415 634 6471 644
rect 6415 5 6471 176
rect 6651 634 6707 644
rect 6651 5 6707 176
rect 6887 634 6943 644
rect 6887 5 6943 176
rect 7123 634 7179 644
rect 7123 5 7179 176
rect 7359 634 7415 644
rect 7359 5 7415 176
rect 7595 634 7651 644
rect 7595 5 7651 176
rect 7831 634 7887 644
rect 7831 5 7887 176
rect 8067 634 8123 644
rect 8067 5 8123 176
rect 2167 -5 8123 5
rect 2167 -107 8123 -97
rect 8391 -238 8447 176
rect 1226 -452 1282 -442
rect 1226 -2006 1282 -1860
rect 1762 -452 1818 -442
rect 1762 -2006 1818 -1860
rect 2298 -452 2354 -442
rect 2298 -2006 2354 -1860
rect 2834 -452 2890 -442
rect 2834 -2006 2890 -1860
rect 3370 -452 3426 -442
rect 3370 -2006 3426 -1860
rect 3906 -452 3962 -442
rect 3906 -2006 3962 -1860
rect 4442 -452 4498 -442
rect 4442 -2006 4498 -1860
rect 4978 -453 5034 -443
rect 4978 -2006 5034 -1861
rect 5514 -452 5570 -442
rect 5514 -2006 5570 -1860
rect 6050 -452 6106 -442
rect 6050 -2006 6106 -1860
rect 6586 -452 6642 -442
rect 6586 -2006 6642 -1860
rect 7122 -452 7178 -442
rect 7122 -1866 7178 -1860
rect 7659 -453 7715 -443
rect 8391 -856 8447 -846
rect 8509 784 8565 794
rect 8509 -238 8565 176
rect 8509 -884 8565 -846
rect 8627 784 8683 822
rect 8627 -238 8683 176
rect 8627 -856 8683 -846
rect 8745 784 8801 794
rect 8745 -238 8801 176
rect 8745 -884 8801 -846
rect 8863 784 8919 822
rect 8863 -238 8919 176
rect 8863 -856 8919 -846
rect 8981 784 9037 794
rect 8981 -238 9037 176
rect 8981 -884 9037 -846
rect 9099 784 9155 822
rect 9099 -238 9155 176
rect 9099 -856 9155 -846
rect 9217 784 9273 794
rect 9217 -238 9273 176
rect 9217 -884 9273 -846
rect 9335 784 9391 822
rect 9335 -238 9391 176
rect 9335 -856 9391 -846
rect 9453 784 9509 794
rect 9453 -238 9509 176
rect 9453 -884 9509 -846
rect 9571 784 9627 822
rect 9571 -238 9627 176
rect 9571 -856 9627 -846
rect 9689 784 9745 794
rect 9689 -238 9745 176
rect 9689 -884 9745 -846
rect 9807 784 9863 822
rect 9807 -238 9863 176
rect 9807 -856 9863 -846
rect 9925 784 9981 794
rect 9925 -238 9981 176
rect 9925 -884 9981 -846
rect 10043 784 10099 822
rect 10043 -238 10099 176
rect 10043 -856 10099 -846
rect 10161 784 10217 794
rect 10161 -238 10217 176
rect 10161 -884 10217 -846
rect 10279 784 10335 822
rect 10279 -238 10335 176
rect 10279 -856 10335 -846
rect 10397 784 10453 794
rect 10397 -238 10453 176
rect 10397 -884 10453 -846
rect 10515 784 10571 822
rect 10515 -238 10571 176
rect 10515 -856 10571 -846
rect 10633 784 10689 794
rect 10633 -238 10689 176
rect 10633 -884 10689 -846
rect 10751 784 10807 822
rect 10751 -238 10807 176
rect 10751 -856 10807 -846
rect 10869 784 10925 794
rect 10869 -238 10925 176
rect 10869 -884 10925 -846
rect 10987 784 11043 822
rect 10987 -238 11043 176
rect 10987 -856 11043 -846
rect 11105 784 11161 794
rect 11105 -238 11161 176
rect 11105 -884 11161 -846
rect 11223 784 11279 822
rect 11223 -238 11279 176
rect 11223 -856 11279 -846
rect 11341 784 11397 794
rect 11341 -238 11397 176
rect 11341 -884 11397 -846
rect 11459 784 11515 822
rect 11459 -238 11515 176
rect 11459 -856 11515 -846
rect 11577 784 11633 794
rect 11577 -238 11633 176
rect 11577 -884 11633 -846
rect 11695 784 11751 822
rect 11695 -238 11751 176
rect 11695 -856 11751 -846
rect 11813 784 11869 794
rect 11813 -238 11869 176
rect 11813 -884 11869 -846
rect 11931 784 11987 822
rect 11931 -238 11987 176
rect 11931 -856 11987 -846
rect 12049 784 12105 794
rect 12049 -238 12105 176
rect 12049 -884 12105 -846
rect 12167 784 12223 822
rect 12167 -238 12223 176
rect 12167 -856 12223 -846
rect 12285 784 12341 794
rect 12285 -238 12341 176
rect 12285 -884 12341 -846
rect 12403 784 12459 822
rect 12403 -238 12459 176
rect 12403 -856 12459 -846
rect 12521 784 12577 794
rect 12521 -238 12577 176
rect 12521 -884 12577 -846
rect 12639 784 12695 822
rect 12639 -238 12695 176
rect 12639 -856 12695 -846
rect 12757 784 12813 794
rect 12757 -238 12813 176
rect 12757 -884 12813 -846
rect 12875 784 12931 822
rect 12875 -238 12931 176
rect 12875 -856 12931 -846
rect 12993 784 13049 794
rect 12993 -238 13049 176
rect 12993 -884 13049 -846
rect 13111 784 13167 822
rect 13111 -238 13167 176
rect 13111 -856 13167 -846
rect 13229 784 13285 794
rect 13229 -238 13285 176
rect 13229 -884 13285 -846
rect 13347 784 13403 822
rect 13347 -238 13403 176
rect 13347 -856 13403 -846
rect 13465 784 13521 794
rect 13465 -238 13521 176
rect 13465 -884 13521 -846
rect 13583 784 13639 822
rect 13583 -238 13639 176
rect 13583 -856 13639 -846
rect 13701 784 13757 794
rect 13701 -238 13757 176
rect 13701 -884 13757 -846
rect 13819 784 13875 822
rect 13819 -238 13875 176
rect 13819 -856 13875 -846
rect 13937 784 13993 794
rect 13937 -238 13993 176
rect 13937 -884 13993 -846
rect 14055 784 14111 822
rect 14292 794 14348 822
rect 14055 -238 14111 176
rect 14055 -856 14111 -846
rect 14173 784 14229 794
rect 14173 -238 14229 176
rect 14291 784 14348 794
rect 14347 176 14348 784
rect 14773 784 14829 822
rect 14291 166 14348 176
rect 14292 -228 14348 166
rect 14173 -884 14229 -846
rect 14291 -238 14348 -228
rect 14347 -239 14348 -238
rect 14416 377 14704 387
rect 14416 308 14704 318
rect 14416 -371 14703 308
rect 14773 -238 14829 176
rect 14416 -381 14704 -371
rect 14416 -445 14704 -435
rect 14416 -447 14703 -445
rect 14291 -856 14347 -846
rect 14773 -856 14829 -846
rect 14891 784 14947 794
rect 14891 -238 14947 176
rect 14891 -884 14947 -846
rect 15009 784 15065 822
rect 15009 -238 15065 176
rect 15009 -856 15065 -846
rect 15127 784 15183 794
rect 15127 -238 15183 176
rect 15127 -884 15183 -846
rect 15245 784 15301 822
rect 15245 -238 15301 176
rect 15245 -856 15301 -846
rect 15363 784 15419 794
rect 15363 -238 15419 176
rect 15363 -884 15419 -846
rect 15481 784 15537 822
rect 15481 -238 15537 176
rect 15481 -856 15537 -846
rect 15599 784 15655 794
rect 15599 -238 15655 176
rect 15599 -884 15655 -846
rect 15717 784 15773 822
rect 15717 -238 15773 176
rect 15717 -856 15773 -846
rect 15835 784 15891 794
rect 15835 -238 15891 176
rect 15835 -884 15891 -846
rect 15953 784 16009 822
rect 15953 -238 16009 176
rect 15953 -856 16009 -846
rect 16071 784 16127 794
rect 16071 -238 16127 176
rect 16071 -884 16127 -846
rect 16189 784 16245 822
rect 16189 -238 16245 176
rect 16189 -856 16245 -846
rect 16307 784 16363 794
rect 16307 -238 16363 176
rect 16307 -884 16363 -846
rect 16425 784 16481 822
rect 16425 -238 16481 176
rect 16425 -856 16481 -846
rect 16543 784 16599 794
rect 16543 -238 16599 176
rect 16543 -884 16599 -846
rect 16661 784 16717 822
rect 16661 -238 16717 176
rect 16661 -856 16717 -846
rect 16779 784 16835 794
rect 16779 -238 16835 176
rect 16779 -884 16835 -846
rect 16897 784 16953 822
rect 16897 -238 16953 176
rect 16897 -856 16953 -846
rect 17015 784 17071 794
rect 17015 -238 17071 176
rect 17015 -884 17071 -846
rect 17133 784 17189 822
rect 17133 -238 17189 176
rect 17133 -856 17189 -846
rect 17251 784 17307 794
rect 17251 -238 17307 176
rect 17251 -884 17307 -846
rect 17369 784 17425 822
rect 17369 -238 17425 176
rect 17369 -856 17425 -846
rect 17487 784 17543 794
rect 17487 -238 17543 176
rect 17487 -884 17543 -846
rect 17605 784 17661 822
rect 17605 -238 17661 176
rect 17605 -856 17661 -846
rect 17723 784 17779 794
rect 17723 -238 17779 176
rect 17723 -884 17779 -846
rect 17841 784 17897 822
rect 17841 -238 17897 176
rect 17841 -856 17897 -846
rect 17959 784 18015 794
rect 17959 -238 18015 176
rect 17959 -884 18015 -846
rect 18077 784 18133 822
rect 18077 -238 18133 176
rect 18077 -856 18133 -846
rect 18195 784 18251 794
rect 18195 -238 18251 176
rect 18195 -884 18251 -846
rect 18313 784 18369 822
rect 18313 -238 18369 176
rect 18313 -856 18369 -846
rect 18431 784 18487 794
rect 18431 -238 18487 176
rect 18431 -884 18487 -846
rect 18549 784 18605 822
rect 18549 -238 18605 176
rect 18549 -856 18605 -846
rect 18667 784 18723 794
rect 18667 -238 18723 176
rect 18667 -884 18723 -846
rect 18785 784 18841 822
rect 18785 -238 18841 176
rect 18785 -856 18841 -846
rect 18903 784 18959 794
rect 18903 -238 18959 176
rect 18903 -884 18959 -846
rect 19021 784 19077 822
rect 19021 -238 19077 176
rect 19021 -856 19077 -846
rect 19139 784 19195 794
rect 19139 -238 19195 176
rect 19139 -884 19195 -846
rect 19257 784 19313 822
rect 19257 -238 19313 176
rect 19257 -856 19313 -846
rect 19375 784 19431 794
rect 19375 -238 19431 176
rect 19375 -884 19431 -846
rect 19493 784 19549 822
rect 19493 -238 19549 176
rect 19493 -856 19549 -846
rect 19611 784 19667 794
rect 19611 -238 19667 176
rect 19611 -884 19667 -846
rect 19729 784 19785 822
rect 19729 -238 19785 176
rect 19729 -856 19785 -846
rect 19847 784 19903 794
rect 19847 -238 19903 176
rect 19847 -884 19903 -846
rect 19965 784 20021 822
rect 19965 -238 20021 176
rect 19965 -856 20021 -846
rect 20083 784 20139 794
rect 20083 -238 20139 176
rect 20083 -884 20139 -846
rect 20201 784 20257 822
rect 20201 -238 20257 176
rect 20201 -856 20257 -846
rect 20319 784 20375 794
rect 20319 -238 20375 176
rect 20319 -884 20375 -846
rect 20437 784 20493 822
rect 20674 794 20730 822
rect 20437 -238 20493 176
rect 20437 -856 20493 -846
rect 20555 784 20611 794
rect 20555 -238 20611 176
rect 20673 784 20730 794
rect 20729 176 20730 784
rect 20673 166 20730 176
rect 20674 -228 20730 166
rect 20555 -884 20611 -846
rect 20673 -238 20730 -228
rect 20729 -239 20730 -238
rect 20673 -856 20729 -846
rect 8509 -967 22770 -884
rect 8509 -972 15310 -967
rect 8509 -1083 9665 -972
rect 14264 -1078 15310 -972
rect 20658 -1078 22770 -967
rect 14264 -1083 22770 -1078
rect 8509 -1183 22770 -1083
rect 7122 -1870 7179 -1866
rect 7123 -2006 7179 -1870
rect 7659 -2006 7715 -1861
rect 8172 -2006 8292 -1996
rect 1226 -2146 8172 -2006
rect 1226 -2292 1282 -2146
rect 1226 -3710 1282 -3700
rect 1762 -2292 1818 -2146
rect 1762 -3710 1818 -3700
rect 2298 -2292 2354 -2146
rect 2298 -3710 2354 -3700
rect 2834 -2292 2890 -2146
rect 2834 -3710 2890 -3700
rect 3370 -2283 3426 -2146
rect 3370 -3711 3426 -3701
rect 3906 -2283 3962 -2146
rect 3906 -3711 3962 -3701
rect 4442 -2283 4498 -2146
rect 4442 -3711 4498 -3701
rect 4978 -2283 5034 -2146
rect 4978 -3711 5034 -3701
rect 5514 -2283 5570 -2146
rect 5514 -3711 5570 -3701
rect 6050 -2283 6106 -2146
rect 6050 -3711 6106 -3701
rect 6586 -2283 6642 -2146
rect 6586 -3711 6642 -3701
rect 7123 -2283 7179 -2146
rect 7123 -3711 7179 -3701
rect 7659 -2284 7715 -2146
rect 8172 -2156 8292 -2146
rect 7659 -3711 7715 -3701
rect 1226 -3981 1282 -3971
rect 1226 -5535 1282 -5389
rect 1762 -3981 1818 -3971
rect 1762 -5535 1818 -5389
rect 2298 -3981 2354 -3971
rect 2298 -5535 2354 -5389
rect 2834 -3981 2890 -3971
rect 2834 -5535 2890 -5389
rect 3370 -3981 3426 -3971
rect 3370 -5535 3426 -5389
rect 3906 -3981 3962 -3971
rect 3906 -5535 3962 -5389
rect 4442 -3981 4498 -3971
rect 4442 -5535 4498 -5389
rect 4978 -3982 5034 -3972
rect 4978 -5535 5034 -5390
rect 5514 -3981 5570 -3971
rect 5514 -5535 5570 -5389
rect 6050 -3981 6106 -3971
rect 6050 -5535 6106 -5389
rect 6586 -3981 6642 -3971
rect 6586 -5535 6642 -5389
rect 7122 -3981 7178 -3971
rect 7122 -5395 7178 -5389
rect 7659 -3982 7715 -3972
rect 7122 -5399 7179 -5395
rect 7123 -5535 7179 -5399
rect 7659 -5535 7715 -5390
rect 1226 -5675 8450 -5535
rect 1226 -5821 1282 -5675
rect 1226 -7239 1282 -7229
rect 1762 -5821 1818 -5675
rect 1762 -7239 1818 -7229
rect 2298 -5821 2354 -5675
rect 2298 -7239 2354 -7229
rect 2834 -5821 2890 -5675
rect 2834 -7239 2890 -7229
rect 3370 -5812 3426 -5675
rect 3370 -7240 3426 -7230
rect 3906 -5812 3962 -5675
rect 3906 -7240 3962 -7230
rect 4442 -5812 4498 -5675
rect 4442 -7240 4498 -7230
rect 4978 -5812 5034 -5675
rect 4978 -7240 5034 -7230
rect 5514 -5812 5570 -5675
rect 5514 -7240 5570 -7230
rect 6050 -5812 6106 -5675
rect 6050 -7240 6106 -7230
rect 6586 -5812 6642 -5675
rect 6586 -7240 6642 -7230
rect 7123 -5812 7179 -5675
rect 7123 -7240 7179 -7230
rect 7659 -5813 7715 -5675
rect 7659 -7240 7715 -7230
rect 8309 -7188 8450 -5675
rect 21166 -6869 22770 -1183
rect 13106 -7150 22770 -6869
rect 12712 -7188 12936 -7187
rect 8309 -7204 12936 -7188
rect 8309 -7557 12726 -7204
rect 6505 -7570 12726 -7557
rect 6505 -7640 10941 -7570
rect 1371 -7776 1427 -7766
rect 1371 -9942 1427 -9884
rect 2247 -7776 2303 -7766
rect 2247 -9942 2303 -9884
rect 3123 -7776 3179 -7766
rect 3123 -9942 3179 -9884
rect 3999 -7776 4055 -7766
rect 3999 -9942 4055 -9884
rect 4875 -7776 4931 -7766
rect 4875 -9942 4931 -9884
rect 5751 -7776 5807 -7766
rect 5751 -9942 5807 -9884
rect 6067 -7776 6123 -7766
rect 6067 -9942 6123 -9884
rect 6505 -7776 6561 -7640
rect 6505 -9894 6561 -9884
rect 6943 -7776 6999 -7766
rect 6943 -9942 6999 -9884
rect 7381 -7776 7437 -7640
rect 7381 -9894 7437 -9884
rect 7819 -7776 7875 -7766
rect 7819 -9942 7875 -9884
rect 8257 -7776 8313 -7640
rect 8257 -9894 8313 -9884
rect 8695 -7776 8751 -7766
rect 8695 -9942 8751 -9884
rect 9133 -7776 9189 -7640
rect 9133 -9894 9189 -9884
rect 9571 -7776 9627 -7766
rect 9571 -9942 9627 -9884
rect 10009 -7776 10065 -7640
rect 10009 -9894 10065 -9884
rect 10447 -7776 10503 -7766
rect 10447 -9942 10503 -9884
rect 10885 -7776 10941 -7640
rect 11219 -7776 11279 -7570
rect 11219 -8094 11279 -8084
rect 11407 -7776 11471 -7570
rect 11407 -8094 11471 -8084
rect 11599 -7776 11663 -7570
rect 11599 -8094 11663 -8084
rect 11791 -7776 11855 -7570
rect 11791 -8094 11855 -8084
rect 11983 -7776 12047 -7570
rect 11983 -8094 12047 -8084
rect 12175 -7776 12239 -7570
rect 12175 -8094 12239 -8084
rect 12367 -7776 12431 -7570
rect 12367 -8094 12431 -8084
rect 12559 -7776 12623 -7570
rect 12559 -8094 12623 -8084
rect 11320 -8138 12512 -8128
rect 11320 -8208 12512 -8198
rect 12712 -9409 12726 -7570
rect 12923 -9409 12936 -7204
rect 12712 -9452 12936 -9409
rect 13106 -9745 13170 -7150
rect 13298 -9746 13362 -7150
rect 13490 -9746 13554 -7150
rect 13682 -9746 13746 -7150
rect 13874 -9746 13938 -7150
rect 14066 -9746 14130 -7150
rect 14258 -9746 14322 -7150
rect 14450 -9746 14514 -7150
rect 14642 -9746 14706 -7150
rect 14834 -9746 14898 -7150
rect 15026 -9746 15090 -7150
rect 15218 -9746 15282 -7150
rect 15410 -9746 15474 -7150
rect 15602 -9746 15666 -7150
rect 15794 -9746 15858 -7150
rect 15986 -9746 16050 -7150
rect 16178 -9746 16242 -7150
rect 16370 -9746 16434 -7150
rect 16562 -9746 16626 -7150
rect 16754 -9746 16818 -7150
rect 16946 -9746 17010 -7150
rect 17138 -9746 17202 -7150
rect 17330 -9746 17394 -7150
rect 17522 -9746 17586 -7150
rect 17714 -9746 17778 -7150
rect 17906 -9746 17970 -7150
rect 18098 -9746 18162 -7150
rect 18290 -9746 18354 -7150
rect 18482 -9746 18546 -7150
rect 18674 -9746 18738 -7150
rect 18866 -9746 18930 -7150
rect 19058 -9746 19122 -7150
rect 19250 -9746 19314 -7150
rect 19442 -9756 19506 -7150
rect 19634 -9756 19698 -7150
rect 19826 -9756 19890 -7150
rect 20018 -9756 20082 -7150
rect 20210 -9756 20274 -7150
rect 20402 -9756 20466 -7150
rect 20594 -9756 20658 -7150
rect 20786 -9756 20850 -7150
rect 20978 -9756 21042 -7150
rect 21170 -9756 21234 -7150
rect 21362 -9756 21426 -7150
rect 21554 -9756 21618 -7150
rect 21746 -9756 21810 -7150
rect 21938 -9756 22002 -7150
rect 22130 -9756 22194 -7150
rect 22322 -9756 22386 -7150
rect 22514 -9756 22578 -7150
rect 22706 -9756 22770 -7150
rect 10885 -9894 10941 -9884
rect 836 -10066 10951 -9942
rect 836 -10132 10951 -10122
<< via2 >>
rect 9665 -1083 14264 -972
rect 15310 -1078 20658 -967
rect 11320 -8141 12512 -8138
rect 11320 -8195 12512 -8141
rect 11320 -8198 12512 -8195
<< metal3 >>
rect 15300 -967 20668 -962
rect 9655 -972 14274 -967
rect 9655 -1083 9665 -972
rect 14264 -1083 14274 -972
rect 15300 -1078 15310 -967
rect 20658 -1078 20668 -967
rect 15300 -1083 20668 -1078
rect 9655 -1088 14274 -1083
rect 8525 -6350 14947 -5755
rect 11716 -8133 12078 -6350
rect 11310 -8138 12522 -8133
rect 11310 -8198 11320 -8138
rect 12512 -8198 12522 -8138
rect 11310 -8203 12522 -8198
<< via3 >>
rect 9665 -1083 14264 -972
rect 15310 -1078 20658 -967
<< metal4 >>
rect 15309 -967 20659 -966
rect 9664 -972 14265 -971
rect 9664 -1083 9665 -972
rect 14264 -1083 14265 -972
rect 15309 -1078 15310 -967
rect 20658 -1078 20659 -967
rect 15309 -1079 20659 -1078
rect 9664 -1084 14265 -1083
rect 9665 -1658 14260 -1084
rect 15310 -1538 20658 -1079
use sky130_fd_pr__pfet_01v8_lvt_7XCYSC  sky130_fd_pr__pfet_01v8_lvt_7XCYSC_1
timestamp 1615997521
transform 1 0 4336 0 1 -6489
box -3517 -884 3517 884
use sky130_fd_pr__pfet_01v8_lvt_RTJWSN  sky130_fd_pr__pfet_01v8_lvt_RTJWSN_1
timestamp 1615997521
transform 1 0 4336 0 1 -4721
box -3517 -884 3517 884
use sky130_fd_pr__nfet_01v8_QVUSYJ  sky130_fd_pr__nfet_01v8_QVUSYJ_0
timestamp 1616176710
transform 1 0 3370 0 1 -8799
box -2576 -1229 2576 1229
use sky130_fd_pr__nfet_01v8_QVUSYJ  sky130_fd_pr__nfet_01v8_QVUSYJ_1
timestamp 1616176710
transform 1 0 8504 0 1 -8799
box -2576 -1229 2576 1229
use sky130_fd_pr__pfet_01v8_lvt_RTJWSN  sky130_fd_pr__pfet_01v8_lvt_RTJWSN_0
timestamp 1615997521
transform 1 0 4336 0 1 -1192
box -3517 -884 3517 884
use sky130_fd_pr__pfet_01v8_lvt_7XCYSC  sky130_fd_pr__pfet_01v8_lvt_7XCYSC_0
timestamp 1615997521
transform 1 0 4336 0 1 -2960
box -3517 -884 3517 884
use sky130_fd_pr__pfet_01v8_65PBSZ  sky130_fd_pr__pfet_01v8_65PBSZ_0
timestamp 1616185029
transform 1 0 11369 0 1 444
box -3117 -484 3117 484
use sky130_fd_pr__pfet_01v8_K4PBSX  sky130_fd_pr__pfet_01v8_K4PBSX_0
timestamp 1616600406
transform 1 0 11369 0 1 -506
box -3117 -484 3117 484
use sky130_fd_pr__pfet_01v8_H98ZZM  sky130_fd_pr__pfet_01v8_H98ZZM_0
timestamp 1615909117
transform 1 0 5145 0 1 369
box -3117 -409 3117 409
use sky130_fd_pr__pfet_01v8_698KZZ  sky130_fd_pr__pfet_01v8_698KZZ_0
timestamp 1619042825
transform 1 0 985 0 1 293
box -1052 -334 1052 334
use sky130_fd_pr__cap_mim_m3_1_XFP5BZ  sky130_fd_pr__cap_mim_m3_1_XFP5BZ_1
timestamp 1616703757
transform -1 0 11666 0 1 -4033
box -3150 -2850 3149 2850
use sky130_fd_pr__pfet_01v8_K4PBSX  sky130_fd_pr__pfet_01v8_K4PBSX_1
timestamp 1616600406
transform 1 0 17751 0 1 -506
box -3117 -484 3117 484
use sky130_fd_pr__cap_mim_m3_1_XFP5BZ  sky130_fd_pr__cap_mim_m3_1_XFP5BZ_0
timestamp 1616703757
transform -1 0 17961 0 1 -4021
box -3150 -2850 3149 2850
use sky130_fd_pr__nfet_01v8_J9MTE9  sky130_fd_pr__nfet_01v8_J9MTE9_0
timestamp 1619042384
transform 1 0 11919 0 1 -7930
box -839 -360 839 360
use sky130_fd_pr__pfet_01v8_65PBSZ  sky130_fd_pr__pfet_01v8_65PBSZ_1
timestamp 1616185029
transform 1 0 17751 0 1 444
box -3117 -484 3117 484
use sky130_fd_pr__nfet_01v8_Z2S3N8  sky130_fd_pr__nfet_01v8_Z2S3N8_0
timestamp 1616876989
transform 1 0 17938 0 1 -9592
box -4967 -360 4967 360
use sky130_fd_pr__nfet_01v8_Z2S3N8  sky130_fd_pr__nfet_01v8_Z2S3N8_1
timestamp 1616876989
transform 1 0 17938 0 1 -8872
box -4967 -360 4967 360
use sky130_fd_pr__nfet_01v8_Z2S3N8  sky130_fd_pr__nfet_01v8_Z2S3N8_2
timestamp 1616876989
transform 1 0 17938 0 1 -8152
box -4967 -360 4967 360
use sky130_fd_pr__nfet_01v8_Z2S3N8  sky130_fd_pr__nfet_01v8_Z2S3N8_3
timestamp 1616876989
transform 1 0 17938 0 1 -7432
box -4967 -360 4967 360
<< labels >>
rlabel nwell 66 973 8178 1089 1 vdd
rlabel pwell 12690 -10122 22854 -9975 1 vss
rlabel metal2 21166 -7150 22770 -884 1 vout
rlabel metal1 796 -344 8133 -97 1 vp
rlabel metal1 63 -425 471 -79 1 iref
rlabel metal1 64 -2249 627 -1903 1 vin_p
rlabel metal1 514 -5778 821 -5432 1 vin_n
<< end >>
