magic
tech sky130A
magscale 1 2
timestamp 1624389981
<< poly >>
rect -78 86 -6 102
rect -78 46 -62 86
rect -22 46 -6 86
rect -78 28 -6 46
rect -56 -99 -26 28
rect 106 -746 174 -730
rect 106 -780 122 -746
rect 156 -780 174 -746
rect 106 -792 174 -780
rect -56 -5074 -26 -4681
rect -74 -5090 -8 -5074
rect -74 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -74 -5140 -8 -5124
<< polycont >>
rect -62 46 -22 86
rect 122 -780 156 -746
rect -58 -5124 -24 -5090
<< locali >>
rect -78 86 -6 102
rect -78 46 -62 86
rect -22 46 -6 86
rect -78 28 -6 46
rect 106 -746 172 -730
rect 106 -780 122 -746
rect 156 -780 172 -746
rect 106 -792 172 -780
rect -74 -5090 -8 -5074
rect -74 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -74 -5140 -8 -5124
<< viali >>
rect -62 46 -22 86
rect 122 -780 156 -746
rect -58 -5124 -24 -5090
<< metal1 >>
rect -2253 6098 -5 6110
rect -2268 6008 -2258 6098
rect -2052 6051 -5 6098
rect -2052 6008 -2042 6051
rect -2654 5184 -114 5196
rect -2664 5040 -2654 5184
rect -2452 5040 -114 5184
rect 2740 4616 2750 4676
rect 2810 4618 2820 4676
rect 2810 4616 2842 4618
rect 11574 4232 11584 4878
rect 13530 4232 13540 4878
rect -2262 4124 -2252 4194
rect -2048 4189 -2038 4194
rect -2048 4130 -5 4189
rect -2048 4124 -2038 4130
rect 6416 3846 6995 3881
rect 11586 3858 12170 4232
rect 1088 3230 1098 3290
rect 1158 3230 1168 3290
rect 6416 2617 6446 3846
rect 6963 2802 6995 3846
rect 12592 3802 13176 4232
rect 6963 2756 7225 2802
rect 6963 2700 7249 2756
rect 6963 2660 7225 2700
rect 16561 2661 17414 2664
rect 6963 2617 7282 2660
rect 15887 2649 17414 2661
rect 6416 2572 7282 2617
rect 14318 1919 14328 2475
rect 15492 1919 15502 2475
rect 15885 2112 15895 2649
rect 17398 2112 17414 2649
rect 15887 2101 17414 2112
rect 14764 1515 14774 1919
rect 15152 1515 15162 1919
rect -536 98 -10 99
rect -546 30 -536 98
rect -336 86 -10 98
rect -336 46 -62 86
rect -22 46 -10 86
rect -336 30 -10 46
rect -186 -216 -176 -18
rect 12 -216 22 -18
rect 7180 -273 7666 368
rect 7840 -273 8326 377
rect 16539 373 17392 376
rect 8554 -273 9166 365
rect 15865 361 17392 373
rect 7180 -337 7192 -273
rect 7182 -514 7192 -337
rect 9157 -514 9167 -273
rect 14318 -322 14328 234
rect 15492 -322 15502 234
rect 15863 -176 15873 361
rect 17376 -176 17392 361
rect 15865 -187 17392 -176
rect 14774 -369 15152 -322
rect 14768 -722 14778 -369
rect 15145 -722 15155 -369
rect 96 -792 106 -730
rect 174 -792 184 -730
rect 14810 -732 14838 -722
rect 52 -1138 118 -1040
rect 52 -1190 62 -1138
rect 114 -1190 124 -1138
rect 52 -1286 118 -1190
rect -2698 -1764 -2688 -1526
rect -2428 -1531 -2418 -1526
rect -1846 -1531 -1836 -1526
rect -2428 -1760 -1836 -1531
rect -2428 -1764 -2418 -1760
rect -1846 -1764 -1836 -1760
rect -1576 -1764 -1566 -1526
rect 16523 -1889 17376 -1886
rect -2288 -2134 -2278 -1896
rect -2018 -1901 -2008 -1896
rect -1836 -1901 -1826 -1894
rect -2018 -2130 -1826 -1901
rect -2018 -2134 -2008 -2130
rect -1836 -2132 -1826 -2130
rect -1566 -2132 -1556 -1894
rect -1842 -2496 -1832 -2258
rect -1572 -2262 -1562 -2258
rect -1572 -2263 -1132 -2262
rect -1572 -2491 -1348 -2263
rect -1572 -2496 -1562 -2491
rect -1358 -2492 -1348 -2491
rect -1119 -2492 -1109 -2263
rect 7158 -2569 7737 -1920
rect 7961 -2569 8270 -1891
rect 15849 -1901 17376 -1889
rect 8549 -2569 9128 -1902
rect -1842 -2888 -1832 -2650
rect -1572 -2659 -1562 -2650
rect -958 -2659 -948 -2657
rect -1572 -2886 -948 -2659
rect -719 -2886 -709 -2657
rect 7143 -2779 7153 -2569
rect 9130 -2779 9140 -2569
rect 14318 -2622 14328 -2066
rect 15492 -2622 15502 -2066
rect 15847 -2438 15857 -1901
rect 17360 -2438 17376 -1901
rect 15849 -2449 17376 -2438
rect 14774 -2800 15152 -2622
rect -1572 -2888 -736 -2886
rect 14764 -3058 14774 -2800
rect 15152 -3058 15162 -2800
rect -1842 -3314 -1832 -3076
rect -1572 -3081 -1562 -3076
rect -1572 -3310 -550 -3081
rect -321 -3310 -311 -3081
rect -1572 -3314 -1562 -3310
rect 52 -3484 118 -3386
rect 52 -3536 64 -3484
rect 116 -3536 126 -3484
rect 52 -3632 118 -3536
rect 16531 -4179 17384 -4176
rect 15857 -4191 17384 -4179
rect 3722 -4712 3732 -4546
rect 3898 -4712 3908 -4546
rect 15855 -4728 15865 -4191
rect 17368 -4728 17384 -4191
rect 15857 -4739 17384 -4728
rect -546 -5140 -536 -5074
rect -336 -5090 -8 -5074
rect -336 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -336 -5140 -8 -5124
rect -2260 -5328 -2250 -5264
rect -2050 -5284 -2040 -5264
rect -2050 -5317 518 -5284
rect -2050 -5328 -2040 -5317
rect 346 -5368 518 -5317
rect 90 -5510 164 -5508
rect -1344 -5562 -1334 -5510
rect -1134 -5562 164 -5510
rect 90 -5564 164 -5562
rect 228 -5564 238 -5508
rect -2664 -6178 -2654 -6118
rect -2454 -6124 -2444 -6118
rect 7577 -6122 7587 -5951
rect -2454 -6170 -104 -6124
rect 7112 -6169 7587 -6122
rect -2454 -6178 -2444 -6170
rect 7577 -6327 7587 -6169
rect 9188 -6327 9198 -5951
rect -942 -6656 -932 -6596
rect -732 -6656 -182 -6596
rect -122 -6656 -112 -6596
rect -2258 -6974 -2248 -6916
rect -2050 -6919 -2040 -6916
rect -2050 -6922 -198 -6919
rect -2050 -6968 -66 -6922
rect -2050 -6970 -198 -6968
rect -2050 -6974 -2040 -6970
<< via1 >>
rect -2258 6008 -2052 6098
rect -2654 5040 -2452 5184
rect 2750 4616 2810 4676
rect 11584 4232 13530 4878
rect -2252 4124 -2048 4194
rect 1098 3230 1158 3290
rect 6446 2617 6963 3846
rect 14328 1919 15492 2475
rect 15895 2112 17398 2649
rect 14774 1515 15152 1919
rect -536 30 -336 98
rect -176 -216 12 -18
rect 7192 -514 9157 -273
rect 14328 -322 15492 234
rect 15873 -176 17376 361
rect 14778 -722 15145 -369
rect 106 -746 174 -730
rect 106 -780 122 -746
rect 122 -780 156 -746
rect 156 -780 174 -746
rect 106 -792 174 -780
rect 62 -1190 114 -1138
rect -2688 -1764 -2428 -1526
rect -1836 -1764 -1576 -1526
rect -2278 -2134 -2018 -1896
rect -1826 -2132 -1566 -1894
rect -1832 -2496 -1572 -2258
rect -1348 -2492 -1119 -2263
rect -1832 -2888 -1572 -2650
rect -948 -2886 -719 -2657
rect 7153 -2779 9130 -2569
rect 14328 -2622 15492 -2066
rect 15857 -2438 17360 -1901
rect 14774 -3058 15152 -2800
rect -1832 -3314 -1572 -3076
rect -550 -3310 -321 -3081
rect 64 -3536 116 -3484
rect 3732 -4712 3898 -4546
rect 15865 -4728 17368 -4191
rect -536 -5140 -336 -5074
rect -2250 -5328 -2050 -5264
rect -1334 -5562 -1134 -5510
rect 164 -5564 228 -5508
rect -2654 -6178 -2454 -6118
rect 7587 -6327 9188 -5951
rect -932 -6656 -732 -6596
rect -182 -6656 -122 -6596
rect -2248 -6974 -2050 -6916
<< metal2 >>
rect -2258 6098 -2052 6108
rect -2652 5194 -2452 6040
rect -2052 6008 -2050 6040
rect -2258 5998 -2050 6008
rect -2654 5184 -2452 5194
rect -2654 5030 -2452 5040
rect -2652 2828 -2452 5030
rect -2250 4204 -2050 5998
rect -1334 6036 -1134 6084
rect -2252 4194 -2048 4204
rect -2252 4114 -2048 4124
rect -2654 2818 -2452 2828
rect -2654 2728 -2452 2738
rect -2652 -20 -2452 2728
rect -2456 -216 -2452 -20
rect -2652 -1516 -2452 -216
rect -2250 1956 -2050 4114
rect -2052 1896 -2050 1956
rect -2688 -1526 -2428 -1516
rect -2688 -1774 -2428 -1764
rect -2652 -6108 -2452 -1774
rect -2250 -1886 -2050 1896
rect -1334 3288 -1134 5964
rect -1334 -1134 -1134 3230
rect -932 4564 -732 6084
rect -536 4712 -336 6056
rect 1494 6026 1560 6036
rect 1494 5958 1560 5968
rect 2812 5888 2872 5898
rect 2786 5828 2812 5886
rect 2786 5818 2872 5828
rect 9648 5836 9906 5846
rect 2786 5712 2846 5818
rect 6110 5752 6170 5762
rect 6110 5682 6170 5692
rect 9906 5600 9910 5836
rect 9648 5598 9910 5600
rect 10239 5834 10499 5844
rect 9648 5590 9906 5598
rect 10239 5592 10499 5602
rect 10791 5832 11074 5842
rect 10791 5596 10800 5832
rect 11058 5596 11074 5832
rect 10791 5587 11074 5596
rect 11584 4878 13530 4888
rect -538 4702 -334 4712
rect -538 4630 -334 4640
rect 232 4708 292 4718
rect 232 4638 292 4648
rect 2750 4676 2810 4686
rect -736 4508 -732 4564
rect -932 2468 -732 4508
rect -940 2458 -732 2468
rect -734 2400 -732 2458
rect -940 2390 -732 2400
rect -932 -720 -732 2390
rect -937 -730 -732 -720
rect -734 -792 -732 -730
rect -937 -802 -732 -792
rect -1836 -1526 -1576 -1516
rect -1836 -1774 -1576 -1764
rect -2278 -1896 -2018 -1886
rect -2278 -2144 -2018 -2134
rect -1826 -1894 -1566 -1884
rect -1826 -2142 -1566 -2132
rect -2654 -6118 -2452 -6108
rect -2454 -6178 -2452 -6118
rect -2654 -6188 -2452 -6178
rect -2652 -6960 -2452 -6188
rect -2250 -4534 -2050 -2144
rect -1832 -2258 -1572 -2248
rect -1334 -2253 -1134 -1194
rect -1832 -2506 -1572 -2496
rect -1348 -2263 -1119 -2253
rect -1348 -2502 -1119 -2492
rect -1832 -2650 -1572 -2640
rect -1832 -2898 -1572 -2888
rect -1832 -3076 -1572 -3066
rect -1832 -3324 -1572 -3314
rect -1334 -3480 -1134 -2502
rect -932 -2647 -732 -802
rect -536 710 -336 4630
rect 2750 4606 2810 4616
rect 6106 4554 6168 4564
rect 2786 4420 2846 4514
rect 6106 4469 6168 4479
rect 2786 4410 2872 4420
rect 2786 4350 2812 4410
rect 2812 4340 2872 4350
rect 11584 4222 13530 4232
rect 16041 4138 16143 4147
rect 3002 4119 3062 4126
rect 2992 4116 6146 4119
rect 2992 4057 3002 4116
rect 3062 4057 6146 4116
rect 3002 4046 3062 4056
rect 5934 4002 5994 4012
rect 2804 3986 2876 3996
rect 2876 3914 5692 3986
rect 2804 3904 2876 3914
rect 1098 3290 1158 3300
rect 1098 3220 1158 3230
rect 2398 3290 2458 3300
rect 2398 3220 2458 3230
rect 5112 3294 5172 3304
rect 5112 3224 5172 3234
rect -120 2810 -60 2820
rect -120 2740 -60 2750
rect 264 2460 324 2470
rect 264 2390 324 2400
rect 5620 2136 5692 3914
rect 5934 3932 5994 3942
rect 5934 3862 6010 3932
rect 5620 2076 5624 2136
rect 5684 2076 5692 2136
rect 5620 2074 5692 2076
rect 5786 3850 5858 3860
rect 5624 2066 5684 2074
rect 2522 1956 2582 1966
rect 2522 1886 2582 1896
rect 2398 1694 2458 1704
rect 2398 1624 2458 1634
rect 5114 1694 5174 1704
rect 5114 1624 5174 1634
rect -536 98 -336 648
rect 2358 708 2418 718
rect 2358 638 2418 648
rect -948 -2657 -719 -2647
rect -948 -2896 -719 -2886
rect -2250 -4544 -2048 -4534
rect -2250 -4712 -2247 -4544
rect -2250 -4722 -2048 -4712
rect -2250 -5264 -2050 -4722
rect -2250 -6916 -2050 -5328
rect -1334 -5510 -1134 -3540
rect -1334 -6916 -1134 -5562
rect -932 -6596 -732 -2896
rect -536 -3071 -336 30
rect -176 -18 12 -8
rect 5786 -154 5858 3778
rect 5786 -214 5794 -154
rect 5854 -214 5858 -154
rect -176 -226 12 -216
rect 5794 -224 5854 -214
rect 106 -730 174 -720
rect 106 -802 174 -792
rect 3042 -766 3102 -756
rect 3042 -836 3102 -826
rect 58 -1134 118 -1124
rect 58 -1204 118 -1194
rect 3046 -1496 3106 -1486
rect 3046 -1566 3106 -1556
rect 5948 -2416 6010 3862
rect 5948 -2488 6010 -2478
rect -550 -3081 -321 -3071
rect 3038 -3106 3110 -3096
rect 3038 -3188 3110 -3178
rect -550 -3320 -321 -3310
rect -932 -6916 -732 -6656
rect -536 -5074 -336 -3320
rect 60 -3480 120 -3470
rect 60 -3550 120 -3540
rect 3044 -3844 3104 -3834
rect 3044 -3914 3104 -3904
rect 3732 -4546 3898 -4536
rect 3732 -4722 3898 -4712
rect 6084 -4702 6146 4057
rect 16041 4057 16050 4138
rect 16134 4057 16143 4138
rect 16041 4054 16143 4057
rect 9671 3991 9888 4001
rect 9671 3913 9888 3923
rect 6446 3846 6963 3856
rect 6250 3294 6310 3302
rect 6248 3292 6310 3294
rect 6248 3232 6250 3292
rect 6248 -2246 6310 3232
rect 16071 3827 16123 4054
rect 17278 3224 17770 3294
rect 17510 3056 17770 3224
rect 6446 2607 6963 2617
rect 15895 2649 17398 2659
rect 6825 2558 6890 2560
rect 7717 2558 7777 2568
rect 12192 2558 12252 2568
rect 6824 2498 7717 2558
rect 7777 2498 12192 2558
rect 6522 2432 6586 2442
rect 6518 2368 6522 2432
rect 6586 2368 6590 2432
rect 6246 -2256 6310 -2246
rect 6308 -2318 6310 -2256
rect 6246 -2323 6310 -2318
rect 6372 1694 6432 1704
rect 6246 -2328 6308 -2323
rect 6372 -4544 6432 1634
rect 6518 -767 6590 2368
rect 6674 142 6734 152
rect 6583 -832 6590 -767
rect 6518 -834 6590 -832
rect 6668 82 6674 140
rect 6734 82 6740 140
rect 6518 -842 6583 -834
rect 6668 -1400 6740 82
rect 6668 -1428 6742 -1400
rect 6670 -1490 6742 -1428
rect 6670 -1572 6742 -1562
rect 6825 -1604 6890 2498
rect 7717 2488 7777 2498
rect 12192 2488 12252 2498
rect 14328 2475 15492 2485
rect 8244 2432 8304 2440
rect 12717 2432 12777 2442
rect 8244 2430 12717 2432
rect 8304 2372 12717 2430
rect 8244 2360 8304 2370
rect 12717 2362 12777 2372
rect 9220 2316 9280 2326
rect 13654 2316 13714 2326
rect 9280 2256 13654 2316
rect 9220 2246 9280 2256
rect 13654 2246 13714 2256
rect 9754 2198 9814 2208
rect 14170 2198 14230 2208
rect 9814 2138 14170 2198
rect 9754 2128 9814 2138
rect 14170 2128 14230 2138
rect 15895 2102 17398 2112
rect 14328 1909 14774 1919
rect 9670 1701 9887 1711
rect 9670 1623 9887 1633
rect 15152 1909 15492 1919
rect 16019 1850 16121 1859
rect 16019 1769 16028 1850
rect 16112 1769 16121 1850
rect 16019 1766 16121 1769
rect 16049 1539 16101 1766
rect 14774 1505 15152 1515
rect 17256 936 17748 1006
rect 17488 768 17748 936
rect 15873 361 17376 371
rect 7694 276 7754 286
rect 12170 276 12230 286
rect 6372 -4614 6432 -4604
rect 6658 -1669 6890 -1604
rect 6968 216 7694 276
rect 7754 216 12170 276
rect 6144 -4762 6146 -4702
rect 6084 -4780 6146 -4762
rect 2768 -5009 2828 -5002
rect 6658 -5009 6723 -1669
rect 6968 -1792 7028 216
rect 7694 206 7754 216
rect 12170 206 12230 216
rect 14328 234 15492 244
rect 8222 144 8282 152
rect 12695 144 12755 154
rect 8222 142 12695 144
rect 8282 84 12695 142
rect 8222 72 8282 82
rect 12695 74 12755 84
rect 9198 28 9258 38
rect 13632 28 13692 38
rect 9258 -32 13632 28
rect 9198 -42 9258 -32
rect 13632 -42 13692 -32
rect 9732 -90 9792 -80
rect 14148 -90 14208 -80
rect 9792 -150 14148 -90
rect 9732 -160 9792 -150
rect 14148 -160 14208 -150
rect 7192 -273 9157 -263
rect 15873 -186 17376 -176
rect 14328 -332 15492 -322
rect 7192 -524 9157 -514
rect 14774 -369 15152 -332
rect 9672 -557 9887 -547
rect 9672 -637 9887 -627
rect 14774 -722 14778 -369
rect 15145 -722 15152 -369
rect 16003 -412 16105 -403
rect 16003 -493 16012 -412
rect 16096 -493 16105 -412
rect 16003 -496 16105 -493
rect 14774 -727 15152 -722
rect 16033 -723 16085 -496
rect 14778 -732 15145 -727
rect 17240 -1428 17732 -1358
rect 17472 -1596 17732 -1428
rect 2766 -5012 6723 -5009
rect 2766 -5072 2768 -5012
rect 2828 -5072 6723 -5012
rect 6802 -1852 7028 -1792
rect 6802 -4998 6870 -1852
rect 15857 -1901 17360 -1891
rect 7679 -1982 7739 -1972
rect 6802 -5058 6806 -4998
rect 6866 -5058 6870 -4998
rect 6802 -5060 6870 -5058
rect 6960 -2042 7679 -1984
rect 12154 -1984 12214 -1974
rect 7739 -2042 12154 -1984
rect 6960 -2044 12154 -2042
rect 6806 -5068 6866 -5060
rect 2766 -5074 6723 -5072
rect 2768 -5082 2828 -5074
rect -536 -5369 -336 -5140
rect 4502 -5134 4562 -5124
rect 6960 -5134 7020 -2044
rect 7679 -2052 7739 -2044
rect 12154 -2054 12214 -2044
rect 14328 -2066 15492 -2056
rect 8206 -2118 8266 -2110
rect 12679 -2118 12739 -2108
rect 8206 -2120 12679 -2118
rect 8266 -2178 12679 -2120
rect 8206 -2190 8266 -2180
rect 12679 -2188 12739 -2178
rect 9182 -2234 9242 -2224
rect 13616 -2234 13676 -2224
rect 9242 -2294 13616 -2234
rect 9182 -2304 9242 -2294
rect 13616 -2304 13676 -2294
rect 9716 -2352 9776 -2342
rect 14132 -2352 14192 -2342
rect 9776 -2412 14132 -2352
rect 9716 -2422 9776 -2412
rect 14132 -2422 14192 -2412
rect 7153 -2569 9130 -2559
rect 15857 -2448 17360 -2438
rect 14328 -2632 15492 -2622
rect 7153 -2789 9130 -2779
rect 14774 -2800 15152 -2632
rect 16020 -2702 16104 -2692
rect 16020 -2793 16104 -2783
rect 9671 -2854 9887 -2844
rect 9671 -2932 9887 -2922
rect 16041 -2982 16093 -2793
rect 14774 -3068 15152 -3058
rect 17250 -3616 17740 -3546
rect 17480 -3784 17740 -3616
rect 15865 -4191 17368 -4181
rect 7687 -4290 7747 -4280
rect 12162 -4290 12222 -4280
rect 7396 -4350 7687 -4290
rect 7747 -4350 12162 -4290
rect 4562 -5194 7020 -5134
rect 7397 -4360 7460 -4350
rect 7687 -4360 7747 -4350
rect 12162 -4360 12222 -4350
rect 4502 -5204 4562 -5194
rect 738 -5256 798 -5246
rect 7397 -5254 7457 -4360
rect 8214 -4408 8274 -4400
rect 12687 -4408 12747 -4398
rect 8214 -4410 12687 -4408
rect 8274 -4468 12687 -4410
rect 8214 -4480 8274 -4470
rect 12687 -4478 12747 -4468
rect 9190 -4524 9250 -4514
rect 13624 -4524 13684 -4514
rect 9250 -4584 13624 -4524
rect 9190 -4594 9250 -4584
rect 13624 -4594 13684 -4584
rect 9724 -4642 9784 -4632
rect 14140 -4642 14200 -4632
rect 9784 -4702 14140 -4642
rect 9724 -4712 9784 -4702
rect 14140 -4712 14200 -4702
rect 15865 -4738 17368 -4728
rect 7396 -5256 7458 -5254
rect 798 -5316 7458 -5256
rect 738 -5326 798 -5316
rect -536 -5397 204 -5369
rect -2250 -6960 -2248 -6916
rect -536 -6944 -336 -5397
rect 164 -5508 228 -5498
rect 164 -5574 228 -5564
rect 738 -5720 798 -5710
rect 738 -5790 798 -5780
rect 4500 -5718 4560 -5708
rect 4500 -5788 4560 -5778
rect 7587 -5951 9188 -5941
rect 7587 -6337 9188 -6327
rect 2768 -6512 2828 -6502
rect 2768 -6582 2828 -6572
rect 6534 -6514 6594 -6504
rect 6534 -6584 6594 -6574
rect -182 -6596 -122 -6586
rect -122 -6640 -30 -6612
rect -182 -6666 -122 -6656
rect -2248 -6984 -2050 -6974
<< via2 >>
rect -1334 5964 -1134 6036
rect -2654 2738 -2452 2818
rect -2652 -216 -2456 -20
rect -2250 1896 -2052 1956
rect -1334 3230 -1134 3288
rect 1494 5968 1560 6026
rect 2812 5828 2872 5888
rect 6110 5692 6170 5752
rect 9648 5600 9906 5836
rect 10239 5602 10499 5834
rect 10800 5596 11058 5832
rect -538 4640 -334 4702
rect 232 4648 292 4708
rect -932 4508 -736 4564
rect -940 2400 -734 2458
rect -937 -792 -734 -730
rect -1334 -1194 -1134 -1134
rect 2750 4616 2810 4676
rect 6106 4479 6168 4554
rect 2812 4350 2872 4410
rect 11584 4232 13530 4878
rect 3002 4056 3062 4116
rect 2804 3914 2876 3986
rect 1098 3230 1158 3290
rect 2398 3230 2458 3290
rect 5112 3234 5172 3294
rect -120 2750 -60 2810
rect 264 2400 324 2460
rect 5934 3942 5994 4002
rect 5624 2076 5684 2136
rect 5786 3778 5858 3850
rect 2522 1896 2582 1956
rect 2398 1634 2458 1694
rect 5114 1634 5174 1694
rect -536 648 -336 710
rect 2358 648 2418 708
rect -1334 -3540 -1134 -3480
rect -2247 -4712 -2048 -4544
rect -176 -216 12 -18
rect 5794 -214 5854 -154
rect 106 -792 174 -730
rect 3042 -826 3102 -766
rect 58 -1138 118 -1134
rect 58 -1190 62 -1138
rect 62 -1190 114 -1138
rect 114 -1190 118 -1138
rect 58 -1194 118 -1190
rect 3046 -1556 3106 -1496
rect 5948 -2478 6010 -2416
rect 3038 -3178 3110 -3106
rect 60 -3484 120 -3480
rect 60 -3536 64 -3484
rect 64 -3536 116 -3484
rect 116 -3536 120 -3484
rect 60 -3540 120 -3536
rect 3044 -3904 3104 -3844
rect 3732 -4712 3898 -4546
rect 16050 4057 16134 4138
rect 9671 3923 9888 3991
rect 6250 3232 6310 3292
rect 6446 2617 6963 3846
rect 7717 2498 7777 2558
rect 12192 2498 12252 2558
rect 6522 2368 6586 2432
rect 6246 -2318 6308 -2256
rect 6372 1634 6432 1694
rect 6518 -832 6583 -767
rect 6674 82 6734 142
rect 6670 -1562 6742 -1490
rect 8244 2370 8304 2430
rect 12717 2372 12777 2432
rect 9220 2256 9280 2316
rect 13654 2256 13714 2316
rect 9754 2138 9814 2198
rect 14170 2138 14230 2198
rect 14328 1919 15492 2475
rect 15895 2112 17398 2649
rect 9670 1633 9887 1701
rect 16028 1769 16112 1850
rect 6372 -4604 6432 -4544
rect 7694 216 7754 276
rect 12170 216 12230 276
rect 6084 -4762 6144 -4702
rect 8222 82 8282 142
rect 12695 84 12755 144
rect 9198 -32 9258 28
rect 13632 -32 13692 28
rect 9732 -150 9792 -90
rect 14148 -150 14208 -90
rect 7192 -514 9157 -280
rect 14328 -322 15492 234
rect 15873 -176 17376 361
rect 9672 -627 9887 -557
rect 16012 -493 16096 -412
rect 2768 -5072 2828 -5012
rect 6806 -5058 6866 -4998
rect 7679 -2042 7739 -1982
rect 12154 -2044 12214 -1984
rect 8206 -2180 8266 -2120
rect 12679 -2178 12739 -2118
rect 9182 -2294 9242 -2234
rect 13616 -2294 13676 -2234
rect 9716 -2412 9776 -2352
rect 14132 -2412 14192 -2352
rect 7153 -2779 9130 -2569
rect 14328 -2622 15492 -2066
rect 15857 -2438 17360 -1901
rect 16020 -2783 16104 -2702
rect 9671 -2922 9887 -2854
rect 7687 -4350 7747 -4290
rect 12162 -4350 12222 -4290
rect 4502 -5194 4562 -5134
rect 8214 -4470 8274 -4410
rect 12687 -4468 12747 -4408
rect 9190 -4584 9250 -4524
rect 13624 -4584 13684 -4524
rect 9724 -4702 9784 -4642
rect 14140 -4702 14200 -4642
rect 15865 -4728 17368 -4191
rect 738 -5316 798 -5256
rect 738 -5780 798 -5720
rect 4500 -5778 4560 -5718
rect 7587 -6327 9188 -5951
rect 2768 -6572 2828 -6512
rect 6534 -6574 6594 -6514
<< metal3 >>
rect -1344 6036 -1124 6041
rect -1344 5964 -1334 6036
rect -1134 6032 -1124 6036
rect -1134 6026 1570 6032
rect -1134 5968 1494 6026
rect 1560 5968 1570 6026
rect -1134 5964 1570 5968
rect -1344 5959 -1124 5964
rect 1484 5963 1570 5964
rect 2802 5888 2882 5893
rect 2802 5828 2812 5888
rect 2872 5828 3062 5888
rect 2802 5823 2882 5828
rect 222 4708 302 4713
rect -548 4702 -324 4707
rect 222 4702 232 4708
rect -548 4640 -538 4702
rect -334 4648 232 4702
rect 292 4648 302 4708
rect -334 4642 302 4648
rect 2740 4676 2820 4681
rect -334 4640 -324 4642
rect -548 4635 -324 4640
rect 2740 4616 2750 4676
rect 2810 4616 2820 4676
rect 2740 4611 2820 4616
rect -942 4568 -726 4569
rect 2740 4568 2810 4611
rect -942 4564 2810 4568
rect -942 4508 -932 4564
rect -736 4508 2810 4564
rect -942 4503 -726 4508
rect 2802 4410 2882 4415
rect 2802 4350 2812 4410
rect 2872 4350 2882 4410
rect 2802 4345 2882 4350
rect 2812 3991 2872 4345
rect 3002 4121 3062 5828
rect 9638 5836 9916 5841
rect 6100 5752 6180 5757
rect 5934 5692 6110 5752
rect 6170 5692 6180 5752
rect 2992 4116 3072 4121
rect 2992 4056 3002 4116
rect 3062 4056 3072 4116
rect 2992 4051 3072 4056
rect 3002 4038 3062 4051
rect 5934 4007 5994 5692
rect 6100 5687 6180 5692
rect 9638 5600 9648 5836
rect 9906 5600 9916 5836
rect 9638 5595 9916 5600
rect 10229 5834 10509 5839
rect 10229 5602 10239 5834
rect 10499 5602 10509 5834
rect 10229 5597 10509 5602
rect 10791 5832 11074 5842
rect 10791 5596 10800 5832
rect 11058 5596 11074 5832
rect 10791 5587 11074 5596
rect 11574 4878 13540 4883
rect 6096 4554 6178 4559
rect 6096 4479 6106 4554
rect 6168 4479 6178 4554
rect 6096 4474 6178 4479
rect 5924 4002 6004 4007
rect 2794 3986 2886 3991
rect 2794 3914 2804 3986
rect 2876 3914 2886 3986
rect 5924 3942 5934 4002
rect 5994 3942 6004 4002
rect 5924 3937 6004 3942
rect 2794 3909 2886 3914
rect 5776 3850 5868 3855
rect 5776 3846 5786 3850
rect 5760 3786 5786 3846
rect 5776 3778 5786 3786
rect 5858 3846 5868 3850
rect 6106 3846 6166 4474
rect 11574 4232 11584 4878
rect 13530 4232 13540 4878
rect 11574 4227 13540 4232
rect 16040 4138 16144 4147
rect 10821 4058 10831 4138
rect 11044 4058 16050 4138
rect 16040 4057 16050 4058
rect 16134 4057 16144 4138
rect 16040 4052 16144 4057
rect 16050 4048 16144 4052
rect 9661 3991 9898 3996
rect 9661 3923 9671 3991
rect 9888 3923 9898 3991
rect 10243 3931 10253 4022
rect 10478 3931 10488 4022
rect 9661 3918 9898 3923
rect 5858 3786 6166 3846
rect 6436 3846 6973 3851
rect 5858 3778 5868 3786
rect 5776 3773 5868 3778
rect -1344 3290 -1124 3293
rect 1088 3290 1168 3295
rect -1344 3288 1098 3290
rect -1344 3230 -1334 3288
rect -1134 3230 1098 3288
rect 1158 3230 1168 3290
rect -1344 3225 -1124 3230
rect 1088 3225 1168 3230
rect 2388 3290 2468 3295
rect 2388 3230 2398 3290
rect 2458 3230 2468 3290
rect 2388 3225 2468 3230
rect 5102 3294 5182 3299
rect 6240 3294 6320 3297
rect 5102 3234 5112 3294
rect 5172 3292 6320 3294
rect 5172 3234 6250 3292
rect 5102 3229 5182 3234
rect 6240 3232 6250 3234
rect 6310 3232 6320 3292
rect 6240 3227 6320 3232
rect -2664 2818 -2442 2823
rect -2664 2738 -2654 2818
rect -2452 2808 -2442 2818
rect -130 2810 -50 2815
rect -130 2808 -120 2810
rect -2452 2750 -120 2808
rect -60 2750 -50 2810
rect -2452 2748 -50 2750
rect -2452 2738 -2442 2748
rect -130 2745 -50 2748
rect -2664 2733 -2442 2738
rect -950 2460 -724 2463
rect 254 2460 334 2465
rect -950 2458 264 2460
rect -950 2400 -940 2458
rect -734 2400 264 2458
rect 324 2400 334 2460
rect -950 2395 -724 2400
rect 254 2395 334 2400
rect 2408 2300 2468 3225
rect 6436 2617 6446 3846
rect 6963 2617 6973 3846
rect 6436 2612 6973 2617
rect 7717 2563 7777 2671
rect 7707 2558 7787 2563
rect 7707 2498 7717 2558
rect 7777 2498 7787 2558
rect 7707 2493 7787 2498
rect 6512 2432 6596 2437
rect 8246 2435 8306 2722
rect 6512 2368 6522 2432
rect 6586 2430 7650 2432
rect 8234 2430 8314 2435
rect 6586 2370 8244 2430
rect 8304 2370 8314 2430
rect 6586 2368 7650 2370
rect 6512 2363 6596 2368
rect 8234 2365 8314 2370
rect 9223 2321 9283 2602
rect 9210 2316 9290 2321
rect 9210 2300 9220 2316
rect 2408 2256 9220 2300
rect 9280 2256 9290 2316
rect 2408 2251 9290 2256
rect 2408 2240 9286 2251
rect 9756 2203 9816 2608
rect 12182 2558 12262 2563
rect 12182 2498 12192 2558
rect 12252 2498 12262 2558
rect 12182 2493 12262 2498
rect 12717 2437 12777 2580
rect 12707 2432 12787 2437
rect 12707 2372 12717 2432
rect 12777 2372 12787 2432
rect 12707 2367 12787 2372
rect 13657 2321 13717 2638
rect 13644 2316 13724 2321
rect 13644 2256 13654 2316
rect 13714 2256 13724 2316
rect 13644 2251 13724 2256
rect 14172 2203 14232 2802
rect 15885 2649 17408 2654
rect 14318 2475 15502 2480
rect 9744 2198 9824 2203
rect 5614 2136 5694 2141
rect 5614 2134 5624 2136
rect 5596 2076 5624 2134
rect 5684 2134 5694 2136
rect 9744 2138 9754 2198
rect 9814 2138 9824 2198
rect 9744 2134 9824 2138
rect 5684 2133 9824 2134
rect 14160 2198 14240 2203
rect 14160 2138 14170 2198
rect 14230 2138 14240 2198
rect 14160 2133 14240 2138
rect 5684 2076 9814 2133
rect 5596 2074 9814 2076
rect 5614 2071 5694 2074
rect -2260 1956 -2042 1961
rect 2512 1956 2592 1961
rect -2260 1896 -2250 1956
rect -2052 1896 2522 1956
rect 2582 1896 2592 1956
rect 14318 1919 14328 2475
rect 15492 1919 15502 2475
rect 15885 2112 15895 2649
rect 17398 2112 17408 2649
rect 15885 2107 17408 2112
rect 14318 1914 15502 1919
rect -2260 1891 -2042 1896
rect 2512 1891 2592 1896
rect 16018 1850 16122 1859
rect 10843 1849 16028 1850
rect 10824 1769 10834 1849
rect 11043 1770 16028 1849
rect 11043 1769 11053 1770
rect 16018 1769 16028 1770
rect 16112 1769 16122 1850
rect 16018 1764 16122 1769
rect 16028 1760 16122 1764
rect 9660 1701 9897 1706
rect 2394 1699 2576 1700
rect 2388 1694 2576 1699
rect 2388 1634 2398 1694
rect 2458 1634 2576 1694
rect 2388 1629 2576 1634
rect 5104 1694 5184 1699
rect 6362 1694 6442 1699
rect 5104 1634 5114 1694
rect 5174 1634 6372 1694
rect 6432 1634 6442 1694
rect 5104 1629 5184 1634
rect 6362 1629 6442 1634
rect 9660 1633 9670 1701
rect 9887 1633 9897 1701
rect 10237 1641 10247 1705
rect 10483 1641 10493 1705
rect 2456 1628 2576 1629
rect 9660 1628 9897 1633
rect -546 710 -326 715
rect -546 648 -536 710
rect -336 708 -326 710
rect 2348 708 2428 713
rect -336 648 2358 708
rect 2418 648 2428 708
rect -546 643 -326 648
rect 2348 643 2428 648
rect 2516 328 2576 1628
rect 2516 268 5292 328
rect 7695 281 7755 428
rect 2516 264 2576 268
rect 5230 244 5292 268
rect 7684 276 7764 281
rect 5230 14 5294 244
rect 7684 216 7694 276
rect 7754 216 7764 276
rect 7684 211 7764 216
rect 8224 148 8284 424
rect 6668 147 8284 148
rect 6664 142 8292 147
rect 6664 82 6674 142
rect 6734 82 8222 142
rect 8282 82 8292 142
rect 6664 77 8292 82
rect 6668 76 8234 77
rect 9201 33 9261 298
rect 9188 28 9268 33
rect 9188 14 9198 28
rect -2662 -20 -2446 -15
rect -186 -18 22 -13
rect -186 -20 -176 -18
rect -2662 -216 -2652 -20
rect -2456 -216 -176 -20
rect 12 -216 22 -18
rect 5230 -32 9198 14
rect 9258 -32 9268 28
rect 5230 -46 9268 -32
rect 5230 -48 5294 -46
rect 9734 -85 9794 296
rect 12160 276 12240 281
rect 12160 216 12170 276
rect 12230 216 12240 276
rect 12160 211 12240 216
rect 12695 149 12755 294
rect 12685 144 12765 149
rect 12685 84 12695 144
rect 12755 84 12765 144
rect 12685 79 12765 84
rect 13635 33 13695 366
rect 13622 28 13702 33
rect 13622 -32 13632 28
rect 13692 -32 13702 28
rect 13622 -37 13702 -32
rect 14150 -85 14210 510
rect 15863 361 17386 366
rect 14318 234 15502 239
rect 9722 -90 9802 -85
rect 5784 -154 5864 -149
rect 9722 -150 9732 -90
rect 9792 -150 9802 -90
rect 9722 -154 9802 -150
rect 5776 -214 5794 -154
rect 5854 -155 9802 -154
rect 14138 -90 14218 -85
rect 14138 -150 14148 -90
rect 14208 -150 14218 -90
rect 14138 -155 14218 -150
rect 5854 -214 9792 -155
rect -2662 -221 -2446 -216
rect -372 -218 22 -216
rect -186 -221 22 -218
rect 5784 -219 5864 -214
rect 7182 -280 9167 -275
rect 7182 -514 7192 -280
rect 9157 -514 9167 -280
rect 14318 -322 14328 234
rect 15492 -322 15502 234
rect 15863 -176 15873 361
rect 17376 -176 17386 361
rect 15863 -181 17386 -176
rect 14318 -327 15502 -322
rect 16002 -412 16106 -403
rect 10842 -413 16012 -412
rect 10832 -492 10842 -413
rect 11044 -492 16012 -413
rect 16002 -493 16012 -492
rect 16096 -493 16106 -412
rect 16002 -498 16106 -493
rect 16012 -502 16106 -498
rect 7182 -519 9167 -514
rect 9662 -557 9897 -552
rect 9662 -627 9672 -557
rect 9887 -627 9897 -557
rect 10237 -621 10247 -557
rect 10483 -621 10493 -557
rect 9662 -632 9897 -627
rect -947 -730 -724 -725
rect 96 -730 184 -725
rect -947 -792 -937 -730
rect -734 -792 106 -730
rect 174 -792 184 -730
rect -947 -797 -724 -792
rect 96 -797 184 -792
rect 3032 -762 3112 -761
rect 3032 -766 6602 -762
rect 3032 -826 3042 -766
rect 3102 -767 6602 -766
rect 3102 -826 6518 -767
rect 3032 -831 6518 -826
rect 3038 -832 6518 -831
rect 6583 -832 6602 -767
rect 3038 -834 6602 -832
rect 6508 -837 6593 -834
rect -1344 -1134 -1124 -1129
rect 48 -1134 128 -1129
rect -1344 -1194 -1334 -1134
rect -1134 -1194 58 -1134
rect 118 -1194 128 -1134
rect -1344 -1199 -1124 -1194
rect 48 -1199 128 -1194
rect 6660 -1490 6752 -1485
rect 3040 -1491 6670 -1490
rect 3036 -1496 6670 -1491
rect 3036 -1556 3046 -1496
rect 3106 -1556 6670 -1496
rect 3036 -1561 6670 -1556
rect 3040 -1562 6670 -1561
rect 6742 -1562 6752 -1490
rect 6660 -1567 6752 -1562
rect 7679 -1977 7739 -1842
rect 7669 -1982 7749 -1977
rect 7669 -2042 7679 -1982
rect 7739 -2042 7749 -1982
rect 7669 -2047 7749 -2042
rect 8208 -2114 8268 -1836
rect 3032 -2115 8268 -2114
rect 3032 -2120 8276 -2115
rect 3032 -2180 8206 -2120
rect 8266 -2180 8276 -2120
rect 3032 -2185 8276 -2180
rect 3032 -2186 8210 -2185
rect 3032 -3101 3104 -2186
rect 9185 -2229 9245 -1956
rect 12144 -1984 12224 -1979
rect 9172 -2234 9252 -2229
rect 9172 -2248 9182 -2234
rect 6222 -2256 9182 -2248
rect 6222 -2308 6246 -2256
rect 6236 -2318 6246 -2308
rect 6308 -2294 9182 -2256
rect 9242 -2294 9252 -2234
rect 6308 -2308 9252 -2294
rect 6308 -2318 6318 -2308
rect 6236 -2323 6318 -2318
rect 9718 -2347 9778 -1994
rect 12144 -2044 12154 -1984
rect 12214 -2044 12224 -1984
rect 12144 -2049 12224 -2044
rect 12679 -2113 12739 -1982
rect 12669 -2118 12749 -2113
rect 12669 -2178 12679 -2118
rect 12739 -2178 12749 -2118
rect 12669 -2183 12749 -2178
rect 13619 -2229 13679 -1906
rect 13606 -2234 13686 -2229
rect 13606 -2294 13616 -2234
rect 13676 -2294 13686 -2234
rect 13606 -2299 13686 -2294
rect 14134 -2347 14194 -1722
rect 15847 -1901 17370 -1896
rect 14318 -2066 15502 -2061
rect 9706 -2352 9786 -2347
rect 5938 -2416 6020 -2411
rect 9706 -2412 9716 -2352
rect 9776 -2412 9786 -2352
rect 9706 -2416 9786 -2412
rect 5905 -2478 5948 -2416
rect 6010 -2417 9786 -2416
rect 14122 -2352 14202 -2347
rect 14122 -2412 14132 -2352
rect 14192 -2412 14202 -2352
rect 14122 -2417 14202 -2412
rect 6010 -2478 9776 -2417
rect 5938 -2483 6020 -2478
rect 7143 -2569 9140 -2564
rect 7137 -2863 7147 -2569
rect 9130 -2863 9140 -2569
rect 14318 -2622 14328 -2066
rect 15492 -2622 15502 -2066
rect 15847 -2438 15857 -1901
rect 17360 -2438 17370 -1901
rect 15847 -2443 17370 -2438
rect 14318 -2627 15502 -2622
rect 16010 -2702 16114 -2697
rect 10816 -2782 10822 -2702
rect 11056 -2782 16020 -2702
rect 16010 -2783 16020 -2782
rect 16104 -2783 16114 -2702
rect 16010 -2788 16114 -2783
rect 9661 -2854 9897 -2849
rect 9661 -2922 9671 -2854
rect 9887 -2922 9897 -2854
rect 9661 -2927 9897 -2922
rect 10129 -2851 10215 -2848
rect 10129 -2917 10251 -2851
rect 10477 -2917 10487 -2851
rect 3028 -3106 3120 -3101
rect 3028 -3178 3038 -3106
rect 3110 -3178 3120 -3106
rect 10129 -3149 10215 -2917
rect 3028 -3183 3120 -3178
rect -1344 -3480 -1124 -3475
rect 50 -3480 130 -3475
rect -1344 -3540 -1334 -3480
rect -1134 -3540 60 -3480
rect 120 -3540 130 -3480
rect -1344 -3545 -1124 -3540
rect 50 -3545 130 -3540
rect 3034 -3844 3114 -3839
rect 3034 -3904 3044 -3844
rect 3104 -3904 3114 -3844
rect 3034 -3909 3114 -3904
rect 3044 -4416 3108 -3909
rect 7687 -4284 7747 -4161
rect 7676 -4285 7747 -4284
rect 7676 -4290 7757 -4285
rect 7676 -4350 7687 -4290
rect 7747 -4350 7757 -4290
rect 7676 -4354 7757 -4350
rect 7677 -4355 7757 -4354
rect 8216 -4405 8276 -4171
rect 8204 -4410 8284 -4405
rect 8204 -4414 8214 -4410
rect 8134 -4416 8214 -4414
rect 3044 -4470 8214 -4416
rect 8274 -4470 8284 -4410
rect 3044 -4475 8284 -4470
rect 3044 -4476 8205 -4475
rect 3044 -4478 3108 -4476
rect 9193 -4519 9253 -4254
rect 9180 -4524 9260 -4519
rect 9180 -4536 9190 -4524
rect -2257 -4544 -2038 -4539
rect -2257 -4712 -2247 -4544
rect -2048 -4546 -2038 -4544
rect 3722 -4546 3908 -4541
rect -2048 -4712 3732 -4546
rect 3898 -4712 3908 -4546
rect 6362 -4544 9190 -4536
rect 6362 -4604 6372 -4544
rect 6432 -4584 9190 -4544
rect 9250 -4584 9260 -4524
rect 6432 -4596 9260 -4584
rect 6432 -4604 6442 -4596
rect 6362 -4609 6442 -4604
rect 9726 -4637 9786 -4254
rect 12152 -4290 12232 -4285
rect 12152 -4350 12162 -4290
rect 12222 -4350 12232 -4290
rect 12152 -4355 12232 -4350
rect 12687 -4403 12747 -4272
rect 12677 -4408 12757 -4403
rect 12677 -4468 12687 -4408
rect 12747 -4468 12757 -4408
rect 12677 -4473 12757 -4468
rect 13627 -4519 13687 -4132
rect 13614 -4524 13694 -4519
rect 13614 -4584 13624 -4524
rect 13684 -4584 13694 -4524
rect 13614 -4589 13694 -4584
rect 14142 -4637 14202 -4009
rect 15855 -4191 17378 -4186
rect 9714 -4642 9794 -4637
rect -2257 -4717 -2038 -4712
rect 3722 -4717 3908 -4712
rect 6074 -4702 6154 -4697
rect 9714 -4702 9724 -4642
rect 9784 -4702 9794 -4642
rect 6074 -4762 6084 -4702
rect 6144 -4707 9794 -4702
rect 14130 -4642 14210 -4637
rect 14130 -4702 14140 -4642
rect 14200 -4702 14210 -4642
rect 14130 -4707 14210 -4702
rect 6144 -4762 9784 -4707
rect 15855 -4728 15865 -4191
rect 17368 -4728 17378 -4191
rect 15855 -4733 17378 -4728
rect 6074 -4767 6154 -4762
rect 6796 -4998 6876 -4993
rect 2758 -5012 2838 -5007
rect 2758 -5072 2768 -5012
rect 2828 -5072 2838 -5012
rect 6796 -5058 6806 -4998
rect 6866 -5058 6876 -4998
rect 6796 -5063 6876 -5058
rect 2758 -5077 2838 -5072
rect 728 -5256 808 -5251
rect 728 -5316 738 -5256
rect 798 -5316 808 -5256
rect 728 -5321 808 -5316
rect 738 -5715 798 -5321
rect 728 -5720 808 -5715
rect 728 -5780 738 -5720
rect 798 -5780 808 -5720
rect 728 -5785 808 -5780
rect 2766 -6507 2831 -5077
rect 4502 -5129 4562 -5118
rect 4492 -5134 4572 -5129
rect 4492 -5194 4502 -5134
rect 4562 -5194 4572 -5134
rect 4492 -5199 4572 -5194
rect 4502 -5713 4562 -5199
rect 4490 -5718 4570 -5713
rect 4490 -5778 4500 -5718
rect 4560 -5778 4570 -5718
rect 4490 -5783 4570 -5778
rect 2758 -6512 2838 -6507
rect 2758 -6572 2768 -6512
rect 2828 -6572 2838 -6512
rect 2758 -6577 2838 -6572
rect 6524 -6510 6604 -6509
rect 6802 -6510 6870 -5063
rect 7577 -5951 9198 -5946
rect 7577 -6327 7587 -5951
rect 9188 -6327 9198 -5951
rect 7577 -6332 9198 -6327
rect 6524 -6514 6870 -6510
rect 6524 -6574 6534 -6514
rect 6594 -6574 6870 -6514
rect 2766 -6578 2831 -6577
rect 6524 -6578 6870 -6574
rect 6524 -6579 6604 -6578
<< via3 >>
rect 9648 5600 9906 5836
rect 10239 5602 10499 5834
rect 10800 5596 11058 5832
rect 11584 4232 13530 4878
rect 10831 4058 11044 4138
rect 9671 3923 9888 3991
rect 10253 3931 10478 4022
rect 6446 2617 6963 3846
rect 14328 1919 15492 2475
rect 15895 2112 17398 2649
rect 10834 1769 11043 1849
rect 9670 1633 9887 1701
rect 10247 1641 10483 1705
rect 7192 -514 9157 -280
rect 14328 -322 15492 234
rect 15873 -176 17376 361
rect 10842 -492 11044 -413
rect 9672 -627 9887 -557
rect 10247 -621 10483 -557
rect 7147 -2779 7153 -2569
rect 7153 -2779 9130 -2569
rect 7147 -2863 9130 -2779
rect 14328 -2622 15492 -2066
rect 15857 -2438 17360 -1901
rect 10822 -2782 11056 -2702
rect 9671 -2922 9887 -2854
rect 10251 -2917 10477 -2851
rect 15865 -4728 17368 -4191
rect 7587 -6327 9188 -5951
<< metal4 >>
rect 9647 5836 9907 5837
rect 9647 5600 9648 5836
rect 9906 5600 9907 5836
rect 10238 5834 10500 5835
rect 10238 5606 10239 5834
rect 9647 5599 9907 5600
rect 10237 5602 10239 5606
rect 10499 5602 10500 5834
rect 10237 5601 10500 5602
rect 10791 5832 11074 5842
rect 9650 5378 9906 5599
rect 6445 3846 6964 3847
rect 6445 2617 6446 3846
rect 6963 3843 6964 3846
rect 7412 3843 9332 4652
rect 6963 2617 9332 3843
rect 6445 2616 6964 2617
rect 7412 -279 9332 2617
rect 7191 -280 9332 -279
rect 7191 -514 7192 -280
rect 9157 -514 9332 -280
rect 7191 -515 9332 -514
rect 7412 -2568 9332 -515
rect 7146 -2569 9332 -2568
rect 7146 -2863 7147 -2569
rect 9130 -2863 9332 -2569
rect 7146 -2864 9332 -2863
rect 7412 -5951 9332 -2864
rect 9669 3991 9891 5378
rect 10237 5366 10497 5601
rect 10791 5596 10800 5832
rect 11058 5596 11074 5832
rect 10791 5587 11074 5596
rect 9669 3923 9671 3991
rect 9888 3923 9891 3991
rect 9669 1701 9891 3923
rect 10247 4022 10483 5366
rect 10800 5362 11070 5587
rect 10247 3931 10253 4022
rect 10478 3931 10483 4022
rect 10247 1706 10483 3931
rect 10821 4138 11055 5362
rect 11583 4878 13531 4879
rect 11583 4596 11584 4878
rect 10821 4058 10831 4138
rect 11044 4058 11055 4138
rect 10821 1849 11055 4058
rect 10821 1769 10834 1849
rect 11043 1769 11055 1849
rect 9669 1633 9670 1701
rect 9887 1633 9891 1701
rect 10246 1705 10484 1706
rect 10246 1641 10247 1705
rect 10483 1641 10484 1705
rect 10246 1640 10484 1641
rect 9669 -557 9891 1633
rect 10247 -556 10483 1640
rect 10821 -413 11055 1769
rect 10821 -492 10842 -413
rect 11044 -492 11055 -413
rect 9669 -627 9672 -557
rect 9887 -627 9891 -557
rect 10246 -557 10484 -556
rect 10246 -621 10247 -557
rect 10483 -621 10484 -557
rect 10246 -622 10484 -621
rect 9669 -2854 9891 -627
rect 9669 -2922 9671 -2854
rect 9887 -2922 9891 -2854
rect 10247 -2851 10483 -622
rect 10821 -2701 11055 -492
rect 11560 4232 11584 4596
rect 13530 4596 13531 4878
rect 13530 4232 13560 4596
rect 11560 2469 13560 4232
rect 15714 2649 17672 4883
rect 14327 2475 15493 2476
rect 14327 2469 14328 2475
rect 11560 1921 14328 2469
rect 11560 228 13560 1921
rect 14327 1919 14328 1921
rect 15492 1919 15493 2475
rect 14327 1918 15493 1919
rect 15714 2112 15895 2649
rect 17398 2112 17672 2649
rect 15714 1872 17672 2112
rect 15714 361 17650 1872
rect 14327 234 15493 235
rect 14327 228 14328 234
rect 11560 -320 14328 228
rect 11560 -2072 13560 -320
rect 14327 -322 14328 -320
rect 15492 -322 15493 234
rect 14327 -323 15493 -322
rect 15714 -176 15873 361
rect 17376 -176 17650 361
rect 15714 -416 17650 -176
rect 15714 -1901 17642 -416
rect 14327 -2066 15493 -2065
rect 14327 -2072 14328 -2066
rect 11560 -2620 14328 -2072
rect 10821 -2702 11057 -2701
rect 10821 -2782 10822 -2702
rect 11056 -2782 11057 -2702
rect 10821 -2784 11057 -2782
rect 10247 -2917 10251 -2851
rect 10477 -2917 10483 -2851
rect 10247 -2920 10483 -2917
rect 9669 -2950 9891 -2922
rect 11560 -5140 13560 -2620
rect 14327 -2622 14328 -2620
rect 15492 -2622 15493 -2066
rect 14327 -2623 15493 -2622
rect 15714 -2438 15857 -1901
rect 17360 -2438 17642 -1901
rect 15714 -2678 17642 -2438
rect 15722 -4191 17642 -2678
rect 15722 -4728 15865 -4191
rect 17368 -4728 17642 -4191
rect 15722 -4968 17642 -4728
rect 7412 -6327 7587 -5951
rect 9188 -6327 9332 -5951
rect 7412 -7058 9332 -6327
use c4b  c4b_0
timestamp 1624338677
transform 1 0 -56 0 1 -2384
box -120 -2346 3972 2370
use contador4bits  contador4bits_0
timestamp 1624338677
transform 1 0 -64 0 1 4130
box -56 0 6948 1980
use 4bitc  4bitc_0
timestamp 1624338677
transform 1 0 -63 0 1 1939
box -107 -1605 5377 1735
use mux_8to1  mux_8to1_3
timestamp 1624381803
transform 1 0 7162 0 1 -5404
box -54 1072 10324 2553
use mux_8to1  mux_8to1_1
timestamp 1624381803
transform 1 0 7170 0 1 -852
box -54 1072 10324 2553
use mux_8to1  mux_8to1_0
timestamp 1624381803
transform 1 0 7192 0 1 1436
box -54 1072 10324 2553
use mux_8to1  mux_8to1_2
timestamp 1624381803
transform 1 0 7154 0 1 -3114
box -54 1072 10324 2553
use contador  contador_0
timestamp 1624388555
transform 1 0 -206 0 1 -6968
box 0 0 7741 1645
<< labels >>
rlabel metal2 -1826 -2132 -1566 -1894 1 VSS
rlabel metal2 -1832 -2890 -1572 -2652 1 CE
rlabel metal2 -1832 -2496 -1572 -2258 1 CLK
rlabel metal2 -1836 -1764 -1576 -1526 1 VDD
rlabel metal2 -1832 -3314 -1572 -3076 1 CLR
rlabel metal2 17488 768 17748 1006 1 Q1
rlabel metal2 17472 -1596 17732 -1358 1 Q2
rlabel metal2 17480 -3784 17740 -3546 1 Q3
rlabel metal2 17510 3056 17770 3294 1 Q0
rlabel metal4 10800 5594 11060 5832 1 reg0
rlabel metal2 10239 5598 10499 5836 1 reg1
rlabel metal2 9650 5598 9910 5836 1 reg2
<< end >>
