magic
tech sky130A
magscale 1 2
timestamp 1615997521
<< nwell >>
rect -6867 -919 6867 919
<< pmoslvt >>
rect -6671 -700 -6461 700
rect -6403 -700 -6193 700
rect -6135 -700 -5925 700
rect -5867 -700 -5657 700
rect -5599 -700 -5389 700
rect -5331 -700 -5121 700
rect -5063 -700 -4853 700
rect -4795 -700 -4585 700
rect -4527 -700 -4317 700
rect -4259 -700 -4049 700
rect -3991 -700 -3781 700
rect -3723 -700 -3513 700
rect -3455 -700 -3245 700
rect -3187 -700 -2977 700
rect -2919 -700 -2709 700
rect -2651 -700 -2441 700
rect -2383 -700 -2173 700
rect -2115 -700 -1905 700
rect -1847 -700 -1637 700
rect -1579 -700 -1369 700
rect -1311 -700 -1101 700
rect -1043 -700 -833 700
rect -775 -700 -565 700
rect -507 -700 -297 700
rect -239 -700 -29 700
rect 29 -700 239 700
rect 297 -700 507 700
rect 565 -700 775 700
rect 833 -700 1043 700
rect 1101 -700 1311 700
rect 1369 -700 1579 700
rect 1637 -700 1847 700
rect 1905 -700 2115 700
rect 2173 -700 2383 700
rect 2441 -700 2651 700
rect 2709 -700 2919 700
rect 2977 -700 3187 700
rect 3245 -700 3455 700
rect 3513 -700 3723 700
rect 3781 -700 3991 700
rect 4049 -700 4259 700
rect 4317 -700 4527 700
rect 4585 -700 4795 700
rect 4853 -700 5063 700
rect 5121 -700 5331 700
rect 5389 -700 5599 700
rect 5657 -700 5867 700
rect 5925 -700 6135 700
rect 6193 -700 6403 700
rect 6461 -700 6671 700
<< pdiff >>
rect -6729 688 -6671 700
rect -6729 -688 -6717 688
rect -6683 -688 -6671 688
rect -6729 -700 -6671 -688
rect -6461 688 -6403 700
rect -6461 -688 -6449 688
rect -6415 -688 -6403 688
rect -6461 -700 -6403 -688
rect -6193 688 -6135 700
rect -6193 -688 -6181 688
rect -6147 -688 -6135 688
rect -6193 -700 -6135 -688
rect -5925 688 -5867 700
rect -5925 -688 -5913 688
rect -5879 -688 -5867 688
rect -5925 -700 -5867 -688
rect -5657 688 -5599 700
rect -5657 -688 -5645 688
rect -5611 -688 -5599 688
rect -5657 -700 -5599 -688
rect -5389 688 -5331 700
rect -5389 -688 -5377 688
rect -5343 -688 -5331 688
rect -5389 -700 -5331 -688
rect -5121 688 -5063 700
rect -5121 -688 -5109 688
rect -5075 -688 -5063 688
rect -5121 -700 -5063 -688
rect -4853 688 -4795 700
rect -4853 -688 -4841 688
rect -4807 -688 -4795 688
rect -4853 -700 -4795 -688
rect -4585 688 -4527 700
rect -4585 -688 -4573 688
rect -4539 -688 -4527 688
rect -4585 -700 -4527 -688
rect -4317 688 -4259 700
rect -4317 -688 -4305 688
rect -4271 -688 -4259 688
rect -4317 -700 -4259 -688
rect -4049 688 -3991 700
rect -4049 -688 -4037 688
rect -4003 -688 -3991 688
rect -4049 -700 -3991 -688
rect -3781 688 -3723 700
rect -3781 -688 -3769 688
rect -3735 -688 -3723 688
rect -3781 -700 -3723 -688
rect -3513 688 -3455 700
rect -3513 -688 -3501 688
rect -3467 -688 -3455 688
rect -3513 -700 -3455 -688
rect -3245 688 -3187 700
rect -3245 -688 -3233 688
rect -3199 -688 -3187 688
rect -3245 -700 -3187 -688
rect -2977 688 -2919 700
rect -2977 -688 -2965 688
rect -2931 -688 -2919 688
rect -2977 -700 -2919 -688
rect -2709 688 -2651 700
rect -2709 -688 -2697 688
rect -2663 -688 -2651 688
rect -2709 -700 -2651 -688
rect -2441 688 -2383 700
rect -2441 -688 -2429 688
rect -2395 -688 -2383 688
rect -2441 -700 -2383 -688
rect -2173 688 -2115 700
rect -2173 -688 -2161 688
rect -2127 -688 -2115 688
rect -2173 -700 -2115 -688
rect -1905 688 -1847 700
rect -1905 -688 -1893 688
rect -1859 -688 -1847 688
rect -1905 -700 -1847 -688
rect -1637 688 -1579 700
rect -1637 -688 -1625 688
rect -1591 -688 -1579 688
rect -1637 -700 -1579 -688
rect -1369 688 -1311 700
rect -1369 -688 -1357 688
rect -1323 -688 -1311 688
rect -1369 -700 -1311 -688
rect -1101 688 -1043 700
rect -1101 -688 -1089 688
rect -1055 -688 -1043 688
rect -1101 -700 -1043 -688
rect -833 688 -775 700
rect -833 -688 -821 688
rect -787 -688 -775 688
rect -833 -700 -775 -688
rect -565 688 -507 700
rect -565 -688 -553 688
rect -519 -688 -507 688
rect -565 -700 -507 -688
rect -297 688 -239 700
rect -297 -688 -285 688
rect -251 -688 -239 688
rect -297 -700 -239 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 239 688 297 700
rect 239 -688 251 688
rect 285 -688 297 688
rect 239 -700 297 -688
rect 507 688 565 700
rect 507 -688 519 688
rect 553 -688 565 688
rect 507 -700 565 -688
rect 775 688 833 700
rect 775 -688 787 688
rect 821 -688 833 688
rect 775 -700 833 -688
rect 1043 688 1101 700
rect 1043 -688 1055 688
rect 1089 -688 1101 688
rect 1043 -700 1101 -688
rect 1311 688 1369 700
rect 1311 -688 1323 688
rect 1357 -688 1369 688
rect 1311 -700 1369 -688
rect 1579 688 1637 700
rect 1579 -688 1591 688
rect 1625 -688 1637 688
rect 1579 -700 1637 -688
rect 1847 688 1905 700
rect 1847 -688 1859 688
rect 1893 -688 1905 688
rect 1847 -700 1905 -688
rect 2115 688 2173 700
rect 2115 -688 2127 688
rect 2161 -688 2173 688
rect 2115 -700 2173 -688
rect 2383 688 2441 700
rect 2383 -688 2395 688
rect 2429 -688 2441 688
rect 2383 -700 2441 -688
rect 2651 688 2709 700
rect 2651 -688 2663 688
rect 2697 -688 2709 688
rect 2651 -700 2709 -688
rect 2919 688 2977 700
rect 2919 -688 2931 688
rect 2965 -688 2977 688
rect 2919 -700 2977 -688
rect 3187 688 3245 700
rect 3187 -688 3199 688
rect 3233 -688 3245 688
rect 3187 -700 3245 -688
rect 3455 688 3513 700
rect 3455 -688 3467 688
rect 3501 -688 3513 688
rect 3455 -700 3513 -688
rect 3723 688 3781 700
rect 3723 -688 3735 688
rect 3769 -688 3781 688
rect 3723 -700 3781 -688
rect 3991 688 4049 700
rect 3991 -688 4003 688
rect 4037 -688 4049 688
rect 3991 -700 4049 -688
rect 4259 688 4317 700
rect 4259 -688 4271 688
rect 4305 -688 4317 688
rect 4259 -700 4317 -688
rect 4527 688 4585 700
rect 4527 -688 4539 688
rect 4573 -688 4585 688
rect 4527 -700 4585 -688
rect 4795 688 4853 700
rect 4795 -688 4807 688
rect 4841 -688 4853 688
rect 4795 -700 4853 -688
rect 5063 688 5121 700
rect 5063 -688 5075 688
rect 5109 -688 5121 688
rect 5063 -700 5121 -688
rect 5331 688 5389 700
rect 5331 -688 5343 688
rect 5377 -688 5389 688
rect 5331 -700 5389 -688
rect 5599 688 5657 700
rect 5599 -688 5611 688
rect 5645 -688 5657 688
rect 5599 -700 5657 -688
rect 5867 688 5925 700
rect 5867 -688 5879 688
rect 5913 -688 5925 688
rect 5867 -700 5925 -688
rect 6135 688 6193 700
rect 6135 -688 6147 688
rect 6181 -688 6193 688
rect 6135 -700 6193 -688
rect 6403 688 6461 700
rect 6403 -688 6415 688
rect 6449 -688 6461 688
rect 6403 -700 6461 -688
rect 6671 688 6729 700
rect 6671 -688 6683 688
rect 6717 -688 6729 688
rect 6671 -700 6729 -688
<< pdiffc >>
rect -6717 -688 -6683 688
rect -6449 -688 -6415 688
rect -6181 -688 -6147 688
rect -5913 -688 -5879 688
rect -5645 -688 -5611 688
rect -5377 -688 -5343 688
rect -5109 -688 -5075 688
rect -4841 -688 -4807 688
rect -4573 -688 -4539 688
rect -4305 -688 -4271 688
rect -4037 -688 -4003 688
rect -3769 -688 -3735 688
rect -3501 -688 -3467 688
rect -3233 -688 -3199 688
rect -2965 -688 -2931 688
rect -2697 -688 -2663 688
rect -2429 -688 -2395 688
rect -2161 -688 -2127 688
rect -1893 -688 -1859 688
rect -1625 -688 -1591 688
rect -1357 -688 -1323 688
rect -1089 -688 -1055 688
rect -821 -688 -787 688
rect -553 -688 -519 688
rect -285 -688 -251 688
rect -17 -688 17 688
rect 251 -688 285 688
rect 519 -688 553 688
rect 787 -688 821 688
rect 1055 -688 1089 688
rect 1323 -688 1357 688
rect 1591 -688 1625 688
rect 1859 -688 1893 688
rect 2127 -688 2161 688
rect 2395 -688 2429 688
rect 2663 -688 2697 688
rect 2931 -688 2965 688
rect 3199 -688 3233 688
rect 3467 -688 3501 688
rect 3735 -688 3769 688
rect 4003 -688 4037 688
rect 4271 -688 4305 688
rect 4539 -688 4573 688
rect 4807 -688 4841 688
rect 5075 -688 5109 688
rect 5343 -688 5377 688
rect 5611 -688 5645 688
rect 5879 -688 5913 688
rect 6147 -688 6181 688
rect 6415 -688 6449 688
rect 6683 -688 6717 688
<< nsubdiff >>
rect -6831 849 -6735 883
rect 6735 849 6831 883
rect -6831 787 -6797 849
rect 6797 787 6831 849
rect -6831 -849 -6797 -787
rect 6797 -849 6831 -787
rect -6831 -883 -6735 -849
rect 6735 -883 6831 -849
<< nsubdiffcont >>
rect -6735 849 6735 883
rect -6831 -787 -6797 787
rect 6797 -787 6831 787
rect -6735 -883 6735 -849
<< poly >>
rect -6671 781 -6461 797
rect -6671 747 -6655 781
rect -6477 747 -6461 781
rect -6671 700 -6461 747
rect -6403 781 -6193 797
rect -6403 747 -6387 781
rect -6209 747 -6193 781
rect -6403 700 -6193 747
rect -6135 781 -5925 797
rect -6135 747 -6119 781
rect -5941 747 -5925 781
rect -6135 700 -5925 747
rect -5867 781 -5657 797
rect -5867 747 -5851 781
rect -5673 747 -5657 781
rect -5867 700 -5657 747
rect -5599 781 -5389 797
rect -5599 747 -5583 781
rect -5405 747 -5389 781
rect -5599 700 -5389 747
rect -5331 781 -5121 797
rect -5331 747 -5315 781
rect -5137 747 -5121 781
rect -5331 700 -5121 747
rect -5063 781 -4853 797
rect -5063 747 -5047 781
rect -4869 747 -4853 781
rect -5063 700 -4853 747
rect -4795 781 -4585 797
rect -4795 747 -4779 781
rect -4601 747 -4585 781
rect -4795 700 -4585 747
rect -4527 781 -4317 797
rect -4527 747 -4511 781
rect -4333 747 -4317 781
rect -4527 700 -4317 747
rect -4259 781 -4049 797
rect -4259 747 -4243 781
rect -4065 747 -4049 781
rect -4259 700 -4049 747
rect -3991 781 -3781 797
rect -3991 747 -3975 781
rect -3797 747 -3781 781
rect -3991 700 -3781 747
rect -3723 781 -3513 797
rect -3723 747 -3707 781
rect -3529 747 -3513 781
rect -3723 700 -3513 747
rect -3455 781 -3245 797
rect -3455 747 -3439 781
rect -3261 747 -3245 781
rect -3455 700 -3245 747
rect -3187 781 -2977 797
rect -3187 747 -3171 781
rect -2993 747 -2977 781
rect -3187 700 -2977 747
rect -2919 781 -2709 797
rect -2919 747 -2903 781
rect -2725 747 -2709 781
rect -2919 700 -2709 747
rect -2651 781 -2441 797
rect -2651 747 -2635 781
rect -2457 747 -2441 781
rect -2651 700 -2441 747
rect -2383 781 -2173 797
rect -2383 747 -2367 781
rect -2189 747 -2173 781
rect -2383 700 -2173 747
rect -2115 781 -1905 797
rect -2115 747 -2099 781
rect -1921 747 -1905 781
rect -2115 700 -1905 747
rect -1847 781 -1637 797
rect -1847 747 -1831 781
rect -1653 747 -1637 781
rect -1847 700 -1637 747
rect -1579 781 -1369 797
rect -1579 747 -1563 781
rect -1385 747 -1369 781
rect -1579 700 -1369 747
rect -1311 781 -1101 797
rect -1311 747 -1295 781
rect -1117 747 -1101 781
rect -1311 700 -1101 747
rect -1043 781 -833 797
rect -1043 747 -1027 781
rect -849 747 -833 781
rect -1043 700 -833 747
rect -775 781 -565 797
rect -775 747 -759 781
rect -581 747 -565 781
rect -775 700 -565 747
rect -507 781 -297 797
rect -507 747 -491 781
rect -313 747 -297 781
rect -507 700 -297 747
rect -239 781 -29 797
rect -239 747 -223 781
rect -45 747 -29 781
rect -239 700 -29 747
rect 29 781 239 797
rect 29 747 45 781
rect 223 747 239 781
rect 29 700 239 747
rect 297 781 507 797
rect 297 747 313 781
rect 491 747 507 781
rect 297 700 507 747
rect 565 781 775 797
rect 565 747 581 781
rect 759 747 775 781
rect 565 700 775 747
rect 833 781 1043 797
rect 833 747 849 781
rect 1027 747 1043 781
rect 833 700 1043 747
rect 1101 781 1311 797
rect 1101 747 1117 781
rect 1295 747 1311 781
rect 1101 700 1311 747
rect 1369 781 1579 797
rect 1369 747 1385 781
rect 1563 747 1579 781
rect 1369 700 1579 747
rect 1637 781 1847 797
rect 1637 747 1653 781
rect 1831 747 1847 781
rect 1637 700 1847 747
rect 1905 781 2115 797
rect 1905 747 1921 781
rect 2099 747 2115 781
rect 1905 700 2115 747
rect 2173 781 2383 797
rect 2173 747 2189 781
rect 2367 747 2383 781
rect 2173 700 2383 747
rect 2441 781 2651 797
rect 2441 747 2457 781
rect 2635 747 2651 781
rect 2441 700 2651 747
rect 2709 781 2919 797
rect 2709 747 2725 781
rect 2903 747 2919 781
rect 2709 700 2919 747
rect 2977 781 3187 797
rect 2977 747 2993 781
rect 3171 747 3187 781
rect 2977 700 3187 747
rect 3245 781 3455 797
rect 3245 747 3261 781
rect 3439 747 3455 781
rect 3245 700 3455 747
rect 3513 781 3723 797
rect 3513 747 3529 781
rect 3707 747 3723 781
rect 3513 700 3723 747
rect 3781 781 3991 797
rect 3781 747 3797 781
rect 3975 747 3991 781
rect 3781 700 3991 747
rect 4049 781 4259 797
rect 4049 747 4065 781
rect 4243 747 4259 781
rect 4049 700 4259 747
rect 4317 781 4527 797
rect 4317 747 4333 781
rect 4511 747 4527 781
rect 4317 700 4527 747
rect 4585 781 4795 797
rect 4585 747 4601 781
rect 4779 747 4795 781
rect 4585 700 4795 747
rect 4853 781 5063 797
rect 4853 747 4869 781
rect 5047 747 5063 781
rect 4853 700 5063 747
rect 5121 781 5331 797
rect 5121 747 5137 781
rect 5315 747 5331 781
rect 5121 700 5331 747
rect 5389 781 5599 797
rect 5389 747 5405 781
rect 5583 747 5599 781
rect 5389 700 5599 747
rect 5657 781 5867 797
rect 5657 747 5673 781
rect 5851 747 5867 781
rect 5657 700 5867 747
rect 5925 781 6135 797
rect 5925 747 5941 781
rect 6119 747 6135 781
rect 5925 700 6135 747
rect 6193 781 6403 797
rect 6193 747 6209 781
rect 6387 747 6403 781
rect 6193 700 6403 747
rect 6461 781 6671 797
rect 6461 747 6477 781
rect 6655 747 6671 781
rect 6461 700 6671 747
rect -6671 -747 -6461 -700
rect -6671 -781 -6655 -747
rect -6477 -781 -6461 -747
rect -6671 -797 -6461 -781
rect -6403 -747 -6193 -700
rect -6403 -781 -6387 -747
rect -6209 -781 -6193 -747
rect -6403 -797 -6193 -781
rect -6135 -747 -5925 -700
rect -6135 -781 -6119 -747
rect -5941 -781 -5925 -747
rect -6135 -797 -5925 -781
rect -5867 -747 -5657 -700
rect -5867 -781 -5851 -747
rect -5673 -781 -5657 -747
rect -5867 -797 -5657 -781
rect -5599 -747 -5389 -700
rect -5599 -781 -5583 -747
rect -5405 -781 -5389 -747
rect -5599 -797 -5389 -781
rect -5331 -747 -5121 -700
rect -5331 -781 -5315 -747
rect -5137 -781 -5121 -747
rect -5331 -797 -5121 -781
rect -5063 -747 -4853 -700
rect -5063 -781 -5047 -747
rect -4869 -781 -4853 -747
rect -5063 -797 -4853 -781
rect -4795 -747 -4585 -700
rect -4795 -781 -4779 -747
rect -4601 -781 -4585 -747
rect -4795 -797 -4585 -781
rect -4527 -747 -4317 -700
rect -4527 -781 -4511 -747
rect -4333 -781 -4317 -747
rect -4527 -797 -4317 -781
rect -4259 -747 -4049 -700
rect -4259 -781 -4243 -747
rect -4065 -781 -4049 -747
rect -4259 -797 -4049 -781
rect -3991 -747 -3781 -700
rect -3991 -781 -3975 -747
rect -3797 -781 -3781 -747
rect -3991 -797 -3781 -781
rect -3723 -747 -3513 -700
rect -3723 -781 -3707 -747
rect -3529 -781 -3513 -747
rect -3723 -797 -3513 -781
rect -3455 -747 -3245 -700
rect -3455 -781 -3439 -747
rect -3261 -781 -3245 -747
rect -3455 -797 -3245 -781
rect -3187 -747 -2977 -700
rect -3187 -781 -3171 -747
rect -2993 -781 -2977 -747
rect -3187 -797 -2977 -781
rect -2919 -747 -2709 -700
rect -2919 -781 -2903 -747
rect -2725 -781 -2709 -747
rect -2919 -797 -2709 -781
rect -2651 -747 -2441 -700
rect -2651 -781 -2635 -747
rect -2457 -781 -2441 -747
rect -2651 -797 -2441 -781
rect -2383 -747 -2173 -700
rect -2383 -781 -2367 -747
rect -2189 -781 -2173 -747
rect -2383 -797 -2173 -781
rect -2115 -747 -1905 -700
rect -2115 -781 -2099 -747
rect -1921 -781 -1905 -747
rect -2115 -797 -1905 -781
rect -1847 -747 -1637 -700
rect -1847 -781 -1831 -747
rect -1653 -781 -1637 -747
rect -1847 -797 -1637 -781
rect -1579 -747 -1369 -700
rect -1579 -781 -1563 -747
rect -1385 -781 -1369 -747
rect -1579 -797 -1369 -781
rect -1311 -747 -1101 -700
rect -1311 -781 -1295 -747
rect -1117 -781 -1101 -747
rect -1311 -797 -1101 -781
rect -1043 -747 -833 -700
rect -1043 -781 -1027 -747
rect -849 -781 -833 -747
rect -1043 -797 -833 -781
rect -775 -747 -565 -700
rect -775 -781 -759 -747
rect -581 -781 -565 -747
rect -775 -797 -565 -781
rect -507 -747 -297 -700
rect -507 -781 -491 -747
rect -313 -781 -297 -747
rect -507 -797 -297 -781
rect -239 -747 -29 -700
rect -239 -781 -223 -747
rect -45 -781 -29 -747
rect -239 -797 -29 -781
rect 29 -747 239 -700
rect 29 -781 45 -747
rect 223 -781 239 -747
rect 29 -797 239 -781
rect 297 -747 507 -700
rect 297 -781 313 -747
rect 491 -781 507 -747
rect 297 -797 507 -781
rect 565 -747 775 -700
rect 565 -781 581 -747
rect 759 -781 775 -747
rect 565 -797 775 -781
rect 833 -747 1043 -700
rect 833 -781 849 -747
rect 1027 -781 1043 -747
rect 833 -797 1043 -781
rect 1101 -747 1311 -700
rect 1101 -781 1117 -747
rect 1295 -781 1311 -747
rect 1101 -797 1311 -781
rect 1369 -747 1579 -700
rect 1369 -781 1385 -747
rect 1563 -781 1579 -747
rect 1369 -797 1579 -781
rect 1637 -747 1847 -700
rect 1637 -781 1653 -747
rect 1831 -781 1847 -747
rect 1637 -797 1847 -781
rect 1905 -747 2115 -700
rect 1905 -781 1921 -747
rect 2099 -781 2115 -747
rect 1905 -797 2115 -781
rect 2173 -747 2383 -700
rect 2173 -781 2189 -747
rect 2367 -781 2383 -747
rect 2173 -797 2383 -781
rect 2441 -747 2651 -700
rect 2441 -781 2457 -747
rect 2635 -781 2651 -747
rect 2441 -797 2651 -781
rect 2709 -747 2919 -700
rect 2709 -781 2725 -747
rect 2903 -781 2919 -747
rect 2709 -797 2919 -781
rect 2977 -747 3187 -700
rect 2977 -781 2993 -747
rect 3171 -781 3187 -747
rect 2977 -797 3187 -781
rect 3245 -747 3455 -700
rect 3245 -781 3261 -747
rect 3439 -781 3455 -747
rect 3245 -797 3455 -781
rect 3513 -747 3723 -700
rect 3513 -781 3529 -747
rect 3707 -781 3723 -747
rect 3513 -797 3723 -781
rect 3781 -747 3991 -700
rect 3781 -781 3797 -747
rect 3975 -781 3991 -747
rect 3781 -797 3991 -781
rect 4049 -747 4259 -700
rect 4049 -781 4065 -747
rect 4243 -781 4259 -747
rect 4049 -797 4259 -781
rect 4317 -747 4527 -700
rect 4317 -781 4333 -747
rect 4511 -781 4527 -747
rect 4317 -797 4527 -781
rect 4585 -747 4795 -700
rect 4585 -781 4601 -747
rect 4779 -781 4795 -747
rect 4585 -797 4795 -781
rect 4853 -747 5063 -700
rect 4853 -781 4869 -747
rect 5047 -781 5063 -747
rect 4853 -797 5063 -781
rect 5121 -747 5331 -700
rect 5121 -781 5137 -747
rect 5315 -781 5331 -747
rect 5121 -797 5331 -781
rect 5389 -747 5599 -700
rect 5389 -781 5405 -747
rect 5583 -781 5599 -747
rect 5389 -797 5599 -781
rect 5657 -747 5867 -700
rect 5657 -781 5673 -747
rect 5851 -781 5867 -747
rect 5657 -797 5867 -781
rect 5925 -747 6135 -700
rect 5925 -781 5941 -747
rect 6119 -781 6135 -747
rect 5925 -797 6135 -781
rect 6193 -747 6403 -700
rect 6193 -781 6209 -747
rect 6387 -781 6403 -747
rect 6193 -797 6403 -781
rect 6461 -747 6671 -700
rect 6461 -781 6477 -747
rect 6655 -781 6671 -747
rect 6461 -797 6671 -781
<< polycont >>
rect -6655 747 -6477 781
rect -6387 747 -6209 781
rect -6119 747 -5941 781
rect -5851 747 -5673 781
rect -5583 747 -5405 781
rect -5315 747 -5137 781
rect -5047 747 -4869 781
rect -4779 747 -4601 781
rect -4511 747 -4333 781
rect -4243 747 -4065 781
rect -3975 747 -3797 781
rect -3707 747 -3529 781
rect -3439 747 -3261 781
rect -3171 747 -2993 781
rect -2903 747 -2725 781
rect -2635 747 -2457 781
rect -2367 747 -2189 781
rect -2099 747 -1921 781
rect -1831 747 -1653 781
rect -1563 747 -1385 781
rect -1295 747 -1117 781
rect -1027 747 -849 781
rect -759 747 -581 781
rect -491 747 -313 781
rect -223 747 -45 781
rect 45 747 223 781
rect 313 747 491 781
rect 581 747 759 781
rect 849 747 1027 781
rect 1117 747 1295 781
rect 1385 747 1563 781
rect 1653 747 1831 781
rect 1921 747 2099 781
rect 2189 747 2367 781
rect 2457 747 2635 781
rect 2725 747 2903 781
rect 2993 747 3171 781
rect 3261 747 3439 781
rect 3529 747 3707 781
rect 3797 747 3975 781
rect 4065 747 4243 781
rect 4333 747 4511 781
rect 4601 747 4779 781
rect 4869 747 5047 781
rect 5137 747 5315 781
rect 5405 747 5583 781
rect 5673 747 5851 781
rect 5941 747 6119 781
rect 6209 747 6387 781
rect 6477 747 6655 781
rect -6655 -781 -6477 -747
rect -6387 -781 -6209 -747
rect -6119 -781 -5941 -747
rect -5851 -781 -5673 -747
rect -5583 -781 -5405 -747
rect -5315 -781 -5137 -747
rect -5047 -781 -4869 -747
rect -4779 -781 -4601 -747
rect -4511 -781 -4333 -747
rect -4243 -781 -4065 -747
rect -3975 -781 -3797 -747
rect -3707 -781 -3529 -747
rect -3439 -781 -3261 -747
rect -3171 -781 -2993 -747
rect -2903 -781 -2725 -747
rect -2635 -781 -2457 -747
rect -2367 -781 -2189 -747
rect -2099 -781 -1921 -747
rect -1831 -781 -1653 -747
rect -1563 -781 -1385 -747
rect -1295 -781 -1117 -747
rect -1027 -781 -849 -747
rect -759 -781 -581 -747
rect -491 -781 -313 -747
rect -223 -781 -45 -747
rect 45 -781 223 -747
rect 313 -781 491 -747
rect 581 -781 759 -747
rect 849 -781 1027 -747
rect 1117 -781 1295 -747
rect 1385 -781 1563 -747
rect 1653 -781 1831 -747
rect 1921 -781 2099 -747
rect 2189 -781 2367 -747
rect 2457 -781 2635 -747
rect 2725 -781 2903 -747
rect 2993 -781 3171 -747
rect 3261 -781 3439 -747
rect 3529 -781 3707 -747
rect 3797 -781 3975 -747
rect 4065 -781 4243 -747
rect 4333 -781 4511 -747
rect 4601 -781 4779 -747
rect 4869 -781 5047 -747
rect 5137 -781 5315 -747
rect 5405 -781 5583 -747
rect 5673 -781 5851 -747
rect 5941 -781 6119 -747
rect 6209 -781 6387 -747
rect 6477 -781 6655 -747
<< locali >>
rect -6831 849 -6735 883
rect 6735 849 6831 883
rect -6831 787 -6797 849
rect 6797 787 6831 849
rect -6671 747 -6655 781
rect -6477 747 -6461 781
rect -6403 747 -6387 781
rect -6209 747 -6193 781
rect -6135 747 -6119 781
rect -5941 747 -5925 781
rect -5867 747 -5851 781
rect -5673 747 -5657 781
rect -5599 747 -5583 781
rect -5405 747 -5389 781
rect -5331 747 -5315 781
rect -5137 747 -5121 781
rect -5063 747 -5047 781
rect -4869 747 -4853 781
rect -4795 747 -4779 781
rect -4601 747 -4585 781
rect -4527 747 -4511 781
rect -4333 747 -4317 781
rect -4259 747 -4243 781
rect -4065 747 -4049 781
rect -3991 747 -3975 781
rect -3797 747 -3781 781
rect -3723 747 -3707 781
rect -3529 747 -3513 781
rect -3455 747 -3439 781
rect -3261 747 -3245 781
rect -3187 747 -3171 781
rect -2993 747 -2977 781
rect -2919 747 -2903 781
rect -2725 747 -2709 781
rect -2651 747 -2635 781
rect -2457 747 -2441 781
rect -2383 747 -2367 781
rect -2189 747 -2173 781
rect -2115 747 -2099 781
rect -1921 747 -1905 781
rect -1847 747 -1831 781
rect -1653 747 -1637 781
rect -1579 747 -1563 781
rect -1385 747 -1369 781
rect -1311 747 -1295 781
rect -1117 747 -1101 781
rect -1043 747 -1027 781
rect -849 747 -833 781
rect -775 747 -759 781
rect -581 747 -565 781
rect -507 747 -491 781
rect -313 747 -297 781
rect -239 747 -223 781
rect -45 747 -29 781
rect 29 747 45 781
rect 223 747 239 781
rect 297 747 313 781
rect 491 747 507 781
rect 565 747 581 781
rect 759 747 775 781
rect 833 747 849 781
rect 1027 747 1043 781
rect 1101 747 1117 781
rect 1295 747 1311 781
rect 1369 747 1385 781
rect 1563 747 1579 781
rect 1637 747 1653 781
rect 1831 747 1847 781
rect 1905 747 1921 781
rect 2099 747 2115 781
rect 2173 747 2189 781
rect 2367 747 2383 781
rect 2441 747 2457 781
rect 2635 747 2651 781
rect 2709 747 2725 781
rect 2903 747 2919 781
rect 2977 747 2993 781
rect 3171 747 3187 781
rect 3245 747 3261 781
rect 3439 747 3455 781
rect 3513 747 3529 781
rect 3707 747 3723 781
rect 3781 747 3797 781
rect 3975 747 3991 781
rect 4049 747 4065 781
rect 4243 747 4259 781
rect 4317 747 4333 781
rect 4511 747 4527 781
rect 4585 747 4601 781
rect 4779 747 4795 781
rect 4853 747 4869 781
rect 5047 747 5063 781
rect 5121 747 5137 781
rect 5315 747 5331 781
rect 5389 747 5405 781
rect 5583 747 5599 781
rect 5657 747 5673 781
rect 5851 747 5867 781
rect 5925 747 5941 781
rect 6119 747 6135 781
rect 6193 747 6209 781
rect 6387 747 6403 781
rect 6461 747 6477 781
rect 6655 747 6671 781
rect -6717 688 -6683 704
rect -6717 -704 -6683 -688
rect -6449 688 -6415 704
rect -6449 -704 -6415 -688
rect -6181 688 -6147 704
rect -6181 -704 -6147 -688
rect -5913 688 -5879 704
rect -5913 -704 -5879 -688
rect -5645 688 -5611 704
rect -5645 -704 -5611 -688
rect -5377 688 -5343 704
rect -5377 -704 -5343 -688
rect -5109 688 -5075 704
rect -5109 -704 -5075 -688
rect -4841 688 -4807 704
rect -4841 -704 -4807 -688
rect -4573 688 -4539 704
rect -4573 -704 -4539 -688
rect -4305 688 -4271 704
rect -4305 -704 -4271 -688
rect -4037 688 -4003 704
rect -4037 -704 -4003 -688
rect -3769 688 -3735 704
rect -3769 -704 -3735 -688
rect -3501 688 -3467 704
rect -3501 -704 -3467 -688
rect -3233 688 -3199 704
rect -3233 -704 -3199 -688
rect -2965 688 -2931 704
rect -2965 -704 -2931 -688
rect -2697 688 -2663 704
rect -2697 -704 -2663 -688
rect -2429 688 -2395 704
rect -2429 -704 -2395 -688
rect -2161 688 -2127 704
rect -2161 -704 -2127 -688
rect -1893 688 -1859 704
rect -1893 -704 -1859 -688
rect -1625 688 -1591 704
rect -1625 -704 -1591 -688
rect -1357 688 -1323 704
rect -1357 -704 -1323 -688
rect -1089 688 -1055 704
rect -1089 -704 -1055 -688
rect -821 688 -787 704
rect -821 -704 -787 -688
rect -553 688 -519 704
rect -553 -704 -519 -688
rect -285 688 -251 704
rect -285 -704 -251 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 251 688 285 704
rect 251 -704 285 -688
rect 519 688 553 704
rect 519 -704 553 -688
rect 787 688 821 704
rect 787 -704 821 -688
rect 1055 688 1089 704
rect 1055 -704 1089 -688
rect 1323 688 1357 704
rect 1323 -704 1357 -688
rect 1591 688 1625 704
rect 1591 -704 1625 -688
rect 1859 688 1893 704
rect 1859 -704 1893 -688
rect 2127 688 2161 704
rect 2127 -704 2161 -688
rect 2395 688 2429 704
rect 2395 -704 2429 -688
rect 2663 688 2697 704
rect 2663 -704 2697 -688
rect 2931 688 2965 704
rect 2931 -704 2965 -688
rect 3199 688 3233 704
rect 3199 -704 3233 -688
rect 3467 688 3501 704
rect 3467 -704 3501 -688
rect 3735 688 3769 704
rect 3735 -704 3769 -688
rect 4003 688 4037 704
rect 4003 -704 4037 -688
rect 4271 688 4305 704
rect 4271 -704 4305 -688
rect 4539 688 4573 704
rect 4539 -704 4573 -688
rect 4807 688 4841 704
rect 4807 -704 4841 -688
rect 5075 688 5109 704
rect 5075 -704 5109 -688
rect 5343 688 5377 704
rect 5343 -704 5377 -688
rect 5611 688 5645 704
rect 5611 -704 5645 -688
rect 5879 688 5913 704
rect 5879 -704 5913 -688
rect 6147 688 6181 704
rect 6147 -704 6181 -688
rect 6415 688 6449 704
rect 6415 -704 6449 -688
rect 6683 688 6717 704
rect 6683 -704 6717 -688
rect -6671 -781 -6655 -747
rect -6477 -781 -6461 -747
rect -6403 -781 -6387 -747
rect -6209 -781 -6193 -747
rect -6135 -781 -6119 -747
rect -5941 -781 -5925 -747
rect -5867 -781 -5851 -747
rect -5673 -781 -5657 -747
rect -5599 -781 -5583 -747
rect -5405 -781 -5389 -747
rect -5331 -781 -5315 -747
rect -5137 -781 -5121 -747
rect -5063 -781 -5047 -747
rect -4869 -781 -4853 -747
rect -4795 -781 -4779 -747
rect -4601 -781 -4585 -747
rect -4527 -781 -4511 -747
rect -4333 -781 -4317 -747
rect -4259 -781 -4243 -747
rect -4065 -781 -4049 -747
rect -3991 -781 -3975 -747
rect -3797 -781 -3781 -747
rect -3723 -781 -3707 -747
rect -3529 -781 -3513 -747
rect -3455 -781 -3439 -747
rect -3261 -781 -3245 -747
rect -3187 -781 -3171 -747
rect -2993 -781 -2977 -747
rect -2919 -781 -2903 -747
rect -2725 -781 -2709 -747
rect -2651 -781 -2635 -747
rect -2457 -781 -2441 -747
rect -2383 -781 -2367 -747
rect -2189 -781 -2173 -747
rect -2115 -781 -2099 -747
rect -1921 -781 -1905 -747
rect -1847 -781 -1831 -747
rect -1653 -781 -1637 -747
rect -1579 -781 -1563 -747
rect -1385 -781 -1369 -747
rect -1311 -781 -1295 -747
rect -1117 -781 -1101 -747
rect -1043 -781 -1027 -747
rect -849 -781 -833 -747
rect -775 -781 -759 -747
rect -581 -781 -565 -747
rect -507 -781 -491 -747
rect -313 -781 -297 -747
rect -239 -781 -223 -747
rect -45 -781 -29 -747
rect 29 -781 45 -747
rect 223 -781 239 -747
rect 297 -781 313 -747
rect 491 -781 507 -747
rect 565 -781 581 -747
rect 759 -781 775 -747
rect 833 -781 849 -747
rect 1027 -781 1043 -747
rect 1101 -781 1117 -747
rect 1295 -781 1311 -747
rect 1369 -781 1385 -747
rect 1563 -781 1579 -747
rect 1637 -781 1653 -747
rect 1831 -781 1847 -747
rect 1905 -781 1921 -747
rect 2099 -781 2115 -747
rect 2173 -781 2189 -747
rect 2367 -781 2383 -747
rect 2441 -781 2457 -747
rect 2635 -781 2651 -747
rect 2709 -781 2725 -747
rect 2903 -781 2919 -747
rect 2977 -781 2993 -747
rect 3171 -781 3187 -747
rect 3245 -781 3261 -747
rect 3439 -781 3455 -747
rect 3513 -781 3529 -747
rect 3707 -781 3723 -747
rect 3781 -781 3797 -747
rect 3975 -781 3991 -747
rect 4049 -781 4065 -747
rect 4243 -781 4259 -747
rect 4317 -781 4333 -747
rect 4511 -781 4527 -747
rect 4585 -781 4601 -747
rect 4779 -781 4795 -747
rect 4853 -781 4869 -747
rect 5047 -781 5063 -747
rect 5121 -781 5137 -747
rect 5315 -781 5331 -747
rect 5389 -781 5405 -747
rect 5583 -781 5599 -747
rect 5657 -781 5673 -747
rect 5851 -781 5867 -747
rect 5925 -781 5941 -747
rect 6119 -781 6135 -747
rect 6193 -781 6209 -747
rect 6387 -781 6403 -747
rect 6461 -781 6477 -747
rect 6655 -781 6671 -747
rect -6831 -849 -6797 -787
rect 6797 -849 6831 -787
rect -6831 -883 -6735 -849
rect 6735 -883 6831 -849
<< viali >>
rect -6655 747 -6477 781
rect -6387 747 -6209 781
rect -6119 747 -5941 781
rect -5851 747 -5673 781
rect -5583 747 -5405 781
rect -5315 747 -5137 781
rect -5047 747 -4869 781
rect -4779 747 -4601 781
rect -4511 747 -4333 781
rect -4243 747 -4065 781
rect -3975 747 -3797 781
rect -3707 747 -3529 781
rect -3439 747 -3261 781
rect -3171 747 -2993 781
rect -2903 747 -2725 781
rect -2635 747 -2457 781
rect -2367 747 -2189 781
rect -2099 747 -1921 781
rect -1831 747 -1653 781
rect -1563 747 -1385 781
rect -1295 747 -1117 781
rect -1027 747 -849 781
rect -759 747 -581 781
rect -491 747 -313 781
rect -223 747 -45 781
rect 45 747 223 781
rect 313 747 491 781
rect 581 747 759 781
rect 849 747 1027 781
rect 1117 747 1295 781
rect 1385 747 1563 781
rect 1653 747 1831 781
rect 1921 747 2099 781
rect 2189 747 2367 781
rect 2457 747 2635 781
rect 2725 747 2903 781
rect 2993 747 3171 781
rect 3261 747 3439 781
rect 3529 747 3707 781
rect 3797 747 3975 781
rect 4065 747 4243 781
rect 4333 747 4511 781
rect 4601 747 4779 781
rect 4869 747 5047 781
rect 5137 747 5315 781
rect 5405 747 5583 781
rect 5673 747 5851 781
rect 5941 747 6119 781
rect 6209 747 6387 781
rect 6477 747 6655 781
rect -6717 -688 -6683 688
rect -6449 -688 -6415 688
rect -6181 -688 -6147 688
rect -5913 -688 -5879 688
rect -5645 -688 -5611 688
rect -5377 -688 -5343 688
rect -5109 -688 -5075 688
rect -4841 -688 -4807 688
rect -4573 -688 -4539 688
rect -4305 -688 -4271 688
rect -4037 -688 -4003 688
rect -3769 -688 -3735 688
rect -3501 -688 -3467 688
rect -3233 -688 -3199 688
rect -2965 -688 -2931 688
rect -2697 -688 -2663 688
rect -2429 -688 -2395 688
rect -2161 -688 -2127 688
rect -1893 -688 -1859 688
rect -1625 -688 -1591 688
rect -1357 -688 -1323 688
rect -1089 -688 -1055 688
rect -821 -688 -787 688
rect -553 -688 -519 688
rect -285 -688 -251 688
rect -17 -688 17 688
rect 251 -688 285 688
rect 519 -688 553 688
rect 787 -688 821 688
rect 1055 -688 1089 688
rect 1323 -688 1357 688
rect 1591 -688 1625 688
rect 1859 -688 1893 688
rect 2127 -688 2161 688
rect 2395 -688 2429 688
rect 2663 -688 2697 688
rect 2931 -688 2965 688
rect 3199 -688 3233 688
rect 3467 -688 3501 688
rect 3735 -688 3769 688
rect 4003 -688 4037 688
rect 4271 -688 4305 688
rect 4539 -688 4573 688
rect 4807 -688 4841 688
rect 5075 -688 5109 688
rect 5343 -688 5377 688
rect 5611 -688 5645 688
rect 5879 -688 5913 688
rect 6147 -688 6181 688
rect 6415 -688 6449 688
rect 6683 -688 6717 688
rect -6655 -781 -6477 -747
rect -6387 -781 -6209 -747
rect -6119 -781 -5941 -747
rect -5851 -781 -5673 -747
rect -5583 -781 -5405 -747
rect -5315 -781 -5137 -747
rect -5047 -781 -4869 -747
rect -4779 -781 -4601 -747
rect -4511 -781 -4333 -747
rect -4243 -781 -4065 -747
rect -3975 -781 -3797 -747
rect -3707 -781 -3529 -747
rect -3439 -781 -3261 -747
rect -3171 -781 -2993 -747
rect -2903 -781 -2725 -747
rect -2635 -781 -2457 -747
rect -2367 -781 -2189 -747
rect -2099 -781 -1921 -747
rect -1831 -781 -1653 -747
rect -1563 -781 -1385 -747
rect -1295 -781 -1117 -747
rect -1027 -781 -849 -747
rect -759 -781 -581 -747
rect -491 -781 -313 -747
rect -223 -781 -45 -747
rect 45 -781 223 -747
rect 313 -781 491 -747
rect 581 -781 759 -747
rect 849 -781 1027 -747
rect 1117 -781 1295 -747
rect 1385 -781 1563 -747
rect 1653 -781 1831 -747
rect 1921 -781 2099 -747
rect 2189 -781 2367 -747
rect 2457 -781 2635 -747
rect 2725 -781 2903 -747
rect 2993 -781 3171 -747
rect 3261 -781 3439 -747
rect 3529 -781 3707 -747
rect 3797 -781 3975 -747
rect 4065 -781 4243 -747
rect 4333 -781 4511 -747
rect 4601 -781 4779 -747
rect 4869 -781 5047 -747
rect 5137 -781 5315 -747
rect 5405 -781 5583 -747
rect 5673 -781 5851 -747
rect 5941 -781 6119 -747
rect 6209 -781 6387 -747
rect 6477 -781 6655 -747
<< metal1 >>
rect -6667 781 -6465 787
rect -6667 747 -6655 781
rect -6477 747 -6465 781
rect -6667 741 -6465 747
rect -6399 781 -6197 787
rect -6399 747 -6387 781
rect -6209 747 -6197 781
rect -6399 741 -6197 747
rect -6131 781 -5929 787
rect -6131 747 -6119 781
rect -5941 747 -5929 781
rect -6131 741 -5929 747
rect -5863 781 -5661 787
rect -5863 747 -5851 781
rect -5673 747 -5661 781
rect -5863 741 -5661 747
rect -5595 781 -5393 787
rect -5595 747 -5583 781
rect -5405 747 -5393 781
rect -5595 741 -5393 747
rect -5327 781 -5125 787
rect -5327 747 -5315 781
rect -5137 747 -5125 781
rect -5327 741 -5125 747
rect -5059 781 -4857 787
rect -5059 747 -5047 781
rect -4869 747 -4857 781
rect -5059 741 -4857 747
rect -4791 781 -4589 787
rect -4791 747 -4779 781
rect -4601 747 -4589 781
rect -4791 741 -4589 747
rect -4523 781 -4321 787
rect -4523 747 -4511 781
rect -4333 747 -4321 781
rect -4523 741 -4321 747
rect -4255 781 -4053 787
rect -4255 747 -4243 781
rect -4065 747 -4053 781
rect -4255 741 -4053 747
rect -3987 781 -3785 787
rect -3987 747 -3975 781
rect -3797 747 -3785 781
rect -3987 741 -3785 747
rect -3719 781 -3517 787
rect -3719 747 -3707 781
rect -3529 747 -3517 781
rect -3719 741 -3517 747
rect -3451 781 -3249 787
rect -3451 747 -3439 781
rect -3261 747 -3249 781
rect -3451 741 -3249 747
rect -3183 781 -2981 787
rect -3183 747 -3171 781
rect -2993 747 -2981 781
rect -3183 741 -2981 747
rect -2915 781 -2713 787
rect -2915 747 -2903 781
rect -2725 747 -2713 781
rect -2915 741 -2713 747
rect -2647 781 -2445 787
rect -2647 747 -2635 781
rect -2457 747 -2445 781
rect -2647 741 -2445 747
rect -2379 781 -2177 787
rect -2379 747 -2367 781
rect -2189 747 -2177 781
rect -2379 741 -2177 747
rect -2111 781 -1909 787
rect -2111 747 -2099 781
rect -1921 747 -1909 781
rect -2111 741 -1909 747
rect -1843 781 -1641 787
rect -1843 747 -1831 781
rect -1653 747 -1641 781
rect -1843 741 -1641 747
rect -1575 781 -1373 787
rect -1575 747 -1563 781
rect -1385 747 -1373 781
rect -1575 741 -1373 747
rect -1307 781 -1105 787
rect -1307 747 -1295 781
rect -1117 747 -1105 781
rect -1307 741 -1105 747
rect -1039 781 -837 787
rect -1039 747 -1027 781
rect -849 747 -837 781
rect -1039 741 -837 747
rect -771 781 -569 787
rect -771 747 -759 781
rect -581 747 -569 781
rect -771 741 -569 747
rect -503 781 -301 787
rect -503 747 -491 781
rect -313 747 -301 781
rect -503 741 -301 747
rect -235 781 -33 787
rect -235 747 -223 781
rect -45 747 -33 781
rect -235 741 -33 747
rect 33 781 235 787
rect 33 747 45 781
rect 223 747 235 781
rect 33 741 235 747
rect 301 781 503 787
rect 301 747 313 781
rect 491 747 503 781
rect 301 741 503 747
rect 569 781 771 787
rect 569 747 581 781
rect 759 747 771 781
rect 569 741 771 747
rect 837 781 1039 787
rect 837 747 849 781
rect 1027 747 1039 781
rect 837 741 1039 747
rect 1105 781 1307 787
rect 1105 747 1117 781
rect 1295 747 1307 781
rect 1105 741 1307 747
rect 1373 781 1575 787
rect 1373 747 1385 781
rect 1563 747 1575 781
rect 1373 741 1575 747
rect 1641 781 1843 787
rect 1641 747 1653 781
rect 1831 747 1843 781
rect 1641 741 1843 747
rect 1909 781 2111 787
rect 1909 747 1921 781
rect 2099 747 2111 781
rect 1909 741 2111 747
rect 2177 781 2379 787
rect 2177 747 2189 781
rect 2367 747 2379 781
rect 2177 741 2379 747
rect 2445 781 2647 787
rect 2445 747 2457 781
rect 2635 747 2647 781
rect 2445 741 2647 747
rect 2713 781 2915 787
rect 2713 747 2725 781
rect 2903 747 2915 781
rect 2713 741 2915 747
rect 2981 781 3183 787
rect 2981 747 2993 781
rect 3171 747 3183 781
rect 2981 741 3183 747
rect 3249 781 3451 787
rect 3249 747 3261 781
rect 3439 747 3451 781
rect 3249 741 3451 747
rect 3517 781 3719 787
rect 3517 747 3529 781
rect 3707 747 3719 781
rect 3517 741 3719 747
rect 3785 781 3987 787
rect 3785 747 3797 781
rect 3975 747 3987 781
rect 3785 741 3987 747
rect 4053 781 4255 787
rect 4053 747 4065 781
rect 4243 747 4255 781
rect 4053 741 4255 747
rect 4321 781 4523 787
rect 4321 747 4333 781
rect 4511 747 4523 781
rect 4321 741 4523 747
rect 4589 781 4791 787
rect 4589 747 4601 781
rect 4779 747 4791 781
rect 4589 741 4791 747
rect 4857 781 5059 787
rect 4857 747 4869 781
rect 5047 747 5059 781
rect 4857 741 5059 747
rect 5125 781 5327 787
rect 5125 747 5137 781
rect 5315 747 5327 781
rect 5125 741 5327 747
rect 5393 781 5595 787
rect 5393 747 5405 781
rect 5583 747 5595 781
rect 5393 741 5595 747
rect 5661 781 5863 787
rect 5661 747 5673 781
rect 5851 747 5863 781
rect 5661 741 5863 747
rect 5929 781 6131 787
rect 5929 747 5941 781
rect 6119 747 6131 781
rect 5929 741 6131 747
rect 6197 781 6399 787
rect 6197 747 6209 781
rect 6387 747 6399 781
rect 6197 741 6399 747
rect 6465 781 6667 787
rect 6465 747 6477 781
rect 6655 747 6667 781
rect 6465 741 6667 747
rect -6723 688 -6677 700
rect -6723 -688 -6717 688
rect -6683 -688 -6677 688
rect -6723 -700 -6677 -688
rect -6455 688 -6409 700
rect -6455 -688 -6449 688
rect -6415 -688 -6409 688
rect -6455 -700 -6409 -688
rect -6187 688 -6141 700
rect -6187 -688 -6181 688
rect -6147 -688 -6141 688
rect -6187 -700 -6141 -688
rect -5919 688 -5873 700
rect -5919 -688 -5913 688
rect -5879 -688 -5873 688
rect -5919 -700 -5873 -688
rect -5651 688 -5605 700
rect -5651 -688 -5645 688
rect -5611 -688 -5605 688
rect -5651 -700 -5605 -688
rect -5383 688 -5337 700
rect -5383 -688 -5377 688
rect -5343 -688 -5337 688
rect -5383 -700 -5337 -688
rect -5115 688 -5069 700
rect -5115 -688 -5109 688
rect -5075 -688 -5069 688
rect -5115 -700 -5069 -688
rect -4847 688 -4801 700
rect -4847 -688 -4841 688
rect -4807 -688 -4801 688
rect -4847 -700 -4801 -688
rect -4579 688 -4533 700
rect -4579 -688 -4573 688
rect -4539 -688 -4533 688
rect -4579 -700 -4533 -688
rect -4311 688 -4265 700
rect -4311 -688 -4305 688
rect -4271 -688 -4265 688
rect -4311 -700 -4265 -688
rect -4043 688 -3997 700
rect -4043 -688 -4037 688
rect -4003 -688 -3997 688
rect -4043 -700 -3997 -688
rect -3775 688 -3729 700
rect -3775 -688 -3769 688
rect -3735 -688 -3729 688
rect -3775 -700 -3729 -688
rect -3507 688 -3461 700
rect -3507 -688 -3501 688
rect -3467 -688 -3461 688
rect -3507 -700 -3461 -688
rect -3239 688 -3193 700
rect -3239 -688 -3233 688
rect -3199 -688 -3193 688
rect -3239 -700 -3193 -688
rect -2971 688 -2925 700
rect -2971 -688 -2965 688
rect -2931 -688 -2925 688
rect -2971 -700 -2925 -688
rect -2703 688 -2657 700
rect -2703 -688 -2697 688
rect -2663 -688 -2657 688
rect -2703 -700 -2657 -688
rect -2435 688 -2389 700
rect -2435 -688 -2429 688
rect -2395 -688 -2389 688
rect -2435 -700 -2389 -688
rect -2167 688 -2121 700
rect -2167 -688 -2161 688
rect -2127 -688 -2121 688
rect -2167 -700 -2121 -688
rect -1899 688 -1853 700
rect -1899 -688 -1893 688
rect -1859 -688 -1853 688
rect -1899 -700 -1853 -688
rect -1631 688 -1585 700
rect -1631 -688 -1625 688
rect -1591 -688 -1585 688
rect -1631 -700 -1585 -688
rect -1363 688 -1317 700
rect -1363 -688 -1357 688
rect -1323 -688 -1317 688
rect -1363 -700 -1317 -688
rect -1095 688 -1049 700
rect -1095 -688 -1089 688
rect -1055 -688 -1049 688
rect -1095 -700 -1049 -688
rect -827 688 -781 700
rect -827 -688 -821 688
rect -787 -688 -781 688
rect -827 -700 -781 -688
rect -559 688 -513 700
rect -559 -688 -553 688
rect -519 -688 -513 688
rect -559 -700 -513 -688
rect -291 688 -245 700
rect -291 -688 -285 688
rect -251 -688 -245 688
rect -291 -700 -245 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 245 688 291 700
rect 245 -688 251 688
rect 285 -688 291 688
rect 245 -700 291 -688
rect 513 688 559 700
rect 513 -688 519 688
rect 553 -688 559 688
rect 513 -700 559 -688
rect 781 688 827 700
rect 781 -688 787 688
rect 821 -688 827 688
rect 781 -700 827 -688
rect 1049 688 1095 700
rect 1049 -688 1055 688
rect 1089 -688 1095 688
rect 1049 -700 1095 -688
rect 1317 688 1363 700
rect 1317 -688 1323 688
rect 1357 -688 1363 688
rect 1317 -700 1363 -688
rect 1585 688 1631 700
rect 1585 -688 1591 688
rect 1625 -688 1631 688
rect 1585 -700 1631 -688
rect 1853 688 1899 700
rect 1853 -688 1859 688
rect 1893 -688 1899 688
rect 1853 -700 1899 -688
rect 2121 688 2167 700
rect 2121 -688 2127 688
rect 2161 -688 2167 688
rect 2121 -700 2167 -688
rect 2389 688 2435 700
rect 2389 -688 2395 688
rect 2429 -688 2435 688
rect 2389 -700 2435 -688
rect 2657 688 2703 700
rect 2657 -688 2663 688
rect 2697 -688 2703 688
rect 2657 -700 2703 -688
rect 2925 688 2971 700
rect 2925 -688 2931 688
rect 2965 -688 2971 688
rect 2925 -700 2971 -688
rect 3193 688 3239 700
rect 3193 -688 3199 688
rect 3233 -688 3239 688
rect 3193 -700 3239 -688
rect 3461 688 3507 700
rect 3461 -688 3467 688
rect 3501 -688 3507 688
rect 3461 -700 3507 -688
rect 3729 688 3775 700
rect 3729 -688 3735 688
rect 3769 -688 3775 688
rect 3729 -700 3775 -688
rect 3997 688 4043 700
rect 3997 -688 4003 688
rect 4037 -688 4043 688
rect 3997 -700 4043 -688
rect 4265 688 4311 700
rect 4265 -688 4271 688
rect 4305 -688 4311 688
rect 4265 -700 4311 -688
rect 4533 688 4579 700
rect 4533 -688 4539 688
rect 4573 -688 4579 688
rect 4533 -700 4579 -688
rect 4801 688 4847 700
rect 4801 -688 4807 688
rect 4841 -688 4847 688
rect 4801 -700 4847 -688
rect 5069 688 5115 700
rect 5069 -688 5075 688
rect 5109 -688 5115 688
rect 5069 -700 5115 -688
rect 5337 688 5383 700
rect 5337 -688 5343 688
rect 5377 -688 5383 688
rect 5337 -700 5383 -688
rect 5605 688 5651 700
rect 5605 -688 5611 688
rect 5645 -688 5651 688
rect 5605 -700 5651 -688
rect 5873 688 5919 700
rect 5873 -688 5879 688
rect 5913 -688 5919 688
rect 5873 -700 5919 -688
rect 6141 688 6187 700
rect 6141 -688 6147 688
rect 6181 -688 6187 688
rect 6141 -700 6187 -688
rect 6409 688 6455 700
rect 6409 -688 6415 688
rect 6449 -688 6455 688
rect 6409 -700 6455 -688
rect 6677 688 6723 700
rect 6677 -688 6683 688
rect 6717 -688 6723 688
rect 6677 -700 6723 -688
rect -6667 -747 -6465 -741
rect -6667 -781 -6655 -747
rect -6477 -781 -6465 -747
rect -6667 -787 -6465 -781
rect -6399 -747 -6197 -741
rect -6399 -781 -6387 -747
rect -6209 -781 -6197 -747
rect -6399 -787 -6197 -781
rect -6131 -747 -5929 -741
rect -6131 -781 -6119 -747
rect -5941 -781 -5929 -747
rect -6131 -787 -5929 -781
rect -5863 -747 -5661 -741
rect -5863 -781 -5851 -747
rect -5673 -781 -5661 -747
rect -5863 -787 -5661 -781
rect -5595 -747 -5393 -741
rect -5595 -781 -5583 -747
rect -5405 -781 -5393 -747
rect -5595 -787 -5393 -781
rect -5327 -747 -5125 -741
rect -5327 -781 -5315 -747
rect -5137 -781 -5125 -747
rect -5327 -787 -5125 -781
rect -5059 -747 -4857 -741
rect -5059 -781 -5047 -747
rect -4869 -781 -4857 -747
rect -5059 -787 -4857 -781
rect -4791 -747 -4589 -741
rect -4791 -781 -4779 -747
rect -4601 -781 -4589 -747
rect -4791 -787 -4589 -781
rect -4523 -747 -4321 -741
rect -4523 -781 -4511 -747
rect -4333 -781 -4321 -747
rect -4523 -787 -4321 -781
rect -4255 -747 -4053 -741
rect -4255 -781 -4243 -747
rect -4065 -781 -4053 -747
rect -4255 -787 -4053 -781
rect -3987 -747 -3785 -741
rect -3987 -781 -3975 -747
rect -3797 -781 -3785 -747
rect -3987 -787 -3785 -781
rect -3719 -747 -3517 -741
rect -3719 -781 -3707 -747
rect -3529 -781 -3517 -747
rect -3719 -787 -3517 -781
rect -3451 -747 -3249 -741
rect -3451 -781 -3439 -747
rect -3261 -781 -3249 -747
rect -3451 -787 -3249 -781
rect -3183 -747 -2981 -741
rect -3183 -781 -3171 -747
rect -2993 -781 -2981 -747
rect -3183 -787 -2981 -781
rect -2915 -747 -2713 -741
rect -2915 -781 -2903 -747
rect -2725 -781 -2713 -747
rect -2915 -787 -2713 -781
rect -2647 -747 -2445 -741
rect -2647 -781 -2635 -747
rect -2457 -781 -2445 -747
rect -2647 -787 -2445 -781
rect -2379 -747 -2177 -741
rect -2379 -781 -2367 -747
rect -2189 -781 -2177 -747
rect -2379 -787 -2177 -781
rect -2111 -747 -1909 -741
rect -2111 -781 -2099 -747
rect -1921 -781 -1909 -747
rect -2111 -787 -1909 -781
rect -1843 -747 -1641 -741
rect -1843 -781 -1831 -747
rect -1653 -781 -1641 -747
rect -1843 -787 -1641 -781
rect -1575 -747 -1373 -741
rect -1575 -781 -1563 -747
rect -1385 -781 -1373 -747
rect -1575 -787 -1373 -781
rect -1307 -747 -1105 -741
rect -1307 -781 -1295 -747
rect -1117 -781 -1105 -747
rect -1307 -787 -1105 -781
rect -1039 -747 -837 -741
rect -1039 -781 -1027 -747
rect -849 -781 -837 -747
rect -1039 -787 -837 -781
rect -771 -747 -569 -741
rect -771 -781 -759 -747
rect -581 -781 -569 -747
rect -771 -787 -569 -781
rect -503 -747 -301 -741
rect -503 -781 -491 -747
rect -313 -781 -301 -747
rect -503 -787 -301 -781
rect -235 -747 -33 -741
rect -235 -781 -223 -747
rect -45 -781 -33 -747
rect -235 -787 -33 -781
rect 33 -747 235 -741
rect 33 -781 45 -747
rect 223 -781 235 -747
rect 33 -787 235 -781
rect 301 -747 503 -741
rect 301 -781 313 -747
rect 491 -781 503 -747
rect 301 -787 503 -781
rect 569 -747 771 -741
rect 569 -781 581 -747
rect 759 -781 771 -747
rect 569 -787 771 -781
rect 837 -747 1039 -741
rect 837 -781 849 -747
rect 1027 -781 1039 -747
rect 837 -787 1039 -781
rect 1105 -747 1307 -741
rect 1105 -781 1117 -747
rect 1295 -781 1307 -747
rect 1105 -787 1307 -781
rect 1373 -747 1575 -741
rect 1373 -781 1385 -747
rect 1563 -781 1575 -747
rect 1373 -787 1575 -781
rect 1641 -747 1843 -741
rect 1641 -781 1653 -747
rect 1831 -781 1843 -747
rect 1641 -787 1843 -781
rect 1909 -747 2111 -741
rect 1909 -781 1921 -747
rect 2099 -781 2111 -747
rect 1909 -787 2111 -781
rect 2177 -747 2379 -741
rect 2177 -781 2189 -747
rect 2367 -781 2379 -747
rect 2177 -787 2379 -781
rect 2445 -747 2647 -741
rect 2445 -781 2457 -747
rect 2635 -781 2647 -747
rect 2445 -787 2647 -781
rect 2713 -747 2915 -741
rect 2713 -781 2725 -747
rect 2903 -781 2915 -747
rect 2713 -787 2915 -781
rect 2981 -747 3183 -741
rect 2981 -781 2993 -747
rect 3171 -781 3183 -747
rect 2981 -787 3183 -781
rect 3249 -747 3451 -741
rect 3249 -781 3261 -747
rect 3439 -781 3451 -747
rect 3249 -787 3451 -781
rect 3517 -747 3719 -741
rect 3517 -781 3529 -747
rect 3707 -781 3719 -747
rect 3517 -787 3719 -781
rect 3785 -747 3987 -741
rect 3785 -781 3797 -747
rect 3975 -781 3987 -747
rect 3785 -787 3987 -781
rect 4053 -747 4255 -741
rect 4053 -781 4065 -747
rect 4243 -781 4255 -747
rect 4053 -787 4255 -781
rect 4321 -747 4523 -741
rect 4321 -781 4333 -747
rect 4511 -781 4523 -747
rect 4321 -787 4523 -781
rect 4589 -747 4791 -741
rect 4589 -781 4601 -747
rect 4779 -781 4791 -747
rect 4589 -787 4791 -781
rect 4857 -747 5059 -741
rect 4857 -781 4869 -747
rect 5047 -781 5059 -747
rect 4857 -787 5059 -781
rect 5125 -747 5327 -741
rect 5125 -781 5137 -747
rect 5315 -781 5327 -747
rect 5125 -787 5327 -781
rect 5393 -747 5595 -741
rect 5393 -781 5405 -747
rect 5583 -781 5595 -747
rect 5393 -787 5595 -781
rect 5661 -747 5863 -741
rect 5661 -781 5673 -747
rect 5851 -781 5863 -747
rect 5661 -787 5863 -781
rect 5929 -747 6131 -741
rect 5929 -781 5941 -747
rect 6119 -781 6131 -747
rect 5929 -787 6131 -781
rect 6197 -747 6399 -741
rect 6197 -781 6209 -747
rect 6387 -781 6399 -747
rect 6197 -787 6399 -781
rect 6465 -747 6667 -741
rect 6465 -781 6477 -747
rect 6655 -781 6667 -747
rect 6465 -787 6667 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -6814 -866 6814 866
string parameters w 7 l 1.05 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
