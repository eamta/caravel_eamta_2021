magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -4781 999 -4723 1005
rect -4589 999 -4531 1005
rect -4397 999 -4339 1005
rect -4205 999 -4147 1005
rect -4013 999 -3955 1005
rect -3821 999 -3763 1005
rect -3629 999 -3571 1005
rect -3437 999 -3379 1005
rect -3245 999 -3187 1005
rect -3053 999 -2995 1005
rect -2861 999 -2803 1005
rect -2669 999 -2611 1005
rect -2477 999 -2419 1005
rect -2285 999 -2227 1005
rect -2093 999 -2035 1005
rect -1901 999 -1843 1005
rect -1709 999 -1651 1005
rect -1517 999 -1459 1005
rect -1325 999 -1267 1005
rect -1133 999 -1075 1005
rect -941 999 -883 1005
rect -749 999 -691 1005
rect -557 999 -499 1005
rect -365 999 -307 1005
rect -173 999 -115 1005
rect 19 999 77 1005
rect 211 999 269 1005
rect 403 999 461 1005
rect 595 999 653 1005
rect 787 999 845 1005
rect 979 999 1037 1005
rect 1171 999 1229 1005
rect 1363 999 1421 1005
rect 1555 999 1613 1005
rect 1747 999 1805 1005
rect 1939 999 1997 1005
rect 2131 999 2189 1005
rect 2323 999 2381 1005
rect 2515 999 2573 1005
rect 2707 999 2765 1005
rect 2899 999 2957 1005
rect 3091 999 3149 1005
rect 3283 999 3341 1005
rect 3475 999 3533 1005
rect 3667 999 3725 1005
rect 3859 999 3917 1005
rect 4051 999 4109 1005
rect 4243 999 4301 1005
rect 4435 999 4493 1005
rect 4627 999 4685 1005
rect -4781 965 -4769 999
rect -4589 965 -4577 999
rect -4397 965 -4385 999
rect -4205 965 -4193 999
rect -4013 965 -4001 999
rect -3821 965 -3809 999
rect -3629 965 -3617 999
rect -3437 965 -3425 999
rect -3245 965 -3233 999
rect -3053 965 -3041 999
rect -2861 965 -2849 999
rect -2669 965 -2657 999
rect -2477 965 -2465 999
rect -2285 965 -2273 999
rect -2093 965 -2081 999
rect -1901 965 -1889 999
rect -1709 965 -1697 999
rect -1517 965 -1505 999
rect -1325 965 -1313 999
rect -1133 965 -1121 999
rect -941 965 -929 999
rect -749 965 -737 999
rect -557 965 -545 999
rect -365 965 -353 999
rect -173 965 -161 999
rect 19 965 31 999
rect 211 965 223 999
rect 403 965 415 999
rect 595 965 607 999
rect 787 965 799 999
rect 979 965 991 999
rect 1171 965 1183 999
rect 1363 965 1375 999
rect 1555 965 1567 999
rect 1747 965 1759 999
rect 1939 965 1951 999
rect 2131 965 2143 999
rect 2323 965 2335 999
rect 2515 965 2527 999
rect 2707 965 2719 999
rect 2899 965 2911 999
rect 3091 965 3103 999
rect 3283 965 3295 999
rect 3475 965 3487 999
rect 3667 965 3679 999
rect 3859 965 3871 999
rect 4051 965 4063 999
rect 4243 965 4255 999
rect 4435 965 4447 999
rect 4627 965 4639 999
rect -4781 959 -4723 965
rect -4589 959 -4531 965
rect -4397 959 -4339 965
rect -4205 959 -4147 965
rect -4013 959 -3955 965
rect -3821 959 -3763 965
rect -3629 959 -3571 965
rect -3437 959 -3379 965
rect -3245 959 -3187 965
rect -3053 959 -2995 965
rect -2861 959 -2803 965
rect -2669 959 -2611 965
rect -2477 959 -2419 965
rect -2285 959 -2227 965
rect -2093 959 -2035 965
rect -1901 959 -1843 965
rect -1709 959 -1651 965
rect -1517 959 -1459 965
rect -1325 959 -1267 965
rect -1133 959 -1075 965
rect -941 959 -883 965
rect -749 959 -691 965
rect -557 959 -499 965
rect -365 959 -307 965
rect -173 959 -115 965
rect 19 959 77 965
rect 211 959 269 965
rect 403 959 461 965
rect 595 959 653 965
rect 787 959 845 965
rect 979 959 1037 965
rect 1171 959 1229 965
rect 1363 959 1421 965
rect 1555 959 1613 965
rect 1747 959 1805 965
rect 1939 959 1997 965
rect 2131 959 2189 965
rect 2323 959 2381 965
rect 2515 959 2573 965
rect 2707 959 2765 965
rect 2899 959 2957 965
rect 3091 959 3149 965
rect 3283 959 3341 965
rect 3475 959 3533 965
rect 3667 959 3725 965
rect 3859 959 3917 965
rect 4051 959 4109 965
rect 4243 959 4301 965
rect 4435 959 4493 965
rect 4627 959 4685 965
rect -4685 589 -4627 595
rect -4493 589 -4435 595
rect -4301 589 -4243 595
rect -4109 589 -4051 595
rect -3917 589 -3859 595
rect -3725 589 -3667 595
rect -3533 589 -3475 595
rect -3341 589 -3283 595
rect -3149 589 -3091 595
rect -2957 589 -2899 595
rect -2765 589 -2707 595
rect -2573 589 -2515 595
rect -2381 589 -2323 595
rect -2189 589 -2131 595
rect -1997 589 -1939 595
rect -1805 589 -1747 595
rect -1613 589 -1555 595
rect -1421 589 -1363 595
rect -1229 589 -1171 595
rect -1037 589 -979 595
rect -845 589 -787 595
rect -653 589 -595 595
rect -461 589 -403 595
rect -269 589 -211 595
rect -77 589 -19 595
rect 115 589 173 595
rect 307 589 365 595
rect 499 589 557 595
rect 691 589 749 595
rect 883 589 941 595
rect 1075 589 1133 595
rect 1267 589 1325 595
rect 1459 589 1517 595
rect 1651 589 1709 595
rect 1843 589 1901 595
rect 2035 589 2093 595
rect 2227 589 2285 595
rect 2419 589 2477 595
rect 2611 589 2669 595
rect 2803 589 2861 595
rect 2995 589 3053 595
rect 3187 589 3245 595
rect 3379 589 3437 595
rect 3571 589 3629 595
rect 3763 589 3821 595
rect 3955 589 4013 595
rect 4147 589 4205 595
rect 4339 589 4397 595
rect 4531 589 4589 595
rect 4723 589 4781 595
rect -4685 555 -4673 589
rect -4493 555 -4481 589
rect -4301 555 -4289 589
rect -4109 555 -4097 589
rect -3917 555 -3905 589
rect -3725 555 -3713 589
rect -3533 555 -3521 589
rect -3341 555 -3329 589
rect -3149 555 -3137 589
rect -2957 555 -2945 589
rect -2765 555 -2753 589
rect -2573 555 -2561 589
rect -2381 555 -2369 589
rect -2189 555 -2177 589
rect -1997 555 -1985 589
rect -1805 555 -1793 589
rect -1613 555 -1601 589
rect -1421 555 -1409 589
rect -1229 555 -1217 589
rect -1037 555 -1025 589
rect -845 555 -833 589
rect -653 555 -641 589
rect -461 555 -449 589
rect -269 555 -257 589
rect -77 555 -65 589
rect 115 555 127 589
rect 307 555 319 589
rect 499 555 511 589
rect 691 555 703 589
rect 883 555 895 589
rect 1075 555 1087 589
rect 1267 555 1279 589
rect 1459 555 1471 589
rect 1651 555 1663 589
rect 1843 555 1855 589
rect 2035 555 2047 589
rect 2227 555 2239 589
rect 2419 555 2431 589
rect 2611 555 2623 589
rect 2803 555 2815 589
rect 2995 555 3007 589
rect 3187 555 3199 589
rect 3379 555 3391 589
rect 3571 555 3583 589
rect 3763 555 3775 589
rect 3955 555 3967 589
rect 4147 555 4159 589
rect 4339 555 4351 589
rect 4531 555 4543 589
rect 4723 555 4735 589
rect -4685 549 -4627 555
rect -4493 549 -4435 555
rect -4301 549 -4243 555
rect -4109 549 -4051 555
rect -3917 549 -3859 555
rect -3725 549 -3667 555
rect -3533 549 -3475 555
rect -3341 549 -3283 555
rect -3149 549 -3091 555
rect -2957 549 -2899 555
rect -2765 549 -2707 555
rect -2573 549 -2515 555
rect -2381 549 -2323 555
rect -2189 549 -2131 555
rect -1997 549 -1939 555
rect -1805 549 -1747 555
rect -1613 549 -1555 555
rect -1421 549 -1363 555
rect -1229 549 -1171 555
rect -1037 549 -979 555
rect -845 549 -787 555
rect -653 549 -595 555
rect -461 549 -403 555
rect -269 549 -211 555
rect -77 549 -19 555
rect 115 549 173 555
rect 307 549 365 555
rect 499 549 557 555
rect 691 549 749 555
rect 883 549 941 555
rect 1075 549 1133 555
rect 1267 549 1325 555
rect 1459 549 1517 555
rect 1651 549 1709 555
rect 1843 549 1901 555
rect 2035 549 2093 555
rect 2227 549 2285 555
rect 2419 549 2477 555
rect 2611 549 2669 555
rect 2803 549 2861 555
rect 2995 549 3053 555
rect 3187 549 3245 555
rect 3379 549 3437 555
rect 3571 549 3629 555
rect 3763 549 3821 555
rect 3955 549 4013 555
rect 4147 549 4205 555
rect 4339 549 4397 555
rect 4531 549 4589 555
rect 4723 549 4781 555
rect -4685 481 -4627 487
rect -4493 481 -4435 487
rect -4301 481 -4243 487
rect -4109 481 -4051 487
rect -3917 481 -3859 487
rect -3725 481 -3667 487
rect -3533 481 -3475 487
rect -3341 481 -3283 487
rect -3149 481 -3091 487
rect -2957 481 -2899 487
rect -2765 481 -2707 487
rect -2573 481 -2515 487
rect -2381 481 -2323 487
rect -2189 481 -2131 487
rect -1997 481 -1939 487
rect -1805 481 -1747 487
rect -1613 481 -1555 487
rect -1421 481 -1363 487
rect -1229 481 -1171 487
rect -1037 481 -979 487
rect -845 481 -787 487
rect -653 481 -595 487
rect -461 481 -403 487
rect -269 481 -211 487
rect -77 481 -19 487
rect 115 481 173 487
rect 307 481 365 487
rect 499 481 557 487
rect 691 481 749 487
rect 883 481 941 487
rect 1075 481 1133 487
rect 1267 481 1325 487
rect 1459 481 1517 487
rect 1651 481 1709 487
rect 1843 481 1901 487
rect 2035 481 2093 487
rect 2227 481 2285 487
rect 2419 481 2477 487
rect 2611 481 2669 487
rect 2803 481 2861 487
rect 2995 481 3053 487
rect 3187 481 3245 487
rect 3379 481 3437 487
rect 3571 481 3629 487
rect 3763 481 3821 487
rect 3955 481 4013 487
rect 4147 481 4205 487
rect 4339 481 4397 487
rect 4531 481 4589 487
rect 4723 481 4781 487
rect -4685 447 -4673 481
rect -4493 447 -4481 481
rect -4301 447 -4289 481
rect -4109 447 -4097 481
rect -3917 447 -3905 481
rect -3725 447 -3713 481
rect -3533 447 -3521 481
rect -3341 447 -3329 481
rect -3149 447 -3137 481
rect -2957 447 -2945 481
rect -2765 447 -2753 481
rect -2573 447 -2561 481
rect -2381 447 -2369 481
rect -2189 447 -2177 481
rect -1997 447 -1985 481
rect -1805 447 -1793 481
rect -1613 447 -1601 481
rect -1421 447 -1409 481
rect -1229 447 -1217 481
rect -1037 447 -1025 481
rect -845 447 -833 481
rect -653 447 -641 481
rect -461 447 -449 481
rect -269 447 -257 481
rect -77 447 -65 481
rect 115 447 127 481
rect 307 447 319 481
rect 499 447 511 481
rect 691 447 703 481
rect 883 447 895 481
rect 1075 447 1087 481
rect 1267 447 1279 481
rect 1459 447 1471 481
rect 1651 447 1663 481
rect 1843 447 1855 481
rect 2035 447 2047 481
rect 2227 447 2239 481
rect 2419 447 2431 481
rect 2611 447 2623 481
rect 2803 447 2815 481
rect 2995 447 3007 481
rect 3187 447 3199 481
rect 3379 447 3391 481
rect 3571 447 3583 481
rect 3763 447 3775 481
rect 3955 447 3967 481
rect 4147 447 4159 481
rect 4339 447 4351 481
rect 4531 447 4543 481
rect 4723 447 4735 481
rect -4685 441 -4627 447
rect -4493 441 -4435 447
rect -4301 441 -4243 447
rect -4109 441 -4051 447
rect -3917 441 -3859 447
rect -3725 441 -3667 447
rect -3533 441 -3475 447
rect -3341 441 -3283 447
rect -3149 441 -3091 447
rect -2957 441 -2899 447
rect -2765 441 -2707 447
rect -2573 441 -2515 447
rect -2381 441 -2323 447
rect -2189 441 -2131 447
rect -1997 441 -1939 447
rect -1805 441 -1747 447
rect -1613 441 -1555 447
rect -1421 441 -1363 447
rect -1229 441 -1171 447
rect -1037 441 -979 447
rect -845 441 -787 447
rect -653 441 -595 447
rect -461 441 -403 447
rect -269 441 -211 447
rect -77 441 -19 447
rect 115 441 173 447
rect 307 441 365 447
rect 499 441 557 447
rect 691 441 749 447
rect 883 441 941 447
rect 1075 441 1133 447
rect 1267 441 1325 447
rect 1459 441 1517 447
rect 1651 441 1709 447
rect 1843 441 1901 447
rect 2035 441 2093 447
rect 2227 441 2285 447
rect 2419 441 2477 447
rect 2611 441 2669 447
rect 2803 441 2861 447
rect 2995 441 3053 447
rect 3187 441 3245 447
rect 3379 441 3437 447
rect 3571 441 3629 447
rect 3763 441 3821 447
rect 3955 441 4013 447
rect 4147 441 4205 447
rect 4339 441 4397 447
rect 4531 441 4589 447
rect 4723 441 4781 447
rect -4781 71 -4723 77
rect -4589 71 -4531 77
rect -4397 71 -4339 77
rect -4205 71 -4147 77
rect -4013 71 -3955 77
rect -3821 71 -3763 77
rect -3629 71 -3571 77
rect -3437 71 -3379 77
rect -3245 71 -3187 77
rect -3053 71 -2995 77
rect -2861 71 -2803 77
rect -2669 71 -2611 77
rect -2477 71 -2419 77
rect -2285 71 -2227 77
rect -2093 71 -2035 77
rect -1901 71 -1843 77
rect -1709 71 -1651 77
rect -1517 71 -1459 77
rect -1325 71 -1267 77
rect -1133 71 -1075 77
rect -941 71 -883 77
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect 979 71 1037 77
rect 1171 71 1229 77
rect 1363 71 1421 77
rect 1555 71 1613 77
rect 1747 71 1805 77
rect 1939 71 1997 77
rect 2131 71 2189 77
rect 2323 71 2381 77
rect 2515 71 2573 77
rect 2707 71 2765 77
rect 2899 71 2957 77
rect 3091 71 3149 77
rect 3283 71 3341 77
rect 3475 71 3533 77
rect 3667 71 3725 77
rect 3859 71 3917 77
rect 4051 71 4109 77
rect 4243 71 4301 77
rect 4435 71 4493 77
rect 4627 71 4685 77
rect -4781 37 -4769 71
rect -4589 37 -4577 71
rect -4397 37 -4385 71
rect -4205 37 -4193 71
rect -4013 37 -4001 71
rect -3821 37 -3809 71
rect -3629 37 -3617 71
rect -3437 37 -3425 71
rect -3245 37 -3233 71
rect -3053 37 -3041 71
rect -2861 37 -2849 71
rect -2669 37 -2657 71
rect -2477 37 -2465 71
rect -2285 37 -2273 71
rect -2093 37 -2081 71
rect -1901 37 -1889 71
rect -1709 37 -1697 71
rect -1517 37 -1505 71
rect -1325 37 -1313 71
rect -1133 37 -1121 71
rect -941 37 -929 71
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect 979 37 991 71
rect 1171 37 1183 71
rect 1363 37 1375 71
rect 1555 37 1567 71
rect 1747 37 1759 71
rect 1939 37 1951 71
rect 2131 37 2143 71
rect 2323 37 2335 71
rect 2515 37 2527 71
rect 2707 37 2719 71
rect 2899 37 2911 71
rect 3091 37 3103 71
rect 3283 37 3295 71
rect 3475 37 3487 71
rect 3667 37 3679 71
rect 3859 37 3871 71
rect 4051 37 4063 71
rect 4243 37 4255 71
rect 4435 37 4447 71
rect 4627 37 4639 71
rect -4781 31 -4723 37
rect -4589 31 -4531 37
rect -4397 31 -4339 37
rect -4205 31 -4147 37
rect -4013 31 -3955 37
rect -3821 31 -3763 37
rect -3629 31 -3571 37
rect -3437 31 -3379 37
rect -3245 31 -3187 37
rect -3053 31 -2995 37
rect -2861 31 -2803 37
rect -2669 31 -2611 37
rect -2477 31 -2419 37
rect -2285 31 -2227 37
rect -2093 31 -2035 37
rect -1901 31 -1843 37
rect -1709 31 -1651 37
rect -1517 31 -1459 37
rect -1325 31 -1267 37
rect -1133 31 -1075 37
rect -941 31 -883 37
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect 979 31 1037 37
rect 1171 31 1229 37
rect 1363 31 1421 37
rect 1555 31 1613 37
rect 1747 31 1805 37
rect 1939 31 1997 37
rect 2131 31 2189 37
rect 2323 31 2381 37
rect 2515 31 2573 37
rect 2707 31 2765 37
rect 2899 31 2957 37
rect 3091 31 3149 37
rect 3283 31 3341 37
rect 3475 31 3533 37
rect 3667 31 3725 37
rect 3859 31 3917 37
rect 4051 31 4109 37
rect 4243 31 4301 37
rect 4435 31 4493 37
rect 4627 31 4685 37
rect -4781 -37 -4723 -31
rect -4589 -37 -4531 -31
rect -4397 -37 -4339 -31
rect -4205 -37 -4147 -31
rect -4013 -37 -3955 -31
rect -3821 -37 -3763 -31
rect -3629 -37 -3571 -31
rect -3437 -37 -3379 -31
rect -3245 -37 -3187 -31
rect -3053 -37 -2995 -31
rect -2861 -37 -2803 -31
rect -2669 -37 -2611 -31
rect -2477 -37 -2419 -31
rect -2285 -37 -2227 -31
rect -2093 -37 -2035 -31
rect -1901 -37 -1843 -31
rect -1709 -37 -1651 -31
rect -1517 -37 -1459 -31
rect -1325 -37 -1267 -31
rect -1133 -37 -1075 -31
rect -941 -37 -883 -31
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect 979 -37 1037 -31
rect 1171 -37 1229 -31
rect 1363 -37 1421 -31
rect 1555 -37 1613 -31
rect 1747 -37 1805 -31
rect 1939 -37 1997 -31
rect 2131 -37 2189 -31
rect 2323 -37 2381 -31
rect 2515 -37 2573 -31
rect 2707 -37 2765 -31
rect 2899 -37 2957 -31
rect 3091 -37 3149 -31
rect 3283 -37 3341 -31
rect 3475 -37 3533 -31
rect 3667 -37 3725 -31
rect 3859 -37 3917 -31
rect 4051 -37 4109 -31
rect 4243 -37 4301 -31
rect 4435 -37 4493 -31
rect 4627 -37 4685 -31
rect -4781 -71 -4769 -37
rect -4589 -71 -4577 -37
rect -4397 -71 -4385 -37
rect -4205 -71 -4193 -37
rect -4013 -71 -4001 -37
rect -3821 -71 -3809 -37
rect -3629 -71 -3617 -37
rect -3437 -71 -3425 -37
rect -3245 -71 -3233 -37
rect -3053 -71 -3041 -37
rect -2861 -71 -2849 -37
rect -2669 -71 -2657 -37
rect -2477 -71 -2465 -37
rect -2285 -71 -2273 -37
rect -2093 -71 -2081 -37
rect -1901 -71 -1889 -37
rect -1709 -71 -1697 -37
rect -1517 -71 -1505 -37
rect -1325 -71 -1313 -37
rect -1133 -71 -1121 -37
rect -941 -71 -929 -37
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect 979 -71 991 -37
rect 1171 -71 1183 -37
rect 1363 -71 1375 -37
rect 1555 -71 1567 -37
rect 1747 -71 1759 -37
rect 1939 -71 1951 -37
rect 2131 -71 2143 -37
rect 2323 -71 2335 -37
rect 2515 -71 2527 -37
rect 2707 -71 2719 -37
rect 2899 -71 2911 -37
rect 3091 -71 3103 -37
rect 3283 -71 3295 -37
rect 3475 -71 3487 -37
rect 3667 -71 3679 -37
rect 3859 -71 3871 -37
rect 4051 -71 4063 -37
rect 4243 -71 4255 -37
rect 4435 -71 4447 -37
rect 4627 -71 4639 -37
rect -4781 -77 -4723 -71
rect -4589 -77 -4531 -71
rect -4397 -77 -4339 -71
rect -4205 -77 -4147 -71
rect -4013 -77 -3955 -71
rect -3821 -77 -3763 -71
rect -3629 -77 -3571 -71
rect -3437 -77 -3379 -71
rect -3245 -77 -3187 -71
rect -3053 -77 -2995 -71
rect -2861 -77 -2803 -71
rect -2669 -77 -2611 -71
rect -2477 -77 -2419 -71
rect -2285 -77 -2227 -71
rect -2093 -77 -2035 -71
rect -1901 -77 -1843 -71
rect -1709 -77 -1651 -71
rect -1517 -77 -1459 -71
rect -1325 -77 -1267 -71
rect -1133 -77 -1075 -71
rect -941 -77 -883 -71
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect 979 -77 1037 -71
rect 1171 -77 1229 -71
rect 1363 -77 1421 -71
rect 1555 -77 1613 -71
rect 1747 -77 1805 -71
rect 1939 -77 1997 -71
rect 2131 -77 2189 -71
rect 2323 -77 2381 -71
rect 2515 -77 2573 -71
rect 2707 -77 2765 -71
rect 2899 -77 2957 -71
rect 3091 -77 3149 -71
rect 3283 -77 3341 -71
rect 3475 -77 3533 -71
rect 3667 -77 3725 -71
rect 3859 -77 3917 -71
rect 4051 -77 4109 -71
rect 4243 -77 4301 -71
rect 4435 -77 4493 -71
rect 4627 -77 4685 -71
rect -4685 -447 -4627 -441
rect -4493 -447 -4435 -441
rect -4301 -447 -4243 -441
rect -4109 -447 -4051 -441
rect -3917 -447 -3859 -441
rect -3725 -447 -3667 -441
rect -3533 -447 -3475 -441
rect -3341 -447 -3283 -441
rect -3149 -447 -3091 -441
rect -2957 -447 -2899 -441
rect -2765 -447 -2707 -441
rect -2573 -447 -2515 -441
rect -2381 -447 -2323 -441
rect -2189 -447 -2131 -441
rect -1997 -447 -1939 -441
rect -1805 -447 -1747 -441
rect -1613 -447 -1555 -441
rect -1421 -447 -1363 -441
rect -1229 -447 -1171 -441
rect -1037 -447 -979 -441
rect -845 -447 -787 -441
rect -653 -447 -595 -441
rect -461 -447 -403 -441
rect -269 -447 -211 -441
rect -77 -447 -19 -441
rect 115 -447 173 -441
rect 307 -447 365 -441
rect 499 -447 557 -441
rect 691 -447 749 -441
rect 883 -447 941 -441
rect 1075 -447 1133 -441
rect 1267 -447 1325 -441
rect 1459 -447 1517 -441
rect 1651 -447 1709 -441
rect 1843 -447 1901 -441
rect 2035 -447 2093 -441
rect 2227 -447 2285 -441
rect 2419 -447 2477 -441
rect 2611 -447 2669 -441
rect 2803 -447 2861 -441
rect 2995 -447 3053 -441
rect 3187 -447 3245 -441
rect 3379 -447 3437 -441
rect 3571 -447 3629 -441
rect 3763 -447 3821 -441
rect 3955 -447 4013 -441
rect 4147 -447 4205 -441
rect 4339 -447 4397 -441
rect 4531 -447 4589 -441
rect 4723 -447 4781 -441
rect -4685 -481 -4673 -447
rect -4493 -481 -4481 -447
rect -4301 -481 -4289 -447
rect -4109 -481 -4097 -447
rect -3917 -481 -3905 -447
rect -3725 -481 -3713 -447
rect -3533 -481 -3521 -447
rect -3341 -481 -3329 -447
rect -3149 -481 -3137 -447
rect -2957 -481 -2945 -447
rect -2765 -481 -2753 -447
rect -2573 -481 -2561 -447
rect -2381 -481 -2369 -447
rect -2189 -481 -2177 -447
rect -1997 -481 -1985 -447
rect -1805 -481 -1793 -447
rect -1613 -481 -1601 -447
rect -1421 -481 -1409 -447
rect -1229 -481 -1217 -447
rect -1037 -481 -1025 -447
rect -845 -481 -833 -447
rect -653 -481 -641 -447
rect -461 -481 -449 -447
rect -269 -481 -257 -447
rect -77 -481 -65 -447
rect 115 -481 127 -447
rect 307 -481 319 -447
rect 499 -481 511 -447
rect 691 -481 703 -447
rect 883 -481 895 -447
rect 1075 -481 1087 -447
rect 1267 -481 1279 -447
rect 1459 -481 1471 -447
rect 1651 -481 1663 -447
rect 1843 -481 1855 -447
rect 2035 -481 2047 -447
rect 2227 -481 2239 -447
rect 2419 -481 2431 -447
rect 2611 -481 2623 -447
rect 2803 -481 2815 -447
rect 2995 -481 3007 -447
rect 3187 -481 3199 -447
rect 3379 -481 3391 -447
rect 3571 -481 3583 -447
rect 3763 -481 3775 -447
rect 3955 -481 3967 -447
rect 4147 -481 4159 -447
rect 4339 -481 4351 -447
rect 4531 -481 4543 -447
rect 4723 -481 4735 -447
rect -4685 -487 -4627 -481
rect -4493 -487 -4435 -481
rect -4301 -487 -4243 -481
rect -4109 -487 -4051 -481
rect -3917 -487 -3859 -481
rect -3725 -487 -3667 -481
rect -3533 -487 -3475 -481
rect -3341 -487 -3283 -481
rect -3149 -487 -3091 -481
rect -2957 -487 -2899 -481
rect -2765 -487 -2707 -481
rect -2573 -487 -2515 -481
rect -2381 -487 -2323 -481
rect -2189 -487 -2131 -481
rect -1997 -487 -1939 -481
rect -1805 -487 -1747 -481
rect -1613 -487 -1555 -481
rect -1421 -487 -1363 -481
rect -1229 -487 -1171 -481
rect -1037 -487 -979 -481
rect -845 -487 -787 -481
rect -653 -487 -595 -481
rect -461 -487 -403 -481
rect -269 -487 -211 -481
rect -77 -487 -19 -481
rect 115 -487 173 -481
rect 307 -487 365 -481
rect 499 -487 557 -481
rect 691 -487 749 -481
rect 883 -487 941 -481
rect 1075 -487 1133 -481
rect 1267 -487 1325 -481
rect 1459 -487 1517 -481
rect 1651 -487 1709 -481
rect 1843 -487 1901 -481
rect 2035 -487 2093 -481
rect 2227 -487 2285 -481
rect 2419 -487 2477 -481
rect 2611 -487 2669 -481
rect 2803 -487 2861 -481
rect 2995 -487 3053 -481
rect 3187 -487 3245 -481
rect 3379 -487 3437 -481
rect 3571 -487 3629 -481
rect 3763 -487 3821 -481
rect 3955 -487 4013 -481
rect 4147 -487 4205 -481
rect 4339 -487 4397 -481
rect 4531 -487 4589 -481
rect 4723 -487 4781 -481
rect -4685 -555 -4627 -549
rect -4493 -555 -4435 -549
rect -4301 -555 -4243 -549
rect -4109 -555 -4051 -549
rect -3917 -555 -3859 -549
rect -3725 -555 -3667 -549
rect -3533 -555 -3475 -549
rect -3341 -555 -3283 -549
rect -3149 -555 -3091 -549
rect -2957 -555 -2899 -549
rect -2765 -555 -2707 -549
rect -2573 -555 -2515 -549
rect -2381 -555 -2323 -549
rect -2189 -555 -2131 -549
rect -1997 -555 -1939 -549
rect -1805 -555 -1747 -549
rect -1613 -555 -1555 -549
rect -1421 -555 -1363 -549
rect -1229 -555 -1171 -549
rect -1037 -555 -979 -549
rect -845 -555 -787 -549
rect -653 -555 -595 -549
rect -461 -555 -403 -549
rect -269 -555 -211 -549
rect -77 -555 -19 -549
rect 115 -555 173 -549
rect 307 -555 365 -549
rect 499 -555 557 -549
rect 691 -555 749 -549
rect 883 -555 941 -549
rect 1075 -555 1133 -549
rect 1267 -555 1325 -549
rect 1459 -555 1517 -549
rect 1651 -555 1709 -549
rect 1843 -555 1901 -549
rect 2035 -555 2093 -549
rect 2227 -555 2285 -549
rect 2419 -555 2477 -549
rect 2611 -555 2669 -549
rect 2803 -555 2861 -549
rect 2995 -555 3053 -549
rect 3187 -555 3245 -549
rect 3379 -555 3437 -549
rect 3571 -555 3629 -549
rect 3763 -555 3821 -549
rect 3955 -555 4013 -549
rect 4147 -555 4205 -549
rect 4339 -555 4397 -549
rect 4531 -555 4589 -549
rect 4723 -555 4781 -549
rect -4685 -589 -4673 -555
rect -4493 -589 -4481 -555
rect -4301 -589 -4289 -555
rect -4109 -589 -4097 -555
rect -3917 -589 -3905 -555
rect -3725 -589 -3713 -555
rect -3533 -589 -3521 -555
rect -3341 -589 -3329 -555
rect -3149 -589 -3137 -555
rect -2957 -589 -2945 -555
rect -2765 -589 -2753 -555
rect -2573 -589 -2561 -555
rect -2381 -589 -2369 -555
rect -2189 -589 -2177 -555
rect -1997 -589 -1985 -555
rect -1805 -589 -1793 -555
rect -1613 -589 -1601 -555
rect -1421 -589 -1409 -555
rect -1229 -589 -1217 -555
rect -1037 -589 -1025 -555
rect -845 -589 -833 -555
rect -653 -589 -641 -555
rect -461 -589 -449 -555
rect -269 -589 -257 -555
rect -77 -589 -65 -555
rect 115 -589 127 -555
rect 307 -589 319 -555
rect 499 -589 511 -555
rect 691 -589 703 -555
rect 883 -589 895 -555
rect 1075 -589 1087 -555
rect 1267 -589 1279 -555
rect 1459 -589 1471 -555
rect 1651 -589 1663 -555
rect 1843 -589 1855 -555
rect 2035 -589 2047 -555
rect 2227 -589 2239 -555
rect 2419 -589 2431 -555
rect 2611 -589 2623 -555
rect 2803 -589 2815 -555
rect 2995 -589 3007 -555
rect 3187 -589 3199 -555
rect 3379 -589 3391 -555
rect 3571 -589 3583 -555
rect 3763 -589 3775 -555
rect 3955 -589 3967 -555
rect 4147 -589 4159 -555
rect 4339 -589 4351 -555
rect 4531 -589 4543 -555
rect 4723 -589 4735 -555
rect -4685 -595 -4627 -589
rect -4493 -595 -4435 -589
rect -4301 -595 -4243 -589
rect -4109 -595 -4051 -589
rect -3917 -595 -3859 -589
rect -3725 -595 -3667 -589
rect -3533 -595 -3475 -589
rect -3341 -595 -3283 -589
rect -3149 -595 -3091 -589
rect -2957 -595 -2899 -589
rect -2765 -595 -2707 -589
rect -2573 -595 -2515 -589
rect -2381 -595 -2323 -589
rect -2189 -595 -2131 -589
rect -1997 -595 -1939 -589
rect -1805 -595 -1747 -589
rect -1613 -595 -1555 -589
rect -1421 -595 -1363 -589
rect -1229 -595 -1171 -589
rect -1037 -595 -979 -589
rect -845 -595 -787 -589
rect -653 -595 -595 -589
rect -461 -595 -403 -589
rect -269 -595 -211 -589
rect -77 -595 -19 -589
rect 115 -595 173 -589
rect 307 -595 365 -589
rect 499 -595 557 -589
rect 691 -595 749 -589
rect 883 -595 941 -589
rect 1075 -595 1133 -589
rect 1267 -595 1325 -589
rect 1459 -595 1517 -589
rect 1651 -595 1709 -589
rect 1843 -595 1901 -589
rect 2035 -595 2093 -589
rect 2227 -595 2285 -589
rect 2419 -595 2477 -589
rect 2611 -595 2669 -589
rect 2803 -595 2861 -589
rect 2995 -595 3053 -589
rect 3187 -595 3245 -589
rect 3379 -595 3437 -589
rect 3571 -595 3629 -589
rect 3763 -595 3821 -589
rect 3955 -595 4013 -589
rect 4147 -595 4205 -589
rect 4339 -595 4397 -589
rect 4531 -595 4589 -589
rect 4723 -595 4781 -589
rect -4781 -965 -4723 -959
rect -4589 -965 -4531 -959
rect -4397 -965 -4339 -959
rect -4205 -965 -4147 -959
rect -4013 -965 -3955 -959
rect -3821 -965 -3763 -959
rect -3629 -965 -3571 -959
rect -3437 -965 -3379 -959
rect -3245 -965 -3187 -959
rect -3053 -965 -2995 -959
rect -2861 -965 -2803 -959
rect -2669 -965 -2611 -959
rect -2477 -965 -2419 -959
rect -2285 -965 -2227 -959
rect -2093 -965 -2035 -959
rect -1901 -965 -1843 -959
rect -1709 -965 -1651 -959
rect -1517 -965 -1459 -959
rect -1325 -965 -1267 -959
rect -1133 -965 -1075 -959
rect -941 -965 -883 -959
rect -749 -965 -691 -959
rect -557 -965 -499 -959
rect -365 -965 -307 -959
rect -173 -965 -115 -959
rect 19 -965 77 -959
rect 211 -965 269 -959
rect 403 -965 461 -959
rect 595 -965 653 -959
rect 787 -965 845 -959
rect 979 -965 1037 -959
rect 1171 -965 1229 -959
rect 1363 -965 1421 -959
rect 1555 -965 1613 -959
rect 1747 -965 1805 -959
rect 1939 -965 1997 -959
rect 2131 -965 2189 -959
rect 2323 -965 2381 -959
rect 2515 -965 2573 -959
rect 2707 -965 2765 -959
rect 2899 -965 2957 -959
rect 3091 -965 3149 -959
rect 3283 -965 3341 -959
rect 3475 -965 3533 -959
rect 3667 -965 3725 -959
rect 3859 -965 3917 -959
rect 4051 -965 4109 -959
rect 4243 -965 4301 -959
rect 4435 -965 4493 -959
rect 4627 -965 4685 -959
rect -4781 -999 -4769 -965
rect -4589 -999 -4577 -965
rect -4397 -999 -4385 -965
rect -4205 -999 -4193 -965
rect -4013 -999 -4001 -965
rect -3821 -999 -3809 -965
rect -3629 -999 -3617 -965
rect -3437 -999 -3425 -965
rect -3245 -999 -3233 -965
rect -3053 -999 -3041 -965
rect -2861 -999 -2849 -965
rect -2669 -999 -2657 -965
rect -2477 -999 -2465 -965
rect -2285 -999 -2273 -965
rect -2093 -999 -2081 -965
rect -1901 -999 -1889 -965
rect -1709 -999 -1697 -965
rect -1517 -999 -1505 -965
rect -1325 -999 -1313 -965
rect -1133 -999 -1121 -965
rect -941 -999 -929 -965
rect -749 -999 -737 -965
rect -557 -999 -545 -965
rect -365 -999 -353 -965
rect -173 -999 -161 -965
rect 19 -999 31 -965
rect 211 -999 223 -965
rect 403 -999 415 -965
rect 595 -999 607 -965
rect 787 -999 799 -965
rect 979 -999 991 -965
rect 1171 -999 1183 -965
rect 1363 -999 1375 -965
rect 1555 -999 1567 -965
rect 1747 -999 1759 -965
rect 1939 -999 1951 -965
rect 2131 -999 2143 -965
rect 2323 -999 2335 -965
rect 2515 -999 2527 -965
rect 2707 -999 2719 -965
rect 2899 -999 2911 -965
rect 3091 -999 3103 -965
rect 3283 -999 3295 -965
rect 3475 -999 3487 -965
rect 3667 -999 3679 -965
rect 3859 -999 3871 -965
rect 4051 -999 4063 -965
rect 4243 -999 4255 -965
rect 4435 -999 4447 -965
rect 4627 -999 4639 -965
rect -4781 -1005 -4723 -999
rect -4589 -1005 -4531 -999
rect -4397 -1005 -4339 -999
rect -4205 -1005 -4147 -999
rect -4013 -1005 -3955 -999
rect -3821 -1005 -3763 -999
rect -3629 -1005 -3571 -999
rect -3437 -1005 -3379 -999
rect -3245 -1005 -3187 -999
rect -3053 -1005 -2995 -999
rect -2861 -1005 -2803 -999
rect -2669 -1005 -2611 -999
rect -2477 -1005 -2419 -999
rect -2285 -1005 -2227 -999
rect -2093 -1005 -2035 -999
rect -1901 -1005 -1843 -999
rect -1709 -1005 -1651 -999
rect -1517 -1005 -1459 -999
rect -1325 -1005 -1267 -999
rect -1133 -1005 -1075 -999
rect -941 -1005 -883 -999
rect -749 -1005 -691 -999
rect -557 -1005 -499 -999
rect -365 -1005 -307 -999
rect -173 -1005 -115 -999
rect 19 -1005 77 -999
rect 211 -1005 269 -999
rect 403 -1005 461 -999
rect 595 -1005 653 -999
rect 787 -1005 845 -999
rect 979 -1005 1037 -999
rect 1171 -1005 1229 -999
rect 1363 -1005 1421 -999
rect 1555 -1005 1613 -999
rect 1747 -1005 1805 -999
rect 1939 -1005 1997 -999
rect 2131 -1005 2189 -999
rect 2323 -1005 2381 -999
rect 2515 -1005 2573 -999
rect 2707 -1005 2765 -999
rect 2899 -1005 2957 -999
rect 3091 -1005 3149 -999
rect 3283 -1005 3341 -999
rect 3475 -1005 3533 -999
rect 3667 -1005 3725 -999
rect 3859 -1005 3917 -999
rect 4051 -1005 4109 -999
rect 4243 -1005 4301 -999
rect 4435 -1005 4493 -999
rect 4627 -1005 4685 -999
<< pwell >>
rect -4967 -1137 4967 1137
<< nmos >>
rect -4767 627 -4737 927
rect -4671 627 -4641 927
rect -4575 627 -4545 927
rect -4479 627 -4449 927
rect -4383 627 -4353 927
rect -4287 627 -4257 927
rect -4191 627 -4161 927
rect -4095 627 -4065 927
rect -3999 627 -3969 927
rect -3903 627 -3873 927
rect -3807 627 -3777 927
rect -3711 627 -3681 927
rect -3615 627 -3585 927
rect -3519 627 -3489 927
rect -3423 627 -3393 927
rect -3327 627 -3297 927
rect -3231 627 -3201 927
rect -3135 627 -3105 927
rect -3039 627 -3009 927
rect -2943 627 -2913 927
rect -2847 627 -2817 927
rect -2751 627 -2721 927
rect -2655 627 -2625 927
rect -2559 627 -2529 927
rect -2463 627 -2433 927
rect -2367 627 -2337 927
rect -2271 627 -2241 927
rect -2175 627 -2145 927
rect -2079 627 -2049 927
rect -1983 627 -1953 927
rect -1887 627 -1857 927
rect -1791 627 -1761 927
rect -1695 627 -1665 927
rect -1599 627 -1569 927
rect -1503 627 -1473 927
rect -1407 627 -1377 927
rect -1311 627 -1281 927
rect -1215 627 -1185 927
rect -1119 627 -1089 927
rect -1023 627 -993 927
rect -927 627 -897 927
rect -831 627 -801 927
rect -735 627 -705 927
rect -639 627 -609 927
rect -543 627 -513 927
rect -447 627 -417 927
rect -351 627 -321 927
rect -255 627 -225 927
rect -159 627 -129 927
rect -63 627 -33 927
rect 33 627 63 927
rect 129 627 159 927
rect 225 627 255 927
rect 321 627 351 927
rect 417 627 447 927
rect 513 627 543 927
rect 609 627 639 927
rect 705 627 735 927
rect 801 627 831 927
rect 897 627 927 927
rect 993 627 1023 927
rect 1089 627 1119 927
rect 1185 627 1215 927
rect 1281 627 1311 927
rect 1377 627 1407 927
rect 1473 627 1503 927
rect 1569 627 1599 927
rect 1665 627 1695 927
rect 1761 627 1791 927
rect 1857 627 1887 927
rect 1953 627 1983 927
rect 2049 627 2079 927
rect 2145 627 2175 927
rect 2241 627 2271 927
rect 2337 627 2367 927
rect 2433 627 2463 927
rect 2529 627 2559 927
rect 2625 627 2655 927
rect 2721 627 2751 927
rect 2817 627 2847 927
rect 2913 627 2943 927
rect 3009 627 3039 927
rect 3105 627 3135 927
rect 3201 627 3231 927
rect 3297 627 3327 927
rect 3393 627 3423 927
rect 3489 627 3519 927
rect 3585 627 3615 927
rect 3681 627 3711 927
rect 3777 627 3807 927
rect 3873 627 3903 927
rect 3969 627 3999 927
rect 4065 627 4095 927
rect 4161 627 4191 927
rect 4257 627 4287 927
rect 4353 627 4383 927
rect 4449 627 4479 927
rect 4545 627 4575 927
rect 4641 627 4671 927
rect 4737 627 4767 927
rect -4767 109 -4737 409
rect -4671 109 -4641 409
rect -4575 109 -4545 409
rect -4479 109 -4449 409
rect -4383 109 -4353 409
rect -4287 109 -4257 409
rect -4191 109 -4161 409
rect -4095 109 -4065 409
rect -3999 109 -3969 409
rect -3903 109 -3873 409
rect -3807 109 -3777 409
rect -3711 109 -3681 409
rect -3615 109 -3585 409
rect -3519 109 -3489 409
rect -3423 109 -3393 409
rect -3327 109 -3297 409
rect -3231 109 -3201 409
rect -3135 109 -3105 409
rect -3039 109 -3009 409
rect -2943 109 -2913 409
rect -2847 109 -2817 409
rect -2751 109 -2721 409
rect -2655 109 -2625 409
rect -2559 109 -2529 409
rect -2463 109 -2433 409
rect -2367 109 -2337 409
rect -2271 109 -2241 409
rect -2175 109 -2145 409
rect -2079 109 -2049 409
rect -1983 109 -1953 409
rect -1887 109 -1857 409
rect -1791 109 -1761 409
rect -1695 109 -1665 409
rect -1599 109 -1569 409
rect -1503 109 -1473 409
rect -1407 109 -1377 409
rect -1311 109 -1281 409
rect -1215 109 -1185 409
rect -1119 109 -1089 409
rect -1023 109 -993 409
rect -927 109 -897 409
rect -831 109 -801 409
rect -735 109 -705 409
rect -639 109 -609 409
rect -543 109 -513 409
rect -447 109 -417 409
rect -351 109 -321 409
rect -255 109 -225 409
rect -159 109 -129 409
rect -63 109 -33 409
rect 33 109 63 409
rect 129 109 159 409
rect 225 109 255 409
rect 321 109 351 409
rect 417 109 447 409
rect 513 109 543 409
rect 609 109 639 409
rect 705 109 735 409
rect 801 109 831 409
rect 897 109 927 409
rect 993 109 1023 409
rect 1089 109 1119 409
rect 1185 109 1215 409
rect 1281 109 1311 409
rect 1377 109 1407 409
rect 1473 109 1503 409
rect 1569 109 1599 409
rect 1665 109 1695 409
rect 1761 109 1791 409
rect 1857 109 1887 409
rect 1953 109 1983 409
rect 2049 109 2079 409
rect 2145 109 2175 409
rect 2241 109 2271 409
rect 2337 109 2367 409
rect 2433 109 2463 409
rect 2529 109 2559 409
rect 2625 109 2655 409
rect 2721 109 2751 409
rect 2817 109 2847 409
rect 2913 109 2943 409
rect 3009 109 3039 409
rect 3105 109 3135 409
rect 3201 109 3231 409
rect 3297 109 3327 409
rect 3393 109 3423 409
rect 3489 109 3519 409
rect 3585 109 3615 409
rect 3681 109 3711 409
rect 3777 109 3807 409
rect 3873 109 3903 409
rect 3969 109 3999 409
rect 4065 109 4095 409
rect 4161 109 4191 409
rect 4257 109 4287 409
rect 4353 109 4383 409
rect 4449 109 4479 409
rect 4545 109 4575 409
rect 4641 109 4671 409
rect 4737 109 4767 409
rect -4767 -409 -4737 -109
rect -4671 -409 -4641 -109
rect -4575 -409 -4545 -109
rect -4479 -409 -4449 -109
rect -4383 -409 -4353 -109
rect -4287 -409 -4257 -109
rect -4191 -409 -4161 -109
rect -4095 -409 -4065 -109
rect -3999 -409 -3969 -109
rect -3903 -409 -3873 -109
rect -3807 -409 -3777 -109
rect -3711 -409 -3681 -109
rect -3615 -409 -3585 -109
rect -3519 -409 -3489 -109
rect -3423 -409 -3393 -109
rect -3327 -409 -3297 -109
rect -3231 -409 -3201 -109
rect -3135 -409 -3105 -109
rect -3039 -409 -3009 -109
rect -2943 -409 -2913 -109
rect -2847 -409 -2817 -109
rect -2751 -409 -2721 -109
rect -2655 -409 -2625 -109
rect -2559 -409 -2529 -109
rect -2463 -409 -2433 -109
rect -2367 -409 -2337 -109
rect -2271 -409 -2241 -109
rect -2175 -409 -2145 -109
rect -2079 -409 -2049 -109
rect -1983 -409 -1953 -109
rect -1887 -409 -1857 -109
rect -1791 -409 -1761 -109
rect -1695 -409 -1665 -109
rect -1599 -409 -1569 -109
rect -1503 -409 -1473 -109
rect -1407 -409 -1377 -109
rect -1311 -409 -1281 -109
rect -1215 -409 -1185 -109
rect -1119 -409 -1089 -109
rect -1023 -409 -993 -109
rect -927 -409 -897 -109
rect -831 -409 -801 -109
rect -735 -409 -705 -109
rect -639 -409 -609 -109
rect -543 -409 -513 -109
rect -447 -409 -417 -109
rect -351 -409 -321 -109
rect -255 -409 -225 -109
rect -159 -409 -129 -109
rect -63 -409 -33 -109
rect 33 -409 63 -109
rect 129 -409 159 -109
rect 225 -409 255 -109
rect 321 -409 351 -109
rect 417 -409 447 -109
rect 513 -409 543 -109
rect 609 -409 639 -109
rect 705 -409 735 -109
rect 801 -409 831 -109
rect 897 -409 927 -109
rect 993 -409 1023 -109
rect 1089 -409 1119 -109
rect 1185 -409 1215 -109
rect 1281 -409 1311 -109
rect 1377 -409 1407 -109
rect 1473 -409 1503 -109
rect 1569 -409 1599 -109
rect 1665 -409 1695 -109
rect 1761 -409 1791 -109
rect 1857 -409 1887 -109
rect 1953 -409 1983 -109
rect 2049 -409 2079 -109
rect 2145 -409 2175 -109
rect 2241 -409 2271 -109
rect 2337 -409 2367 -109
rect 2433 -409 2463 -109
rect 2529 -409 2559 -109
rect 2625 -409 2655 -109
rect 2721 -409 2751 -109
rect 2817 -409 2847 -109
rect 2913 -409 2943 -109
rect 3009 -409 3039 -109
rect 3105 -409 3135 -109
rect 3201 -409 3231 -109
rect 3297 -409 3327 -109
rect 3393 -409 3423 -109
rect 3489 -409 3519 -109
rect 3585 -409 3615 -109
rect 3681 -409 3711 -109
rect 3777 -409 3807 -109
rect 3873 -409 3903 -109
rect 3969 -409 3999 -109
rect 4065 -409 4095 -109
rect 4161 -409 4191 -109
rect 4257 -409 4287 -109
rect 4353 -409 4383 -109
rect 4449 -409 4479 -109
rect 4545 -409 4575 -109
rect 4641 -409 4671 -109
rect 4737 -409 4767 -109
rect -4767 -927 -4737 -627
rect -4671 -927 -4641 -627
rect -4575 -927 -4545 -627
rect -4479 -927 -4449 -627
rect -4383 -927 -4353 -627
rect -4287 -927 -4257 -627
rect -4191 -927 -4161 -627
rect -4095 -927 -4065 -627
rect -3999 -927 -3969 -627
rect -3903 -927 -3873 -627
rect -3807 -927 -3777 -627
rect -3711 -927 -3681 -627
rect -3615 -927 -3585 -627
rect -3519 -927 -3489 -627
rect -3423 -927 -3393 -627
rect -3327 -927 -3297 -627
rect -3231 -927 -3201 -627
rect -3135 -927 -3105 -627
rect -3039 -927 -3009 -627
rect -2943 -927 -2913 -627
rect -2847 -927 -2817 -627
rect -2751 -927 -2721 -627
rect -2655 -927 -2625 -627
rect -2559 -927 -2529 -627
rect -2463 -927 -2433 -627
rect -2367 -927 -2337 -627
rect -2271 -927 -2241 -627
rect -2175 -927 -2145 -627
rect -2079 -927 -2049 -627
rect -1983 -927 -1953 -627
rect -1887 -927 -1857 -627
rect -1791 -927 -1761 -627
rect -1695 -927 -1665 -627
rect -1599 -927 -1569 -627
rect -1503 -927 -1473 -627
rect -1407 -927 -1377 -627
rect -1311 -927 -1281 -627
rect -1215 -927 -1185 -627
rect -1119 -927 -1089 -627
rect -1023 -927 -993 -627
rect -927 -927 -897 -627
rect -831 -927 -801 -627
rect -735 -927 -705 -627
rect -639 -927 -609 -627
rect -543 -927 -513 -627
rect -447 -927 -417 -627
rect -351 -927 -321 -627
rect -255 -927 -225 -627
rect -159 -927 -129 -627
rect -63 -927 -33 -627
rect 33 -927 63 -627
rect 129 -927 159 -627
rect 225 -927 255 -627
rect 321 -927 351 -627
rect 417 -927 447 -627
rect 513 -927 543 -627
rect 609 -927 639 -627
rect 705 -927 735 -627
rect 801 -927 831 -627
rect 897 -927 927 -627
rect 993 -927 1023 -627
rect 1089 -927 1119 -627
rect 1185 -927 1215 -627
rect 1281 -927 1311 -627
rect 1377 -927 1407 -627
rect 1473 -927 1503 -627
rect 1569 -927 1599 -627
rect 1665 -927 1695 -627
rect 1761 -927 1791 -627
rect 1857 -927 1887 -627
rect 1953 -927 1983 -627
rect 2049 -927 2079 -627
rect 2145 -927 2175 -627
rect 2241 -927 2271 -627
rect 2337 -927 2367 -627
rect 2433 -927 2463 -627
rect 2529 -927 2559 -627
rect 2625 -927 2655 -627
rect 2721 -927 2751 -627
rect 2817 -927 2847 -627
rect 2913 -927 2943 -627
rect 3009 -927 3039 -627
rect 3105 -927 3135 -627
rect 3201 -927 3231 -627
rect 3297 -927 3327 -627
rect 3393 -927 3423 -627
rect 3489 -927 3519 -627
rect 3585 -927 3615 -627
rect 3681 -927 3711 -627
rect 3777 -927 3807 -627
rect 3873 -927 3903 -627
rect 3969 -927 3999 -627
rect 4065 -927 4095 -627
rect 4161 -927 4191 -627
rect 4257 -927 4287 -627
rect 4353 -927 4383 -627
rect 4449 -927 4479 -627
rect 4545 -927 4575 -627
rect 4641 -927 4671 -627
rect 4737 -927 4767 -627
<< ndiff >>
rect -4829 915 -4767 927
rect -4829 639 -4817 915
rect -4783 639 -4767 915
rect -4829 627 -4767 639
rect -4737 915 -4671 927
rect -4737 639 -4721 915
rect -4687 639 -4671 915
rect -4737 627 -4671 639
rect -4641 915 -4575 927
rect -4641 639 -4625 915
rect -4591 639 -4575 915
rect -4641 627 -4575 639
rect -4545 915 -4479 927
rect -4545 639 -4529 915
rect -4495 639 -4479 915
rect -4545 627 -4479 639
rect -4449 915 -4383 927
rect -4449 639 -4433 915
rect -4399 639 -4383 915
rect -4449 627 -4383 639
rect -4353 915 -4287 927
rect -4353 639 -4337 915
rect -4303 639 -4287 915
rect -4353 627 -4287 639
rect -4257 915 -4191 927
rect -4257 639 -4241 915
rect -4207 639 -4191 915
rect -4257 627 -4191 639
rect -4161 915 -4095 927
rect -4161 639 -4145 915
rect -4111 639 -4095 915
rect -4161 627 -4095 639
rect -4065 915 -3999 927
rect -4065 639 -4049 915
rect -4015 639 -3999 915
rect -4065 627 -3999 639
rect -3969 915 -3903 927
rect -3969 639 -3953 915
rect -3919 639 -3903 915
rect -3969 627 -3903 639
rect -3873 915 -3807 927
rect -3873 639 -3857 915
rect -3823 639 -3807 915
rect -3873 627 -3807 639
rect -3777 915 -3711 927
rect -3777 639 -3761 915
rect -3727 639 -3711 915
rect -3777 627 -3711 639
rect -3681 915 -3615 927
rect -3681 639 -3665 915
rect -3631 639 -3615 915
rect -3681 627 -3615 639
rect -3585 915 -3519 927
rect -3585 639 -3569 915
rect -3535 639 -3519 915
rect -3585 627 -3519 639
rect -3489 915 -3423 927
rect -3489 639 -3473 915
rect -3439 639 -3423 915
rect -3489 627 -3423 639
rect -3393 915 -3327 927
rect -3393 639 -3377 915
rect -3343 639 -3327 915
rect -3393 627 -3327 639
rect -3297 915 -3231 927
rect -3297 639 -3281 915
rect -3247 639 -3231 915
rect -3297 627 -3231 639
rect -3201 915 -3135 927
rect -3201 639 -3185 915
rect -3151 639 -3135 915
rect -3201 627 -3135 639
rect -3105 915 -3039 927
rect -3105 639 -3089 915
rect -3055 639 -3039 915
rect -3105 627 -3039 639
rect -3009 915 -2943 927
rect -3009 639 -2993 915
rect -2959 639 -2943 915
rect -3009 627 -2943 639
rect -2913 915 -2847 927
rect -2913 639 -2897 915
rect -2863 639 -2847 915
rect -2913 627 -2847 639
rect -2817 915 -2751 927
rect -2817 639 -2801 915
rect -2767 639 -2751 915
rect -2817 627 -2751 639
rect -2721 915 -2655 927
rect -2721 639 -2705 915
rect -2671 639 -2655 915
rect -2721 627 -2655 639
rect -2625 915 -2559 927
rect -2625 639 -2609 915
rect -2575 639 -2559 915
rect -2625 627 -2559 639
rect -2529 915 -2463 927
rect -2529 639 -2513 915
rect -2479 639 -2463 915
rect -2529 627 -2463 639
rect -2433 915 -2367 927
rect -2433 639 -2417 915
rect -2383 639 -2367 915
rect -2433 627 -2367 639
rect -2337 915 -2271 927
rect -2337 639 -2321 915
rect -2287 639 -2271 915
rect -2337 627 -2271 639
rect -2241 915 -2175 927
rect -2241 639 -2225 915
rect -2191 639 -2175 915
rect -2241 627 -2175 639
rect -2145 915 -2079 927
rect -2145 639 -2129 915
rect -2095 639 -2079 915
rect -2145 627 -2079 639
rect -2049 915 -1983 927
rect -2049 639 -2033 915
rect -1999 639 -1983 915
rect -2049 627 -1983 639
rect -1953 915 -1887 927
rect -1953 639 -1937 915
rect -1903 639 -1887 915
rect -1953 627 -1887 639
rect -1857 915 -1791 927
rect -1857 639 -1841 915
rect -1807 639 -1791 915
rect -1857 627 -1791 639
rect -1761 915 -1695 927
rect -1761 639 -1745 915
rect -1711 639 -1695 915
rect -1761 627 -1695 639
rect -1665 915 -1599 927
rect -1665 639 -1649 915
rect -1615 639 -1599 915
rect -1665 627 -1599 639
rect -1569 915 -1503 927
rect -1569 639 -1553 915
rect -1519 639 -1503 915
rect -1569 627 -1503 639
rect -1473 915 -1407 927
rect -1473 639 -1457 915
rect -1423 639 -1407 915
rect -1473 627 -1407 639
rect -1377 915 -1311 927
rect -1377 639 -1361 915
rect -1327 639 -1311 915
rect -1377 627 -1311 639
rect -1281 915 -1215 927
rect -1281 639 -1265 915
rect -1231 639 -1215 915
rect -1281 627 -1215 639
rect -1185 915 -1119 927
rect -1185 639 -1169 915
rect -1135 639 -1119 915
rect -1185 627 -1119 639
rect -1089 915 -1023 927
rect -1089 639 -1073 915
rect -1039 639 -1023 915
rect -1089 627 -1023 639
rect -993 915 -927 927
rect -993 639 -977 915
rect -943 639 -927 915
rect -993 627 -927 639
rect -897 915 -831 927
rect -897 639 -881 915
rect -847 639 -831 915
rect -897 627 -831 639
rect -801 915 -735 927
rect -801 639 -785 915
rect -751 639 -735 915
rect -801 627 -735 639
rect -705 915 -639 927
rect -705 639 -689 915
rect -655 639 -639 915
rect -705 627 -639 639
rect -609 915 -543 927
rect -609 639 -593 915
rect -559 639 -543 915
rect -609 627 -543 639
rect -513 915 -447 927
rect -513 639 -497 915
rect -463 639 -447 915
rect -513 627 -447 639
rect -417 915 -351 927
rect -417 639 -401 915
rect -367 639 -351 915
rect -417 627 -351 639
rect -321 915 -255 927
rect -321 639 -305 915
rect -271 639 -255 915
rect -321 627 -255 639
rect -225 915 -159 927
rect -225 639 -209 915
rect -175 639 -159 915
rect -225 627 -159 639
rect -129 915 -63 927
rect -129 639 -113 915
rect -79 639 -63 915
rect -129 627 -63 639
rect -33 915 33 927
rect -33 639 -17 915
rect 17 639 33 915
rect -33 627 33 639
rect 63 915 129 927
rect 63 639 79 915
rect 113 639 129 915
rect 63 627 129 639
rect 159 915 225 927
rect 159 639 175 915
rect 209 639 225 915
rect 159 627 225 639
rect 255 915 321 927
rect 255 639 271 915
rect 305 639 321 915
rect 255 627 321 639
rect 351 915 417 927
rect 351 639 367 915
rect 401 639 417 915
rect 351 627 417 639
rect 447 915 513 927
rect 447 639 463 915
rect 497 639 513 915
rect 447 627 513 639
rect 543 915 609 927
rect 543 639 559 915
rect 593 639 609 915
rect 543 627 609 639
rect 639 915 705 927
rect 639 639 655 915
rect 689 639 705 915
rect 639 627 705 639
rect 735 915 801 927
rect 735 639 751 915
rect 785 639 801 915
rect 735 627 801 639
rect 831 915 897 927
rect 831 639 847 915
rect 881 639 897 915
rect 831 627 897 639
rect 927 915 993 927
rect 927 639 943 915
rect 977 639 993 915
rect 927 627 993 639
rect 1023 915 1089 927
rect 1023 639 1039 915
rect 1073 639 1089 915
rect 1023 627 1089 639
rect 1119 915 1185 927
rect 1119 639 1135 915
rect 1169 639 1185 915
rect 1119 627 1185 639
rect 1215 915 1281 927
rect 1215 639 1231 915
rect 1265 639 1281 915
rect 1215 627 1281 639
rect 1311 915 1377 927
rect 1311 639 1327 915
rect 1361 639 1377 915
rect 1311 627 1377 639
rect 1407 915 1473 927
rect 1407 639 1423 915
rect 1457 639 1473 915
rect 1407 627 1473 639
rect 1503 915 1569 927
rect 1503 639 1519 915
rect 1553 639 1569 915
rect 1503 627 1569 639
rect 1599 915 1665 927
rect 1599 639 1615 915
rect 1649 639 1665 915
rect 1599 627 1665 639
rect 1695 915 1761 927
rect 1695 639 1711 915
rect 1745 639 1761 915
rect 1695 627 1761 639
rect 1791 915 1857 927
rect 1791 639 1807 915
rect 1841 639 1857 915
rect 1791 627 1857 639
rect 1887 915 1953 927
rect 1887 639 1903 915
rect 1937 639 1953 915
rect 1887 627 1953 639
rect 1983 915 2049 927
rect 1983 639 1999 915
rect 2033 639 2049 915
rect 1983 627 2049 639
rect 2079 915 2145 927
rect 2079 639 2095 915
rect 2129 639 2145 915
rect 2079 627 2145 639
rect 2175 915 2241 927
rect 2175 639 2191 915
rect 2225 639 2241 915
rect 2175 627 2241 639
rect 2271 915 2337 927
rect 2271 639 2287 915
rect 2321 639 2337 915
rect 2271 627 2337 639
rect 2367 915 2433 927
rect 2367 639 2383 915
rect 2417 639 2433 915
rect 2367 627 2433 639
rect 2463 915 2529 927
rect 2463 639 2479 915
rect 2513 639 2529 915
rect 2463 627 2529 639
rect 2559 915 2625 927
rect 2559 639 2575 915
rect 2609 639 2625 915
rect 2559 627 2625 639
rect 2655 915 2721 927
rect 2655 639 2671 915
rect 2705 639 2721 915
rect 2655 627 2721 639
rect 2751 915 2817 927
rect 2751 639 2767 915
rect 2801 639 2817 915
rect 2751 627 2817 639
rect 2847 915 2913 927
rect 2847 639 2863 915
rect 2897 639 2913 915
rect 2847 627 2913 639
rect 2943 915 3009 927
rect 2943 639 2959 915
rect 2993 639 3009 915
rect 2943 627 3009 639
rect 3039 915 3105 927
rect 3039 639 3055 915
rect 3089 639 3105 915
rect 3039 627 3105 639
rect 3135 915 3201 927
rect 3135 639 3151 915
rect 3185 639 3201 915
rect 3135 627 3201 639
rect 3231 915 3297 927
rect 3231 639 3247 915
rect 3281 639 3297 915
rect 3231 627 3297 639
rect 3327 915 3393 927
rect 3327 639 3343 915
rect 3377 639 3393 915
rect 3327 627 3393 639
rect 3423 915 3489 927
rect 3423 639 3439 915
rect 3473 639 3489 915
rect 3423 627 3489 639
rect 3519 915 3585 927
rect 3519 639 3535 915
rect 3569 639 3585 915
rect 3519 627 3585 639
rect 3615 915 3681 927
rect 3615 639 3631 915
rect 3665 639 3681 915
rect 3615 627 3681 639
rect 3711 915 3777 927
rect 3711 639 3727 915
rect 3761 639 3777 915
rect 3711 627 3777 639
rect 3807 915 3873 927
rect 3807 639 3823 915
rect 3857 639 3873 915
rect 3807 627 3873 639
rect 3903 915 3969 927
rect 3903 639 3919 915
rect 3953 639 3969 915
rect 3903 627 3969 639
rect 3999 915 4065 927
rect 3999 639 4015 915
rect 4049 639 4065 915
rect 3999 627 4065 639
rect 4095 915 4161 927
rect 4095 639 4111 915
rect 4145 639 4161 915
rect 4095 627 4161 639
rect 4191 915 4257 927
rect 4191 639 4207 915
rect 4241 639 4257 915
rect 4191 627 4257 639
rect 4287 915 4353 927
rect 4287 639 4303 915
rect 4337 639 4353 915
rect 4287 627 4353 639
rect 4383 915 4449 927
rect 4383 639 4399 915
rect 4433 639 4449 915
rect 4383 627 4449 639
rect 4479 915 4545 927
rect 4479 639 4495 915
rect 4529 639 4545 915
rect 4479 627 4545 639
rect 4575 915 4641 927
rect 4575 639 4591 915
rect 4625 639 4641 915
rect 4575 627 4641 639
rect 4671 915 4737 927
rect 4671 639 4687 915
rect 4721 639 4737 915
rect 4671 627 4737 639
rect 4767 915 4829 927
rect 4767 639 4783 915
rect 4817 639 4829 915
rect 4767 627 4829 639
rect -4829 397 -4767 409
rect -4829 121 -4817 397
rect -4783 121 -4767 397
rect -4829 109 -4767 121
rect -4737 397 -4671 409
rect -4737 121 -4721 397
rect -4687 121 -4671 397
rect -4737 109 -4671 121
rect -4641 397 -4575 409
rect -4641 121 -4625 397
rect -4591 121 -4575 397
rect -4641 109 -4575 121
rect -4545 397 -4479 409
rect -4545 121 -4529 397
rect -4495 121 -4479 397
rect -4545 109 -4479 121
rect -4449 397 -4383 409
rect -4449 121 -4433 397
rect -4399 121 -4383 397
rect -4449 109 -4383 121
rect -4353 397 -4287 409
rect -4353 121 -4337 397
rect -4303 121 -4287 397
rect -4353 109 -4287 121
rect -4257 397 -4191 409
rect -4257 121 -4241 397
rect -4207 121 -4191 397
rect -4257 109 -4191 121
rect -4161 397 -4095 409
rect -4161 121 -4145 397
rect -4111 121 -4095 397
rect -4161 109 -4095 121
rect -4065 397 -3999 409
rect -4065 121 -4049 397
rect -4015 121 -3999 397
rect -4065 109 -3999 121
rect -3969 397 -3903 409
rect -3969 121 -3953 397
rect -3919 121 -3903 397
rect -3969 109 -3903 121
rect -3873 397 -3807 409
rect -3873 121 -3857 397
rect -3823 121 -3807 397
rect -3873 109 -3807 121
rect -3777 397 -3711 409
rect -3777 121 -3761 397
rect -3727 121 -3711 397
rect -3777 109 -3711 121
rect -3681 397 -3615 409
rect -3681 121 -3665 397
rect -3631 121 -3615 397
rect -3681 109 -3615 121
rect -3585 397 -3519 409
rect -3585 121 -3569 397
rect -3535 121 -3519 397
rect -3585 109 -3519 121
rect -3489 397 -3423 409
rect -3489 121 -3473 397
rect -3439 121 -3423 397
rect -3489 109 -3423 121
rect -3393 397 -3327 409
rect -3393 121 -3377 397
rect -3343 121 -3327 397
rect -3393 109 -3327 121
rect -3297 397 -3231 409
rect -3297 121 -3281 397
rect -3247 121 -3231 397
rect -3297 109 -3231 121
rect -3201 397 -3135 409
rect -3201 121 -3185 397
rect -3151 121 -3135 397
rect -3201 109 -3135 121
rect -3105 397 -3039 409
rect -3105 121 -3089 397
rect -3055 121 -3039 397
rect -3105 109 -3039 121
rect -3009 397 -2943 409
rect -3009 121 -2993 397
rect -2959 121 -2943 397
rect -3009 109 -2943 121
rect -2913 397 -2847 409
rect -2913 121 -2897 397
rect -2863 121 -2847 397
rect -2913 109 -2847 121
rect -2817 397 -2751 409
rect -2817 121 -2801 397
rect -2767 121 -2751 397
rect -2817 109 -2751 121
rect -2721 397 -2655 409
rect -2721 121 -2705 397
rect -2671 121 -2655 397
rect -2721 109 -2655 121
rect -2625 397 -2559 409
rect -2625 121 -2609 397
rect -2575 121 -2559 397
rect -2625 109 -2559 121
rect -2529 397 -2463 409
rect -2529 121 -2513 397
rect -2479 121 -2463 397
rect -2529 109 -2463 121
rect -2433 397 -2367 409
rect -2433 121 -2417 397
rect -2383 121 -2367 397
rect -2433 109 -2367 121
rect -2337 397 -2271 409
rect -2337 121 -2321 397
rect -2287 121 -2271 397
rect -2337 109 -2271 121
rect -2241 397 -2175 409
rect -2241 121 -2225 397
rect -2191 121 -2175 397
rect -2241 109 -2175 121
rect -2145 397 -2079 409
rect -2145 121 -2129 397
rect -2095 121 -2079 397
rect -2145 109 -2079 121
rect -2049 397 -1983 409
rect -2049 121 -2033 397
rect -1999 121 -1983 397
rect -2049 109 -1983 121
rect -1953 397 -1887 409
rect -1953 121 -1937 397
rect -1903 121 -1887 397
rect -1953 109 -1887 121
rect -1857 397 -1791 409
rect -1857 121 -1841 397
rect -1807 121 -1791 397
rect -1857 109 -1791 121
rect -1761 397 -1695 409
rect -1761 121 -1745 397
rect -1711 121 -1695 397
rect -1761 109 -1695 121
rect -1665 397 -1599 409
rect -1665 121 -1649 397
rect -1615 121 -1599 397
rect -1665 109 -1599 121
rect -1569 397 -1503 409
rect -1569 121 -1553 397
rect -1519 121 -1503 397
rect -1569 109 -1503 121
rect -1473 397 -1407 409
rect -1473 121 -1457 397
rect -1423 121 -1407 397
rect -1473 109 -1407 121
rect -1377 397 -1311 409
rect -1377 121 -1361 397
rect -1327 121 -1311 397
rect -1377 109 -1311 121
rect -1281 397 -1215 409
rect -1281 121 -1265 397
rect -1231 121 -1215 397
rect -1281 109 -1215 121
rect -1185 397 -1119 409
rect -1185 121 -1169 397
rect -1135 121 -1119 397
rect -1185 109 -1119 121
rect -1089 397 -1023 409
rect -1089 121 -1073 397
rect -1039 121 -1023 397
rect -1089 109 -1023 121
rect -993 397 -927 409
rect -993 121 -977 397
rect -943 121 -927 397
rect -993 109 -927 121
rect -897 397 -831 409
rect -897 121 -881 397
rect -847 121 -831 397
rect -897 109 -831 121
rect -801 397 -735 409
rect -801 121 -785 397
rect -751 121 -735 397
rect -801 109 -735 121
rect -705 397 -639 409
rect -705 121 -689 397
rect -655 121 -639 397
rect -705 109 -639 121
rect -609 397 -543 409
rect -609 121 -593 397
rect -559 121 -543 397
rect -609 109 -543 121
rect -513 397 -447 409
rect -513 121 -497 397
rect -463 121 -447 397
rect -513 109 -447 121
rect -417 397 -351 409
rect -417 121 -401 397
rect -367 121 -351 397
rect -417 109 -351 121
rect -321 397 -255 409
rect -321 121 -305 397
rect -271 121 -255 397
rect -321 109 -255 121
rect -225 397 -159 409
rect -225 121 -209 397
rect -175 121 -159 397
rect -225 109 -159 121
rect -129 397 -63 409
rect -129 121 -113 397
rect -79 121 -63 397
rect -129 109 -63 121
rect -33 397 33 409
rect -33 121 -17 397
rect 17 121 33 397
rect -33 109 33 121
rect 63 397 129 409
rect 63 121 79 397
rect 113 121 129 397
rect 63 109 129 121
rect 159 397 225 409
rect 159 121 175 397
rect 209 121 225 397
rect 159 109 225 121
rect 255 397 321 409
rect 255 121 271 397
rect 305 121 321 397
rect 255 109 321 121
rect 351 397 417 409
rect 351 121 367 397
rect 401 121 417 397
rect 351 109 417 121
rect 447 397 513 409
rect 447 121 463 397
rect 497 121 513 397
rect 447 109 513 121
rect 543 397 609 409
rect 543 121 559 397
rect 593 121 609 397
rect 543 109 609 121
rect 639 397 705 409
rect 639 121 655 397
rect 689 121 705 397
rect 639 109 705 121
rect 735 397 801 409
rect 735 121 751 397
rect 785 121 801 397
rect 735 109 801 121
rect 831 397 897 409
rect 831 121 847 397
rect 881 121 897 397
rect 831 109 897 121
rect 927 397 993 409
rect 927 121 943 397
rect 977 121 993 397
rect 927 109 993 121
rect 1023 397 1089 409
rect 1023 121 1039 397
rect 1073 121 1089 397
rect 1023 109 1089 121
rect 1119 397 1185 409
rect 1119 121 1135 397
rect 1169 121 1185 397
rect 1119 109 1185 121
rect 1215 397 1281 409
rect 1215 121 1231 397
rect 1265 121 1281 397
rect 1215 109 1281 121
rect 1311 397 1377 409
rect 1311 121 1327 397
rect 1361 121 1377 397
rect 1311 109 1377 121
rect 1407 397 1473 409
rect 1407 121 1423 397
rect 1457 121 1473 397
rect 1407 109 1473 121
rect 1503 397 1569 409
rect 1503 121 1519 397
rect 1553 121 1569 397
rect 1503 109 1569 121
rect 1599 397 1665 409
rect 1599 121 1615 397
rect 1649 121 1665 397
rect 1599 109 1665 121
rect 1695 397 1761 409
rect 1695 121 1711 397
rect 1745 121 1761 397
rect 1695 109 1761 121
rect 1791 397 1857 409
rect 1791 121 1807 397
rect 1841 121 1857 397
rect 1791 109 1857 121
rect 1887 397 1953 409
rect 1887 121 1903 397
rect 1937 121 1953 397
rect 1887 109 1953 121
rect 1983 397 2049 409
rect 1983 121 1999 397
rect 2033 121 2049 397
rect 1983 109 2049 121
rect 2079 397 2145 409
rect 2079 121 2095 397
rect 2129 121 2145 397
rect 2079 109 2145 121
rect 2175 397 2241 409
rect 2175 121 2191 397
rect 2225 121 2241 397
rect 2175 109 2241 121
rect 2271 397 2337 409
rect 2271 121 2287 397
rect 2321 121 2337 397
rect 2271 109 2337 121
rect 2367 397 2433 409
rect 2367 121 2383 397
rect 2417 121 2433 397
rect 2367 109 2433 121
rect 2463 397 2529 409
rect 2463 121 2479 397
rect 2513 121 2529 397
rect 2463 109 2529 121
rect 2559 397 2625 409
rect 2559 121 2575 397
rect 2609 121 2625 397
rect 2559 109 2625 121
rect 2655 397 2721 409
rect 2655 121 2671 397
rect 2705 121 2721 397
rect 2655 109 2721 121
rect 2751 397 2817 409
rect 2751 121 2767 397
rect 2801 121 2817 397
rect 2751 109 2817 121
rect 2847 397 2913 409
rect 2847 121 2863 397
rect 2897 121 2913 397
rect 2847 109 2913 121
rect 2943 397 3009 409
rect 2943 121 2959 397
rect 2993 121 3009 397
rect 2943 109 3009 121
rect 3039 397 3105 409
rect 3039 121 3055 397
rect 3089 121 3105 397
rect 3039 109 3105 121
rect 3135 397 3201 409
rect 3135 121 3151 397
rect 3185 121 3201 397
rect 3135 109 3201 121
rect 3231 397 3297 409
rect 3231 121 3247 397
rect 3281 121 3297 397
rect 3231 109 3297 121
rect 3327 397 3393 409
rect 3327 121 3343 397
rect 3377 121 3393 397
rect 3327 109 3393 121
rect 3423 397 3489 409
rect 3423 121 3439 397
rect 3473 121 3489 397
rect 3423 109 3489 121
rect 3519 397 3585 409
rect 3519 121 3535 397
rect 3569 121 3585 397
rect 3519 109 3585 121
rect 3615 397 3681 409
rect 3615 121 3631 397
rect 3665 121 3681 397
rect 3615 109 3681 121
rect 3711 397 3777 409
rect 3711 121 3727 397
rect 3761 121 3777 397
rect 3711 109 3777 121
rect 3807 397 3873 409
rect 3807 121 3823 397
rect 3857 121 3873 397
rect 3807 109 3873 121
rect 3903 397 3969 409
rect 3903 121 3919 397
rect 3953 121 3969 397
rect 3903 109 3969 121
rect 3999 397 4065 409
rect 3999 121 4015 397
rect 4049 121 4065 397
rect 3999 109 4065 121
rect 4095 397 4161 409
rect 4095 121 4111 397
rect 4145 121 4161 397
rect 4095 109 4161 121
rect 4191 397 4257 409
rect 4191 121 4207 397
rect 4241 121 4257 397
rect 4191 109 4257 121
rect 4287 397 4353 409
rect 4287 121 4303 397
rect 4337 121 4353 397
rect 4287 109 4353 121
rect 4383 397 4449 409
rect 4383 121 4399 397
rect 4433 121 4449 397
rect 4383 109 4449 121
rect 4479 397 4545 409
rect 4479 121 4495 397
rect 4529 121 4545 397
rect 4479 109 4545 121
rect 4575 397 4641 409
rect 4575 121 4591 397
rect 4625 121 4641 397
rect 4575 109 4641 121
rect 4671 397 4737 409
rect 4671 121 4687 397
rect 4721 121 4737 397
rect 4671 109 4737 121
rect 4767 397 4829 409
rect 4767 121 4783 397
rect 4817 121 4829 397
rect 4767 109 4829 121
rect -4829 -121 -4767 -109
rect -4829 -397 -4817 -121
rect -4783 -397 -4767 -121
rect -4829 -409 -4767 -397
rect -4737 -121 -4671 -109
rect -4737 -397 -4721 -121
rect -4687 -397 -4671 -121
rect -4737 -409 -4671 -397
rect -4641 -121 -4575 -109
rect -4641 -397 -4625 -121
rect -4591 -397 -4575 -121
rect -4641 -409 -4575 -397
rect -4545 -121 -4479 -109
rect -4545 -397 -4529 -121
rect -4495 -397 -4479 -121
rect -4545 -409 -4479 -397
rect -4449 -121 -4383 -109
rect -4449 -397 -4433 -121
rect -4399 -397 -4383 -121
rect -4449 -409 -4383 -397
rect -4353 -121 -4287 -109
rect -4353 -397 -4337 -121
rect -4303 -397 -4287 -121
rect -4353 -409 -4287 -397
rect -4257 -121 -4191 -109
rect -4257 -397 -4241 -121
rect -4207 -397 -4191 -121
rect -4257 -409 -4191 -397
rect -4161 -121 -4095 -109
rect -4161 -397 -4145 -121
rect -4111 -397 -4095 -121
rect -4161 -409 -4095 -397
rect -4065 -121 -3999 -109
rect -4065 -397 -4049 -121
rect -4015 -397 -3999 -121
rect -4065 -409 -3999 -397
rect -3969 -121 -3903 -109
rect -3969 -397 -3953 -121
rect -3919 -397 -3903 -121
rect -3969 -409 -3903 -397
rect -3873 -121 -3807 -109
rect -3873 -397 -3857 -121
rect -3823 -397 -3807 -121
rect -3873 -409 -3807 -397
rect -3777 -121 -3711 -109
rect -3777 -397 -3761 -121
rect -3727 -397 -3711 -121
rect -3777 -409 -3711 -397
rect -3681 -121 -3615 -109
rect -3681 -397 -3665 -121
rect -3631 -397 -3615 -121
rect -3681 -409 -3615 -397
rect -3585 -121 -3519 -109
rect -3585 -397 -3569 -121
rect -3535 -397 -3519 -121
rect -3585 -409 -3519 -397
rect -3489 -121 -3423 -109
rect -3489 -397 -3473 -121
rect -3439 -397 -3423 -121
rect -3489 -409 -3423 -397
rect -3393 -121 -3327 -109
rect -3393 -397 -3377 -121
rect -3343 -397 -3327 -121
rect -3393 -409 -3327 -397
rect -3297 -121 -3231 -109
rect -3297 -397 -3281 -121
rect -3247 -397 -3231 -121
rect -3297 -409 -3231 -397
rect -3201 -121 -3135 -109
rect -3201 -397 -3185 -121
rect -3151 -397 -3135 -121
rect -3201 -409 -3135 -397
rect -3105 -121 -3039 -109
rect -3105 -397 -3089 -121
rect -3055 -397 -3039 -121
rect -3105 -409 -3039 -397
rect -3009 -121 -2943 -109
rect -3009 -397 -2993 -121
rect -2959 -397 -2943 -121
rect -3009 -409 -2943 -397
rect -2913 -121 -2847 -109
rect -2913 -397 -2897 -121
rect -2863 -397 -2847 -121
rect -2913 -409 -2847 -397
rect -2817 -121 -2751 -109
rect -2817 -397 -2801 -121
rect -2767 -397 -2751 -121
rect -2817 -409 -2751 -397
rect -2721 -121 -2655 -109
rect -2721 -397 -2705 -121
rect -2671 -397 -2655 -121
rect -2721 -409 -2655 -397
rect -2625 -121 -2559 -109
rect -2625 -397 -2609 -121
rect -2575 -397 -2559 -121
rect -2625 -409 -2559 -397
rect -2529 -121 -2463 -109
rect -2529 -397 -2513 -121
rect -2479 -397 -2463 -121
rect -2529 -409 -2463 -397
rect -2433 -121 -2367 -109
rect -2433 -397 -2417 -121
rect -2383 -397 -2367 -121
rect -2433 -409 -2367 -397
rect -2337 -121 -2271 -109
rect -2337 -397 -2321 -121
rect -2287 -397 -2271 -121
rect -2337 -409 -2271 -397
rect -2241 -121 -2175 -109
rect -2241 -397 -2225 -121
rect -2191 -397 -2175 -121
rect -2241 -409 -2175 -397
rect -2145 -121 -2079 -109
rect -2145 -397 -2129 -121
rect -2095 -397 -2079 -121
rect -2145 -409 -2079 -397
rect -2049 -121 -1983 -109
rect -2049 -397 -2033 -121
rect -1999 -397 -1983 -121
rect -2049 -409 -1983 -397
rect -1953 -121 -1887 -109
rect -1953 -397 -1937 -121
rect -1903 -397 -1887 -121
rect -1953 -409 -1887 -397
rect -1857 -121 -1791 -109
rect -1857 -397 -1841 -121
rect -1807 -397 -1791 -121
rect -1857 -409 -1791 -397
rect -1761 -121 -1695 -109
rect -1761 -397 -1745 -121
rect -1711 -397 -1695 -121
rect -1761 -409 -1695 -397
rect -1665 -121 -1599 -109
rect -1665 -397 -1649 -121
rect -1615 -397 -1599 -121
rect -1665 -409 -1599 -397
rect -1569 -121 -1503 -109
rect -1569 -397 -1553 -121
rect -1519 -397 -1503 -121
rect -1569 -409 -1503 -397
rect -1473 -121 -1407 -109
rect -1473 -397 -1457 -121
rect -1423 -397 -1407 -121
rect -1473 -409 -1407 -397
rect -1377 -121 -1311 -109
rect -1377 -397 -1361 -121
rect -1327 -397 -1311 -121
rect -1377 -409 -1311 -397
rect -1281 -121 -1215 -109
rect -1281 -397 -1265 -121
rect -1231 -397 -1215 -121
rect -1281 -409 -1215 -397
rect -1185 -121 -1119 -109
rect -1185 -397 -1169 -121
rect -1135 -397 -1119 -121
rect -1185 -409 -1119 -397
rect -1089 -121 -1023 -109
rect -1089 -397 -1073 -121
rect -1039 -397 -1023 -121
rect -1089 -409 -1023 -397
rect -993 -121 -927 -109
rect -993 -397 -977 -121
rect -943 -397 -927 -121
rect -993 -409 -927 -397
rect -897 -121 -831 -109
rect -897 -397 -881 -121
rect -847 -397 -831 -121
rect -897 -409 -831 -397
rect -801 -121 -735 -109
rect -801 -397 -785 -121
rect -751 -397 -735 -121
rect -801 -409 -735 -397
rect -705 -121 -639 -109
rect -705 -397 -689 -121
rect -655 -397 -639 -121
rect -705 -409 -639 -397
rect -609 -121 -543 -109
rect -609 -397 -593 -121
rect -559 -397 -543 -121
rect -609 -409 -543 -397
rect -513 -121 -447 -109
rect -513 -397 -497 -121
rect -463 -397 -447 -121
rect -513 -409 -447 -397
rect -417 -121 -351 -109
rect -417 -397 -401 -121
rect -367 -397 -351 -121
rect -417 -409 -351 -397
rect -321 -121 -255 -109
rect -321 -397 -305 -121
rect -271 -397 -255 -121
rect -321 -409 -255 -397
rect -225 -121 -159 -109
rect -225 -397 -209 -121
rect -175 -397 -159 -121
rect -225 -409 -159 -397
rect -129 -121 -63 -109
rect -129 -397 -113 -121
rect -79 -397 -63 -121
rect -129 -409 -63 -397
rect -33 -121 33 -109
rect -33 -397 -17 -121
rect 17 -397 33 -121
rect -33 -409 33 -397
rect 63 -121 129 -109
rect 63 -397 79 -121
rect 113 -397 129 -121
rect 63 -409 129 -397
rect 159 -121 225 -109
rect 159 -397 175 -121
rect 209 -397 225 -121
rect 159 -409 225 -397
rect 255 -121 321 -109
rect 255 -397 271 -121
rect 305 -397 321 -121
rect 255 -409 321 -397
rect 351 -121 417 -109
rect 351 -397 367 -121
rect 401 -397 417 -121
rect 351 -409 417 -397
rect 447 -121 513 -109
rect 447 -397 463 -121
rect 497 -397 513 -121
rect 447 -409 513 -397
rect 543 -121 609 -109
rect 543 -397 559 -121
rect 593 -397 609 -121
rect 543 -409 609 -397
rect 639 -121 705 -109
rect 639 -397 655 -121
rect 689 -397 705 -121
rect 639 -409 705 -397
rect 735 -121 801 -109
rect 735 -397 751 -121
rect 785 -397 801 -121
rect 735 -409 801 -397
rect 831 -121 897 -109
rect 831 -397 847 -121
rect 881 -397 897 -121
rect 831 -409 897 -397
rect 927 -121 993 -109
rect 927 -397 943 -121
rect 977 -397 993 -121
rect 927 -409 993 -397
rect 1023 -121 1089 -109
rect 1023 -397 1039 -121
rect 1073 -397 1089 -121
rect 1023 -409 1089 -397
rect 1119 -121 1185 -109
rect 1119 -397 1135 -121
rect 1169 -397 1185 -121
rect 1119 -409 1185 -397
rect 1215 -121 1281 -109
rect 1215 -397 1231 -121
rect 1265 -397 1281 -121
rect 1215 -409 1281 -397
rect 1311 -121 1377 -109
rect 1311 -397 1327 -121
rect 1361 -397 1377 -121
rect 1311 -409 1377 -397
rect 1407 -121 1473 -109
rect 1407 -397 1423 -121
rect 1457 -397 1473 -121
rect 1407 -409 1473 -397
rect 1503 -121 1569 -109
rect 1503 -397 1519 -121
rect 1553 -397 1569 -121
rect 1503 -409 1569 -397
rect 1599 -121 1665 -109
rect 1599 -397 1615 -121
rect 1649 -397 1665 -121
rect 1599 -409 1665 -397
rect 1695 -121 1761 -109
rect 1695 -397 1711 -121
rect 1745 -397 1761 -121
rect 1695 -409 1761 -397
rect 1791 -121 1857 -109
rect 1791 -397 1807 -121
rect 1841 -397 1857 -121
rect 1791 -409 1857 -397
rect 1887 -121 1953 -109
rect 1887 -397 1903 -121
rect 1937 -397 1953 -121
rect 1887 -409 1953 -397
rect 1983 -121 2049 -109
rect 1983 -397 1999 -121
rect 2033 -397 2049 -121
rect 1983 -409 2049 -397
rect 2079 -121 2145 -109
rect 2079 -397 2095 -121
rect 2129 -397 2145 -121
rect 2079 -409 2145 -397
rect 2175 -121 2241 -109
rect 2175 -397 2191 -121
rect 2225 -397 2241 -121
rect 2175 -409 2241 -397
rect 2271 -121 2337 -109
rect 2271 -397 2287 -121
rect 2321 -397 2337 -121
rect 2271 -409 2337 -397
rect 2367 -121 2433 -109
rect 2367 -397 2383 -121
rect 2417 -397 2433 -121
rect 2367 -409 2433 -397
rect 2463 -121 2529 -109
rect 2463 -397 2479 -121
rect 2513 -397 2529 -121
rect 2463 -409 2529 -397
rect 2559 -121 2625 -109
rect 2559 -397 2575 -121
rect 2609 -397 2625 -121
rect 2559 -409 2625 -397
rect 2655 -121 2721 -109
rect 2655 -397 2671 -121
rect 2705 -397 2721 -121
rect 2655 -409 2721 -397
rect 2751 -121 2817 -109
rect 2751 -397 2767 -121
rect 2801 -397 2817 -121
rect 2751 -409 2817 -397
rect 2847 -121 2913 -109
rect 2847 -397 2863 -121
rect 2897 -397 2913 -121
rect 2847 -409 2913 -397
rect 2943 -121 3009 -109
rect 2943 -397 2959 -121
rect 2993 -397 3009 -121
rect 2943 -409 3009 -397
rect 3039 -121 3105 -109
rect 3039 -397 3055 -121
rect 3089 -397 3105 -121
rect 3039 -409 3105 -397
rect 3135 -121 3201 -109
rect 3135 -397 3151 -121
rect 3185 -397 3201 -121
rect 3135 -409 3201 -397
rect 3231 -121 3297 -109
rect 3231 -397 3247 -121
rect 3281 -397 3297 -121
rect 3231 -409 3297 -397
rect 3327 -121 3393 -109
rect 3327 -397 3343 -121
rect 3377 -397 3393 -121
rect 3327 -409 3393 -397
rect 3423 -121 3489 -109
rect 3423 -397 3439 -121
rect 3473 -397 3489 -121
rect 3423 -409 3489 -397
rect 3519 -121 3585 -109
rect 3519 -397 3535 -121
rect 3569 -397 3585 -121
rect 3519 -409 3585 -397
rect 3615 -121 3681 -109
rect 3615 -397 3631 -121
rect 3665 -397 3681 -121
rect 3615 -409 3681 -397
rect 3711 -121 3777 -109
rect 3711 -397 3727 -121
rect 3761 -397 3777 -121
rect 3711 -409 3777 -397
rect 3807 -121 3873 -109
rect 3807 -397 3823 -121
rect 3857 -397 3873 -121
rect 3807 -409 3873 -397
rect 3903 -121 3969 -109
rect 3903 -397 3919 -121
rect 3953 -397 3969 -121
rect 3903 -409 3969 -397
rect 3999 -121 4065 -109
rect 3999 -397 4015 -121
rect 4049 -397 4065 -121
rect 3999 -409 4065 -397
rect 4095 -121 4161 -109
rect 4095 -397 4111 -121
rect 4145 -397 4161 -121
rect 4095 -409 4161 -397
rect 4191 -121 4257 -109
rect 4191 -397 4207 -121
rect 4241 -397 4257 -121
rect 4191 -409 4257 -397
rect 4287 -121 4353 -109
rect 4287 -397 4303 -121
rect 4337 -397 4353 -121
rect 4287 -409 4353 -397
rect 4383 -121 4449 -109
rect 4383 -397 4399 -121
rect 4433 -397 4449 -121
rect 4383 -409 4449 -397
rect 4479 -121 4545 -109
rect 4479 -397 4495 -121
rect 4529 -397 4545 -121
rect 4479 -409 4545 -397
rect 4575 -121 4641 -109
rect 4575 -397 4591 -121
rect 4625 -397 4641 -121
rect 4575 -409 4641 -397
rect 4671 -121 4737 -109
rect 4671 -397 4687 -121
rect 4721 -397 4737 -121
rect 4671 -409 4737 -397
rect 4767 -121 4829 -109
rect 4767 -397 4783 -121
rect 4817 -397 4829 -121
rect 4767 -409 4829 -397
rect -4829 -639 -4767 -627
rect -4829 -915 -4817 -639
rect -4783 -915 -4767 -639
rect -4829 -927 -4767 -915
rect -4737 -639 -4671 -627
rect -4737 -915 -4721 -639
rect -4687 -915 -4671 -639
rect -4737 -927 -4671 -915
rect -4641 -639 -4575 -627
rect -4641 -915 -4625 -639
rect -4591 -915 -4575 -639
rect -4641 -927 -4575 -915
rect -4545 -639 -4479 -627
rect -4545 -915 -4529 -639
rect -4495 -915 -4479 -639
rect -4545 -927 -4479 -915
rect -4449 -639 -4383 -627
rect -4449 -915 -4433 -639
rect -4399 -915 -4383 -639
rect -4449 -927 -4383 -915
rect -4353 -639 -4287 -627
rect -4353 -915 -4337 -639
rect -4303 -915 -4287 -639
rect -4353 -927 -4287 -915
rect -4257 -639 -4191 -627
rect -4257 -915 -4241 -639
rect -4207 -915 -4191 -639
rect -4257 -927 -4191 -915
rect -4161 -639 -4095 -627
rect -4161 -915 -4145 -639
rect -4111 -915 -4095 -639
rect -4161 -927 -4095 -915
rect -4065 -639 -3999 -627
rect -4065 -915 -4049 -639
rect -4015 -915 -3999 -639
rect -4065 -927 -3999 -915
rect -3969 -639 -3903 -627
rect -3969 -915 -3953 -639
rect -3919 -915 -3903 -639
rect -3969 -927 -3903 -915
rect -3873 -639 -3807 -627
rect -3873 -915 -3857 -639
rect -3823 -915 -3807 -639
rect -3873 -927 -3807 -915
rect -3777 -639 -3711 -627
rect -3777 -915 -3761 -639
rect -3727 -915 -3711 -639
rect -3777 -927 -3711 -915
rect -3681 -639 -3615 -627
rect -3681 -915 -3665 -639
rect -3631 -915 -3615 -639
rect -3681 -927 -3615 -915
rect -3585 -639 -3519 -627
rect -3585 -915 -3569 -639
rect -3535 -915 -3519 -639
rect -3585 -927 -3519 -915
rect -3489 -639 -3423 -627
rect -3489 -915 -3473 -639
rect -3439 -915 -3423 -639
rect -3489 -927 -3423 -915
rect -3393 -639 -3327 -627
rect -3393 -915 -3377 -639
rect -3343 -915 -3327 -639
rect -3393 -927 -3327 -915
rect -3297 -639 -3231 -627
rect -3297 -915 -3281 -639
rect -3247 -915 -3231 -639
rect -3297 -927 -3231 -915
rect -3201 -639 -3135 -627
rect -3201 -915 -3185 -639
rect -3151 -915 -3135 -639
rect -3201 -927 -3135 -915
rect -3105 -639 -3039 -627
rect -3105 -915 -3089 -639
rect -3055 -915 -3039 -639
rect -3105 -927 -3039 -915
rect -3009 -639 -2943 -627
rect -3009 -915 -2993 -639
rect -2959 -915 -2943 -639
rect -3009 -927 -2943 -915
rect -2913 -639 -2847 -627
rect -2913 -915 -2897 -639
rect -2863 -915 -2847 -639
rect -2913 -927 -2847 -915
rect -2817 -639 -2751 -627
rect -2817 -915 -2801 -639
rect -2767 -915 -2751 -639
rect -2817 -927 -2751 -915
rect -2721 -639 -2655 -627
rect -2721 -915 -2705 -639
rect -2671 -915 -2655 -639
rect -2721 -927 -2655 -915
rect -2625 -639 -2559 -627
rect -2625 -915 -2609 -639
rect -2575 -915 -2559 -639
rect -2625 -927 -2559 -915
rect -2529 -639 -2463 -627
rect -2529 -915 -2513 -639
rect -2479 -915 -2463 -639
rect -2529 -927 -2463 -915
rect -2433 -639 -2367 -627
rect -2433 -915 -2417 -639
rect -2383 -915 -2367 -639
rect -2433 -927 -2367 -915
rect -2337 -639 -2271 -627
rect -2337 -915 -2321 -639
rect -2287 -915 -2271 -639
rect -2337 -927 -2271 -915
rect -2241 -639 -2175 -627
rect -2241 -915 -2225 -639
rect -2191 -915 -2175 -639
rect -2241 -927 -2175 -915
rect -2145 -639 -2079 -627
rect -2145 -915 -2129 -639
rect -2095 -915 -2079 -639
rect -2145 -927 -2079 -915
rect -2049 -639 -1983 -627
rect -2049 -915 -2033 -639
rect -1999 -915 -1983 -639
rect -2049 -927 -1983 -915
rect -1953 -639 -1887 -627
rect -1953 -915 -1937 -639
rect -1903 -915 -1887 -639
rect -1953 -927 -1887 -915
rect -1857 -639 -1791 -627
rect -1857 -915 -1841 -639
rect -1807 -915 -1791 -639
rect -1857 -927 -1791 -915
rect -1761 -639 -1695 -627
rect -1761 -915 -1745 -639
rect -1711 -915 -1695 -639
rect -1761 -927 -1695 -915
rect -1665 -639 -1599 -627
rect -1665 -915 -1649 -639
rect -1615 -915 -1599 -639
rect -1665 -927 -1599 -915
rect -1569 -639 -1503 -627
rect -1569 -915 -1553 -639
rect -1519 -915 -1503 -639
rect -1569 -927 -1503 -915
rect -1473 -639 -1407 -627
rect -1473 -915 -1457 -639
rect -1423 -915 -1407 -639
rect -1473 -927 -1407 -915
rect -1377 -639 -1311 -627
rect -1377 -915 -1361 -639
rect -1327 -915 -1311 -639
rect -1377 -927 -1311 -915
rect -1281 -639 -1215 -627
rect -1281 -915 -1265 -639
rect -1231 -915 -1215 -639
rect -1281 -927 -1215 -915
rect -1185 -639 -1119 -627
rect -1185 -915 -1169 -639
rect -1135 -915 -1119 -639
rect -1185 -927 -1119 -915
rect -1089 -639 -1023 -627
rect -1089 -915 -1073 -639
rect -1039 -915 -1023 -639
rect -1089 -927 -1023 -915
rect -993 -639 -927 -627
rect -993 -915 -977 -639
rect -943 -915 -927 -639
rect -993 -927 -927 -915
rect -897 -639 -831 -627
rect -897 -915 -881 -639
rect -847 -915 -831 -639
rect -897 -927 -831 -915
rect -801 -639 -735 -627
rect -801 -915 -785 -639
rect -751 -915 -735 -639
rect -801 -927 -735 -915
rect -705 -639 -639 -627
rect -705 -915 -689 -639
rect -655 -915 -639 -639
rect -705 -927 -639 -915
rect -609 -639 -543 -627
rect -609 -915 -593 -639
rect -559 -915 -543 -639
rect -609 -927 -543 -915
rect -513 -639 -447 -627
rect -513 -915 -497 -639
rect -463 -915 -447 -639
rect -513 -927 -447 -915
rect -417 -639 -351 -627
rect -417 -915 -401 -639
rect -367 -915 -351 -639
rect -417 -927 -351 -915
rect -321 -639 -255 -627
rect -321 -915 -305 -639
rect -271 -915 -255 -639
rect -321 -927 -255 -915
rect -225 -639 -159 -627
rect -225 -915 -209 -639
rect -175 -915 -159 -639
rect -225 -927 -159 -915
rect -129 -639 -63 -627
rect -129 -915 -113 -639
rect -79 -915 -63 -639
rect -129 -927 -63 -915
rect -33 -639 33 -627
rect -33 -915 -17 -639
rect 17 -915 33 -639
rect -33 -927 33 -915
rect 63 -639 129 -627
rect 63 -915 79 -639
rect 113 -915 129 -639
rect 63 -927 129 -915
rect 159 -639 225 -627
rect 159 -915 175 -639
rect 209 -915 225 -639
rect 159 -927 225 -915
rect 255 -639 321 -627
rect 255 -915 271 -639
rect 305 -915 321 -639
rect 255 -927 321 -915
rect 351 -639 417 -627
rect 351 -915 367 -639
rect 401 -915 417 -639
rect 351 -927 417 -915
rect 447 -639 513 -627
rect 447 -915 463 -639
rect 497 -915 513 -639
rect 447 -927 513 -915
rect 543 -639 609 -627
rect 543 -915 559 -639
rect 593 -915 609 -639
rect 543 -927 609 -915
rect 639 -639 705 -627
rect 639 -915 655 -639
rect 689 -915 705 -639
rect 639 -927 705 -915
rect 735 -639 801 -627
rect 735 -915 751 -639
rect 785 -915 801 -639
rect 735 -927 801 -915
rect 831 -639 897 -627
rect 831 -915 847 -639
rect 881 -915 897 -639
rect 831 -927 897 -915
rect 927 -639 993 -627
rect 927 -915 943 -639
rect 977 -915 993 -639
rect 927 -927 993 -915
rect 1023 -639 1089 -627
rect 1023 -915 1039 -639
rect 1073 -915 1089 -639
rect 1023 -927 1089 -915
rect 1119 -639 1185 -627
rect 1119 -915 1135 -639
rect 1169 -915 1185 -639
rect 1119 -927 1185 -915
rect 1215 -639 1281 -627
rect 1215 -915 1231 -639
rect 1265 -915 1281 -639
rect 1215 -927 1281 -915
rect 1311 -639 1377 -627
rect 1311 -915 1327 -639
rect 1361 -915 1377 -639
rect 1311 -927 1377 -915
rect 1407 -639 1473 -627
rect 1407 -915 1423 -639
rect 1457 -915 1473 -639
rect 1407 -927 1473 -915
rect 1503 -639 1569 -627
rect 1503 -915 1519 -639
rect 1553 -915 1569 -639
rect 1503 -927 1569 -915
rect 1599 -639 1665 -627
rect 1599 -915 1615 -639
rect 1649 -915 1665 -639
rect 1599 -927 1665 -915
rect 1695 -639 1761 -627
rect 1695 -915 1711 -639
rect 1745 -915 1761 -639
rect 1695 -927 1761 -915
rect 1791 -639 1857 -627
rect 1791 -915 1807 -639
rect 1841 -915 1857 -639
rect 1791 -927 1857 -915
rect 1887 -639 1953 -627
rect 1887 -915 1903 -639
rect 1937 -915 1953 -639
rect 1887 -927 1953 -915
rect 1983 -639 2049 -627
rect 1983 -915 1999 -639
rect 2033 -915 2049 -639
rect 1983 -927 2049 -915
rect 2079 -639 2145 -627
rect 2079 -915 2095 -639
rect 2129 -915 2145 -639
rect 2079 -927 2145 -915
rect 2175 -639 2241 -627
rect 2175 -915 2191 -639
rect 2225 -915 2241 -639
rect 2175 -927 2241 -915
rect 2271 -639 2337 -627
rect 2271 -915 2287 -639
rect 2321 -915 2337 -639
rect 2271 -927 2337 -915
rect 2367 -639 2433 -627
rect 2367 -915 2383 -639
rect 2417 -915 2433 -639
rect 2367 -927 2433 -915
rect 2463 -639 2529 -627
rect 2463 -915 2479 -639
rect 2513 -915 2529 -639
rect 2463 -927 2529 -915
rect 2559 -639 2625 -627
rect 2559 -915 2575 -639
rect 2609 -915 2625 -639
rect 2559 -927 2625 -915
rect 2655 -639 2721 -627
rect 2655 -915 2671 -639
rect 2705 -915 2721 -639
rect 2655 -927 2721 -915
rect 2751 -639 2817 -627
rect 2751 -915 2767 -639
rect 2801 -915 2817 -639
rect 2751 -927 2817 -915
rect 2847 -639 2913 -627
rect 2847 -915 2863 -639
rect 2897 -915 2913 -639
rect 2847 -927 2913 -915
rect 2943 -639 3009 -627
rect 2943 -915 2959 -639
rect 2993 -915 3009 -639
rect 2943 -927 3009 -915
rect 3039 -639 3105 -627
rect 3039 -915 3055 -639
rect 3089 -915 3105 -639
rect 3039 -927 3105 -915
rect 3135 -639 3201 -627
rect 3135 -915 3151 -639
rect 3185 -915 3201 -639
rect 3135 -927 3201 -915
rect 3231 -639 3297 -627
rect 3231 -915 3247 -639
rect 3281 -915 3297 -639
rect 3231 -927 3297 -915
rect 3327 -639 3393 -627
rect 3327 -915 3343 -639
rect 3377 -915 3393 -639
rect 3327 -927 3393 -915
rect 3423 -639 3489 -627
rect 3423 -915 3439 -639
rect 3473 -915 3489 -639
rect 3423 -927 3489 -915
rect 3519 -639 3585 -627
rect 3519 -915 3535 -639
rect 3569 -915 3585 -639
rect 3519 -927 3585 -915
rect 3615 -639 3681 -627
rect 3615 -915 3631 -639
rect 3665 -915 3681 -639
rect 3615 -927 3681 -915
rect 3711 -639 3777 -627
rect 3711 -915 3727 -639
rect 3761 -915 3777 -639
rect 3711 -927 3777 -915
rect 3807 -639 3873 -627
rect 3807 -915 3823 -639
rect 3857 -915 3873 -639
rect 3807 -927 3873 -915
rect 3903 -639 3969 -627
rect 3903 -915 3919 -639
rect 3953 -915 3969 -639
rect 3903 -927 3969 -915
rect 3999 -639 4065 -627
rect 3999 -915 4015 -639
rect 4049 -915 4065 -639
rect 3999 -927 4065 -915
rect 4095 -639 4161 -627
rect 4095 -915 4111 -639
rect 4145 -915 4161 -639
rect 4095 -927 4161 -915
rect 4191 -639 4257 -627
rect 4191 -915 4207 -639
rect 4241 -915 4257 -639
rect 4191 -927 4257 -915
rect 4287 -639 4353 -627
rect 4287 -915 4303 -639
rect 4337 -915 4353 -639
rect 4287 -927 4353 -915
rect 4383 -639 4449 -627
rect 4383 -915 4399 -639
rect 4433 -915 4449 -639
rect 4383 -927 4449 -915
rect 4479 -639 4545 -627
rect 4479 -915 4495 -639
rect 4529 -915 4545 -639
rect 4479 -927 4545 -915
rect 4575 -639 4641 -627
rect 4575 -915 4591 -639
rect 4625 -915 4641 -639
rect 4575 -927 4641 -915
rect 4671 -639 4737 -627
rect 4671 -915 4687 -639
rect 4721 -915 4737 -639
rect 4671 -927 4737 -915
rect 4767 -639 4829 -627
rect 4767 -915 4783 -639
rect 4817 -915 4829 -639
rect 4767 -927 4829 -915
<< ndiffc >>
rect -4817 639 -4783 915
rect -4721 639 -4687 915
rect -4625 639 -4591 915
rect -4529 639 -4495 915
rect -4433 639 -4399 915
rect -4337 639 -4303 915
rect -4241 639 -4207 915
rect -4145 639 -4111 915
rect -4049 639 -4015 915
rect -3953 639 -3919 915
rect -3857 639 -3823 915
rect -3761 639 -3727 915
rect -3665 639 -3631 915
rect -3569 639 -3535 915
rect -3473 639 -3439 915
rect -3377 639 -3343 915
rect -3281 639 -3247 915
rect -3185 639 -3151 915
rect -3089 639 -3055 915
rect -2993 639 -2959 915
rect -2897 639 -2863 915
rect -2801 639 -2767 915
rect -2705 639 -2671 915
rect -2609 639 -2575 915
rect -2513 639 -2479 915
rect -2417 639 -2383 915
rect -2321 639 -2287 915
rect -2225 639 -2191 915
rect -2129 639 -2095 915
rect -2033 639 -1999 915
rect -1937 639 -1903 915
rect -1841 639 -1807 915
rect -1745 639 -1711 915
rect -1649 639 -1615 915
rect -1553 639 -1519 915
rect -1457 639 -1423 915
rect -1361 639 -1327 915
rect -1265 639 -1231 915
rect -1169 639 -1135 915
rect -1073 639 -1039 915
rect -977 639 -943 915
rect -881 639 -847 915
rect -785 639 -751 915
rect -689 639 -655 915
rect -593 639 -559 915
rect -497 639 -463 915
rect -401 639 -367 915
rect -305 639 -271 915
rect -209 639 -175 915
rect -113 639 -79 915
rect -17 639 17 915
rect 79 639 113 915
rect 175 639 209 915
rect 271 639 305 915
rect 367 639 401 915
rect 463 639 497 915
rect 559 639 593 915
rect 655 639 689 915
rect 751 639 785 915
rect 847 639 881 915
rect 943 639 977 915
rect 1039 639 1073 915
rect 1135 639 1169 915
rect 1231 639 1265 915
rect 1327 639 1361 915
rect 1423 639 1457 915
rect 1519 639 1553 915
rect 1615 639 1649 915
rect 1711 639 1745 915
rect 1807 639 1841 915
rect 1903 639 1937 915
rect 1999 639 2033 915
rect 2095 639 2129 915
rect 2191 639 2225 915
rect 2287 639 2321 915
rect 2383 639 2417 915
rect 2479 639 2513 915
rect 2575 639 2609 915
rect 2671 639 2705 915
rect 2767 639 2801 915
rect 2863 639 2897 915
rect 2959 639 2993 915
rect 3055 639 3089 915
rect 3151 639 3185 915
rect 3247 639 3281 915
rect 3343 639 3377 915
rect 3439 639 3473 915
rect 3535 639 3569 915
rect 3631 639 3665 915
rect 3727 639 3761 915
rect 3823 639 3857 915
rect 3919 639 3953 915
rect 4015 639 4049 915
rect 4111 639 4145 915
rect 4207 639 4241 915
rect 4303 639 4337 915
rect 4399 639 4433 915
rect 4495 639 4529 915
rect 4591 639 4625 915
rect 4687 639 4721 915
rect 4783 639 4817 915
rect -4817 121 -4783 397
rect -4721 121 -4687 397
rect -4625 121 -4591 397
rect -4529 121 -4495 397
rect -4433 121 -4399 397
rect -4337 121 -4303 397
rect -4241 121 -4207 397
rect -4145 121 -4111 397
rect -4049 121 -4015 397
rect -3953 121 -3919 397
rect -3857 121 -3823 397
rect -3761 121 -3727 397
rect -3665 121 -3631 397
rect -3569 121 -3535 397
rect -3473 121 -3439 397
rect -3377 121 -3343 397
rect -3281 121 -3247 397
rect -3185 121 -3151 397
rect -3089 121 -3055 397
rect -2993 121 -2959 397
rect -2897 121 -2863 397
rect -2801 121 -2767 397
rect -2705 121 -2671 397
rect -2609 121 -2575 397
rect -2513 121 -2479 397
rect -2417 121 -2383 397
rect -2321 121 -2287 397
rect -2225 121 -2191 397
rect -2129 121 -2095 397
rect -2033 121 -1999 397
rect -1937 121 -1903 397
rect -1841 121 -1807 397
rect -1745 121 -1711 397
rect -1649 121 -1615 397
rect -1553 121 -1519 397
rect -1457 121 -1423 397
rect -1361 121 -1327 397
rect -1265 121 -1231 397
rect -1169 121 -1135 397
rect -1073 121 -1039 397
rect -977 121 -943 397
rect -881 121 -847 397
rect -785 121 -751 397
rect -689 121 -655 397
rect -593 121 -559 397
rect -497 121 -463 397
rect -401 121 -367 397
rect -305 121 -271 397
rect -209 121 -175 397
rect -113 121 -79 397
rect -17 121 17 397
rect 79 121 113 397
rect 175 121 209 397
rect 271 121 305 397
rect 367 121 401 397
rect 463 121 497 397
rect 559 121 593 397
rect 655 121 689 397
rect 751 121 785 397
rect 847 121 881 397
rect 943 121 977 397
rect 1039 121 1073 397
rect 1135 121 1169 397
rect 1231 121 1265 397
rect 1327 121 1361 397
rect 1423 121 1457 397
rect 1519 121 1553 397
rect 1615 121 1649 397
rect 1711 121 1745 397
rect 1807 121 1841 397
rect 1903 121 1937 397
rect 1999 121 2033 397
rect 2095 121 2129 397
rect 2191 121 2225 397
rect 2287 121 2321 397
rect 2383 121 2417 397
rect 2479 121 2513 397
rect 2575 121 2609 397
rect 2671 121 2705 397
rect 2767 121 2801 397
rect 2863 121 2897 397
rect 2959 121 2993 397
rect 3055 121 3089 397
rect 3151 121 3185 397
rect 3247 121 3281 397
rect 3343 121 3377 397
rect 3439 121 3473 397
rect 3535 121 3569 397
rect 3631 121 3665 397
rect 3727 121 3761 397
rect 3823 121 3857 397
rect 3919 121 3953 397
rect 4015 121 4049 397
rect 4111 121 4145 397
rect 4207 121 4241 397
rect 4303 121 4337 397
rect 4399 121 4433 397
rect 4495 121 4529 397
rect 4591 121 4625 397
rect 4687 121 4721 397
rect 4783 121 4817 397
rect -4817 -397 -4783 -121
rect -4721 -397 -4687 -121
rect -4625 -397 -4591 -121
rect -4529 -397 -4495 -121
rect -4433 -397 -4399 -121
rect -4337 -397 -4303 -121
rect -4241 -397 -4207 -121
rect -4145 -397 -4111 -121
rect -4049 -397 -4015 -121
rect -3953 -397 -3919 -121
rect -3857 -397 -3823 -121
rect -3761 -397 -3727 -121
rect -3665 -397 -3631 -121
rect -3569 -397 -3535 -121
rect -3473 -397 -3439 -121
rect -3377 -397 -3343 -121
rect -3281 -397 -3247 -121
rect -3185 -397 -3151 -121
rect -3089 -397 -3055 -121
rect -2993 -397 -2959 -121
rect -2897 -397 -2863 -121
rect -2801 -397 -2767 -121
rect -2705 -397 -2671 -121
rect -2609 -397 -2575 -121
rect -2513 -397 -2479 -121
rect -2417 -397 -2383 -121
rect -2321 -397 -2287 -121
rect -2225 -397 -2191 -121
rect -2129 -397 -2095 -121
rect -2033 -397 -1999 -121
rect -1937 -397 -1903 -121
rect -1841 -397 -1807 -121
rect -1745 -397 -1711 -121
rect -1649 -397 -1615 -121
rect -1553 -397 -1519 -121
rect -1457 -397 -1423 -121
rect -1361 -397 -1327 -121
rect -1265 -397 -1231 -121
rect -1169 -397 -1135 -121
rect -1073 -397 -1039 -121
rect -977 -397 -943 -121
rect -881 -397 -847 -121
rect -785 -397 -751 -121
rect -689 -397 -655 -121
rect -593 -397 -559 -121
rect -497 -397 -463 -121
rect -401 -397 -367 -121
rect -305 -397 -271 -121
rect -209 -397 -175 -121
rect -113 -397 -79 -121
rect -17 -397 17 -121
rect 79 -397 113 -121
rect 175 -397 209 -121
rect 271 -397 305 -121
rect 367 -397 401 -121
rect 463 -397 497 -121
rect 559 -397 593 -121
rect 655 -397 689 -121
rect 751 -397 785 -121
rect 847 -397 881 -121
rect 943 -397 977 -121
rect 1039 -397 1073 -121
rect 1135 -397 1169 -121
rect 1231 -397 1265 -121
rect 1327 -397 1361 -121
rect 1423 -397 1457 -121
rect 1519 -397 1553 -121
rect 1615 -397 1649 -121
rect 1711 -397 1745 -121
rect 1807 -397 1841 -121
rect 1903 -397 1937 -121
rect 1999 -397 2033 -121
rect 2095 -397 2129 -121
rect 2191 -397 2225 -121
rect 2287 -397 2321 -121
rect 2383 -397 2417 -121
rect 2479 -397 2513 -121
rect 2575 -397 2609 -121
rect 2671 -397 2705 -121
rect 2767 -397 2801 -121
rect 2863 -397 2897 -121
rect 2959 -397 2993 -121
rect 3055 -397 3089 -121
rect 3151 -397 3185 -121
rect 3247 -397 3281 -121
rect 3343 -397 3377 -121
rect 3439 -397 3473 -121
rect 3535 -397 3569 -121
rect 3631 -397 3665 -121
rect 3727 -397 3761 -121
rect 3823 -397 3857 -121
rect 3919 -397 3953 -121
rect 4015 -397 4049 -121
rect 4111 -397 4145 -121
rect 4207 -397 4241 -121
rect 4303 -397 4337 -121
rect 4399 -397 4433 -121
rect 4495 -397 4529 -121
rect 4591 -397 4625 -121
rect 4687 -397 4721 -121
rect 4783 -397 4817 -121
rect -4817 -915 -4783 -639
rect -4721 -915 -4687 -639
rect -4625 -915 -4591 -639
rect -4529 -915 -4495 -639
rect -4433 -915 -4399 -639
rect -4337 -915 -4303 -639
rect -4241 -915 -4207 -639
rect -4145 -915 -4111 -639
rect -4049 -915 -4015 -639
rect -3953 -915 -3919 -639
rect -3857 -915 -3823 -639
rect -3761 -915 -3727 -639
rect -3665 -915 -3631 -639
rect -3569 -915 -3535 -639
rect -3473 -915 -3439 -639
rect -3377 -915 -3343 -639
rect -3281 -915 -3247 -639
rect -3185 -915 -3151 -639
rect -3089 -915 -3055 -639
rect -2993 -915 -2959 -639
rect -2897 -915 -2863 -639
rect -2801 -915 -2767 -639
rect -2705 -915 -2671 -639
rect -2609 -915 -2575 -639
rect -2513 -915 -2479 -639
rect -2417 -915 -2383 -639
rect -2321 -915 -2287 -639
rect -2225 -915 -2191 -639
rect -2129 -915 -2095 -639
rect -2033 -915 -1999 -639
rect -1937 -915 -1903 -639
rect -1841 -915 -1807 -639
rect -1745 -915 -1711 -639
rect -1649 -915 -1615 -639
rect -1553 -915 -1519 -639
rect -1457 -915 -1423 -639
rect -1361 -915 -1327 -639
rect -1265 -915 -1231 -639
rect -1169 -915 -1135 -639
rect -1073 -915 -1039 -639
rect -977 -915 -943 -639
rect -881 -915 -847 -639
rect -785 -915 -751 -639
rect -689 -915 -655 -639
rect -593 -915 -559 -639
rect -497 -915 -463 -639
rect -401 -915 -367 -639
rect -305 -915 -271 -639
rect -209 -915 -175 -639
rect -113 -915 -79 -639
rect -17 -915 17 -639
rect 79 -915 113 -639
rect 175 -915 209 -639
rect 271 -915 305 -639
rect 367 -915 401 -639
rect 463 -915 497 -639
rect 559 -915 593 -639
rect 655 -915 689 -639
rect 751 -915 785 -639
rect 847 -915 881 -639
rect 943 -915 977 -639
rect 1039 -915 1073 -639
rect 1135 -915 1169 -639
rect 1231 -915 1265 -639
rect 1327 -915 1361 -639
rect 1423 -915 1457 -639
rect 1519 -915 1553 -639
rect 1615 -915 1649 -639
rect 1711 -915 1745 -639
rect 1807 -915 1841 -639
rect 1903 -915 1937 -639
rect 1999 -915 2033 -639
rect 2095 -915 2129 -639
rect 2191 -915 2225 -639
rect 2287 -915 2321 -639
rect 2383 -915 2417 -639
rect 2479 -915 2513 -639
rect 2575 -915 2609 -639
rect 2671 -915 2705 -639
rect 2767 -915 2801 -639
rect 2863 -915 2897 -639
rect 2959 -915 2993 -639
rect 3055 -915 3089 -639
rect 3151 -915 3185 -639
rect 3247 -915 3281 -639
rect 3343 -915 3377 -639
rect 3439 -915 3473 -639
rect 3535 -915 3569 -639
rect 3631 -915 3665 -639
rect 3727 -915 3761 -639
rect 3823 -915 3857 -639
rect 3919 -915 3953 -639
rect 4015 -915 4049 -639
rect 4111 -915 4145 -639
rect 4207 -915 4241 -639
rect 4303 -915 4337 -639
rect 4399 -915 4433 -639
rect 4495 -915 4529 -639
rect 4591 -915 4625 -639
rect 4687 -915 4721 -639
rect 4783 -915 4817 -639
<< psubdiff >>
rect -4931 1067 -4835 1101
rect 4835 1067 4931 1101
rect -4931 1005 -4897 1067
rect 4897 1005 4931 1067
rect -4931 -1067 -4897 -1005
rect 4897 -1067 4931 -1005
rect -4931 -1101 -4835 -1067
rect 4835 -1101 4931 -1067
<< psubdiffcont >>
rect -4835 1067 4835 1101
rect -4931 -1005 -4897 1005
rect 4897 -1005 4931 1005
rect -4835 -1101 4835 -1067
<< poly >>
rect -4785 999 -4719 1015
rect -4785 965 -4769 999
rect -4735 965 -4719 999
rect -4785 949 -4719 965
rect -4593 999 -4527 1015
rect -4593 965 -4577 999
rect -4543 965 -4527 999
rect -4767 927 -4737 949
rect -4671 927 -4641 953
rect -4593 949 -4527 965
rect -4401 999 -4335 1015
rect -4401 965 -4385 999
rect -4351 965 -4335 999
rect -4575 927 -4545 949
rect -4479 927 -4449 953
rect -4401 949 -4335 965
rect -4209 999 -4143 1015
rect -4209 965 -4193 999
rect -4159 965 -4143 999
rect -4383 927 -4353 949
rect -4287 927 -4257 953
rect -4209 949 -4143 965
rect -4017 999 -3951 1015
rect -4017 965 -4001 999
rect -3967 965 -3951 999
rect -4191 927 -4161 949
rect -4095 927 -4065 953
rect -4017 949 -3951 965
rect -3825 999 -3759 1015
rect -3825 965 -3809 999
rect -3775 965 -3759 999
rect -3999 927 -3969 949
rect -3903 927 -3873 953
rect -3825 949 -3759 965
rect -3633 999 -3567 1015
rect -3633 965 -3617 999
rect -3583 965 -3567 999
rect -3807 927 -3777 949
rect -3711 927 -3681 953
rect -3633 949 -3567 965
rect -3441 999 -3375 1015
rect -3441 965 -3425 999
rect -3391 965 -3375 999
rect -3615 927 -3585 949
rect -3519 927 -3489 953
rect -3441 949 -3375 965
rect -3249 999 -3183 1015
rect -3249 965 -3233 999
rect -3199 965 -3183 999
rect -3423 927 -3393 949
rect -3327 927 -3297 953
rect -3249 949 -3183 965
rect -3057 999 -2991 1015
rect -3057 965 -3041 999
rect -3007 965 -2991 999
rect -3231 927 -3201 949
rect -3135 927 -3105 953
rect -3057 949 -2991 965
rect -2865 999 -2799 1015
rect -2865 965 -2849 999
rect -2815 965 -2799 999
rect -3039 927 -3009 949
rect -2943 927 -2913 953
rect -2865 949 -2799 965
rect -2673 999 -2607 1015
rect -2673 965 -2657 999
rect -2623 965 -2607 999
rect -2847 927 -2817 949
rect -2751 927 -2721 953
rect -2673 949 -2607 965
rect -2481 999 -2415 1015
rect -2481 965 -2465 999
rect -2431 965 -2415 999
rect -2655 927 -2625 949
rect -2559 927 -2529 953
rect -2481 949 -2415 965
rect -2289 999 -2223 1015
rect -2289 965 -2273 999
rect -2239 965 -2223 999
rect -2463 927 -2433 949
rect -2367 927 -2337 953
rect -2289 949 -2223 965
rect -2097 999 -2031 1015
rect -2097 965 -2081 999
rect -2047 965 -2031 999
rect -2271 927 -2241 949
rect -2175 927 -2145 953
rect -2097 949 -2031 965
rect -1905 999 -1839 1015
rect -1905 965 -1889 999
rect -1855 965 -1839 999
rect -2079 927 -2049 949
rect -1983 927 -1953 953
rect -1905 949 -1839 965
rect -1713 999 -1647 1015
rect -1713 965 -1697 999
rect -1663 965 -1647 999
rect -1887 927 -1857 949
rect -1791 927 -1761 953
rect -1713 949 -1647 965
rect -1521 999 -1455 1015
rect -1521 965 -1505 999
rect -1471 965 -1455 999
rect -1695 927 -1665 949
rect -1599 927 -1569 953
rect -1521 949 -1455 965
rect -1329 999 -1263 1015
rect -1329 965 -1313 999
rect -1279 965 -1263 999
rect -1503 927 -1473 949
rect -1407 927 -1377 953
rect -1329 949 -1263 965
rect -1137 999 -1071 1015
rect -1137 965 -1121 999
rect -1087 965 -1071 999
rect -1311 927 -1281 949
rect -1215 927 -1185 953
rect -1137 949 -1071 965
rect -945 999 -879 1015
rect -945 965 -929 999
rect -895 965 -879 999
rect -1119 927 -1089 949
rect -1023 927 -993 953
rect -945 949 -879 965
rect -753 999 -687 1015
rect -753 965 -737 999
rect -703 965 -687 999
rect -927 927 -897 949
rect -831 927 -801 953
rect -753 949 -687 965
rect -561 999 -495 1015
rect -561 965 -545 999
rect -511 965 -495 999
rect -735 927 -705 949
rect -639 927 -609 953
rect -561 949 -495 965
rect -369 999 -303 1015
rect -369 965 -353 999
rect -319 965 -303 999
rect -543 927 -513 949
rect -447 927 -417 953
rect -369 949 -303 965
rect -177 999 -111 1015
rect -177 965 -161 999
rect -127 965 -111 999
rect -351 927 -321 949
rect -255 927 -225 953
rect -177 949 -111 965
rect 15 999 81 1015
rect 15 965 31 999
rect 65 965 81 999
rect -159 927 -129 949
rect -63 927 -33 953
rect 15 949 81 965
rect 207 999 273 1015
rect 207 965 223 999
rect 257 965 273 999
rect 33 927 63 949
rect 129 927 159 953
rect 207 949 273 965
rect 399 999 465 1015
rect 399 965 415 999
rect 449 965 465 999
rect 225 927 255 949
rect 321 927 351 953
rect 399 949 465 965
rect 591 999 657 1015
rect 591 965 607 999
rect 641 965 657 999
rect 417 927 447 949
rect 513 927 543 953
rect 591 949 657 965
rect 783 999 849 1015
rect 783 965 799 999
rect 833 965 849 999
rect 609 927 639 949
rect 705 927 735 953
rect 783 949 849 965
rect 975 999 1041 1015
rect 975 965 991 999
rect 1025 965 1041 999
rect 801 927 831 949
rect 897 927 927 953
rect 975 949 1041 965
rect 1167 999 1233 1015
rect 1167 965 1183 999
rect 1217 965 1233 999
rect 993 927 1023 949
rect 1089 927 1119 953
rect 1167 949 1233 965
rect 1359 999 1425 1015
rect 1359 965 1375 999
rect 1409 965 1425 999
rect 1185 927 1215 949
rect 1281 927 1311 953
rect 1359 949 1425 965
rect 1551 999 1617 1015
rect 1551 965 1567 999
rect 1601 965 1617 999
rect 1377 927 1407 949
rect 1473 927 1503 953
rect 1551 949 1617 965
rect 1743 999 1809 1015
rect 1743 965 1759 999
rect 1793 965 1809 999
rect 1569 927 1599 949
rect 1665 927 1695 953
rect 1743 949 1809 965
rect 1935 999 2001 1015
rect 1935 965 1951 999
rect 1985 965 2001 999
rect 1761 927 1791 949
rect 1857 927 1887 953
rect 1935 949 2001 965
rect 2127 999 2193 1015
rect 2127 965 2143 999
rect 2177 965 2193 999
rect 1953 927 1983 949
rect 2049 927 2079 953
rect 2127 949 2193 965
rect 2319 999 2385 1015
rect 2319 965 2335 999
rect 2369 965 2385 999
rect 2145 927 2175 949
rect 2241 927 2271 953
rect 2319 949 2385 965
rect 2511 999 2577 1015
rect 2511 965 2527 999
rect 2561 965 2577 999
rect 2337 927 2367 949
rect 2433 927 2463 953
rect 2511 949 2577 965
rect 2703 999 2769 1015
rect 2703 965 2719 999
rect 2753 965 2769 999
rect 2529 927 2559 949
rect 2625 927 2655 953
rect 2703 949 2769 965
rect 2895 999 2961 1015
rect 2895 965 2911 999
rect 2945 965 2961 999
rect 2721 927 2751 949
rect 2817 927 2847 953
rect 2895 949 2961 965
rect 3087 999 3153 1015
rect 3087 965 3103 999
rect 3137 965 3153 999
rect 2913 927 2943 949
rect 3009 927 3039 953
rect 3087 949 3153 965
rect 3279 999 3345 1015
rect 3279 965 3295 999
rect 3329 965 3345 999
rect 3105 927 3135 949
rect 3201 927 3231 953
rect 3279 949 3345 965
rect 3471 999 3537 1015
rect 3471 965 3487 999
rect 3521 965 3537 999
rect 3297 927 3327 949
rect 3393 927 3423 953
rect 3471 949 3537 965
rect 3663 999 3729 1015
rect 3663 965 3679 999
rect 3713 965 3729 999
rect 3489 927 3519 949
rect 3585 927 3615 953
rect 3663 949 3729 965
rect 3855 999 3921 1015
rect 3855 965 3871 999
rect 3905 965 3921 999
rect 3681 927 3711 949
rect 3777 927 3807 953
rect 3855 949 3921 965
rect 4047 999 4113 1015
rect 4047 965 4063 999
rect 4097 965 4113 999
rect 3873 927 3903 949
rect 3969 927 3999 953
rect 4047 949 4113 965
rect 4239 999 4305 1015
rect 4239 965 4255 999
rect 4289 965 4305 999
rect 4065 927 4095 949
rect 4161 927 4191 953
rect 4239 949 4305 965
rect 4431 999 4497 1015
rect 4431 965 4447 999
rect 4481 965 4497 999
rect 4257 927 4287 949
rect 4353 927 4383 953
rect 4431 949 4497 965
rect 4623 999 4689 1015
rect 4623 965 4639 999
rect 4673 965 4689 999
rect 4449 927 4479 949
rect 4545 927 4575 953
rect 4623 949 4689 965
rect 4641 927 4671 949
rect 4737 927 4767 953
rect -4767 601 -4737 627
rect -4671 605 -4641 627
rect -4689 589 -4623 605
rect -4575 601 -4545 627
rect -4479 605 -4449 627
rect -4689 555 -4673 589
rect -4639 555 -4623 589
rect -4689 539 -4623 555
rect -4497 589 -4431 605
rect -4383 601 -4353 627
rect -4287 605 -4257 627
rect -4497 555 -4481 589
rect -4447 555 -4431 589
rect -4497 539 -4431 555
rect -4305 589 -4239 605
rect -4191 601 -4161 627
rect -4095 605 -4065 627
rect -4305 555 -4289 589
rect -4255 555 -4239 589
rect -4305 539 -4239 555
rect -4113 589 -4047 605
rect -3999 601 -3969 627
rect -3903 605 -3873 627
rect -4113 555 -4097 589
rect -4063 555 -4047 589
rect -4113 539 -4047 555
rect -3921 589 -3855 605
rect -3807 601 -3777 627
rect -3711 605 -3681 627
rect -3921 555 -3905 589
rect -3871 555 -3855 589
rect -3921 539 -3855 555
rect -3729 589 -3663 605
rect -3615 601 -3585 627
rect -3519 605 -3489 627
rect -3729 555 -3713 589
rect -3679 555 -3663 589
rect -3729 539 -3663 555
rect -3537 589 -3471 605
rect -3423 601 -3393 627
rect -3327 605 -3297 627
rect -3537 555 -3521 589
rect -3487 555 -3471 589
rect -3537 539 -3471 555
rect -3345 589 -3279 605
rect -3231 601 -3201 627
rect -3135 605 -3105 627
rect -3345 555 -3329 589
rect -3295 555 -3279 589
rect -3345 539 -3279 555
rect -3153 589 -3087 605
rect -3039 601 -3009 627
rect -2943 605 -2913 627
rect -3153 555 -3137 589
rect -3103 555 -3087 589
rect -3153 539 -3087 555
rect -2961 589 -2895 605
rect -2847 601 -2817 627
rect -2751 605 -2721 627
rect -2961 555 -2945 589
rect -2911 555 -2895 589
rect -2961 539 -2895 555
rect -2769 589 -2703 605
rect -2655 601 -2625 627
rect -2559 605 -2529 627
rect -2769 555 -2753 589
rect -2719 555 -2703 589
rect -2769 539 -2703 555
rect -2577 589 -2511 605
rect -2463 601 -2433 627
rect -2367 605 -2337 627
rect -2577 555 -2561 589
rect -2527 555 -2511 589
rect -2577 539 -2511 555
rect -2385 589 -2319 605
rect -2271 601 -2241 627
rect -2175 605 -2145 627
rect -2385 555 -2369 589
rect -2335 555 -2319 589
rect -2385 539 -2319 555
rect -2193 589 -2127 605
rect -2079 601 -2049 627
rect -1983 605 -1953 627
rect -2193 555 -2177 589
rect -2143 555 -2127 589
rect -2193 539 -2127 555
rect -2001 589 -1935 605
rect -1887 601 -1857 627
rect -1791 605 -1761 627
rect -2001 555 -1985 589
rect -1951 555 -1935 589
rect -2001 539 -1935 555
rect -1809 589 -1743 605
rect -1695 601 -1665 627
rect -1599 605 -1569 627
rect -1809 555 -1793 589
rect -1759 555 -1743 589
rect -1809 539 -1743 555
rect -1617 589 -1551 605
rect -1503 601 -1473 627
rect -1407 605 -1377 627
rect -1617 555 -1601 589
rect -1567 555 -1551 589
rect -1617 539 -1551 555
rect -1425 589 -1359 605
rect -1311 601 -1281 627
rect -1215 605 -1185 627
rect -1425 555 -1409 589
rect -1375 555 -1359 589
rect -1425 539 -1359 555
rect -1233 589 -1167 605
rect -1119 601 -1089 627
rect -1023 605 -993 627
rect -1233 555 -1217 589
rect -1183 555 -1167 589
rect -1233 539 -1167 555
rect -1041 589 -975 605
rect -927 601 -897 627
rect -831 605 -801 627
rect -1041 555 -1025 589
rect -991 555 -975 589
rect -1041 539 -975 555
rect -849 589 -783 605
rect -735 601 -705 627
rect -639 605 -609 627
rect -849 555 -833 589
rect -799 555 -783 589
rect -849 539 -783 555
rect -657 589 -591 605
rect -543 601 -513 627
rect -447 605 -417 627
rect -657 555 -641 589
rect -607 555 -591 589
rect -657 539 -591 555
rect -465 589 -399 605
rect -351 601 -321 627
rect -255 605 -225 627
rect -465 555 -449 589
rect -415 555 -399 589
rect -465 539 -399 555
rect -273 589 -207 605
rect -159 601 -129 627
rect -63 605 -33 627
rect -273 555 -257 589
rect -223 555 -207 589
rect -273 539 -207 555
rect -81 589 -15 605
rect 33 601 63 627
rect 129 605 159 627
rect -81 555 -65 589
rect -31 555 -15 589
rect -81 539 -15 555
rect 111 589 177 605
rect 225 601 255 627
rect 321 605 351 627
rect 111 555 127 589
rect 161 555 177 589
rect 111 539 177 555
rect 303 589 369 605
rect 417 601 447 627
rect 513 605 543 627
rect 303 555 319 589
rect 353 555 369 589
rect 303 539 369 555
rect 495 589 561 605
rect 609 601 639 627
rect 705 605 735 627
rect 495 555 511 589
rect 545 555 561 589
rect 495 539 561 555
rect 687 589 753 605
rect 801 601 831 627
rect 897 605 927 627
rect 687 555 703 589
rect 737 555 753 589
rect 687 539 753 555
rect 879 589 945 605
rect 993 601 1023 627
rect 1089 605 1119 627
rect 879 555 895 589
rect 929 555 945 589
rect 879 539 945 555
rect 1071 589 1137 605
rect 1185 601 1215 627
rect 1281 605 1311 627
rect 1071 555 1087 589
rect 1121 555 1137 589
rect 1071 539 1137 555
rect 1263 589 1329 605
rect 1377 601 1407 627
rect 1473 605 1503 627
rect 1263 555 1279 589
rect 1313 555 1329 589
rect 1263 539 1329 555
rect 1455 589 1521 605
rect 1569 601 1599 627
rect 1665 605 1695 627
rect 1455 555 1471 589
rect 1505 555 1521 589
rect 1455 539 1521 555
rect 1647 589 1713 605
rect 1761 601 1791 627
rect 1857 605 1887 627
rect 1647 555 1663 589
rect 1697 555 1713 589
rect 1647 539 1713 555
rect 1839 589 1905 605
rect 1953 601 1983 627
rect 2049 605 2079 627
rect 1839 555 1855 589
rect 1889 555 1905 589
rect 1839 539 1905 555
rect 2031 589 2097 605
rect 2145 601 2175 627
rect 2241 605 2271 627
rect 2031 555 2047 589
rect 2081 555 2097 589
rect 2031 539 2097 555
rect 2223 589 2289 605
rect 2337 601 2367 627
rect 2433 605 2463 627
rect 2223 555 2239 589
rect 2273 555 2289 589
rect 2223 539 2289 555
rect 2415 589 2481 605
rect 2529 601 2559 627
rect 2625 605 2655 627
rect 2415 555 2431 589
rect 2465 555 2481 589
rect 2415 539 2481 555
rect 2607 589 2673 605
rect 2721 601 2751 627
rect 2817 605 2847 627
rect 2607 555 2623 589
rect 2657 555 2673 589
rect 2607 539 2673 555
rect 2799 589 2865 605
rect 2913 601 2943 627
rect 3009 605 3039 627
rect 2799 555 2815 589
rect 2849 555 2865 589
rect 2799 539 2865 555
rect 2991 589 3057 605
rect 3105 601 3135 627
rect 3201 605 3231 627
rect 2991 555 3007 589
rect 3041 555 3057 589
rect 2991 539 3057 555
rect 3183 589 3249 605
rect 3297 601 3327 627
rect 3393 605 3423 627
rect 3183 555 3199 589
rect 3233 555 3249 589
rect 3183 539 3249 555
rect 3375 589 3441 605
rect 3489 601 3519 627
rect 3585 605 3615 627
rect 3375 555 3391 589
rect 3425 555 3441 589
rect 3375 539 3441 555
rect 3567 589 3633 605
rect 3681 601 3711 627
rect 3777 605 3807 627
rect 3567 555 3583 589
rect 3617 555 3633 589
rect 3567 539 3633 555
rect 3759 589 3825 605
rect 3873 601 3903 627
rect 3969 605 3999 627
rect 3759 555 3775 589
rect 3809 555 3825 589
rect 3759 539 3825 555
rect 3951 589 4017 605
rect 4065 601 4095 627
rect 4161 605 4191 627
rect 3951 555 3967 589
rect 4001 555 4017 589
rect 3951 539 4017 555
rect 4143 589 4209 605
rect 4257 601 4287 627
rect 4353 605 4383 627
rect 4143 555 4159 589
rect 4193 555 4209 589
rect 4143 539 4209 555
rect 4335 589 4401 605
rect 4449 601 4479 627
rect 4545 605 4575 627
rect 4335 555 4351 589
rect 4385 555 4401 589
rect 4335 539 4401 555
rect 4527 589 4593 605
rect 4641 601 4671 627
rect 4737 605 4767 627
rect 4527 555 4543 589
rect 4577 555 4593 589
rect 4527 539 4593 555
rect 4719 589 4785 605
rect 4719 555 4735 589
rect 4769 555 4785 589
rect 4719 539 4785 555
rect -4689 481 -4623 497
rect -4689 447 -4673 481
rect -4639 447 -4623 481
rect -4767 409 -4737 435
rect -4689 431 -4623 447
rect -4497 481 -4431 497
rect -4497 447 -4481 481
rect -4447 447 -4431 481
rect -4671 409 -4641 431
rect -4575 409 -4545 435
rect -4497 431 -4431 447
rect -4305 481 -4239 497
rect -4305 447 -4289 481
rect -4255 447 -4239 481
rect -4479 409 -4449 431
rect -4383 409 -4353 435
rect -4305 431 -4239 447
rect -4113 481 -4047 497
rect -4113 447 -4097 481
rect -4063 447 -4047 481
rect -4287 409 -4257 431
rect -4191 409 -4161 435
rect -4113 431 -4047 447
rect -3921 481 -3855 497
rect -3921 447 -3905 481
rect -3871 447 -3855 481
rect -4095 409 -4065 431
rect -3999 409 -3969 435
rect -3921 431 -3855 447
rect -3729 481 -3663 497
rect -3729 447 -3713 481
rect -3679 447 -3663 481
rect -3903 409 -3873 431
rect -3807 409 -3777 435
rect -3729 431 -3663 447
rect -3537 481 -3471 497
rect -3537 447 -3521 481
rect -3487 447 -3471 481
rect -3711 409 -3681 431
rect -3615 409 -3585 435
rect -3537 431 -3471 447
rect -3345 481 -3279 497
rect -3345 447 -3329 481
rect -3295 447 -3279 481
rect -3519 409 -3489 431
rect -3423 409 -3393 435
rect -3345 431 -3279 447
rect -3153 481 -3087 497
rect -3153 447 -3137 481
rect -3103 447 -3087 481
rect -3327 409 -3297 431
rect -3231 409 -3201 435
rect -3153 431 -3087 447
rect -2961 481 -2895 497
rect -2961 447 -2945 481
rect -2911 447 -2895 481
rect -3135 409 -3105 431
rect -3039 409 -3009 435
rect -2961 431 -2895 447
rect -2769 481 -2703 497
rect -2769 447 -2753 481
rect -2719 447 -2703 481
rect -2943 409 -2913 431
rect -2847 409 -2817 435
rect -2769 431 -2703 447
rect -2577 481 -2511 497
rect -2577 447 -2561 481
rect -2527 447 -2511 481
rect -2751 409 -2721 431
rect -2655 409 -2625 435
rect -2577 431 -2511 447
rect -2385 481 -2319 497
rect -2385 447 -2369 481
rect -2335 447 -2319 481
rect -2559 409 -2529 431
rect -2463 409 -2433 435
rect -2385 431 -2319 447
rect -2193 481 -2127 497
rect -2193 447 -2177 481
rect -2143 447 -2127 481
rect -2367 409 -2337 431
rect -2271 409 -2241 435
rect -2193 431 -2127 447
rect -2001 481 -1935 497
rect -2001 447 -1985 481
rect -1951 447 -1935 481
rect -2175 409 -2145 431
rect -2079 409 -2049 435
rect -2001 431 -1935 447
rect -1809 481 -1743 497
rect -1809 447 -1793 481
rect -1759 447 -1743 481
rect -1983 409 -1953 431
rect -1887 409 -1857 435
rect -1809 431 -1743 447
rect -1617 481 -1551 497
rect -1617 447 -1601 481
rect -1567 447 -1551 481
rect -1791 409 -1761 431
rect -1695 409 -1665 435
rect -1617 431 -1551 447
rect -1425 481 -1359 497
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1599 409 -1569 431
rect -1503 409 -1473 435
rect -1425 431 -1359 447
rect -1233 481 -1167 497
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1407 409 -1377 431
rect -1311 409 -1281 435
rect -1233 431 -1167 447
rect -1041 481 -975 497
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -1215 409 -1185 431
rect -1119 409 -1089 435
rect -1041 431 -975 447
rect -849 481 -783 497
rect -849 447 -833 481
rect -799 447 -783 481
rect -1023 409 -993 431
rect -927 409 -897 435
rect -849 431 -783 447
rect -657 481 -591 497
rect -657 447 -641 481
rect -607 447 -591 481
rect -831 409 -801 431
rect -735 409 -705 435
rect -657 431 -591 447
rect -465 481 -399 497
rect -465 447 -449 481
rect -415 447 -399 481
rect -639 409 -609 431
rect -543 409 -513 435
rect -465 431 -399 447
rect -273 481 -207 497
rect -273 447 -257 481
rect -223 447 -207 481
rect -447 409 -417 431
rect -351 409 -321 435
rect -273 431 -207 447
rect -81 481 -15 497
rect -81 447 -65 481
rect -31 447 -15 481
rect -255 409 -225 431
rect -159 409 -129 435
rect -81 431 -15 447
rect 111 481 177 497
rect 111 447 127 481
rect 161 447 177 481
rect -63 409 -33 431
rect 33 409 63 435
rect 111 431 177 447
rect 303 481 369 497
rect 303 447 319 481
rect 353 447 369 481
rect 129 409 159 431
rect 225 409 255 435
rect 303 431 369 447
rect 495 481 561 497
rect 495 447 511 481
rect 545 447 561 481
rect 321 409 351 431
rect 417 409 447 435
rect 495 431 561 447
rect 687 481 753 497
rect 687 447 703 481
rect 737 447 753 481
rect 513 409 543 431
rect 609 409 639 435
rect 687 431 753 447
rect 879 481 945 497
rect 879 447 895 481
rect 929 447 945 481
rect 705 409 735 431
rect 801 409 831 435
rect 879 431 945 447
rect 1071 481 1137 497
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 897 409 927 431
rect 993 409 1023 435
rect 1071 431 1137 447
rect 1263 481 1329 497
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1089 409 1119 431
rect 1185 409 1215 435
rect 1263 431 1329 447
rect 1455 481 1521 497
rect 1455 447 1471 481
rect 1505 447 1521 481
rect 1281 409 1311 431
rect 1377 409 1407 435
rect 1455 431 1521 447
rect 1647 481 1713 497
rect 1647 447 1663 481
rect 1697 447 1713 481
rect 1473 409 1503 431
rect 1569 409 1599 435
rect 1647 431 1713 447
rect 1839 481 1905 497
rect 1839 447 1855 481
rect 1889 447 1905 481
rect 1665 409 1695 431
rect 1761 409 1791 435
rect 1839 431 1905 447
rect 2031 481 2097 497
rect 2031 447 2047 481
rect 2081 447 2097 481
rect 1857 409 1887 431
rect 1953 409 1983 435
rect 2031 431 2097 447
rect 2223 481 2289 497
rect 2223 447 2239 481
rect 2273 447 2289 481
rect 2049 409 2079 431
rect 2145 409 2175 435
rect 2223 431 2289 447
rect 2415 481 2481 497
rect 2415 447 2431 481
rect 2465 447 2481 481
rect 2241 409 2271 431
rect 2337 409 2367 435
rect 2415 431 2481 447
rect 2607 481 2673 497
rect 2607 447 2623 481
rect 2657 447 2673 481
rect 2433 409 2463 431
rect 2529 409 2559 435
rect 2607 431 2673 447
rect 2799 481 2865 497
rect 2799 447 2815 481
rect 2849 447 2865 481
rect 2625 409 2655 431
rect 2721 409 2751 435
rect 2799 431 2865 447
rect 2991 481 3057 497
rect 2991 447 3007 481
rect 3041 447 3057 481
rect 2817 409 2847 431
rect 2913 409 2943 435
rect 2991 431 3057 447
rect 3183 481 3249 497
rect 3183 447 3199 481
rect 3233 447 3249 481
rect 3009 409 3039 431
rect 3105 409 3135 435
rect 3183 431 3249 447
rect 3375 481 3441 497
rect 3375 447 3391 481
rect 3425 447 3441 481
rect 3201 409 3231 431
rect 3297 409 3327 435
rect 3375 431 3441 447
rect 3567 481 3633 497
rect 3567 447 3583 481
rect 3617 447 3633 481
rect 3393 409 3423 431
rect 3489 409 3519 435
rect 3567 431 3633 447
rect 3759 481 3825 497
rect 3759 447 3775 481
rect 3809 447 3825 481
rect 3585 409 3615 431
rect 3681 409 3711 435
rect 3759 431 3825 447
rect 3951 481 4017 497
rect 3951 447 3967 481
rect 4001 447 4017 481
rect 3777 409 3807 431
rect 3873 409 3903 435
rect 3951 431 4017 447
rect 4143 481 4209 497
rect 4143 447 4159 481
rect 4193 447 4209 481
rect 3969 409 3999 431
rect 4065 409 4095 435
rect 4143 431 4209 447
rect 4335 481 4401 497
rect 4335 447 4351 481
rect 4385 447 4401 481
rect 4161 409 4191 431
rect 4257 409 4287 435
rect 4335 431 4401 447
rect 4527 481 4593 497
rect 4527 447 4543 481
rect 4577 447 4593 481
rect 4353 409 4383 431
rect 4449 409 4479 435
rect 4527 431 4593 447
rect 4719 481 4785 497
rect 4719 447 4735 481
rect 4769 447 4785 481
rect 4545 409 4575 431
rect 4641 409 4671 435
rect 4719 431 4785 447
rect 4737 409 4767 431
rect -4767 87 -4737 109
rect -4785 71 -4719 87
rect -4671 83 -4641 109
rect -4575 87 -4545 109
rect -4785 37 -4769 71
rect -4735 37 -4719 71
rect -4785 21 -4719 37
rect -4593 71 -4527 87
rect -4479 83 -4449 109
rect -4383 87 -4353 109
rect -4593 37 -4577 71
rect -4543 37 -4527 71
rect -4593 21 -4527 37
rect -4401 71 -4335 87
rect -4287 83 -4257 109
rect -4191 87 -4161 109
rect -4401 37 -4385 71
rect -4351 37 -4335 71
rect -4401 21 -4335 37
rect -4209 71 -4143 87
rect -4095 83 -4065 109
rect -3999 87 -3969 109
rect -4209 37 -4193 71
rect -4159 37 -4143 71
rect -4209 21 -4143 37
rect -4017 71 -3951 87
rect -3903 83 -3873 109
rect -3807 87 -3777 109
rect -4017 37 -4001 71
rect -3967 37 -3951 71
rect -4017 21 -3951 37
rect -3825 71 -3759 87
rect -3711 83 -3681 109
rect -3615 87 -3585 109
rect -3825 37 -3809 71
rect -3775 37 -3759 71
rect -3825 21 -3759 37
rect -3633 71 -3567 87
rect -3519 83 -3489 109
rect -3423 87 -3393 109
rect -3633 37 -3617 71
rect -3583 37 -3567 71
rect -3633 21 -3567 37
rect -3441 71 -3375 87
rect -3327 83 -3297 109
rect -3231 87 -3201 109
rect -3441 37 -3425 71
rect -3391 37 -3375 71
rect -3441 21 -3375 37
rect -3249 71 -3183 87
rect -3135 83 -3105 109
rect -3039 87 -3009 109
rect -3249 37 -3233 71
rect -3199 37 -3183 71
rect -3249 21 -3183 37
rect -3057 71 -2991 87
rect -2943 83 -2913 109
rect -2847 87 -2817 109
rect -3057 37 -3041 71
rect -3007 37 -2991 71
rect -3057 21 -2991 37
rect -2865 71 -2799 87
rect -2751 83 -2721 109
rect -2655 87 -2625 109
rect -2865 37 -2849 71
rect -2815 37 -2799 71
rect -2865 21 -2799 37
rect -2673 71 -2607 87
rect -2559 83 -2529 109
rect -2463 87 -2433 109
rect -2673 37 -2657 71
rect -2623 37 -2607 71
rect -2673 21 -2607 37
rect -2481 71 -2415 87
rect -2367 83 -2337 109
rect -2271 87 -2241 109
rect -2481 37 -2465 71
rect -2431 37 -2415 71
rect -2481 21 -2415 37
rect -2289 71 -2223 87
rect -2175 83 -2145 109
rect -2079 87 -2049 109
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2289 21 -2223 37
rect -2097 71 -2031 87
rect -1983 83 -1953 109
rect -1887 87 -1857 109
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -2097 21 -2031 37
rect -1905 71 -1839 87
rect -1791 83 -1761 109
rect -1695 87 -1665 109
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1905 21 -1839 37
rect -1713 71 -1647 87
rect -1599 83 -1569 109
rect -1503 87 -1473 109
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1713 21 -1647 37
rect -1521 71 -1455 87
rect -1407 83 -1377 109
rect -1311 87 -1281 109
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1521 21 -1455 37
rect -1329 71 -1263 87
rect -1215 83 -1185 109
rect -1119 87 -1089 109
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1329 21 -1263 37
rect -1137 71 -1071 87
rect -1023 83 -993 109
rect -927 87 -897 109
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -1137 21 -1071 37
rect -945 71 -879 87
rect -831 83 -801 109
rect -735 87 -705 109
rect -945 37 -929 71
rect -895 37 -879 71
rect -945 21 -879 37
rect -753 71 -687 87
rect -639 83 -609 109
rect -543 87 -513 109
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 609 87 639 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 705 83 735 109
rect 801 87 831 109
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 897 83 927 109
rect 993 87 1023 109
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect 975 71 1041 87
rect 1089 83 1119 109
rect 1185 87 1215 109
rect 975 37 991 71
rect 1025 37 1041 71
rect 975 21 1041 37
rect 1167 71 1233 87
rect 1281 83 1311 109
rect 1377 87 1407 109
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1167 21 1233 37
rect 1359 71 1425 87
rect 1473 83 1503 109
rect 1569 87 1599 109
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1359 21 1425 37
rect 1551 71 1617 87
rect 1665 83 1695 109
rect 1761 87 1791 109
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1551 21 1617 37
rect 1743 71 1809 87
rect 1857 83 1887 109
rect 1953 87 1983 109
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1743 21 1809 37
rect 1935 71 2001 87
rect 2049 83 2079 109
rect 2145 87 2175 109
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 1935 21 2001 37
rect 2127 71 2193 87
rect 2241 83 2271 109
rect 2337 87 2367 109
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2127 21 2193 37
rect 2319 71 2385 87
rect 2433 83 2463 109
rect 2529 87 2559 109
rect 2319 37 2335 71
rect 2369 37 2385 71
rect 2319 21 2385 37
rect 2511 71 2577 87
rect 2625 83 2655 109
rect 2721 87 2751 109
rect 2511 37 2527 71
rect 2561 37 2577 71
rect 2511 21 2577 37
rect 2703 71 2769 87
rect 2817 83 2847 109
rect 2913 87 2943 109
rect 2703 37 2719 71
rect 2753 37 2769 71
rect 2703 21 2769 37
rect 2895 71 2961 87
rect 3009 83 3039 109
rect 3105 87 3135 109
rect 2895 37 2911 71
rect 2945 37 2961 71
rect 2895 21 2961 37
rect 3087 71 3153 87
rect 3201 83 3231 109
rect 3297 87 3327 109
rect 3087 37 3103 71
rect 3137 37 3153 71
rect 3087 21 3153 37
rect 3279 71 3345 87
rect 3393 83 3423 109
rect 3489 87 3519 109
rect 3279 37 3295 71
rect 3329 37 3345 71
rect 3279 21 3345 37
rect 3471 71 3537 87
rect 3585 83 3615 109
rect 3681 87 3711 109
rect 3471 37 3487 71
rect 3521 37 3537 71
rect 3471 21 3537 37
rect 3663 71 3729 87
rect 3777 83 3807 109
rect 3873 87 3903 109
rect 3663 37 3679 71
rect 3713 37 3729 71
rect 3663 21 3729 37
rect 3855 71 3921 87
rect 3969 83 3999 109
rect 4065 87 4095 109
rect 3855 37 3871 71
rect 3905 37 3921 71
rect 3855 21 3921 37
rect 4047 71 4113 87
rect 4161 83 4191 109
rect 4257 87 4287 109
rect 4047 37 4063 71
rect 4097 37 4113 71
rect 4047 21 4113 37
rect 4239 71 4305 87
rect 4353 83 4383 109
rect 4449 87 4479 109
rect 4239 37 4255 71
rect 4289 37 4305 71
rect 4239 21 4305 37
rect 4431 71 4497 87
rect 4545 83 4575 109
rect 4641 87 4671 109
rect 4431 37 4447 71
rect 4481 37 4497 71
rect 4431 21 4497 37
rect 4623 71 4689 87
rect 4737 83 4767 109
rect 4623 37 4639 71
rect 4673 37 4689 71
rect 4623 21 4689 37
rect -4785 -37 -4719 -21
rect -4785 -71 -4769 -37
rect -4735 -71 -4719 -37
rect -4785 -87 -4719 -71
rect -4593 -37 -4527 -21
rect -4593 -71 -4577 -37
rect -4543 -71 -4527 -37
rect -4767 -109 -4737 -87
rect -4671 -109 -4641 -83
rect -4593 -87 -4527 -71
rect -4401 -37 -4335 -21
rect -4401 -71 -4385 -37
rect -4351 -71 -4335 -37
rect -4575 -109 -4545 -87
rect -4479 -109 -4449 -83
rect -4401 -87 -4335 -71
rect -4209 -37 -4143 -21
rect -4209 -71 -4193 -37
rect -4159 -71 -4143 -37
rect -4383 -109 -4353 -87
rect -4287 -109 -4257 -83
rect -4209 -87 -4143 -71
rect -4017 -37 -3951 -21
rect -4017 -71 -4001 -37
rect -3967 -71 -3951 -37
rect -4191 -109 -4161 -87
rect -4095 -109 -4065 -83
rect -4017 -87 -3951 -71
rect -3825 -37 -3759 -21
rect -3825 -71 -3809 -37
rect -3775 -71 -3759 -37
rect -3999 -109 -3969 -87
rect -3903 -109 -3873 -83
rect -3825 -87 -3759 -71
rect -3633 -37 -3567 -21
rect -3633 -71 -3617 -37
rect -3583 -71 -3567 -37
rect -3807 -109 -3777 -87
rect -3711 -109 -3681 -83
rect -3633 -87 -3567 -71
rect -3441 -37 -3375 -21
rect -3441 -71 -3425 -37
rect -3391 -71 -3375 -37
rect -3615 -109 -3585 -87
rect -3519 -109 -3489 -83
rect -3441 -87 -3375 -71
rect -3249 -37 -3183 -21
rect -3249 -71 -3233 -37
rect -3199 -71 -3183 -37
rect -3423 -109 -3393 -87
rect -3327 -109 -3297 -83
rect -3249 -87 -3183 -71
rect -3057 -37 -2991 -21
rect -3057 -71 -3041 -37
rect -3007 -71 -2991 -37
rect -3231 -109 -3201 -87
rect -3135 -109 -3105 -83
rect -3057 -87 -2991 -71
rect -2865 -37 -2799 -21
rect -2865 -71 -2849 -37
rect -2815 -71 -2799 -37
rect -3039 -109 -3009 -87
rect -2943 -109 -2913 -83
rect -2865 -87 -2799 -71
rect -2673 -37 -2607 -21
rect -2673 -71 -2657 -37
rect -2623 -71 -2607 -37
rect -2847 -109 -2817 -87
rect -2751 -109 -2721 -83
rect -2673 -87 -2607 -71
rect -2481 -37 -2415 -21
rect -2481 -71 -2465 -37
rect -2431 -71 -2415 -37
rect -2655 -109 -2625 -87
rect -2559 -109 -2529 -83
rect -2481 -87 -2415 -71
rect -2289 -37 -2223 -21
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2463 -109 -2433 -87
rect -2367 -109 -2337 -83
rect -2289 -87 -2223 -71
rect -2097 -37 -2031 -21
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -2271 -109 -2241 -87
rect -2175 -109 -2145 -83
rect -2097 -87 -2031 -71
rect -1905 -37 -1839 -21
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -2079 -109 -2049 -87
rect -1983 -109 -1953 -83
rect -1905 -87 -1839 -71
rect -1713 -37 -1647 -21
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1887 -109 -1857 -87
rect -1791 -109 -1761 -83
rect -1713 -87 -1647 -71
rect -1521 -37 -1455 -21
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1695 -109 -1665 -87
rect -1599 -109 -1569 -83
rect -1521 -87 -1455 -71
rect -1329 -37 -1263 -21
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1503 -109 -1473 -87
rect -1407 -109 -1377 -83
rect -1329 -87 -1263 -71
rect -1137 -37 -1071 -21
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -1311 -109 -1281 -87
rect -1215 -109 -1185 -83
rect -1137 -87 -1071 -71
rect -945 -37 -879 -21
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -1119 -109 -1089 -87
rect -1023 -109 -993 -83
rect -945 -87 -879 -71
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -927 -109 -897 -87
rect -831 -109 -801 -83
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -735 -109 -705 -87
rect -639 -109 -609 -83
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 417 -109 447 -87
rect 513 -109 543 -83
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 609 -109 639 -87
rect 705 -109 735 -83
rect 783 -87 849 -71
rect 975 -37 1041 -21
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 801 -109 831 -87
rect 897 -109 927 -83
rect 975 -87 1041 -71
rect 1167 -37 1233 -21
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 993 -109 1023 -87
rect 1089 -109 1119 -83
rect 1167 -87 1233 -71
rect 1359 -37 1425 -21
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1185 -109 1215 -87
rect 1281 -109 1311 -83
rect 1359 -87 1425 -71
rect 1551 -37 1617 -21
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1377 -109 1407 -87
rect 1473 -109 1503 -83
rect 1551 -87 1617 -71
rect 1743 -37 1809 -21
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1569 -109 1599 -87
rect 1665 -109 1695 -83
rect 1743 -87 1809 -71
rect 1935 -37 2001 -21
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 1761 -109 1791 -87
rect 1857 -109 1887 -83
rect 1935 -87 2001 -71
rect 2127 -37 2193 -21
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 1953 -109 1983 -87
rect 2049 -109 2079 -83
rect 2127 -87 2193 -71
rect 2319 -37 2385 -21
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect 2145 -109 2175 -87
rect 2241 -109 2271 -83
rect 2319 -87 2385 -71
rect 2511 -37 2577 -21
rect 2511 -71 2527 -37
rect 2561 -71 2577 -37
rect 2337 -109 2367 -87
rect 2433 -109 2463 -83
rect 2511 -87 2577 -71
rect 2703 -37 2769 -21
rect 2703 -71 2719 -37
rect 2753 -71 2769 -37
rect 2529 -109 2559 -87
rect 2625 -109 2655 -83
rect 2703 -87 2769 -71
rect 2895 -37 2961 -21
rect 2895 -71 2911 -37
rect 2945 -71 2961 -37
rect 2721 -109 2751 -87
rect 2817 -109 2847 -83
rect 2895 -87 2961 -71
rect 3087 -37 3153 -21
rect 3087 -71 3103 -37
rect 3137 -71 3153 -37
rect 2913 -109 2943 -87
rect 3009 -109 3039 -83
rect 3087 -87 3153 -71
rect 3279 -37 3345 -21
rect 3279 -71 3295 -37
rect 3329 -71 3345 -37
rect 3105 -109 3135 -87
rect 3201 -109 3231 -83
rect 3279 -87 3345 -71
rect 3471 -37 3537 -21
rect 3471 -71 3487 -37
rect 3521 -71 3537 -37
rect 3297 -109 3327 -87
rect 3393 -109 3423 -83
rect 3471 -87 3537 -71
rect 3663 -37 3729 -21
rect 3663 -71 3679 -37
rect 3713 -71 3729 -37
rect 3489 -109 3519 -87
rect 3585 -109 3615 -83
rect 3663 -87 3729 -71
rect 3855 -37 3921 -21
rect 3855 -71 3871 -37
rect 3905 -71 3921 -37
rect 3681 -109 3711 -87
rect 3777 -109 3807 -83
rect 3855 -87 3921 -71
rect 4047 -37 4113 -21
rect 4047 -71 4063 -37
rect 4097 -71 4113 -37
rect 3873 -109 3903 -87
rect 3969 -109 3999 -83
rect 4047 -87 4113 -71
rect 4239 -37 4305 -21
rect 4239 -71 4255 -37
rect 4289 -71 4305 -37
rect 4065 -109 4095 -87
rect 4161 -109 4191 -83
rect 4239 -87 4305 -71
rect 4431 -37 4497 -21
rect 4431 -71 4447 -37
rect 4481 -71 4497 -37
rect 4257 -109 4287 -87
rect 4353 -109 4383 -83
rect 4431 -87 4497 -71
rect 4623 -37 4689 -21
rect 4623 -71 4639 -37
rect 4673 -71 4689 -37
rect 4449 -109 4479 -87
rect 4545 -109 4575 -83
rect 4623 -87 4689 -71
rect 4641 -109 4671 -87
rect 4737 -109 4767 -83
rect -4767 -435 -4737 -409
rect -4671 -431 -4641 -409
rect -4689 -447 -4623 -431
rect -4575 -435 -4545 -409
rect -4479 -431 -4449 -409
rect -4689 -481 -4673 -447
rect -4639 -481 -4623 -447
rect -4689 -497 -4623 -481
rect -4497 -447 -4431 -431
rect -4383 -435 -4353 -409
rect -4287 -431 -4257 -409
rect -4497 -481 -4481 -447
rect -4447 -481 -4431 -447
rect -4497 -497 -4431 -481
rect -4305 -447 -4239 -431
rect -4191 -435 -4161 -409
rect -4095 -431 -4065 -409
rect -4305 -481 -4289 -447
rect -4255 -481 -4239 -447
rect -4305 -497 -4239 -481
rect -4113 -447 -4047 -431
rect -3999 -435 -3969 -409
rect -3903 -431 -3873 -409
rect -4113 -481 -4097 -447
rect -4063 -481 -4047 -447
rect -4113 -497 -4047 -481
rect -3921 -447 -3855 -431
rect -3807 -435 -3777 -409
rect -3711 -431 -3681 -409
rect -3921 -481 -3905 -447
rect -3871 -481 -3855 -447
rect -3921 -497 -3855 -481
rect -3729 -447 -3663 -431
rect -3615 -435 -3585 -409
rect -3519 -431 -3489 -409
rect -3729 -481 -3713 -447
rect -3679 -481 -3663 -447
rect -3729 -497 -3663 -481
rect -3537 -447 -3471 -431
rect -3423 -435 -3393 -409
rect -3327 -431 -3297 -409
rect -3537 -481 -3521 -447
rect -3487 -481 -3471 -447
rect -3537 -497 -3471 -481
rect -3345 -447 -3279 -431
rect -3231 -435 -3201 -409
rect -3135 -431 -3105 -409
rect -3345 -481 -3329 -447
rect -3295 -481 -3279 -447
rect -3345 -497 -3279 -481
rect -3153 -447 -3087 -431
rect -3039 -435 -3009 -409
rect -2943 -431 -2913 -409
rect -3153 -481 -3137 -447
rect -3103 -481 -3087 -447
rect -3153 -497 -3087 -481
rect -2961 -447 -2895 -431
rect -2847 -435 -2817 -409
rect -2751 -431 -2721 -409
rect -2961 -481 -2945 -447
rect -2911 -481 -2895 -447
rect -2961 -497 -2895 -481
rect -2769 -447 -2703 -431
rect -2655 -435 -2625 -409
rect -2559 -431 -2529 -409
rect -2769 -481 -2753 -447
rect -2719 -481 -2703 -447
rect -2769 -497 -2703 -481
rect -2577 -447 -2511 -431
rect -2463 -435 -2433 -409
rect -2367 -431 -2337 -409
rect -2577 -481 -2561 -447
rect -2527 -481 -2511 -447
rect -2577 -497 -2511 -481
rect -2385 -447 -2319 -431
rect -2271 -435 -2241 -409
rect -2175 -431 -2145 -409
rect -2385 -481 -2369 -447
rect -2335 -481 -2319 -447
rect -2385 -497 -2319 -481
rect -2193 -447 -2127 -431
rect -2079 -435 -2049 -409
rect -1983 -431 -1953 -409
rect -2193 -481 -2177 -447
rect -2143 -481 -2127 -447
rect -2193 -497 -2127 -481
rect -2001 -447 -1935 -431
rect -1887 -435 -1857 -409
rect -1791 -431 -1761 -409
rect -2001 -481 -1985 -447
rect -1951 -481 -1935 -447
rect -2001 -497 -1935 -481
rect -1809 -447 -1743 -431
rect -1695 -435 -1665 -409
rect -1599 -431 -1569 -409
rect -1809 -481 -1793 -447
rect -1759 -481 -1743 -447
rect -1809 -497 -1743 -481
rect -1617 -447 -1551 -431
rect -1503 -435 -1473 -409
rect -1407 -431 -1377 -409
rect -1617 -481 -1601 -447
rect -1567 -481 -1551 -447
rect -1617 -497 -1551 -481
rect -1425 -447 -1359 -431
rect -1311 -435 -1281 -409
rect -1215 -431 -1185 -409
rect -1425 -481 -1409 -447
rect -1375 -481 -1359 -447
rect -1425 -497 -1359 -481
rect -1233 -447 -1167 -431
rect -1119 -435 -1089 -409
rect -1023 -431 -993 -409
rect -1233 -481 -1217 -447
rect -1183 -481 -1167 -447
rect -1233 -497 -1167 -481
rect -1041 -447 -975 -431
rect -927 -435 -897 -409
rect -831 -431 -801 -409
rect -1041 -481 -1025 -447
rect -991 -481 -975 -447
rect -1041 -497 -975 -481
rect -849 -447 -783 -431
rect -735 -435 -705 -409
rect -639 -431 -609 -409
rect -849 -481 -833 -447
rect -799 -481 -783 -447
rect -849 -497 -783 -481
rect -657 -447 -591 -431
rect -543 -435 -513 -409
rect -447 -431 -417 -409
rect -657 -481 -641 -447
rect -607 -481 -591 -447
rect -657 -497 -591 -481
rect -465 -447 -399 -431
rect -351 -435 -321 -409
rect -255 -431 -225 -409
rect -465 -481 -449 -447
rect -415 -481 -399 -447
rect -465 -497 -399 -481
rect -273 -447 -207 -431
rect -159 -435 -129 -409
rect -63 -431 -33 -409
rect -273 -481 -257 -447
rect -223 -481 -207 -447
rect -273 -497 -207 -481
rect -81 -447 -15 -431
rect 33 -435 63 -409
rect 129 -431 159 -409
rect -81 -481 -65 -447
rect -31 -481 -15 -447
rect -81 -497 -15 -481
rect 111 -447 177 -431
rect 225 -435 255 -409
rect 321 -431 351 -409
rect 111 -481 127 -447
rect 161 -481 177 -447
rect 111 -497 177 -481
rect 303 -447 369 -431
rect 417 -435 447 -409
rect 513 -431 543 -409
rect 303 -481 319 -447
rect 353 -481 369 -447
rect 303 -497 369 -481
rect 495 -447 561 -431
rect 609 -435 639 -409
rect 705 -431 735 -409
rect 495 -481 511 -447
rect 545 -481 561 -447
rect 495 -497 561 -481
rect 687 -447 753 -431
rect 801 -435 831 -409
rect 897 -431 927 -409
rect 687 -481 703 -447
rect 737 -481 753 -447
rect 687 -497 753 -481
rect 879 -447 945 -431
rect 993 -435 1023 -409
rect 1089 -431 1119 -409
rect 879 -481 895 -447
rect 929 -481 945 -447
rect 879 -497 945 -481
rect 1071 -447 1137 -431
rect 1185 -435 1215 -409
rect 1281 -431 1311 -409
rect 1071 -481 1087 -447
rect 1121 -481 1137 -447
rect 1071 -497 1137 -481
rect 1263 -447 1329 -431
rect 1377 -435 1407 -409
rect 1473 -431 1503 -409
rect 1263 -481 1279 -447
rect 1313 -481 1329 -447
rect 1263 -497 1329 -481
rect 1455 -447 1521 -431
rect 1569 -435 1599 -409
rect 1665 -431 1695 -409
rect 1455 -481 1471 -447
rect 1505 -481 1521 -447
rect 1455 -497 1521 -481
rect 1647 -447 1713 -431
rect 1761 -435 1791 -409
rect 1857 -431 1887 -409
rect 1647 -481 1663 -447
rect 1697 -481 1713 -447
rect 1647 -497 1713 -481
rect 1839 -447 1905 -431
rect 1953 -435 1983 -409
rect 2049 -431 2079 -409
rect 1839 -481 1855 -447
rect 1889 -481 1905 -447
rect 1839 -497 1905 -481
rect 2031 -447 2097 -431
rect 2145 -435 2175 -409
rect 2241 -431 2271 -409
rect 2031 -481 2047 -447
rect 2081 -481 2097 -447
rect 2031 -497 2097 -481
rect 2223 -447 2289 -431
rect 2337 -435 2367 -409
rect 2433 -431 2463 -409
rect 2223 -481 2239 -447
rect 2273 -481 2289 -447
rect 2223 -497 2289 -481
rect 2415 -447 2481 -431
rect 2529 -435 2559 -409
rect 2625 -431 2655 -409
rect 2415 -481 2431 -447
rect 2465 -481 2481 -447
rect 2415 -497 2481 -481
rect 2607 -447 2673 -431
rect 2721 -435 2751 -409
rect 2817 -431 2847 -409
rect 2607 -481 2623 -447
rect 2657 -481 2673 -447
rect 2607 -497 2673 -481
rect 2799 -447 2865 -431
rect 2913 -435 2943 -409
rect 3009 -431 3039 -409
rect 2799 -481 2815 -447
rect 2849 -481 2865 -447
rect 2799 -497 2865 -481
rect 2991 -447 3057 -431
rect 3105 -435 3135 -409
rect 3201 -431 3231 -409
rect 2991 -481 3007 -447
rect 3041 -481 3057 -447
rect 2991 -497 3057 -481
rect 3183 -447 3249 -431
rect 3297 -435 3327 -409
rect 3393 -431 3423 -409
rect 3183 -481 3199 -447
rect 3233 -481 3249 -447
rect 3183 -497 3249 -481
rect 3375 -447 3441 -431
rect 3489 -435 3519 -409
rect 3585 -431 3615 -409
rect 3375 -481 3391 -447
rect 3425 -481 3441 -447
rect 3375 -497 3441 -481
rect 3567 -447 3633 -431
rect 3681 -435 3711 -409
rect 3777 -431 3807 -409
rect 3567 -481 3583 -447
rect 3617 -481 3633 -447
rect 3567 -497 3633 -481
rect 3759 -447 3825 -431
rect 3873 -435 3903 -409
rect 3969 -431 3999 -409
rect 3759 -481 3775 -447
rect 3809 -481 3825 -447
rect 3759 -497 3825 -481
rect 3951 -447 4017 -431
rect 4065 -435 4095 -409
rect 4161 -431 4191 -409
rect 3951 -481 3967 -447
rect 4001 -481 4017 -447
rect 3951 -497 4017 -481
rect 4143 -447 4209 -431
rect 4257 -435 4287 -409
rect 4353 -431 4383 -409
rect 4143 -481 4159 -447
rect 4193 -481 4209 -447
rect 4143 -497 4209 -481
rect 4335 -447 4401 -431
rect 4449 -435 4479 -409
rect 4545 -431 4575 -409
rect 4335 -481 4351 -447
rect 4385 -481 4401 -447
rect 4335 -497 4401 -481
rect 4527 -447 4593 -431
rect 4641 -435 4671 -409
rect 4737 -431 4767 -409
rect 4527 -481 4543 -447
rect 4577 -481 4593 -447
rect 4527 -497 4593 -481
rect 4719 -447 4785 -431
rect 4719 -481 4735 -447
rect 4769 -481 4785 -447
rect 4719 -497 4785 -481
rect -4689 -555 -4623 -539
rect -4689 -589 -4673 -555
rect -4639 -589 -4623 -555
rect -4767 -627 -4737 -601
rect -4689 -605 -4623 -589
rect -4497 -555 -4431 -539
rect -4497 -589 -4481 -555
rect -4447 -589 -4431 -555
rect -4671 -627 -4641 -605
rect -4575 -627 -4545 -601
rect -4497 -605 -4431 -589
rect -4305 -555 -4239 -539
rect -4305 -589 -4289 -555
rect -4255 -589 -4239 -555
rect -4479 -627 -4449 -605
rect -4383 -627 -4353 -601
rect -4305 -605 -4239 -589
rect -4113 -555 -4047 -539
rect -4113 -589 -4097 -555
rect -4063 -589 -4047 -555
rect -4287 -627 -4257 -605
rect -4191 -627 -4161 -601
rect -4113 -605 -4047 -589
rect -3921 -555 -3855 -539
rect -3921 -589 -3905 -555
rect -3871 -589 -3855 -555
rect -4095 -627 -4065 -605
rect -3999 -627 -3969 -601
rect -3921 -605 -3855 -589
rect -3729 -555 -3663 -539
rect -3729 -589 -3713 -555
rect -3679 -589 -3663 -555
rect -3903 -627 -3873 -605
rect -3807 -627 -3777 -601
rect -3729 -605 -3663 -589
rect -3537 -555 -3471 -539
rect -3537 -589 -3521 -555
rect -3487 -589 -3471 -555
rect -3711 -627 -3681 -605
rect -3615 -627 -3585 -601
rect -3537 -605 -3471 -589
rect -3345 -555 -3279 -539
rect -3345 -589 -3329 -555
rect -3295 -589 -3279 -555
rect -3519 -627 -3489 -605
rect -3423 -627 -3393 -601
rect -3345 -605 -3279 -589
rect -3153 -555 -3087 -539
rect -3153 -589 -3137 -555
rect -3103 -589 -3087 -555
rect -3327 -627 -3297 -605
rect -3231 -627 -3201 -601
rect -3153 -605 -3087 -589
rect -2961 -555 -2895 -539
rect -2961 -589 -2945 -555
rect -2911 -589 -2895 -555
rect -3135 -627 -3105 -605
rect -3039 -627 -3009 -601
rect -2961 -605 -2895 -589
rect -2769 -555 -2703 -539
rect -2769 -589 -2753 -555
rect -2719 -589 -2703 -555
rect -2943 -627 -2913 -605
rect -2847 -627 -2817 -601
rect -2769 -605 -2703 -589
rect -2577 -555 -2511 -539
rect -2577 -589 -2561 -555
rect -2527 -589 -2511 -555
rect -2751 -627 -2721 -605
rect -2655 -627 -2625 -601
rect -2577 -605 -2511 -589
rect -2385 -555 -2319 -539
rect -2385 -589 -2369 -555
rect -2335 -589 -2319 -555
rect -2559 -627 -2529 -605
rect -2463 -627 -2433 -601
rect -2385 -605 -2319 -589
rect -2193 -555 -2127 -539
rect -2193 -589 -2177 -555
rect -2143 -589 -2127 -555
rect -2367 -627 -2337 -605
rect -2271 -627 -2241 -601
rect -2193 -605 -2127 -589
rect -2001 -555 -1935 -539
rect -2001 -589 -1985 -555
rect -1951 -589 -1935 -555
rect -2175 -627 -2145 -605
rect -2079 -627 -2049 -601
rect -2001 -605 -1935 -589
rect -1809 -555 -1743 -539
rect -1809 -589 -1793 -555
rect -1759 -589 -1743 -555
rect -1983 -627 -1953 -605
rect -1887 -627 -1857 -601
rect -1809 -605 -1743 -589
rect -1617 -555 -1551 -539
rect -1617 -589 -1601 -555
rect -1567 -589 -1551 -555
rect -1791 -627 -1761 -605
rect -1695 -627 -1665 -601
rect -1617 -605 -1551 -589
rect -1425 -555 -1359 -539
rect -1425 -589 -1409 -555
rect -1375 -589 -1359 -555
rect -1599 -627 -1569 -605
rect -1503 -627 -1473 -601
rect -1425 -605 -1359 -589
rect -1233 -555 -1167 -539
rect -1233 -589 -1217 -555
rect -1183 -589 -1167 -555
rect -1407 -627 -1377 -605
rect -1311 -627 -1281 -601
rect -1233 -605 -1167 -589
rect -1041 -555 -975 -539
rect -1041 -589 -1025 -555
rect -991 -589 -975 -555
rect -1215 -627 -1185 -605
rect -1119 -627 -1089 -601
rect -1041 -605 -975 -589
rect -849 -555 -783 -539
rect -849 -589 -833 -555
rect -799 -589 -783 -555
rect -1023 -627 -993 -605
rect -927 -627 -897 -601
rect -849 -605 -783 -589
rect -657 -555 -591 -539
rect -657 -589 -641 -555
rect -607 -589 -591 -555
rect -831 -627 -801 -605
rect -735 -627 -705 -601
rect -657 -605 -591 -589
rect -465 -555 -399 -539
rect -465 -589 -449 -555
rect -415 -589 -399 -555
rect -639 -627 -609 -605
rect -543 -627 -513 -601
rect -465 -605 -399 -589
rect -273 -555 -207 -539
rect -273 -589 -257 -555
rect -223 -589 -207 -555
rect -447 -627 -417 -605
rect -351 -627 -321 -601
rect -273 -605 -207 -589
rect -81 -555 -15 -539
rect -81 -589 -65 -555
rect -31 -589 -15 -555
rect -255 -627 -225 -605
rect -159 -627 -129 -601
rect -81 -605 -15 -589
rect 111 -555 177 -539
rect 111 -589 127 -555
rect 161 -589 177 -555
rect -63 -627 -33 -605
rect 33 -627 63 -601
rect 111 -605 177 -589
rect 303 -555 369 -539
rect 303 -589 319 -555
rect 353 -589 369 -555
rect 129 -627 159 -605
rect 225 -627 255 -601
rect 303 -605 369 -589
rect 495 -555 561 -539
rect 495 -589 511 -555
rect 545 -589 561 -555
rect 321 -627 351 -605
rect 417 -627 447 -601
rect 495 -605 561 -589
rect 687 -555 753 -539
rect 687 -589 703 -555
rect 737 -589 753 -555
rect 513 -627 543 -605
rect 609 -627 639 -601
rect 687 -605 753 -589
rect 879 -555 945 -539
rect 879 -589 895 -555
rect 929 -589 945 -555
rect 705 -627 735 -605
rect 801 -627 831 -601
rect 879 -605 945 -589
rect 1071 -555 1137 -539
rect 1071 -589 1087 -555
rect 1121 -589 1137 -555
rect 897 -627 927 -605
rect 993 -627 1023 -601
rect 1071 -605 1137 -589
rect 1263 -555 1329 -539
rect 1263 -589 1279 -555
rect 1313 -589 1329 -555
rect 1089 -627 1119 -605
rect 1185 -627 1215 -601
rect 1263 -605 1329 -589
rect 1455 -555 1521 -539
rect 1455 -589 1471 -555
rect 1505 -589 1521 -555
rect 1281 -627 1311 -605
rect 1377 -627 1407 -601
rect 1455 -605 1521 -589
rect 1647 -555 1713 -539
rect 1647 -589 1663 -555
rect 1697 -589 1713 -555
rect 1473 -627 1503 -605
rect 1569 -627 1599 -601
rect 1647 -605 1713 -589
rect 1839 -555 1905 -539
rect 1839 -589 1855 -555
rect 1889 -589 1905 -555
rect 1665 -627 1695 -605
rect 1761 -627 1791 -601
rect 1839 -605 1905 -589
rect 2031 -555 2097 -539
rect 2031 -589 2047 -555
rect 2081 -589 2097 -555
rect 1857 -627 1887 -605
rect 1953 -627 1983 -601
rect 2031 -605 2097 -589
rect 2223 -555 2289 -539
rect 2223 -589 2239 -555
rect 2273 -589 2289 -555
rect 2049 -627 2079 -605
rect 2145 -627 2175 -601
rect 2223 -605 2289 -589
rect 2415 -555 2481 -539
rect 2415 -589 2431 -555
rect 2465 -589 2481 -555
rect 2241 -627 2271 -605
rect 2337 -627 2367 -601
rect 2415 -605 2481 -589
rect 2607 -555 2673 -539
rect 2607 -589 2623 -555
rect 2657 -589 2673 -555
rect 2433 -627 2463 -605
rect 2529 -627 2559 -601
rect 2607 -605 2673 -589
rect 2799 -555 2865 -539
rect 2799 -589 2815 -555
rect 2849 -589 2865 -555
rect 2625 -627 2655 -605
rect 2721 -627 2751 -601
rect 2799 -605 2865 -589
rect 2991 -555 3057 -539
rect 2991 -589 3007 -555
rect 3041 -589 3057 -555
rect 2817 -627 2847 -605
rect 2913 -627 2943 -601
rect 2991 -605 3057 -589
rect 3183 -555 3249 -539
rect 3183 -589 3199 -555
rect 3233 -589 3249 -555
rect 3009 -627 3039 -605
rect 3105 -627 3135 -601
rect 3183 -605 3249 -589
rect 3375 -555 3441 -539
rect 3375 -589 3391 -555
rect 3425 -589 3441 -555
rect 3201 -627 3231 -605
rect 3297 -627 3327 -601
rect 3375 -605 3441 -589
rect 3567 -555 3633 -539
rect 3567 -589 3583 -555
rect 3617 -589 3633 -555
rect 3393 -627 3423 -605
rect 3489 -627 3519 -601
rect 3567 -605 3633 -589
rect 3759 -555 3825 -539
rect 3759 -589 3775 -555
rect 3809 -589 3825 -555
rect 3585 -627 3615 -605
rect 3681 -627 3711 -601
rect 3759 -605 3825 -589
rect 3951 -555 4017 -539
rect 3951 -589 3967 -555
rect 4001 -589 4017 -555
rect 3777 -627 3807 -605
rect 3873 -627 3903 -601
rect 3951 -605 4017 -589
rect 4143 -555 4209 -539
rect 4143 -589 4159 -555
rect 4193 -589 4209 -555
rect 3969 -627 3999 -605
rect 4065 -627 4095 -601
rect 4143 -605 4209 -589
rect 4335 -555 4401 -539
rect 4335 -589 4351 -555
rect 4385 -589 4401 -555
rect 4161 -627 4191 -605
rect 4257 -627 4287 -601
rect 4335 -605 4401 -589
rect 4527 -555 4593 -539
rect 4527 -589 4543 -555
rect 4577 -589 4593 -555
rect 4353 -627 4383 -605
rect 4449 -627 4479 -601
rect 4527 -605 4593 -589
rect 4719 -555 4785 -539
rect 4719 -589 4735 -555
rect 4769 -589 4785 -555
rect 4545 -627 4575 -605
rect 4641 -627 4671 -601
rect 4719 -605 4785 -589
rect 4737 -627 4767 -605
rect -4767 -949 -4737 -927
rect -4785 -965 -4719 -949
rect -4671 -953 -4641 -927
rect -4575 -949 -4545 -927
rect -4785 -999 -4769 -965
rect -4735 -999 -4719 -965
rect -4785 -1015 -4719 -999
rect -4593 -965 -4527 -949
rect -4479 -953 -4449 -927
rect -4383 -949 -4353 -927
rect -4593 -999 -4577 -965
rect -4543 -999 -4527 -965
rect -4593 -1015 -4527 -999
rect -4401 -965 -4335 -949
rect -4287 -953 -4257 -927
rect -4191 -949 -4161 -927
rect -4401 -999 -4385 -965
rect -4351 -999 -4335 -965
rect -4401 -1015 -4335 -999
rect -4209 -965 -4143 -949
rect -4095 -953 -4065 -927
rect -3999 -949 -3969 -927
rect -4209 -999 -4193 -965
rect -4159 -999 -4143 -965
rect -4209 -1015 -4143 -999
rect -4017 -965 -3951 -949
rect -3903 -953 -3873 -927
rect -3807 -949 -3777 -927
rect -4017 -999 -4001 -965
rect -3967 -999 -3951 -965
rect -4017 -1015 -3951 -999
rect -3825 -965 -3759 -949
rect -3711 -953 -3681 -927
rect -3615 -949 -3585 -927
rect -3825 -999 -3809 -965
rect -3775 -999 -3759 -965
rect -3825 -1015 -3759 -999
rect -3633 -965 -3567 -949
rect -3519 -953 -3489 -927
rect -3423 -949 -3393 -927
rect -3633 -999 -3617 -965
rect -3583 -999 -3567 -965
rect -3633 -1015 -3567 -999
rect -3441 -965 -3375 -949
rect -3327 -953 -3297 -927
rect -3231 -949 -3201 -927
rect -3441 -999 -3425 -965
rect -3391 -999 -3375 -965
rect -3441 -1015 -3375 -999
rect -3249 -965 -3183 -949
rect -3135 -953 -3105 -927
rect -3039 -949 -3009 -927
rect -3249 -999 -3233 -965
rect -3199 -999 -3183 -965
rect -3249 -1015 -3183 -999
rect -3057 -965 -2991 -949
rect -2943 -953 -2913 -927
rect -2847 -949 -2817 -927
rect -3057 -999 -3041 -965
rect -3007 -999 -2991 -965
rect -3057 -1015 -2991 -999
rect -2865 -965 -2799 -949
rect -2751 -953 -2721 -927
rect -2655 -949 -2625 -927
rect -2865 -999 -2849 -965
rect -2815 -999 -2799 -965
rect -2865 -1015 -2799 -999
rect -2673 -965 -2607 -949
rect -2559 -953 -2529 -927
rect -2463 -949 -2433 -927
rect -2673 -999 -2657 -965
rect -2623 -999 -2607 -965
rect -2673 -1015 -2607 -999
rect -2481 -965 -2415 -949
rect -2367 -953 -2337 -927
rect -2271 -949 -2241 -927
rect -2481 -999 -2465 -965
rect -2431 -999 -2415 -965
rect -2481 -1015 -2415 -999
rect -2289 -965 -2223 -949
rect -2175 -953 -2145 -927
rect -2079 -949 -2049 -927
rect -2289 -999 -2273 -965
rect -2239 -999 -2223 -965
rect -2289 -1015 -2223 -999
rect -2097 -965 -2031 -949
rect -1983 -953 -1953 -927
rect -1887 -949 -1857 -927
rect -2097 -999 -2081 -965
rect -2047 -999 -2031 -965
rect -2097 -1015 -2031 -999
rect -1905 -965 -1839 -949
rect -1791 -953 -1761 -927
rect -1695 -949 -1665 -927
rect -1905 -999 -1889 -965
rect -1855 -999 -1839 -965
rect -1905 -1015 -1839 -999
rect -1713 -965 -1647 -949
rect -1599 -953 -1569 -927
rect -1503 -949 -1473 -927
rect -1713 -999 -1697 -965
rect -1663 -999 -1647 -965
rect -1713 -1015 -1647 -999
rect -1521 -965 -1455 -949
rect -1407 -953 -1377 -927
rect -1311 -949 -1281 -927
rect -1521 -999 -1505 -965
rect -1471 -999 -1455 -965
rect -1521 -1015 -1455 -999
rect -1329 -965 -1263 -949
rect -1215 -953 -1185 -927
rect -1119 -949 -1089 -927
rect -1329 -999 -1313 -965
rect -1279 -999 -1263 -965
rect -1329 -1015 -1263 -999
rect -1137 -965 -1071 -949
rect -1023 -953 -993 -927
rect -927 -949 -897 -927
rect -1137 -999 -1121 -965
rect -1087 -999 -1071 -965
rect -1137 -1015 -1071 -999
rect -945 -965 -879 -949
rect -831 -953 -801 -927
rect -735 -949 -705 -927
rect -945 -999 -929 -965
rect -895 -999 -879 -965
rect -945 -1015 -879 -999
rect -753 -965 -687 -949
rect -639 -953 -609 -927
rect -543 -949 -513 -927
rect -753 -999 -737 -965
rect -703 -999 -687 -965
rect -753 -1015 -687 -999
rect -561 -965 -495 -949
rect -447 -953 -417 -927
rect -351 -949 -321 -927
rect -561 -999 -545 -965
rect -511 -999 -495 -965
rect -561 -1015 -495 -999
rect -369 -965 -303 -949
rect -255 -953 -225 -927
rect -159 -949 -129 -927
rect -369 -999 -353 -965
rect -319 -999 -303 -965
rect -369 -1015 -303 -999
rect -177 -965 -111 -949
rect -63 -953 -33 -927
rect 33 -949 63 -927
rect -177 -999 -161 -965
rect -127 -999 -111 -965
rect -177 -1015 -111 -999
rect 15 -965 81 -949
rect 129 -953 159 -927
rect 225 -949 255 -927
rect 15 -999 31 -965
rect 65 -999 81 -965
rect 15 -1015 81 -999
rect 207 -965 273 -949
rect 321 -953 351 -927
rect 417 -949 447 -927
rect 207 -999 223 -965
rect 257 -999 273 -965
rect 207 -1015 273 -999
rect 399 -965 465 -949
rect 513 -953 543 -927
rect 609 -949 639 -927
rect 399 -999 415 -965
rect 449 -999 465 -965
rect 399 -1015 465 -999
rect 591 -965 657 -949
rect 705 -953 735 -927
rect 801 -949 831 -927
rect 591 -999 607 -965
rect 641 -999 657 -965
rect 591 -1015 657 -999
rect 783 -965 849 -949
rect 897 -953 927 -927
rect 993 -949 1023 -927
rect 783 -999 799 -965
rect 833 -999 849 -965
rect 783 -1015 849 -999
rect 975 -965 1041 -949
rect 1089 -953 1119 -927
rect 1185 -949 1215 -927
rect 975 -999 991 -965
rect 1025 -999 1041 -965
rect 975 -1015 1041 -999
rect 1167 -965 1233 -949
rect 1281 -953 1311 -927
rect 1377 -949 1407 -927
rect 1167 -999 1183 -965
rect 1217 -999 1233 -965
rect 1167 -1015 1233 -999
rect 1359 -965 1425 -949
rect 1473 -953 1503 -927
rect 1569 -949 1599 -927
rect 1359 -999 1375 -965
rect 1409 -999 1425 -965
rect 1359 -1015 1425 -999
rect 1551 -965 1617 -949
rect 1665 -953 1695 -927
rect 1761 -949 1791 -927
rect 1551 -999 1567 -965
rect 1601 -999 1617 -965
rect 1551 -1015 1617 -999
rect 1743 -965 1809 -949
rect 1857 -953 1887 -927
rect 1953 -949 1983 -927
rect 1743 -999 1759 -965
rect 1793 -999 1809 -965
rect 1743 -1015 1809 -999
rect 1935 -965 2001 -949
rect 2049 -953 2079 -927
rect 2145 -949 2175 -927
rect 1935 -999 1951 -965
rect 1985 -999 2001 -965
rect 1935 -1015 2001 -999
rect 2127 -965 2193 -949
rect 2241 -953 2271 -927
rect 2337 -949 2367 -927
rect 2127 -999 2143 -965
rect 2177 -999 2193 -965
rect 2127 -1015 2193 -999
rect 2319 -965 2385 -949
rect 2433 -953 2463 -927
rect 2529 -949 2559 -927
rect 2319 -999 2335 -965
rect 2369 -999 2385 -965
rect 2319 -1015 2385 -999
rect 2511 -965 2577 -949
rect 2625 -953 2655 -927
rect 2721 -949 2751 -927
rect 2511 -999 2527 -965
rect 2561 -999 2577 -965
rect 2511 -1015 2577 -999
rect 2703 -965 2769 -949
rect 2817 -953 2847 -927
rect 2913 -949 2943 -927
rect 2703 -999 2719 -965
rect 2753 -999 2769 -965
rect 2703 -1015 2769 -999
rect 2895 -965 2961 -949
rect 3009 -953 3039 -927
rect 3105 -949 3135 -927
rect 2895 -999 2911 -965
rect 2945 -999 2961 -965
rect 2895 -1015 2961 -999
rect 3087 -965 3153 -949
rect 3201 -953 3231 -927
rect 3297 -949 3327 -927
rect 3087 -999 3103 -965
rect 3137 -999 3153 -965
rect 3087 -1015 3153 -999
rect 3279 -965 3345 -949
rect 3393 -953 3423 -927
rect 3489 -949 3519 -927
rect 3279 -999 3295 -965
rect 3329 -999 3345 -965
rect 3279 -1015 3345 -999
rect 3471 -965 3537 -949
rect 3585 -953 3615 -927
rect 3681 -949 3711 -927
rect 3471 -999 3487 -965
rect 3521 -999 3537 -965
rect 3471 -1015 3537 -999
rect 3663 -965 3729 -949
rect 3777 -953 3807 -927
rect 3873 -949 3903 -927
rect 3663 -999 3679 -965
rect 3713 -999 3729 -965
rect 3663 -1015 3729 -999
rect 3855 -965 3921 -949
rect 3969 -953 3999 -927
rect 4065 -949 4095 -927
rect 3855 -999 3871 -965
rect 3905 -999 3921 -965
rect 3855 -1015 3921 -999
rect 4047 -965 4113 -949
rect 4161 -953 4191 -927
rect 4257 -949 4287 -927
rect 4047 -999 4063 -965
rect 4097 -999 4113 -965
rect 4047 -1015 4113 -999
rect 4239 -965 4305 -949
rect 4353 -953 4383 -927
rect 4449 -949 4479 -927
rect 4239 -999 4255 -965
rect 4289 -999 4305 -965
rect 4239 -1015 4305 -999
rect 4431 -965 4497 -949
rect 4545 -953 4575 -927
rect 4641 -949 4671 -927
rect 4431 -999 4447 -965
rect 4481 -999 4497 -965
rect 4431 -1015 4497 -999
rect 4623 -965 4689 -949
rect 4737 -953 4767 -927
rect 4623 -999 4639 -965
rect 4673 -999 4689 -965
rect 4623 -1015 4689 -999
<< polycont >>
rect -4769 965 -4735 999
rect -4577 965 -4543 999
rect -4385 965 -4351 999
rect -4193 965 -4159 999
rect -4001 965 -3967 999
rect -3809 965 -3775 999
rect -3617 965 -3583 999
rect -3425 965 -3391 999
rect -3233 965 -3199 999
rect -3041 965 -3007 999
rect -2849 965 -2815 999
rect -2657 965 -2623 999
rect -2465 965 -2431 999
rect -2273 965 -2239 999
rect -2081 965 -2047 999
rect -1889 965 -1855 999
rect -1697 965 -1663 999
rect -1505 965 -1471 999
rect -1313 965 -1279 999
rect -1121 965 -1087 999
rect -929 965 -895 999
rect -737 965 -703 999
rect -545 965 -511 999
rect -353 965 -319 999
rect -161 965 -127 999
rect 31 965 65 999
rect 223 965 257 999
rect 415 965 449 999
rect 607 965 641 999
rect 799 965 833 999
rect 991 965 1025 999
rect 1183 965 1217 999
rect 1375 965 1409 999
rect 1567 965 1601 999
rect 1759 965 1793 999
rect 1951 965 1985 999
rect 2143 965 2177 999
rect 2335 965 2369 999
rect 2527 965 2561 999
rect 2719 965 2753 999
rect 2911 965 2945 999
rect 3103 965 3137 999
rect 3295 965 3329 999
rect 3487 965 3521 999
rect 3679 965 3713 999
rect 3871 965 3905 999
rect 4063 965 4097 999
rect 4255 965 4289 999
rect 4447 965 4481 999
rect 4639 965 4673 999
rect -4673 555 -4639 589
rect -4481 555 -4447 589
rect -4289 555 -4255 589
rect -4097 555 -4063 589
rect -3905 555 -3871 589
rect -3713 555 -3679 589
rect -3521 555 -3487 589
rect -3329 555 -3295 589
rect -3137 555 -3103 589
rect -2945 555 -2911 589
rect -2753 555 -2719 589
rect -2561 555 -2527 589
rect -2369 555 -2335 589
rect -2177 555 -2143 589
rect -1985 555 -1951 589
rect -1793 555 -1759 589
rect -1601 555 -1567 589
rect -1409 555 -1375 589
rect -1217 555 -1183 589
rect -1025 555 -991 589
rect -833 555 -799 589
rect -641 555 -607 589
rect -449 555 -415 589
rect -257 555 -223 589
rect -65 555 -31 589
rect 127 555 161 589
rect 319 555 353 589
rect 511 555 545 589
rect 703 555 737 589
rect 895 555 929 589
rect 1087 555 1121 589
rect 1279 555 1313 589
rect 1471 555 1505 589
rect 1663 555 1697 589
rect 1855 555 1889 589
rect 2047 555 2081 589
rect 2239 555 2273 589
rect 2431 555 2465 589
rect 2623 555 2657 589
rect 2815 555 2849 589
rect 3007 555 3041 589
rect 3199 555 3233 589
rect 3391 555 3425 589
rect 3583 555 3617 589
rect 3775 555 3809 589
rect 3967 555 4001 589
rect 4159 555 4193 589
rect 4351 555 4385 589
rect 4543 555 4577 589
rect 4735 555 4769 589
rect -4673 447 -4639 481
rect -4481 447 -4447 481
rect -4289 447 -4255 481
rect -4097 447 -4063 481
rect -3905 447 -3871 481
rect -3713 447 -3679 481
rect -3521 447 -3487 481
rect -3329 447 -3295 481
rect -3137 447 -3103 481
rect -2945 447 -2911 481
rect -2753 447 -2719 481
rect -2561 447 -2527 481
rect -2369 447 -2335 481
rect -2177 447 -2143 481
rect -1985 447 -1951 481
rect -1793 447 -1759 481
rect -1601 447 -1567 481
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect 1663 447 1697 481
rect 1855 447 1889 481
rect 2047 447 2081 481
rect 2239 447 2273 481
rect 2431 447 2465 481
rect 2623 447 2657 481
rect 2815 447 2849 481
rect 3007 447 3041 481
rect 3199 447 3233 481
rect 3391 447 3425 481
rect 3583 447 3617 481
rect 3775 447 3809 481
rect 3967 447 4001 481
rect 4159 447 4193 481
rect 4351 447 4385 481
rect 4543 447 4577 481
rect 4735 447 4769 481
rect -4769 37 -4735 71
rect -4577 37 -4543 71
rect -4385 37 -4351 71
rect -4193 37 -4159 71
rect -4001 37 -3967 71
rect -3809 37 -3775 71
rect -3617 37 -3583 71
rect -3425 37 -3391 71
rect -3233 37 -3199 71
rect -3041 37 -3007 71
rect -2849 37 -2815 71
rect -2657 37 -2623 71
rect -2465 37 -2431 71
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect 2527 37 2561 71
rect 2719 37 2753 71
rect 2911 37 2945 71
rect 3103 37 3137 71
rect 3295 37 3329 71
rect 3487 37 3521 71
rect 3679 37 3713 71
rect 3871 37 3905 71
rect 4063 37 4097 71
rect 4255 37 4289 71
rect 4447 37 4481 71
rect 4639 37 4673 71
rect -4769 -71 -4735 -37
rect -4577 -71 -4543 -37
rect -4385 -71 -4351 -37
rect -4193 -71 -4159 -37
rect -4001 -71 -3967 -37
rect -3809 -71 -3775 -37
rect -3617 -71 -3583 -37
rect -3425 -71 -3391 -37
rect -3233 -71 -3199 -37
rect -3041 -71 -3007 -37
rect -2849 -71 -2815 -37
rect -2657 -71 -2623 -37
rect -2465 -71 -2431 -37
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect 2527 -71 2561 -37
rect 2719 -71 2753 -37
rect 2911 -71 2945 -37
rect 3103 -71 3137 -37
rect 3295 -71 3329 -37
rect 3487 -71 3521 -37
rect 3679 -71 3713 -37
rect 3871 -71 3905 -37
rect 4063 -71 4097 -37
rect 4255 -71 4289 -37
rect 4447 -71 4481 -37
rect 4639 -71 4673 -37
rect -4673 -481 -4639 -447
rect -4481 -481 -4447 -447
rect -4289 -481 -4255 -447
rect -4097 -481 -4063 -447
rect -3905 -481 -3871 -447
rect -3713 -481 -3679 -447
rect -3521 -481 -3487 -447
rect -3329 -481 -3295 -447
rect -3137 -481 -3103 -447
rect -2945 -481 -2911 -447
rect -2753 -481 -2719 -447
rect -2561 -481 -2527 -447
rect -2369 -481 -2335 -447
rect -2177 -481 -2143 -447
rect -1985 -481 -1951 -447
rect -1793 -481 -1759 -447
rect -1601 -481 -1567 -447
rect -1409 -481 -1375 -447
rect -1217 -481 -1183 -447
rect -1025 -481 -991 -447
rect -833 -481 -799 -447
rect -641 -481 -607 -447
rect -449 -481 -415 -447
rect -257 -481 -223 -447
rect -65 -481 -31 -447
rect 127 -481 161 -447
rect 319 -481 353 -447
rect 511 -481 545 -447
rect 703 -481 737 -447
rect 895 -481 929 -447
rect 1087 -481 1121 -447
rect 1279 -481 1313 -447
rect 1471 -481 1505 -447
rect 1663 -481 1697 -447
rect 1855 -481 1889 -447
rect 2047 -481 2081 -447
rect 2239 -481 2273 -447
rect 2431 -481 2465 -447
rect 2623 -481 2657 -447
rect 2815 -481 2849 -447
rect 3007 -481 3041 -447
rect 3199 -481 3233 -447
rect 3391 -481 3425 -447
rect 3583 -481 3617 -447
rect 3775 -481 3809 -447
rect 3967 -481 4001 -447
rect 4159 -481 4193 -447
rect 4351 -481 4385 -447
rect 4543 -481 4577 -447
rect 4735 -481 4769 -447
rect -4673 -589 -4639 -555
rect -4481 -589 -4447 -555
rect -4289 -589 -4255 -555
rect -4097 -589 -4063 -555
rect -3905 -589 -3871 -555
rect -3713 -589 -3679 -555
rect -3521 -589 -3487 -555
rect -3329 -589 -3295 -555
rect -3137 -589 -3103 -555
rect -2945 -589 -2911 -555
rect -2753 -589 -2719 -555
rect -2561 -589 -2527 -555
rect -2369 -589 -2335 -555
rect -2177 -589 -2143 -555
rect -1985 -589 -1951 -555
rect -1793 -589 -1759 -555
rect -1601 -589 -1567 -555
rect -1409 -589 -1375 -555
rect -1217 -589 -1183 -555
rect -1025 -589 -991 -555
rect -833 -589 -799 -555
rect -641 -589 -607 -555
rect -449 -589 -415 -555
rect -257 -589 -223 -555
rect -65 -589 -31 -555
rect 127 -589 161 -555
rect 319 -589 353 -555
rect 511 -589 545 -555
rect 703 -589 737 -555
rect 895 -589 929 -555
rect 1087 -589 1121 -555
rect 1279 -589 1313 -555
rect 1471 -589 1505 -555
rect 1663 -589 1697 -555
rect 1855 -589 1889 -555
rect 2047 -589 2081 -555
rect 2239 -589 2273 -555
rect 2431 -589 2465 -555
rect 2623 -589 2657 -555
rect 2815 -589 2849 -555
rect 3007 -589 3041 -555
rect 3199 -589 3233 -555
rect 3391 -589 3425 -555
rect 3583 -589 3617 -555
rect 3775 -589 3809 -555
rect 3967 -589 4001 -555
rect 4159 -589 4193 -555
rect 4351 -589 4385 -555
rect 4543 -589 4577 -555
rect 4735 -589 4769 -555
rect -4769 -999 -4735 -965
rect -4577 -999 -4543 -965
rect -4385 -999 -4351 -965
rect -4193 -999 -4159 -965
rect -4001 -999 -3967 -965
rect -3809 -999 -3775 -965
rect -3617 -999 -3583 -965
rect -3425 -999 -3391 -965
rect -3233 -999 -3199 -965
rect -3041 -999 -3007 -965
rect -2849 -999 -2815 -965
rect -2657 -999 -2623 -965
rect -2465 -999 -2431 -965
rect -2273 -999 -2239 -965
rect -2081 -999 -2047 -965
rect -1889 -999 -1855 -965
rect -1697 -999 -1663 -965
rect -1505 -999 -1471 -965
rect -1313 -999 -1279 -965
rect -1121 -999 -1087 -965
rect -929 -999 -895 -965
rect -737 -999 -703 -965
rect -545 -999 -511 -965
rect -353 -999 -319 -965
rect -161 -999 -127 -965
rect 31 -999 65 -965
rect 223 -999 257 -965
rect 415 -999 449 -965
rect 607 -999 641 -965
rect 799 -999 833 -965
rect 991 -999 1025 -965
rect 1183 -999 1217 -965
rect 1375 -999 1409 -965
rect 1567 -999 1601 -965
rect 1759 -999 1793 -965
rect 1951 -999 1985 -965
rect 2143 -999 2177 -965
rect 2335 -999 2369 -965
rect 2527 -999 2561 -965
rect 2719 -999 2753 -965
rect 2911 -999 2945 -965
rect 3103 -999 3137 -965
rect 3295 -999 3329 -965
rect 3487 -999 3521 -965
rect 3679 -999 3713 -965
rect 3871 -999 3905 -965
rect 4063 -999 4097 -965
rect 4255 -999 4289 -965
rect 4447 -999 4481 -965
rect 4639 -999 4673 -965
<< locali >>
rect -4931 1067 -4835 1101
rect 4835 1067 4931 1101
rect -4931 1005 -4897 1067
rect 4897 1005 4931 1067
rect -4785 965 -4769 999
rect -4735 965 -4719 999
rect -4593 965 -4577 999
rect -4543 965 -4527 999
rect -4401 965 -4385 999
rect -4351 965 -4335 999
rect -4209 965 -4193 999
rect -4159 965 -4143 999
rect -4017 965 -4001 999
rect -3967 965 -3951 999
rect -3825 965 -3809 999
rect -3775 965 -3759 999
rect -3633 965 -3617 999
rect -3583 965 -3567 999
rect -3441 965 -3425 999
rect -3391 965 -3375 999
rect -3249 965 -3233 999
rect -3199 965 -3183 999
rect -3057 965 -3041 999
rect -3007 965 -2991 999
rect -2865 965 -2849 999
rect -2815 965 -2799 999
rect -2673 965 -2657 999
rect -2623 965 -2607 999
rect -2481 965 -2465 999
rect -2431 965 -2415 999
rect -2289 965 -2273 999
rect -2239 965 -2223 999
rect -2097 965 -2081 999
rect -2047 965 -2031 999
rect -1905 965 -1889 999
rect -1855 965 -1839 999
rect -1713 965 -1697 999
rect -1663 965 -1647 999
rect -1521 965 -1505 999
rect -1471 965 -1455 999
rect -1329 965 -1313 999
rect -1279 965 -1263 999
rect -1137 965 -1121 999
rect -1087 965 -1071 999
rect -945 965 -929 999
rect -895 965 -879 999
rect -753 965 -737 999
rect -703 965 -687 999
rect -561 965 -545 999
rect -511 965 -495 999
rect -369 965 -353 999
rect -319 965 -303 999
rect -177 965 -161 999
rect -127 965 -111 999
rect 15 965 31 999
rect 65 965 81 999
rect 207 965 223 999
rect 257 965 273 999
rect 399 965 415 999
rect 449 965 465 999
rect 591 965 607 999
rect 641 965 657 999
rect 783 965 799 999
rect 833 965 849 999
rect 975 965 991 999
rect 1025 965 1041 999
rect 1167 965 1183 999
rect 1217 965 1233 999
rect 1359 965 1375 999
rect 1409 965 1425 999
rect 1551 965 1567 999
rect 1601 965 1617 999
rect 1743 965 1759 999
rect 1793 965 1809 999
rect 1935 965 1951 999
rect 1985 965 2001 999
rect 2127 965 2143 999
rect 2177 965 2193 999
rect 2319 965 2335 999
rect 2369 965 2385 999
rect 2511 965 2527 999
rect 2561 965 2577 999
rect 2703 965 2719 999
rect 2753 965 2769 999
rect 2895 965 2911 999
rect 2945 965 2961 999
rect 3087 965 3103 999
rect 3137 965 3153 999
rect 3279 965 3295 999
rect 3329 965 3345 999
rect 3471 965 3487 999
rect 3521 965 3537 999
rect 3663 965 3679 999
rect 3713 965 3729 999
rect 3855 965 3871 999
rect 3905 965 3921 999
rect 4047 965 4063 999
rect 4097 965 4113 999
rect 4239 965 4255 999
rect 4289 965 4305 999
rect 4431 965 4447 999
rect 4481 965 4497 999
rect 4623 965 4639 999
rect 4673 965 4689 999
rect -4817 915 -4783 931
rect -4817 623 -4783 639
rect -4721 915 -4687 931
rect -4721 623 -4687 639
rect -4625 915 -4591 931
rect -4625 623 -4591 639
rect -4529 915 -4495 931
rect -4529 623 -4495 639
rect -4433 915 -4399 931
rect -4433 623 -4399 639
rect -4337 915 -4303 931
rect -4337 623 -4303 639
rect -4241 915 -4207 931
rect -4241 623 -4207 639
rect -4145 915 -4111 931
rect -4145 623 -4111 639
rect -4049 915 -4015 931
rect -4049 623 -4015 639
rect -3953 915 -3919 931
rect -3953 623 -3919 639
rect -3857 915 -3823 931
rect -3857 623 -3823 639
rect -3761 915 -3727 931
rect -3761 623 -3727 639
rect -3665 915 -3631 931
rect -3665 623 -3631 639
rect -3569 915 -3535 931
rect -3569 623 -3535 639
rect -3473 915 -3439 931
rect -3473 623 -3439 639
rect -3377 915 -3343 931
rect -3377 623 -3343 639
rect -3281 915 -3247 931
rect -3281 623 -3247 639
rect -3185 915 -3151 931
rect -3185 623 -3151 639
rect -3089 915 -3055 931
rect -3089 623 -3055 639
rect -2993 915 -2959 931
rect -2993 623 -2959 639
rect -2897 915 -2863 931
rect -2897 623 -2863 639
rect -2801 915 -2767 931
rect -2801 623 -2767 639
rect -2705 915 -2671 931
rect -2705 623 -2671 639
rect -2609 915 -2575 931
rect -2609 623 -2575 639
rect -2513 915 -2479 931
rect -2513 623 -2479 639
rect -2417 915 -2383 931
rect -2417 623 -2383 639
rect -2321 915 -2287 931
rect -2321 623 -2287 639
rect -2225 915 -2191 931
rect -2225 623 -2191 639
rect -2129 915 -2095 931
rect -2129 623 -2095 639
rect -2033 915 -1999 931
rect -2033 623 -1999 639
rect -1937 915 -1903 931
rect -1937 623 -1903 639
rect -1841 915 -1807 931
rect -1841 623 -1807 639
rect -1745 915 -1711 931
rect -1745 623 -1711 639
rect -1649 915 -1615 931
rect -1649 623 -1615 639
rect -1553 915 -1519 931
rect -1553 623 -1519 639
rect -1457 915 -1423 931
rect -1457 623 -1423 639
rect -1361 915 -1327 931
rect -1361 623 -1327 639
rect -1265 915 -1231 931
rect -1265 623 -1231 639
rect -1169 915 -1135 931
rect -1169 623 -1135 639
rect -1073 915 -1039 931
rect -1073 623 -1039 639
rect -977 915 -943 931
rect -977 623 -943 639
rect -881 915 -847 931
rect -881 623 -847 639
rect -785 915 -751 931
rect -785 623 -751 639
rect -689 915 -655 931
rect -689 623 -655 639
rect -593 915 -559 931
rect -593 623 -559 639
rect -497 915 -463 931
rect -497 623 -463 639
rect -401 915 -367 931
rect -401 623 -367 639
rect -305 915 -271 931
rect -305 623 -271 639
rect -209 915 -175 931
rect -209 623 -175 639
rect -113 915 -79 931
rect -113 623 -79 639
rect -17 915 17 931
rect -17 623 17 639
rect 79 915 113 931
rect 79 623 113 639
rect 175 915 209 931
rect 175 623 209 639
rect 271 915 305 931
rect 271 623 305 639
rect 367 915 401 931
rect 367 623 401 639
rect 463 915 497 931
rect 463 623 497 639
rect 559 915 593 931
rect 559 623 593 639
rect 655 915 689 931
rect 655 623 689 639
rect 751 915 785 931
rect 751 623 785 639
rect 847 915 881 931
rect 847 623 881 639
rect 943 915 977 931
rect 943 623 977 639
rect 1039 915 1073 931
rect 1039 623 1073 639
rect 1135 915 1169 931
rect 1135 623 1169 639
rect 1231 915 1265 931
rect 1231 623 1265 639
rect 1327 915 1361 931
rect 1327 623 1361 639
rect 1423 915 1457 931
rect 1423 623 1457 639
rect 1519 915 1553 931
rect 1519 623 1553 639
rect 1615 915 1649 931
rect 1615 623 1649 639
rect 1711 915 1745 931
rect 1711 623 1745 639
rect 1807 915 1841 931
rect 1807 623 1841 639
rect 1903 915 1937 931
rect 1903 623 1937 639
rect 1999 915 2033 931
rect 1999 623 2033 639
rect 2095 915 2129 931
rect 2095 623 2129 639
rect 2191 915 2225 931
rect 2191 623 2225 639
rect 2287 915 2321 931
rect 2287 623 2321 639
rect 2383 915 2417 931
rect 2383 623 2417 639
rect 2479 915 2513 931
rect 2479 623 2513 639
rect 2575 915 2609 931
rect 2575 623 2609 639
rect 2671 915 2705 931
rect 2671 623 2705 639
rect 2767 915 2801 931
rect 2767 623 2801 639
rect 2863 915 2897 931
rect 2863 623 2897 639
rect 2959 915 2993 931
rect 2959 623 2993 639
rect 3055 915 3089 931
rect 3055 623 3089 639
rect 3151 915 3185 931
rect 3151 623 3185 639
rect 3247 915 3281 931
rect 3247 623 3281 639
rect 3343 915 3377 931
rect 3343 623 3377 639
rect 3439 915 3473 931
rect 3439 623 3473 639
rect 3535 915 3569 931
rect 3535 623 3569 639
rect 3631 915 3665 931
rect 3631 623 3665 639
rect 3727 915 3761 931
rect 3727 623 3761 639
rect 3823 915 3857 931
rect 3823 623 3857 639
rect 3919 915 3953 931
rect 3919 623 3953 639
rect 4015 915 4049 931
rect 4015 623 4049 639
rect 4111 915 4145 931
rect 4111 623 4145 639
rect 4207 915 4241 931
rect 4207 623 4241 639
rect 4303 915 4337 931
rect 4303 623 4337 639
rect 4399 915 4433 931
rect 4399 623 4433 639
rect 4495 915 4529 931
rect 4495 623 4529 639
rect 4591 915 4625 931
rect 4591 623 4625 639
rect 4687 915 4721 931
rect 4687 623 4721 639
rect 4783 915 4817 931
rect 4783 623 4817 639
rect -4689 555 -4673 589
rect -4639 555 -4623 589
rect -4497 555 -4481 589
rect -4447 555 -4431 589
rect -4305 555 -4289 589
rect -4255 555 -4239 589
rect -4113 555 -4097 589
rect -4063 555 -4047 589
rect -3921 555 -3905 589
rect -3871 555 -3855 589
rect -3729 555 -3713 589
rect -3679 555 -3663 589
rect -3537 555 -3521 589
rect -3487 555 -3471 589
rect -3345 555 -3329 589
rect -3295 555 -3279 589
rect -3153 555 -3137 589
rect -3103 555 -3087 589
rect -2961 555 -2945 589
rect -2911 555 -2895 589
rect -2769 555 -2753 589
rect -2719 555 -2703 589
rect -2577 555 -2561 589
rect -2527 555 -2511 589
rect -2385 555 -2369 589
rect -2335 555 -2319 589
rect -2193 555 -2177 589
rect -2143 555 -2127 589
rect -2001 555 -1985 589
rect -1951 555 -1935 589
rect -1809 555 -1793 589
rect -1759 555 -1743 589
rect -1617 555 -1601 589
rect -1567 555 -1551 589
rect -1425 555 -1409 589
rect -1375 555 -1359 589
rect -1233 555 -1217 589
rect -1183 555 -1167 589
rect -1041 555 -1025 589
rect -991 555 -975 589
rect -849 555 -833 589
rect -799 555 -783 589
rect -657 555 -641 589
rect -607 555 -591 589
rect -465 555 -449 589
rect -415 555 -399 589
rect -273 555 -257 589
rect -223 555 -207 589
rect -81 555 -65 589
rect -31 555 -15 589
rect 111 555 127 589
rect 161 555 177 589
rect 303 555 319 589
rect 353 555 369 589
rect 495 555 511 589
rect 545 555 561 589
rect 687 555 703 589
rect 737 555 753 589
rect 879 555 895 589
rect 929 555 945 589
rect 1071 555 1087 589
rect 1121 555 1137 589
rect 1263 555 1279 589
rect 1313 555 1329 589
rect 1455 555 1471 589
rect 1505 555 1521 589
rect 1647 555 1663 589
rect 1697 555 1713 589
rect 1839 555 1855 589
rect 1889 555 1905 589
rect 2031 555 2047 589
rect 2081 555 2097 589
rect 2223 555 2239 589
rect 2273 555 2289 589
rect 2415 555 2431 589
rect 2465 555 2481 589
rect 2607 555 2623 589
rect 2657 555 2673 589
rect 2799 555 2815 589
rect 2849 555 2865 589
rect 2991 555 3007 589
rect 3041 555 3057 589
rect 3183 555 3199 589
rect 3233 555 3249 589
rect 3375 555 3391 589
rect 3425 555 3441 589
rect 3567 555 3583 589
rect 3617 555 3633 589
rect 3759 555 3775 589
rect 3809 555 3825 589
rect 3951 555 3967 589
rect 4001 555 4017 589
rect 4143 555 4159 589
rect 4193 555 4209 589
rect 4335 555 4351 589
rect 4385 555 4401 589
rect 4527 555 4543 589
rect 4577 555 4593 589
rect 4719 555 4735 589
rect 4769 555 4785 589
rect -4689 447 -4673 481
rect -4639 447 -4623 481
rect -4497 447 -4481 481
rect -4447 447 -4431 481
rect -4305 447 -4289 481
rect -4255 447 -4239 481
rect -4113 447 -4097 481
rect -4063 447 -4047 481
rect -3921 447 -3905 481
rect -3871 447 -3855 481
rect -3729 447 -3713 481
rect -3679 447 -3663 481
rect -3537 447 -3521 481
rect -3487 447 -3471 481
rect -3345 447 -3329 481
rect -3295 447 -3279 481
rect -3153 447 -3137 481
rect -3103 447 -3087 481
rect -2961 447 -2945 481
rect -2911 447 -2895 481
rect -2769 447 -2753 481
rect -2719 447 -2703 481
rect -2577 447 -2561 481
rect -2527 447 -2511 481
rect -2385 447 -2369 481
rect -2335 447 -2319 481
rect -2193 447 -2177 481
rect -2143 447 -2127 481
rect -2001 447 -1985 481
rect -1951 447 -1935 481
rect -1809 447 -1793 481
rect -1759 447 -1743 481
rect -1617 447 -1601 481
rect -1567 447 -1551 481
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -849 447 -833 481
rect -799 447 -783 481
rect -657 447 -641 481
rect -607 447 -591 481
rect -465 447 -449 481
rect -415 447 -399 481
rect -273 447 -257 481
rect -223 447 -207 481
rect -81 447 -65 481
rect -31 447 -15 481
rect 111 447 127 481
rect 161 447 177 481
rect 303 447 319 481
rect 353 447 369 481
rect 495 447 511 481
rect 545 447 561 481
rect 687 447 703 481
rect 737 447 753 481
rect 879 447 895 481
rect 929 447 945 481
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1455 447 1471 481
rect 1505 447 1521 481
rect 1647 447 1663 481
rect 1697 447 1713 481
rect 1839 447 1855 481
rect 1889 447 1905 481
rect 2031 447 2047 481
rect 2081 447 2097 481
rect 2223 447 2239 481
rect 2273 447 2289 481
rect 2415 447 2431 481
rect 2465 447 2481 481
rect 2607 447 2623 481
rect 2657 447 2673 481
rect 2799 447 2815 481
rect 2849 447 2865 481
rect 2991 447 3007 481
rect 3041 447 3057 481
rect 3183 447 3199 481
rect 3233 447 3249 481
rect 3375 447 3391 481
rect 3425 447 3441 481
rect 3567 447 3583 481
rect 3617 447 3633 481
rect 3759 447 3775 481
rect 3809 447 3825 481
rect 3951 447 3967 481
rect 4001 447 4017 481
rect 4143 447 4159 481
rect 4193 447 4209 481
rect 4335 447 4351 481
rect 4385 447 4401 481
rect 4527 447 4543 481
rect 4577 447 4593 481
rect 4719 447 4735 481
rect 4769 447 4785 481
rect -4817 397 -4783 413
rect -4817 105 -4783 121
rect -4721 397 -4687 413
rect -4721 105 -4687 121
rect -4625 397 -4591 413
rect -4625 105 -4591 121
rect -4529 397 -4495 413
rect -4529 105 -4495 121
rect -4433 397 -4399 413
rect -4433 105 -4399 121
rect -4337 397 -4303 413
rect -4337 105 -4303 121
rect -4241 397 -4207 413
rect -4241 105 -4207 121
rect -4145 397 -4111 413
rect -4145 105 -4111 121
rect -4049 397 -4015 413
rect -4049 105 -4015 121
rect -3953 397 -3919 413
rect -3953 105 -3919 121
rect -3857 397 -3823 413
rect -3857 105 -3823 121
rect -3761 397 -3727 413
rect -3761 105 -3727 121
rect -3665 397 -3631 413
rect -3665 105 -3631 121
rect -3569 397 -3535 413
rect -3569 105 -3535 121
rect -3473 397 -3439 413
rect -3473 105 -3439 121
rect -3377 397 -3343 413
rect -3377 105 -3343 121
rect -3281 397 -3247 413
rect -3281 105 -3247 121
rect -3185 397 -3151 413
rect -3185 105 -3151 121
rect -3089 397 -3055 413
rect -3089 105 -3055 121
rect -2993 397 -2959 413
rect -2993 105 -2959 121
rect -2897 397 -2863 413
rect -2897 105 -2863 121
rect -2801 397 -2767 413
rect -2801 105 -2767 121
rect -2705 397 -2671 413
rect -2705 105 -2671 121
rect -2609 397 -2575 413
rect -2609 105 -2575 121
rect -2513 397 -2479 413
rect -2513 105 -2479 121
rect -2417 397 -2383 413
rect -2417 105 -2383 121
rect -2321 397 -2287 413
rect -2321 105 -2287 121
rect -2225 397 -2191 413
rect -2225 105 -2191 121
rect -2129 397 -2095 413
rect -2129 105 -2095 121
rect -2033 397 -1999 413
rect -2033 105 -1999 121
rect -1937 397 -1903 413
rect -1937 105 -1903 121
rect -1841 397 -1807 413
rect -1841 105 -1807 121
rect -1745 397 -1711 413
rect -1745 105 -1711 121
rect -1649 397 -1615 413
rect -1649 105 -1615 121
rect -1553 397 -1519 413
rect -1553 105 -1519 121
rect -1457 397 -1423 413
rect -1457 105 -1423 121
rect -1361 397 -1327 413
rect -1361 105 -1327 121
rect -1265 397 -1231 413
rect -1265 105 -1231 121
rect -1169 397 -1135 413
rect -1169 105 -1135 121
rect -1073 397 -1039 413
rect -1073 105 -1039 121
rect -977 397 -943 413
rect -977 105 -943 121
rect -881 397 -847 413
rect -881 105 -847 121
rect -785 397 -751 413
rect -785 105 -751 121
rect -689 397 -655 413
rect -689 105 -655 121
rect -593 397 -559 413
rect -593 105 -559 121
rect -497 397 -463 413
rect -497 105 -463 121
rect -401 397 -367 413
rect -401 105 -367 121
rect -305 397 -271 413
rect -305 105 -271 121
rect -209 397 -175 413
rect -209 105 -175 121
rect -113 397 -79 413
rect -113 105 -79 121
rect -17 397 17 413
rect -17 105 17 121
rect 79 397 113 413
rect 79 105 113 121
rect 175 397 209 413
rect 175 105 209 121
rect 271 397 305 413
rect 271 105 305 121
rect 367 397 401 413
rect 367 105 401 121
rect 463 397 497 413
rect 463 105 497 121
rect 559 397 593 413
rect 559 105 593 121
rect 655 397 689 413
rect 655 105 689 121
rect 751 397 785 413
rect 751 105 785 121
rect 847 397 881 413
rect 847 105 881 121
rect 943 397 977 413
rect 943 105 977 121
rect 1039 397 1073 413
rect 1039 105 1073 121
rect 1135 397 1169 413
rect 1135 105 1169 121
rect 1231 397 1265 413
rect 1231 105 1265 121
rect 1327 397 1361 413
rect 1327 105 1361 121
rect 1423 397 1457 413
rect 1423 105 1457 121
rect 1519 397 1553 413
rect 1519 105 1553 121
rect 1615 397 1649 413
rect 1615 105 1649 121
rect 1711 397 1745 413
rect 1711 105 1745 121
rect 1807 397 1841 413
rect 1807 105 1841 121
rect 1903 397 1937 413
rect 1903 105 1937 121
rect 1999 397 2033 413
rect 1999 105 2033 121
rect 2095 397 2129 413
rect 2095 105 2129 121
rect 2191 397 2225 413
rect 2191 105 2225 121
rect 2287 397 2321 413
rect 2287 105 2321 121
rect 2383 397 2417 413
rect 2383 105 2417 121
rect 2479 397 2513 413
rect 2479 105 2513 121
rect 2575 397 2609 413
rect 2575 105 2609 121
rect 2671 397 2705 413
rect 2671 105 2705 121
rect 2767 397 2801 413
rect 2767 105 2801 121
rect 2863 397 2897 413
rect 2863 105 2897 121
rect 2959 397 2993 413
rect 2959 105 2993 121
rect 3055 397 3089 413
rect 3055 105 3089 121
rect 3151 397 3185 413
rect 3151 105 3185 121
rect 3247 397 3281 413
rect 3247 105 3281 121
rect 3343 397 3377 413
rect 3343 105 3377 121
rect 3439 397 3473 413
rect 3439 105 3473 121
rect 3535 397 3569 413
rect 3535 105 3569 121
rect 3631 397 3665 413
rect 3631 105 3665 121
rect 3727 397 3761 413
rect 3727 105 3761 121
rect 3823 397 3857 413
rect 3823 105 3857 121
rect 3919 397 3953 413
rect 3919 105 3953 121
rect 4015 397 4049 413
rect 4015 105 4049 121
rect 4111 397 4145 413
rect 4111 105 4145 121
rect 4207 397 4241 413
rect 4207 105 4241 121
rect 4303 397 4337 413
rect 4303 105 4337 121
rect 4399 397 4433 413
rect 4399 105 4433 121
rect 4495 397 4529 413
rect 4495 105 4529 121
rect 4591 397 4625 413
rect 4591 105 4625 121
rect 4687 397 4721 413
rect 4687 105 4721 121
rect 4783 397 4817 413
rect 4783 105 4817 121
rect -4785 37 -4769 71
rect -4735 37 -4719 71
rect -4593 37 -4577 71
rect -4543 37 -4527 71
rect -4401 37 -4385 71
rect -4351 37 -4335 71
rect -4209 37 -4193 71
rect -4159 37 -4143 71
rect -4017 37 -4001 71
rect -3967 37 -3951 71
rect -3825 37 -3809 71
rect -3775 37 -3759 71
rect -3633 37 -3617 71
rect -3583 37 -3567 71
rect -3441 37 -3425 71
rect -3391 37 -3375 71
rect -3249 37 -3233 71
rect -3199 37 -3183 71
rect -3057 37 -3041 71
rect -3007 37 -2991 71
rect -2865 37 -2849 71
rect -2815 37 -2799 71
rect -2673 37 -2657 71
rect -2623 37 -2607 71
rect -2481 37 -2465 71
rect -2431 37 -2415 71
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -945 37 -929 71
rect -895 37 -879 71
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect 975 37 991 71
rect 1025 37 1041 71
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2319 37 2335 71
rect 2369 37 2385 71
rect 2511 37 2527 71
rect 2561 37 2577 71
rect 2703 37 2719 71
rect 2753 37 2769 71
rect 2895 37 2911 71
rect 2945 37 2961 71
rect 3087 37 3103 71
rect 3137 37 3153 71
rect 3279 37 3295 71
rect 3329 37 3345 71
rect 3471 37 3487 71
rect 3521 37 3537 71
rect 3663 37 3679 71
rect 3713 37 3729 71
rect 3855 37 3871 71
rect 3905 37 3921 71
rect 4047 37 4063 71
rect 4097 37 4113 71
rect 4239 37 4255 71
rect 4289 37 4305 71
rect 4431 37 4447 71
rect 4481 37 4497 71
rect 4623 37 4639 71
rect 4673 37 4689 71
rect -4785 -71 -4769 -37
rect -4735 -71 -4719 -37
rect -4593 -71 -4577 -37
rect -4543 -71 -4527 -37
rect -4401 -71 -4385 -37
rect -4351 -71 -4335 -37
rect -4209 -71 -4193 -37
rect -4159 -71 -4143 -37
rect -4017 -71 -4001 -37
rect -3967 -71 -3951 -37
rect -3825 -71 -3809 -37
rect -3775 -71 -3759 -37
rect -3633 -71 -3617 -37
rect -3583 -71 -3567 -37
rect -3441 -71 -3425 -37
rect -3391 -71 -3375 -37
rect -3249 -71 -3233 -37
rect -3199 -71 -3183 -37
rect -3057 -71 -3041 -37
rect -3007 -71 -2991 -37
rect -2865 -71 -2849 -37
rect -2815 -71 -2799 -37
rect -2673 -71 -2657 -37
rect -2623 -71 -2607 -37
rect -2481 -71 -2465 -37
rect -2431 -71 -2415 -37
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect 2511 -71 2527 -37
rect 2561 -71 2577 -37
rect 2703 -71 2719 -37
rect 2753 -71 2769 -37
rect 2895 -71 2911 -37
rect 2945 -71 2961 -37
rect 3087 -71 3103 -37
rect 3137 -71 3153 -37
rect 3279 -71 3295 -37
rect 3329 -71 3345 -37
rect 3471 -71 3487 -37
rect 3521 -71 3537 -37
rect 3663 -71 3679 -37
rect 3713 -71 3729 -37
rect 3855 -71 3871 -37
rect 3905 -71 3921 -37
rect 4047 -71 4063 -37
rect 4097 -71 4113 -37
rect 4239 -71 4255 -37
rect 4289 -71 4305 -37
rect 4431 -71 4447 -37
rect 4481 -71 4497 -37
rect 4623 -71 4639 -37
rect 4673 -71 4689 -37
rect -4817 -121 -4783 -105
rect -4817 -413 -4783 -397
rect -4721 -121 -4687 -105
rect -4721 -413 -4687 -397
rect -4625 -121 -4591 -105
rect -4625 -413 -4591 -397
rect -4529 -121 -4495 -105
rect -4529 -413 -4495 -397
rect -4433 -121 -4399 -105
rect -4433 -413 -4399 -397
rect -4337 -121 -4303 -105
rect -4337 -413 -4303 -397
rect -4241 -121 -4207 -105
rect -4241 -413 -4207 -397
rect -4145 -121 -4111 -105
rect -4145 -413 -4111 -397
rect -4049 -121 -4015 -105
rect -4049 -413 -4015 -397
rect -3953 -121 -3919 -105
rect -3953 -413 -3919 -397
rect -3857 -121 -3823 -105
rect -3857 -413 -3823 -397
rect -3761 -121 -3727 -105
rect -3761 -413 -3727 -397
rect -3665 -121 -3631 -105
rect -3665 -413 -3631 -397
rect -3569 -121 -3535 -105
rect -3569 -413 -3535 -397
rect -3473 -121 -3439 -105
rect -3473 -413 -3439 -397
rect -3377 -121 -3343 -105
rect -3377 -413 -3343 -397
rect -3281 -121 -3247 -105
rect -3281 -413 -3247 -397
rect -3185 -121 -3151 -105
rect -3185 -413 -3151 -397
rect -3089 -121 -3055 -105
rect -3089 -413 -3055 -397
rect -2993 -121 -2959 -105
rect -2993 -413 -2959 -397
rect -2897 -121 -2863 -105
rect -2897 -413 -2863 -397
rect -2801 -121 -2767 -105
rect -2801 -413 -2767 -397
rect -2705 -121 -2671 -105
rect -2705 -413 -2671 -397
rect -2609 -121 -2575 -105
rect -2609 -413 -2575 -397
rect -2513 -121 -2479 -105
rect -2513 -413 -2479 -397
rect -2417 -121 -2383 -105
rect -2417 -413 -2383 -397
rect -2321 -121 -2287 -105
rect -2321 -413 -2287 -397
rect -2225 -121 -2191 -105
rect -2225 -413 -2191 -397
rect -2129 -121 -2095 -105
rect -2129 -413 -2095 -397
rect -2033 -121 -1999 -105
rect -2033 -413 -1999 -397
rect -1937 -121 -1903 -105
rect -1937 -413 -1903 -397
rect -1841 -121 -1807 -105
rect -1841 -413 -1807 -397
rect -1745 -121 -1711 -105
rect -1745 -413 -1711 -397
rect -1649 -121 -1615 -105
rect -1649 -413 -1615 -397
rect -1553 -121 -1519 -105
rect -1553 -413 -1519 -397
rect -1457 -121 -1423 -105
rect -1457 -413 -1423 -397
rect -1361 -121 -1327 -105
rect -1361 -413 -1327 -397
rect -1265 -121 -1231 -105
rect -1265 -413 -1231 -397
rect -1169 -121 -1135 -105
rect -1169 -413 -1135 -397
rect -1073 -121 -1039 -105
rect -1073 -413 -1039 -397
rect -977 -121 -943 -105
rect -977 -413 -943 -397
rect -881 -121 -847 -105
rect -881 -413 -847 -397
rect -785 -121 -751 -105
rect -785 -413 -751 -397
rect -689 -121 -655 -105
rect -689 -413 -655 -397
rect -593 -121 -559 -105
rect -593 -413 -559 -397
rect -497 -121 -463 -105
rect -497 -413 -463 -397
rect -401 -121 -367 -105
rect -401 -413 -367 -397
rect -305 -121 -271 -105
rect -305 -413 -271 -397
rect -209 -121 -175 -105
rect -209 -413 -175 -397
rect -113 -121 -79 -105
rect -113 -413 -79 -397
rect -17 -121 17 -105
rect -17 -413 17 -397
rect 79 -121 113 -105
rect 79 -413 113 -397
rect 175 -121 209 -105
rect 175 -413 209 -397
rect 271 -121 305 -105
rect 271 -413 305 -397
rect 367 -121 401 -105
rect 367 -413 401 -397
rect 463 -121 497 -105
rect 463 -413 497 -397
rect 559 -121 593 -105
rect 559 -413 593 -397
rect 655 -121 689 -105
rect 655 -413 689 -397
rect 751 -121 785 -105
rect 751 -413 785 -397
rect 847 -121 881 -105
rect 847 -413 881 -397
rect 943 -121 977 -105
rect 943 -413 977 -397
rect 1039 -121 1073 -105
rect 1039 -413 1073 -397
rect 1135 -121 1169 -105
rect 1135 -413 1169 -397
rect 1231 -121 1265 -105
rect 1231 -413 1265 -397
rect 1327 -121 1361 -105
rect 1327 -413 1361 -397
rect 1423 -121 1457 -105
rect 1423 -413 1457 -397
rect 1519 -121 1553 -105
rect 1519 -413 1553 -397
rect 1615 -121 1649 -105
rect 1615 -413 1649 -397
rect 1711 -121 1745 -105
rect 1711 -413 1745 -397
rect 1807 -121 1841 -105
rect 1807 -413 1841 -397
rect 1903 -121 1937 -105
rect 1903 -413 1937 -397
rect 1999 -121 2033 -105
rect 1999 -413 2033 -397
rect 2095 -121 2129 -105
rect 2095 -413 2129 -397
rect 2191 -121 2225 -105
rect 2191 -413 2225 -397
rect 2287 -121 2321 -105
rect 2287 -413 2321 -397
rect 2383 -121 2417 -105
rect 2383 -413 2417 -397
rect 2479 -121 2513 -105
rect 2479 -413 2513 -397
rect 2575 -121 2609 -105
rect 2575 -413 2609 -397
rect 2671 -121 2705 -105
rect 2671 -413 2705 -397
rect 2767 -121 2801 -105
rect 2767 -413 2801 -397
rect 2863 -121 2897 -105
rect 2863 -413 2897 -397
rect 2959 -121 2993 -105
rect 2959 -413 2993 -397
rect 3055 -121 3089 -105
rect 3055 -413 3089 -397
rect 3151 -121 3185 -105
rect 3151 -413 3185 -397
rect 3247 -121 3281 -105
rect 3247 -413 3281 -397
rect 3343 -121 3377 -105
rect 3343 -413 3377 -397
rect 3439 -121 3473 -105
rect 3439 -413 3473 -397
rect 3535 -121 3569 -105
rect 3535 -413 3569 -397
rect 3631 -121 3665 -105
rect 3631 -413 3665 -397
rect 3727 -121 3761 -105
rect 3727 -413 3761 -397
rect 3823 -121 3857 -105
rect 3823 -413 3857 -397
rect 3919 -121 3953 -105
rect 3919 -413 3953 -397
rect 4015 -121 4049 -105
rect 4015 -413 4049 -397
rect 4111 -121 4145 -105
rect 4111 -413 4145 -397
rect 4207 -121 4241 -105
rect 4207 -413 4241 -397
rect 4303 -121 4337 -105
rect 4303 -413 4337 -397
rect 4399 -121 4433 -105
rect 4399 -413 4433 -397
rect 4495 -121 4529 -105
rect 4495 -413 4529 -397
rect 4591 -121 4625 -105
rect 4591 -413 4625 -397
rect 4687 -121 4721 -105
rect 4687 -413 4721 -397
rect 4783 -121 4817 -105
rect 4783 -413 4817 -397
rect -4689 -481 -4673 -447
rect -4639 -481 -4623 -447
rect -4497 -481 -4481 -447
rect -4447 -481 -4431 -447
rect -4305 -481 -4289 -447
rect -4255 -481 -4239 -447
rect -4113 -481 -4097 -447
rect -4063 -481 -4047 -447
rect -3921 -481 -3905 -447
rect -3871 -481 -3855 -447
rect -3729 -481 -3713 -447
rect -3679 -481 -3663 -447
rect -3537 -481 -3521 -447
rect -3487 -481 -3471 -447
rect -3345 -481 -3329 -447
rect -3295 -481 -3279 -447
rect -3153 -481 -3137 -447
rect -3103 -481 -3087 -447
rect -2961 -481 -2945 -447
rect -2911 -481 -2895 -447
rect -2769 -481 -2753 -447
rect -2719 -481 -2703 -447
rect -2577 -481 -2561 -447
rect -2527 -481 -2511 -447
rect -2385 -481 -2369 -447
rect -2335 -481 -2319 -447
rect -2193 -481 -2177 -447
rect -2143 -481 -2127 -447
rect -2001 -481 -1985 -447
rect -1951 -481 -1935 -447
rect -1809 -481 -1793 -447
rect -1759 -481 -1743 -447
rect -1617 -481 -1601 -447
rect -1567 -481 -1551 -447
rect -1425 -481 -1409 -447
rect -1375 -481 -1359 -447
rect -1233 -481 -1217 -447
rect -1183 -481 -1167 -447
rect -1041 -481 -1025 -447
rect -991 -481 -975 -447
rect -849 -481 -833 -447
rect -799 -481 -783 -447
rect -657 -481 -641 -447
rect -607 -481 -591 -447
rect -465 -481 -449 -447
rect -415 -481 -399 -447
rect -273 -481 -257 -447
rect -223 -481 -207 -447
rect -81 -481 -65 -447
rect -31 -481 -15 -447
rect 111 -481 127 -447
rect 161 -481 177 -447
rect 303 -481 319 -447
rect 353 -481 369 -447
rect 495 -481 511 -447
rect 545 -481 561 -447
rect 687 -481 703 -447
rect 737 -481 753 -447
rect 879 -481 895 -447
rect 929 -481 945 -447
rect 1071 -481 1087 -447
rect 1121 -481 1137 -447
rect 1263 -481 1279 -447
rect 1313 -481 1329 -447
rect 1455 -481 1471 -447
rect 1505 -481 1521 -447
rect 1647 -481 1663 -447
rect 1697 -481 1713 -447
rect 1839 -481 1855 -447
rect 1889 -481 1905 -447
rect 2031 -481 2047 -447
rect 2081 -481 2097 -447
rect 2223 -481 2239 -447
rect 2273 -481 2289 -447
rect 2415 -481 2431 -447
rect 2465 -481 2481 -447
rect 2607 -481 2623 -447
rect 2657 -481 2673 -447
rect 2799 -481 2815 -447
rect 2849 -481 2865 -447
rect 2991 -481 3007 -447
rect 3041 -481 3057 -447
rect 3183 -481 3199 -447
rect 3233 -481 3249 -447
rect 3375 -481 3391 -447
rect 3425 -481 3441 -447
rect 3567 -481 3583 -447
rect 3617 -481 3633 -447
rect 3759 -481 3775 -447
rect 3809 -481 3825 -447
rect 3951 -481 3967 -447
rect 4001 -481 4017 -447
rect 4143 -481 4159 -447
rect 4193 -481 4209 -447
rect 4335 -481 4351 -447
rect 4385 -481 4401 -447
rect 4527 -481 4543 -447
rect 4577 -481 4593 -447
rect 4719 -481 4735 -447
rect 4769 -481 4785 -447
rect -4689 -589 -4673 -555
rect -4639 -589 -4623 -555
rect -4497 -589 -4481 -555
rect -4447 -589 -4431 -555
rect -4305 -589 -4289 -555
rect -4255 -589 -4239 -555
rect -4113 -589 -4097 -555
rect -4063 -589 -4047 -555
rect -3921 -589 -3905 -555
rect -3871 -589 -3855 -555
rect -3729 -589 -3713 -555
rect -3679 -589 -3663 -555
rect -3537 -589 -3521 -555
rect -3487 -589 -3471 -555
rect -3345 -589 -3329 -555
rect -3295 -589 -3279 -555
rect -3153 -589 -3137 -555
rect -3103 -589 -3087 -555
rect -2961 -589 -2945 -555
rect -2911 -589 -2895 -555
rect -2769 -589 -2753 -555
rect -2719 -589 -2703 -555
rect -2577 -589 -2561 -555
rect -2527 -589 -2511 -555
rect -2385 -589 -2369 -555
rect -2335 -589 -2319 -555
rect -2193 -589 -2177 -555
rect -2143 -589 -2127 -555
rect -2001 -589 -1985 -555
rect -1951 -589 -1935 -555
rect -1809 -589 -1793 -555
rect -1759 -589 -1743 -555
rect -1617 -589 -1601 -555
rect -1567 -589 -1551 -555
rect -1425 -589 -1409 -555
rect -1375 -589 -1359 -555
rect -1233 -589 -1217 -555
rect -1183 -589 -1167 -555
rect -1041 -589 -1025 -555
rect -991 -589 -975 -555
rect -849 -589 -833 -555
rect -799 -589 -783 -555
rect -657 -589 -641 -555
rect -607 -589 -591 -555
rect -465 -589 -449 -555
rect -415 -589 -399 -555
rect -273 -589 -257 -555
rect -223 -589 -207 -555
rect -81 -589 -65 -555
rect -31 -589 -15 -555
rect 111 -589 127 -555
rect 161 -589 177 -555
rect 303 -589 319 -555
rect 353 -589 369 -555
rect 495 -589 511 -555
rect 545 -589 561 -555
rect 687 -589 703 -555
rect 737 -589 753 -555
rect 879 -589 895 -555
rect 929 -589 945 -555
rect 1071 -589 1087 -555
rect 1121 -589 1137 -555
rect 1263 -589 1279 -555
rect 1313 -589 1329 -555
rect 1455 -589 1471 -555
rect 1505 -589 1521 -555
rect 1647 -589 1663 -555
rect 1697 -589 1713 -555
rect 1839 -589 1855 -555
rect 1889 -589 1905 -555
rect 2031 -589 2047 -555
rect 2081 -589 2097 -555
rect 2223 -589 2239 -555
rect 2273 -589 2289 -555
rect 2415 -589 2431 -555
rect 2465 -589 2481 -555
rect 2607 -589 2623 -555
rect 2657 -589 2673 -555
rect 2799 -589 2815 -555
rect 2849 -589 2865 -555
rect 2991 -589 3007 -555
rect 3041 -589 3057 -555
rect 3183 -589 3199 -555
rect 3233 -589 3249 -555
rect 3375 -589 3391 -555
rect 3425 -589 3441 -555
rect 3567 -589 3583 -555
rect 3617 -589 3633 -555
rect 3759 -589 3775 -555
rect 3809 -589 3825 -555
rect 3951 -589 3967 -555
rect 4001 -589 4017 -555
rect 4143 -589 4159 -555
rect 4193 -589 4209 -555
rect 4335 -589 4351 -555
rect 4385 -589 4401 -555
rect 4527 -589 4543 -555
rect 4577 -589 4593 -555
rect 4719 -589 4735 -555
rect 4769 -589 4785 -555
rect -4817 -639 -4783 -623
rect -4817 -931 -4783 -915
rect -4721 -639 -4687 -623
rect -4721 -931 -4687 -915
rect -4625 -639 -4591 -623
rect -4625 -931 -4591 -915
rect -4529 -639 -4495 -623
rect -4529 -931 -4495 -915
rect -4433 -639 -4399 -623
rect -4433 -931 -4399 -915
rect -4337 -639 -4303 -623
rect -4337 -931 -4303 -915
rect -4241 -639 -4207 -623
rect -4241 -931 -4207 -915
rect -4145 -639 -4111 -623
rect -4145 -931 -4111 -915
rect -4049 -639 -4015 -623
rect -4049 -931 -4015 -915
rect -3953 -639 -3919 -623
rect -3953 -931 -3919 -915
rect -3857 -639 -3823 -623
rect -3857 -931 -3823 -915
rect -3761 -639 -3727 -623
rect -3761 -931 -3727 -915
rect -3665 -639 -3631 -623
rect -3665 -931 -3631 -915
rect -3569 -639 -3535 -623
rect -3569 -931 -3535 -915
rect -3473 -639 -3439 -623
rect -3473 -931 -3439 -915
rect -3377 -639 -3343 -623
rect -3377 -931 -3343 -915
rect -3281 -639 -3247 -623
rect -3281 -931 -3247 -915
rect -3185 -639 -3151 -623
rect -3185 -931 -3151 -915
rect -3089 -639 -3055 -623
rect -3089 -931 -3055 -915
rect -2993 -639 -2959 -623
rect -2993 -931 -2959 -915
rect -2897 -639 -2863 -623
rect -2897 -931 -2863 -915
rect -2801 -639 -2767 -623
rect -2801 -931 -2767 -915
rect -2705 -639 -2671 -623
rect -2705 -931 -2671 -915
rect -2609 -639 -2575 -623
rect -2609 -931 -2575 -915
rect -2513 -639 -2479 -623
rect -2513 -931 -2479 -915
rect -2417 -639 -2383 -623
rect -2417 -931 -2383 -915
rect -2321 -639 -2287 -623
rect -2321 -931 -2287 -915
rect -2225 -639 -2191 -623
rect -2225 -931 -2191 -915
rect -2129 -639 -2095 -623
rect -2129 -931 -2095 -915
rect -2033 -639 -1999 -623
rect -2033 -931 -1999 -915
rect -1937 -639 -1903 -623
rect -1937 -931 -1903 -915
rect -1841 -639 -1807 -623
rect -1841 -931 -1807 -915
rect -1745 -639 -1711 -623
rect -1745 -931 -1711 -915
rect -1649 -639 -1615 -623
rect -1649 -931 -1615 -915
rect -1553 -639 -1519 -623
rect -1553 -931 -1519 -915
rect -1457 -639 -1423 -623
rect -1457 -931 -1423 -915
rect -1361 -639 -1327 -623
rect -1361 -931 -1327 -915
rect -1265 -639 -1231 -623
rect -1265 -931 -1231 -915
rect -1169 -639 -1135 -623
rect -1169 -931 -1135 -915
rect -1073 -639 -1039 -623
rect -1073 -931 -1039 -915
rect -977 -639 -943 -623
rect -977 -931 -943 -915
rect -881 -639 -847 -623
rect -881 -931 -847 -915
rect -785 -639 -751 -623
rect -785 -931 -751 -915
rect -689 -639 -655 -623
rect -689 -931 -655 -915
rect -593 -639 -559 -623
rect -593 -931 -559 -915
rect -497 -639 -463 -623
rect -497 -931 -463 -915
rect -401 -639 -367 -623
rect -401 -931 -367 -915
rect -305 -639 -271 -623
rect -305 -931 -271 -915
rect -209 -639 -175 -623
rect -209 -931 -175 -915
rect -113 -639 -79 -623
rect -113 -931 -79 -915
rect -17 -639 17 -623
rect -17 -931 17 -915
rect 79 -639 113 -623
rect 79 -931 113 -915
rect 175 -639 209 -623
rect 175 -931 209 -915
rect 271 -639 305 -623
rect 271 -931 305 -915
rect 367 -639 401 -623
rect 367 -931 401 -915
rect 463 -639 497 -623
rect 463 -931 497 -915
rect 559 -639 593 -623
rect 559 -931 593 -915
rect 655 -639 689 -623
rect 655 -931 689 -915
rect 751 -639 785 -623
rect 751 -931 785 -915
rect 847 -639 881 -623
rect 847 -931 881 -915
rect 943 -639 977 -623
rect 943 -931 977 -915
rect 1039 -639 1073 -623
rect 1039 -931 1073 -915
rect 1135 -639 1169 -623
rect 1135 -931 1169 -915
rect 1231 -639 1265 -623
rect 1231 -931 1265 -915
rect 1327 -639 1361 -623
rect 1327 -931 1361 -915
rect 1423 -639 1457 -623
rect 1423 -931 1457 -915
rect 1519 -639 1553 -623
rect 1519 -931 1553 -915
rect 1615 -639 1649 -623
rect 1615 -931 1649 -915
rect 1711 -639 1745 -623
rect 1711 -931 1745 -915
rect 1807 -639 1841 -623
rect 1807 -931 1841 -915
rect 1903 -639 1937 -623
rect 1903 -931 1937 -915
rect 1999 -639 2033 -623
rect 1999 -931 2033 -915
rect 2095 -639 2129 -623
rect 2095 -931 2129 -915
rect 2191 -639 2225 -623
rect 2191 -931 2225 -915
rect 2287 -639 2321 -623
rect 2287 -931 2321 -915
rect 2383 -639 2417 -623
rect 2383 -931 2417 -915
rect 2479 -639 2513 -623
rect 2479 -931 2513 -915
rect 2575 -639 2609 -623
rect 2575 -931 2609 -915
rect 2671 -639 2705 -623
rect 2671 -931 2705 -915
rect 2767 -639 2801 -623
rect 2767 -931 2801 -915
rect 2863 -639 2897 -623
rect 2863 -931 2897 -915
rect 2959 -639 2993 -623
rect 2959 -931 2993 -915
rect 3055 -639 3089 -623
rect 3055 -931 3089 -915
rect 3151 -639 3185 -623
rect 3151 -931 3185 -915
rect 3247 -639 3281 -623
rect 3247 -931 3281 -915
rect 3343 -639 3377 -623
rect 3343 -931 3377 -915
rect 3439 -639 3473 -623
rect 3439 -931 3473 -915
rect 3535 -639 3569 -623
rect 3535 -931 3569 -915
rect 3631 -639 3665 -623
rect 3631 -931 3665 -915
rect 3727 -639 3761 -623
rect 3727 -931 3761 -915
rect 3823 -639 3857 -623
rect 3823 -931 3857 -915
rect 3919 -639 3953 -623
rect 3919 -931 3953 -915
rect 4015 -639 4049 -623
rect 4015 -931 4049 -915
rect 4111 -639 4145 -623
rect 4111 -931 4145 -915
rect 4207 -639 4241 -623
rect 4207 -931 4241 -915
rect 4303 -639 4337 -623
rect 4303 -931 4337 -915
rect 4399 -639 4433 -623
rect 4399 -931 4433 -915
rect 4495 -639 4529 -623
rect 4495 -931 4529 -915
rect 4591 -639 4625 -623
rect 4591 -931 4625 -915
rect 4687 -639 4721 -623
rect 4687 -931 4721 -915
rect 4783 -639 4817 -623
rect 4783 -931 4817 -915
rect -4785 -999 -4769 -965
rect -4735 -999 -4719 -965
rect -4593 -999 -4577 -965
rect -4543 -999 -4527 -965
rect -4401 -999 -4385 -965
rect -4351 -999 -4335 -965
rect -4209 -999 -4193 -965
rect -4159 -999 -4143 -965
rect -4017 -999 -4001 -965
rect -3967 -999 -3951 -965
rect -3825 -999 -3809 -965
rect -3775 -999 -3759 -965
rect -3633 -999 -3617 -965
rect -3583 -999 -3567 -965
rect -3441 -999 -3425 -965
rect -3391 -999 -3375 -965
rect -3249 -999 -3233 -965
rect -3199 -999 -3183 -965
rect -3057 -999 -3041 -965
rect -3007 -999 -2991 -965
rect -2865 -999 -2849 -965
rect -2815 -999 -2799 -965
rect -2673 -999 -2657 -965
rect -2623 -999 -2607 -965
rect -2481 -999 -2465 -965
rect -2431 -999 -2415 -965
rect -2289 -999 -2273 -965
rect -2239 -999 -2223 -965
rect -2097 -999 -2081 -965
rect -2047 -999 -2031 -965
rect -1905 -999 -1889 -965
rect -1855 -999 -1839 -965
rect -1713 -999 -1697 -965
rect -1663 -999 -1647 -965
rect -1521 -999 -1505 -965
rect -1471 -999 -1455 -965
rect -1329 -999 -1313 -965
rect -1279 -999 -1263 -965
rect -1137 -999 -1121 -965
rect -1087 -999 -1071 -965
rect -945 -999 -929 -965
rect -895 -999 -879 -965
rect -753 -999 -737 -965
rect -703 -999 -687 -965
rect -561 -999 -545 -965
rect -511 -999 -495 -965
rect -369 -999 -353 -965
rect -319 -999 -303 -965
rect -177 -999 -161 -965
rect -127 -999 -111 -965
rect 15 -999 31 -965
rect 65 -999 81 -965
rect 207 -999 223 -965
rect 257 -999 273 -965
rect 399 -999 415 -965
rect 449 -999 465 -965
rect 591 -999 607 -965
rect 641 -999 657 -965
rect 783 -999 799 -965
rect 833 -999 849 -965
rect 975 -999 991 -965
rect 1025 -999 1041 -965
rect 1167 -999 1183 -965
rect 1217 -999 1233 -965
rect 1359 -999 1375 -965
rect 1409 -999 1425 -965
rect 1551 -999 1567 -965
rect 1601 -999 1617 -965
rect 1743 -999 1759 -965
rect 1793 -999 1809 -965
rect 1935 -999 1951 -965
rect 1985 -999 2001 -965
rect 2127 -999 2143 -965
rect 2177 -999 2193 -965
rect 2319 -999 2335 -965
rect 2369 -999 2385 -965
rect 2511 -999 2527 -965
rect 2561 -999 2577 -965
rect 2703 -999 2719 -965
rect 2753 -999 2769 -965
rect 2895 -999 2911 -965
rect 2945 -999 2961 -965
rect 3087 -999 3103 -965
rect 3137 -999 3153 -965
rect 3279 -999 3295 -965
rect 3329 -999 3345 -965
rect 3471 -999 3487 -965
rect 3521 -999 3537 -965
rect 3663 -999 3679 -965
rect 3713 -999 3729 -965
rect 3855 -999 3871 -965
rect 3905 -999 3921 -965
rect 4047 -999 4063 -965
rect 4097 -999 4113 -965
rect 4239 -999 4255 -965
rect 4289 -999 4305 -965
rect 4431 -999 4447 -965
rect 4481 -999 4497 -965
rect 4623 -999 4639 -965
rect 4673 -999 4689 -965
rect -4931 -1067 -4897 -1005
rect 4897 -1067 4931 -1005
rect -4931 -1101 -4835 -1067
rect 4835 -1101 4931 -1067
<< viali >>
rect -4769 965 -4735 999
rect -4577 965 -4543 999
rect -4385 965 -4351 999
rect -4193 965 -4159 999
rect -4001 965 -3967 999
rect -3809 965 -3775 999
rect -3617 965 -3583 999
rect -3425 965 -3391 999
rect -3233 965 -3199 999
rect -3041 965 -3007 999
rect -2849 965 -2815 999
rect -2657 965 -2623 999
rect -2465 965 -2431 999
rect -2273 965 -2239 999
rect -2081 965 -2047 999
rect -1889 965 -1855 999
rect -1697 965 -1663 999
rect -1505 965 -1471 999
rect -1313 965 -1279 999
rect -1121 965 -1087 999
rect -929 965 -895 999
rect -737 965 -703 999
rect -545 965 -511 999
rect -353 965 -319 999
rect -161 965 -127 999
rect 31 965 65 999
rect 223 965 257 999
rect 415 965 449 999
rect 607 965 641 999
rect 799 965 833 999
rect 991 965 1025 999
rect 1183 965 1217 999
rect 1375 965 1409 999
rect 1567 965 1601 999
rect 1759 965 1793 999
rect 1951 965 1985 999
rect 2143 965 2177 999
rect 2335 965 2369 999
rect 2527 965 2561 999
rect 2719 965 2753 999
rect 2911 965 2945 999
rect 3103 965 3137 999
rect 3295 965 3329 999
rect 3487 965 3521 999
rect 3679 965 3713 999
rect 3871 965 3905 999
rect 4063 965 4097 999
rect 4255 965 4289 999
rect 4447 965 4481 999
rect 4639 965 4673 999
rect -4817 639 -4783 915
rect -4721 639 -4687 915
rect -4625 639 -4591 915
rect -4529 639 -4495 915
rect -4433 639 -4399 915
rect -4337 639 -4303 915
rect -4241 639 -4207 915
rect -4145 639 -4111 915
rect -4049 639 -4015 915
rect -3953 639 -3919 915
rect -3857 639 -3823 915
rect -3761 639 -3727 915
rect -3665 639 -3631 915
rect -3569 639 -3535 915
rect -3473 639 -3439 915
rect -3377 639 -3343 915
rect -3281 639 -3247 915
rect -3185 639 -3151 915
rect -3089 639 -3055 915
rect -2993 639 -2959 915
rect -2897 639 -2863 915
rect -2801 639 -2767 915
rect -2705 639 -2671 915
rect -2609 639 -2575 915
rect -2513 639 -2479 915
rect -2417 639 -2383 915
rect -2321 639 -2287 915
rect -2225 639 -2191 915
rect -2129 639 -2095 915
rect -2033 639 -1999 915
rect -1937 639 -1903 915
rect -1841 639 -1807 915
rect -1745 639 -1711 915
rect -1649 639 -1615 915
rect -1553 639 -1519 915
rect -1457 639 -1423 915
rect -1361 639 -1327 915
rect -1265 639 -1231 915
rect -1169 639 -1135 915
rect -1073 639 -1039 915
rect -977 639 -943 915
rect -881 639 -847 915
rect -785 639 -751 915
rect -689 639 -655 915
rect -593 639 -559 915
rect -497 639 -463 915
rect -401 639 -367 915
rect -305 639 -271 915
rect -209 639 -175 915
rect -113 639 -79 915
rect -17 639 17 915
rect 79 639 113 915
rect 175 639 209 915
rect 271 639 305 915
rect 367 639 401 915
rect 463 639 497 915
rect 559 639 593 915
rect 655 639 689 915
rect 751 639 785 915
rect 847 639 881 915
rect 943 639 977 915
rect 1039 639 1073 915
rect 1135 639 1169 915
rect 1231 639 1265 915
rect 1327 639 1361 915
rect 1423 639 1457 915
rect 1519 639 1553 915
rect 1615 639 1649 915
rect 1711 639 1745 915
rect 1807 639 1841 915
rect 1903 639 1937 915
rect 1999 639 2033 915
rect 2095 639 2129 915
rect 2191 639 2225 915
rect 2287 639 2321 915
rect 2383 639 2417 915
rect 2479 639 2513 915
rect 2575 639 2609 915
rect 2671 639 2705 915
rect 2767 639 2801 915
rect 2863 639 2897 915
rect 2959 639 2993 915
rect 3055 639 3089 915
rect 3151 639 3185 915
rect 3247 639 3281 915
rect 3343 639 3377 915
rect 3439 639 3473 915
rect 3535 639 3569 915
rect 3631 639 3665 915
rect 3727 639 3761 915
rect 3823 639 3857 915
rect 3919 639 3953 915
rect 4015 639 4049 915
rect 4111 639 4145 915
rect 4207 639 4241 915
rect 4303 639 4337 915
rect 4399 639 4433 915
rect 4495 639 4529 915
rect 4591 639 4625 915
rect 4687 639 4721 915
rect 4783 639 4817 915
rect -4673 555 -4639 589
rect -4481 555 -4447 589
rect -4289 555 -4255 589
rect -4097 555 -4063 589
rect -3905 555 -3871 589
rect -3713 555 -3679 589
rect -3521 555 -3487 589
rect -3329 555 -3295 589
rect -3137 555 -3103 589
rect -2945 555 -2911 589
rect -2753 555 -2719 589
rect -2561 555 -2527 589
rect -2369 555 -2335 589
rect -2177 555 -2143 589
rect -1985 555 -1951 589
rect -1793 555 -1759 589
rect -1601 555 -1567 589
rect -1409 555 -1375 589
rect -1217 555 -1183 589
rect -1025 555 -991 589
rect -833 555 -799 589
rect -641 555 -607 589
rect -449 555 -415 589
rect -257 555 -223 589
rect -65 555 -31 589
rect 127 555 161 589
rect 319 555 353 589
rect 511 555 545 589
rect 703 555 737 589
rect 895 555 929 589
rect 1087 555 1121 589
rect 1279 555 1313 589
rect 1471 555 1505 589
rect 1663 555 1697 589
rect 1855 555 1889 589
rect 2047 555 2081 589
rect 2239 555 2273 589
rect 2431 555 2465 589
rect 2623 555 2657 589
rect 2815 555 2849 589
rect 3007 555 3041 589
rect 3199 555 3233 589
rect 3391 555 3425 589
rect 3583 555 3617 589
rect 3775 555 3809 589
rect 3967 555 4001 589
rect 4159 555 4193 589
rect 4351 555 4385 589
rect 4543 555 4577 589
rect 4735 555 4769 589
rect -4673 447 -4639 481
rect -4481 447 -4447 481
rect -4289 447 -4255 481
rect -4097 447 -4063 481
rect -3905 447 -3871 481
rect -3713 447 -3679 481
rect -3521 447 -3487 481
rect -3329 447 -3295 481
rect -3137 447 -3103 481
rect -2945 447 -2911 481
rect -2753 447 -2719 481
rect -2561 447 -2527 481
rect -2369 447 -2335 481
rect -2177 447 -2143 481
rect -1985 447 -1951 481
rect -1793 447 -1759 481
rect -1601 447 -1567 481
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect 1663 447 1697 481
rect 1855 447 1889 481
rect 2047 447 2081 481
rect 2239 447 2273 481
rect 2431 447 2465 481
rect 2623 447 2657 481
rect 2815 447 2849 481
rect 3007 447 3041 481
rect 3199 447 3233 481
rect 3391 447 3425 481
rect 3583 447 3617 481
rect 3775 447 3809 481
rect 3967 447 4001 481
rect 4159 447 4193 481
rect 4351 447 4385 481
rect 4543 447 4577 481
rect 4735 447 4769 481
rect -4817 121 -4783 397
rect -4721 121 -4687 397
rect -4625 121 -4591 397
rect -4529 121 -4495 397
rect -4433 121 -4399 397
rect -4337 121 -4303 397
rect -4241 121 -4207 397
rect -4145 121 -4111 397
rect -4049 121 -4015 397
rect -3953 121 -3919 397
rect -3857 121 -3823 397
rect -3761 121 -3727 397
rect -3665 121 -3631 397
rect -3569 121 -3535 397
rect -3473 121 -3439 397
rect -3377 121 -3343 397
rect -3281 121 -3247 397
rect -3185 121 -3151 397
rect -3089 121 -3055 397
rect -2993 121 -2959 397
rect -2897 121 -2863 397
rect -2801 121 -2767 397
rect -2705 121 -2671 397
rect -2609 121 -2575 397
rect -2513 121 -2479 397
rect -2417 121 -2383 397
rect -2321 121 -2287 397
rect -2225 121 -2191 397
rect -2129 121 -2095 397
rect -2033 121 -1999 397
rect -1937 121 -1903 397
rect -1841 121 -1807 397
rect -1745 121 -1711 397
rect -1649 121 -1615 397
rect -1553 121 -1519 397
rect -1457 121 -1423 397
rect -1361 121 -1327 397
rect -1265 121 -1231 397
rect -1169 121 -1135 397
rect -1073 121 -1039 397
rect -977 121 -943 397
rect -881 121 -847 397
rect -785 121 -751 397
rect -689 121 -655 397
rect -593 121 -559 397
rect -497 121 -463 397
rect -401 121 -367 397
rect -305 121 -271 397
rect -209 121 -175 397
rect -113 121 -79 397
rect -17 121 17 397
rect 79 121 113 397
rect 175 121 209 397
rect 271 121 305 397
rect 367 121 401 397
rect 463 121 497 397
rect 559 121 593 397
rect 655 121 689 397
rect 751 121 785 397
rect 847 121 881 397
rect 943 121 977 397
rect 1039 121 1073 397
rect 1135 121 1169 397
rect 1231 121 1265 397
rect 1327 121 1361 397
rect 1423 121 1457 397
rect 1519 121 1553 397
rect 1615 121 1649 397
rect 1711 121 1745 397
rect 1807 121 1841 397
rect 1903 121 1937 397
rect 1999 121 2033 397
rect 2095 121 2129 397
rect 2191 121 2225 397
rect 2287 121 2321 397
rect 2383 121 2417 397
rect 2479 121 2513 397
rect 2575 121 2609 397
rect 2671 121 2705 397
rect 2767 121 2801 397
rect 2863 121 2897 397
rect 2959 121 2993 397
rect 3055 121 3089 397
rect 3151 121 3185 397
rect 3247 121 3281 397
rect 3343 121 3377 397
rect 3439 121 3473 397
rect 3535 121 3569 397
rect 3631 121 3665 397
rect 3727 121 3761 397
rect 3823 121 3857 397
rect 3919 121 3953 397
rect 4015 121 4049 397
rect 4111 121 4145 397
rect 4207 121 4241 397
rect 4303 121 4337 397
rect 4399 121 4433 397
rect 4495 121 4529 397
rect 4591 121 4625 397
rect 4687 121 4721 397
rect 4783 121 4817 397
rect -4769 37 -4735 71
rect -4577 37 -4543 71
rect -4385 37 -4351 71
rect -4193 37 -4159 71
rect -4001 37 -3967 71
rect -3809 37 -3775 71
rect -3617 37 -3583 71
rect -3425 37 -3391 71
rect -3233 37 -3199 71
rect -3041 37 -3007 71
rect -2849 37 -2815 71
rect -2657 37 -2623 71
rect -2465 37 -2431 71
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect 2527 37 2561 71
rect 2719 37 2753 71
rect 2911 37 2945 71
rect 3103 37 3137 71
rect 3295 37 3329 71
rect 3487 37 3521 71
rect 3679 37 3713 71
rect 3871 37 3905 71
rect 4063 37 4097 71
rect 4255 37 4289 71
rect 4447 37 4481 71
rect 4639 37 4673 71
rect -4769 -71 -4735 -37
rect -4577 -71 -4543 -37
rect -4385 -71 -4351 -37
rect -4193 -71 -4159 -37
rect -4001 -71 -3967 -37
rect -3809 -71 -3775 -37
rect -3617 -71 -3583 -37
rect -3425 -71 -3391 -37
rect -3233 -71 -3199 -37
rect -3041 -71 -3007 -37
rect -2849 -71 -2815 -37
rect -2657 -71 -2623 -37
rect -2465 -71 -2431 -37
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect 2527 -71 2561 -37
rect 2719 -71 2753 -37
rect 2911 -71 2945 -37
rect 3103 -71 3137 -37
rect 3295 -71 3329 -37
rect 3487 -71 3521 -37
rect 3679 -71 3713 -37
rect 3871 -71 3905 -37
rect 4063 -71 4097 -37
rect 4255 -71 4289 -37
rect 4447 -71 4481 -37
rect 4639 -71 4673 -37
rect -4817 -397 -4783 -121
rect -4721 -397 -4687 -121
rect -4625 -397 -4591 -121
rect -4529 -397 -4495 -121
rect -4433 -397 -4399 -121
rect -4337 -397 -4303 -121
rect -4241 -397 -4207 -121
rect -4145 -397 -4111 -121
rect -4049 -397 -4015 -121
rect -3953 -397 -3919 -121
rect -3857 -397 -3823 -121
rect -3761 -397 -3727 -121
rect -3665 -397 -3631 -121
rect -3569 -397 -3535 -121
rect -3473 -397 -3439 -121
rect -3377 -397 -3343 -121
rect -3281 -397 -3247 -121
rect -3185 -397 -3151 -121
rect -3089 -397 -3055 -121
rect -2993 -397 -2959 -121
rect -2897 -397 -2863 -121
rect -2801 -397 -2767 -121
rect -2705 -397 -2671 -121
rect -2609 -397 -2575 -121
rect -2513 -397 -2479 -121
rect -2417 -397 -2383 -121
rect -2321 -397 -2287 -121
rect -2225 -397 -2191 -121
rect -2129 -397 -2095 -121
rect -2033 -397 -1999 -121
rect -1937 -397 -1903 -121
rect -1841 -397 -1807 -121
rect -1745 -397 -1711 -121
rect -1649 -397 -1615 -121
rect -1553 -397 -1519 -121
rect -1457 -397 -1423 -121
rect -1361 -397 -1327 -121
rect -1265 -397 -1231 -121
rect -1169 -397 -1135 -121
rect -1073 -397 -1039 -121
rect -977 -397 -943 -121
rect -881 -397 -847 -121
rect -785 -397 -751 -121
rect -689 -397 -655 -121
rect -593 -397 -559 -121
rect -497 -397 -463 -121
rect -401 -397 -367 -121
rect -305 -397 -271 -121
rect -209 -397 -175 -121
rect -113 -397 -79 -121
rect -17 -397 17 -121
rect 79 -397 113 -121
rect 175 -397 209 -121
rect 271 -397 305 -121
rect 367 -397 401 -121
rect 463 -397 497 -121
rect 559 -397 593 -121
rect 655 -397 689 -121
rect 751 -397 785 -121
rect 847 -397 881 -121
rect 943 -397 977 -121
rect 1039 -397 1073 -121
rect 1135 -397 1169 -121
rect 1231 -397 1265 -121
rect 1327 -397 1361 -121
rect 1423 -397 1457 -121
rect 1519 -397 1553 -121
rect 1615 -397 1649 -121
rect 1711 -397 1745 -121
rect 1807 -397 1841 -121
rect 1903 -397 1937 -121
rect 1999 -397 2033 -121
rect 2095 -397 2129 -121
rect 2191 -397 2225 -121
rect 2287 -397 2321 -121
rect 2383 -397 2417 -121
rect 2479 -397 2513 -121
rect 2575 -397 2609 -121
rect 2671 -397 2705 -121
rect 2767 -397 2801 -121
rect 2863 -397 2897 -121
rect 2959 -397 2993 -121
rect 3055 -397 3089 -121
rect 3151 -397 3185 -121
rect 3247 -397 3281 -121
rect 3343 -397 3377 -121
rect 3439 -397 3473 -121
rect 3535 -397 3569 -121
rect 3631 -397 3665 -121
rect 3727 -397 3761 -121
rect 3823 -397 3857 -121
rect 3919 -397 3953 -121
rect 4015 -397 4049 -121
rect 4111 -397 4145 -121
rect 4207 -397 4241 -121
rect 4303 -397 4337 -121
rect 4399 -397 4433 -121
rect 4495 -397 4529 -121
rect 4591 -397 4625 -121
rect 4687 -397 4721 -121
rect 4783 -397 4817 -121
rect -4673 -481 -4639 -447
rect -4481 -481 -4447 -447
rect -4289 -481 -4255 -447
rect -4097 -481 -4063 -447
rect -3905 -481 -3871 -447
rect -3713 -481 -3679 -447
rect -3521 -481 -3487 -447
rect -3329 -481 -3295 -447
rect -3137 -481 -3103 -447
rect -2945 -481 -2911 -447
rect -2753 -481 -2719 -447
rect -2561 -481 -2527 -447
rect -2369 -481 -2335 -447
rect -2177 -481 -2143 -447
rect -1985 -481 -1951 -447
rect -1793 -481 -1759 -447
rect -1601 -481 -1567 -447
rect -1409 -481 -1375 -447
rect -1217 -481 -1183 -447
rect -1025 -481 -991 -447
rect -833 -481 -799 -447
rect -641 -481 -607 -447
rect -449 -481 -415 -447
rect -257 -481 -223 -447
rect -65 -481 -31 -447
rect 127 -481 161 -447
rect 319 -481 353 -447
rect 511 -481 545 -447
rect 703 -481 737 -447
rect 895 -481 929 -447
rect 1087 -481 1121 -447
rect 1279 -481 1313 -447
rect 1471 -481 1505 -447
rect 1663 -481 1697 -447
rect 1855 -481 1889 -447
rect 2047 -481 2081 -447
rect 2239 -481 2273 -447
rect 2431 -481 2465 -447
rect 2623 -481 2657 -447
rect 2815 -481 2849 -447
rect 3007 -481 3041 -447
rect 3199 -481 3233 -447
rect 3391 -481 3425 -447
rect 3583 -481 3617 -447
rect 3775 -481 3809 -447
rect 3967 -481 4001 -447
rect 4159 -481 4193 -447
rect 4351 -481 4385 -447
rect 4543 -481 4577 -447
rect 4735 -481 4769 -447
rect -4673 -589 -4639 -555
rect -4481 -589 -4447 -555
rect -4289 -589 -4255 -555
rect -4097 -589 -4063 -555
rect -3905 -589 -3871 -555
rect -3713 -589 -3679 -555
rect -3521 -589 -3487 -555
rect -3329 -589 -3295 -555
rect -3137 -589 -3103 -555
rect -2945 -589 -2911 -555
rect -2753 -589 -2719 -555
rect -2561 -589 -2527 -555
rect -2369 -589 -2335 -555
rect -2177 -589 -2143 -555
rect -1985 -589 -1951 -555
rect -1793 -589 -1759 -555
rect -1601 -589 -1567 -555
rect -1409 -589 -1375 -555
rect -1217 -589 -1183 -555
rect -1025 -589 -991 -555
rect -833 -589 -799 -555
rect -641 -589 -607 -555
rect -449 -589 -415 -555
rect -257 -589 -223 -555
rect -65 -589 -31 -555
rect 127 -589 161 -555
rect 319 -589 353 -555
rect 511 -589 545 -555
rect 703 -589 737 -555
rect 895 -589 929 -555
rect 1087 -589 1121 -555
rect 1279 -589 1313 -555
rect 1471 -589 1505 -555
rect 1663 -589 1697 -555
rect 1855 -589 1889 -555
rect 2047 -589 2081 -555
rect 2239 -589 2273 -555
rect 2431 -589 2465 -555
rect 2623 -589 2657 -555
rect 2815 -589 2849 -555
rect 3007 -589 3041 -555
rect 3199 -589 3233 -555
rect 3391 -589 3425 -555
rect 3583 -589 3617 -555
rect 3775 -589 3809 -555
rect 3967 -589 4001 -555
rect 4159 -589 4193 -555
rect 4351 -589 4385 -555
rect 4543 -589 4577 -555
rect 4735 -589 4769 -555
rect -4817 -915 -4783 -639
rect -4721 -915 -4687 -639
rect -4625 -915 -4591 -639
rect -4529 -915 -4495 -639
rect -4433 -915 -4399 -639
rect -4337 -915 -4303 -639
rect -4241 -915 -4207 -639
rect -4145 -915 -4111 -639
rect -4049 -915 -4015 -639
rect -3953 -915 -3919 -639
rect -3857 -915 -3823 -639
rect -3761 -915 -3727 -639
rect -3665 -915 -3631 -639
rect -3569 -915 -3535 -639
rect -3473 -915 -3439 -639
rect -3377 -915 -3343 -639
rect -3281 -915 -3247 -639
rect -3185 -915 -3151 -639
rect -3089 -915 -3055 -639
rect -2993 -915 -2959 -639
rect -2897 -915 -2863 -639
rect -2801 -915 -2767 -639
rect -2705 -915 -2671 -639
rect -2609 -915 -2575 -639
rect -2513 -915 -2479 -639
rect -2417 -915 -2383 -639
rect -2321 -915 -2287 -639
rect -2225 -915 -2191 -639
rect -2129 -915 -2095 -639
rect -2033 -915 -1999 -639
rect -1937 -915 -1903 -639
rect -1841 -915 -1807 -639
rect -1745 -915 -1711 -639
rect -1649 -915 -1615 -639
rect -1553 -915 -1519 -639
rect -1457 -915 -1423 -639
rect -1361 -915 -1327 -639
rect -1265 -915 -1231 -639
rect -1169 -915 -1135 -639
rect -1073 -915 -1039 -639
rect -977 -915 -943 -639
rect -881 -915 -847 -639
rect -785 -915 -751 -639
rect -689 -915 -655 -639
rect -593 -915 -559 -639
rect -497 -915 -463 -639
rect -401 -915 -367 -639
rect -305 -915 -271 -639
rect -209 -915 -175 -639
rect -113 -915 -79 -639
rect -17 -915 17 -639
rect 79 -915 113 -639
rect 175 -915 209 -639
rect 271 -915 305 -639
rect 367 -915 401 -639
rect 463 -915 497 -639
rect 559 -915 593 -639
rect 655 -915 689 -639
rect 751 -915 785 -639
rect 847 -915 881 -639
rect 943 -915 977 -639
rect 1039 -915 1073 -639
rect 1135 -915 1169 -639
rect 1231 -915 1265 -639
rect 1327 -915 1361 -639
rect 1423 -915 1457 -639
rect 1519 -915 1553 -639
rect 1615 -915 1649 -639
rect 1711 -915 1745 -639
rect 1807 -915 1841 -639
rect 1903 -915 1937 -639
rect 1999 -915 2033 -639
rect 2095 -915 2129 -639
rect 2191 -915 2225 -639
rect 2287 -915 2321 -639
rect 2383 -915 2417 -639
rect 2479 -915 2513 -639
rect 2575 -915 2609 -639
rect 2671 -915 2705 -639
rect 2767 -915 2801 -639
rect 2863 -915 2897 -639
rect 2959 -915 2993 -639
rect 3055 -915 3089 -639
rect 3151 -915 3185 -639
rect 3247 -915 3281 -639
rect 3343 -915 3377 -639
rect 3439 -915 3473 -639
rect 3535 -915 3569 -639
rect 3631 -915 3665 -639
rect 3727 -915 3761 -639
rect 3823 -915 3857 -639
rect 3919 -915 3953 -639
rect 4015 -915 4049 -639
rect 4111 -915 4145 -639
rect 4207 -915 4241 -639
rect 4303 -915 4337 -639
rect 4399 -915 4433 -639
rect 4495 -915 4529 -639
rect 4591 -915 4625 -639
rect 4687 -915 4721 -639
rect 4783 -915 4817 -639
rect -4769 -999 -4735 -965
rect -4577 -999 -4543 -965
rect -4385 -999 -4351 -965
rect -4193 -999 -4159 -965
rect -4001 -999 -3967 -965
rect -3809 -999 -3775 -965
rect -3617 -999 -3583 -965
rect -3425 -999 -3391 -965
rect -3233 -999 -3199 -965
rect -3041 -999 -3007 -965
rect -2849 -999 -2815 -965
rect -2657 -999 -2623 -965
rect -2465 -999 -2431 -965
rect -2273 -999 -2239 -965
rect -2081 -999 -2047 -965
rect -1889 -999 -1855 -965
rect -1697 -999 -1663 -965
rect -1505 -999 -1471 -965
rect -1313 -999 -1279 -965
rect -1121 -999 -1087 -965
rect -929 -999 -895 -965
rect -737 -999 -703 -965
rect -545 -999 -511 -965
rect -353 -999 -319 -965
rect -161 -999 -127 -965
rect 31 -999 65 -965
rect 223 -999 257 -965
rect 415 -999 449 -965
rect 607 -999 641 -965
rect 799 -999 833 -965
rect 991 -999 1025 -965
rect 1183 -999 1217 -965
rect 1375 -999 1409 -965
rect 1567 -999 1601 -965
rect 1759 -999 1793 -965
rect 1951 -999 1985 -965
rect 2143 -999 2177 -965
rect 2335 -999 2369 -965
rect 2527 -999 2561 -965
rect 2719 -999 2753 -965
rect 2911 -999 2945 -965
rect 3103 -999 3137 -965
rect 3295 -999 3329 -965
rect 3487 -999 3521 -965
rect 3679 -999 3713 -965
rect 3871 -999 3905 -965
rect 4063 -999 4097 -965
rect 4255 -999 4289 -965
rect 4447 -999 4481 -965
rect 4639 -999 4673 -965
<< metal1 >>
rect -4781 999 -4723 1005
rect -4781 965 -4769 999
rect -4735 965 -4723 999
rect -4781 959 -4723 965
rect -4589 999 -4531 1005
rect -4589 965 -4577 999
rect -4543 965 -4531 999
rect -4589 959 -4531 965
rect -4397 999 -4339 1005
rect -4397 965 -4385 999
rect -4351 965 -4339 999
rect -4397 959 -4339 965
rect -4205 999 -4147 1005
rect -4205 965 -4193 999
rect -4159 965 -4147 999
rect -4205 959 -4147 965
rect -4013 999 -3955 1005
rect -4013 965 -4001 999
rect -3967 965 -3955 999
rect -4013 959 -3955 965
rect -3821 999 -3763 1005
rect -3821 965 -3809 999
rect -3775 965 -3763 999
rect -3821 959 -3763 965
rect -3629 999 -3571 1005
rect -3629 965 -3617 999
rect -3583 965 -3571 999
rect -3629 959 -3571 965
rect -3437 999 -3379 1005
rect -3437 965 -3425 999
rect -3391 965 -3379 999
rect -3437 959 -3379 965
rect -3245 999 -3187 1005
rect -3245 965 -3233 999
rect -3199 965 -3187 999
rect -3245 959 -3187 965
rect -3053 999 -2995 1005
rect -3053 965 -3041 999
rect -3007 965 -2995 999
rect -3053 959 -2995 965
rect -2861 999 -2803 1005
rect -2861 965 -2849 999
rect -2815 965 -2803 999
rect -2861 959 -2803 965
rect -2669 999 -2611 1005
rect -2669 965 -2657 999
rect -2623 965 -2611 999
rect -2669 959 -2611 965
rect -2477 999 -2419 1005
rect -2477 965 -2465 999
rect -2431 965 -2419 999
rect -2477 959 -2419 965
rect -2285 999 -2227 1005
rect -2285 965 -2273 999
rect -2239 965 -2227 999
rect -2285 959 -2227 965
rect -2093 999 -2035 1005
rect -2093 965 -2081 999
rect -2047 965 -2035 999
rect -2093 959 -2035 965
rect -1901 999 -1843 1005
rect -1901 965 -1889 999
rect -1855 965 -1843 999
rect -1901 959 -1843 965
rect -1709 999 -1651 1005
rect -1709 965 -1697 999
rect -1663 965 -1651 999
rect -1709 959 -1651 965
rect -1517 999 -1459 1005
rect -1517 965 -1505 999
rect -1471 965 -1459 999
rect -1517 959 -1459 965
rect -1325 999 -1267 1005
rect -1325 965 -1313 999
rect -1279 965 -1267 999
rect -1325 959 -1267 965
rect -1133 999 -1075 1005
rect -1133 965 -1121 999
rect -1087 965 -1075 999
rect -1133 959 -1075 965
rect -941 999 -883 1005
rect -941 965 -929 999
rect -895 965 -883 999
rect -941 959 -883 965
rect -749 999 -691 1005
rect -749 965 -737 999
rect -703 965 -691 999
rect -749 959 -691 965
rect -557 999 -499 1005
rect -557 965 -545 999
rect -511 965 -499 999
rect -557 959 -499 965
rect -365 999 -307 1005
rect -365 965 -353 999
rect -319 965 -307 999
rect -365 959 -307 965
rect -173 999 -115 1005
rect -173 965 -161 999
rect -127 965 -115 999
rect -173 959 -115 965
rect 19 999 77 1005
rect 19 965 31 999
rect 65 965 77 999
rect 19 959 77 965
rect 211 999 269 1005
rect 211 965 223 999
rect 257 965 269 999
rect 211 959 269 965
rect 403 999 461 1005
rect 403 965 415 999
rect 449 965 461 999
rect 403 959 461 965
rect 595 999 653 1005
rect 595 965 607 999
rect 641 965 653 999
rect 595 959 653 965
rect 787 999 845 1005
rect 787 965 799 999
rect 833 965 845 999
rect 787 959 845 965
rect 979 999 1037 1005
rect 979 965 991 999
rect 1025 965 1037 999
rect 979 959 1037 965
rect 1171 999 1229 1005
rect 1171 965 1183 999
rect 1217 965 1229 999
rect 1171 959 1229 965
rect 1363 999 1421 1005
rect 1363 965 1375 999
rect 1409 965 1421 999
rect 1363 959 1421 965
rect 1555 999 1613 1005
rect 1555 965 1567 999
rect 1601 965 1613 999
rect 1555 959 1613 965
rect 1747 999 1805 1005
rect 1747 965 1759 999
rect 1793 965 1805 999
rect 1747 959 1805 965
rect 1939 999 1997 1005
rect 1939 965 1951 999
rect 1985 965 1997 999
rect 1939 959 1997 965
rect 2131 999 2189 1005
rect 2131 965 2143 999
rect 2177 965 2189 999
rect 2131 959 2189 965
rect 2323 999 2381 1005
rect 2323 965 2335 999
rect 2369 965 2381 999
rect 2323 959 2381 965
rect 2515 999 2573 1005
rect 2515 965 2527 999
rect 2561 965 2573 999
rect 2515 959 2573 965
rect 2707 999 2765 1005
rect 2707 965 2719 999
rect 2753 965 2765 999
rect 2707 959 2765 965
rect 2899 999 2957 1005
rect 2899 965 2911 999
rect 2945 965 2957 999
rect 2899 959 2957 965
rect 3091 999 3149 1005
rect 3091 965 3103 999
rect 3137 965 3149 999
rect 3091 959 3149 965
rect 3283 999 3341 1005
rect 3283 965 3295 999
rect 3329 965 3341 999
rect 3283 959 3341 965
rect 3475 999 3533 1005
rect 3475 965 3487 999
rect 3521 965 3533 999
rect 3475 959 3533 965
rect 3667 999 3725 1005
rect 3667 965 3679 999
rect 3713 965 3725 999
rect 3667 959 3725 965
rect 3859 999 3917 1005
rect 3859 965 3871 999
rect 3905 965 3917 999
rect 3859 959 3917 965
rect 4051 999 4109 1005
rect 4051 965 4063 999
rect 4097 965 4109 999
rect 4051 959 4109 965
rect 4243 999 4301 1005
rect 4243 965 4255 999
rect 4289 965 4301 999
rect 4243 959 4301 965
rect 4435 999 4493 1005
rect 4435 965 4447 999
rect 4481 965 4493 999
rect 4435 959 4493 965
rect 4627 999 4685 1005
rect 4627 965 4639 999
rect 4673 965 4685 999
rect 4627 959 4685 965
rect -4823 915 -4777 927
rect -4823 639 -4817 915
rect -4783 639 -4777 915
rect -4823 627 -4777 639
rect -4727 915 -4681 927
rect -4727 639 -4721 915
rect -4687 639 -4681 915
rect -4727 627 -4681 639
rect -4631 915 -4585 927
rect -4631 639 -4625 915
rect -4591 639 -4585 915
rect -4631 627 -4585 639
rect -4535 915 -4489 927
rect -4535 639 -4529 915
rect -4495 639 -4489 915
rect -4535 627 -4489 639
rect -4439 915 -4393 927
rect -4439 639 -4433 915
rect -4399 639 -4393 915
rect -4439 627 -4393 639
rect -4343 915 -4297 927
rect -4343 639 -4337 915
rect -4303 639 -4297 915
rect -4343 627 -4297 639
rect -4247 915 -4201 927
rect -4247 639 -4241 915
rect -4207 639 -4201 915
rect -4247 627 -4201 639
rect -4151 915 -4105 927
rect -4151 639 -4145 915
rect -4111 639 -4105 915
rect -4151 627 -4105 639
rect -4055 915 -4009 927
rect -4055 639 -4049 915
rect -4015 639 -4009 915
rect -4055 627 -4009 639
rect -3959 915 -3913 927
rect -3959 639 -3953 915
rect -3919 639 -3913 915
rect -3959 627 -3913 639
rect -3863 915 -3817 927
rect -3863 639 -3857 915
rect -3823 639 -3817 915
rect -3863 627 -3817 639
rect -3767 915 -3721 927
rect -3767 639 -3761 915
rect -3727 639 -3721 915
rect -3767 627 -3721 639
rect -3671 915 -3625 927
rect -3671 639 -3665 915
rect -3631 639 -3625 915
rect -3671 627 -3625 639
rect -3575 915 -3529 927
rect -3575 639 -3569 915
rect -3535 639 -3529 915
rect -3575 627 -3529 639
rect -3479 915 -3433 927
rect -3479 639 -3473 915
rect -3439 639 -3433 915
rect -3479 627 -3433 639
rect -3383 915 -3337 927
rect -3383 639 -3377 915
rect -3343 639 -3337 915
rect -3383 627 -3337 639
rect -3287 915 -3241 927
rect -3287 639 -3281 915
rect -3247 639 -3241 915
rect -3287 627 -3241 639
rect -3191 915 -3145 927
rect -3191 639 -3185 915
rect -3151 639 -3145 915
rect -3191 627 -3145 639
rect -3095 915 -3049 927
rect -3095 639 -3089 915
rect -3055 639 -3049 915
rect -3095 627 -3049 639
rect -2999 915 -2953 927
rect -2999 639 -2993 915
rect -2959 639 -2953 915
rect -2999 627 -2953 639
rect -2903 915 -2857 927
rect -2903 639 -2897 915
rect -2863 639 -2857 915
rect -2903 627 -2857 639
rect -2807 915 -2761 927
rect -2807 639 -2801 915
rect -2767 639 -2761 915
rect -2807 627 -2761 639
rect -2711 915 -2665 927
rect -2711 639 -2705 915
rect -2671 639 -2665 915
rect -2711 627 -2665 639
rect -2615 915 -2569 927
rect -2615 639 -2609 915
rect -2575 639 -2569 915
rect -2615 627 -2569 639
rect -2519 915 -2473 927
rect -2519 639 -2513 915
rect -2479 639 -2473 915
rect -2519 627 -2473 639
rect -2423 915 -2377 927
rect -2423 639 -2417 915
rect -2383 639 -2377 915
rect -2423 627 -2377 639
rect -2327 915 -2281 927
rect -2327 639 -2321 915
rect -2287 639 -2281 915
rect -2327 627 -2281 639
rect -2231 915 -2185 927
rect -2231 639 -2225 915
rect -2191 639 -2185 915
rect -2231 627 -2185 639
rect -2135 915 -2089 927
rect -2135 639 -2129 915
rect -2095 639 -2089 915
rect -2135 627 -2089 639
rect -2039 915 -1993 927
rect -2039 639 -2033 915
rect -1999 639 -1993 915
rect -2039 627 -1993 639
rect -1943 915 -1897 927
rect -1943 639 -1937 915
rect -1903 639 -1897 915
rect -1943 627 -1897 639
rect -1847 915 -1801 927
rect -1847 639 -1841 915
rect -1807 639 -1801 915
rect -1847 627 -1801 639
rect -1751 915 -1705 927
rect -1751 639 -1745 915
rect -1711 639 -1705 915
rect -1751 627 -1705 639
rect -1655 915 -1609 927
rect -1655 639 -1649 915
rect -1615 639 -1609 915
rect -1655 627 -1609 639
rect -1559 915 -1513 927
rect -1559 639 -1553 915
rect -1519 639 -1513 915
rect -1559 627 -1513 639
rect -1463 915 -1417 927
rect -1463 639 -1457 915
rect -1423 639 -1417 915
rect -1463 627 -1417 639
rect -1367 915 -1321 927
rect -1367 639 -1361 915
rect -1327 639 -1321 915
rect -1367 627 -1321 639
rect -1271 915 -1225 927
rect -1271 639 -1265 915
rect -1231 639 -1225 915
rect -1271 627 -1225 639
rect -1175 915 -1129 927
rect -1175 639 -1169 915
rect -1135 639 -1129 915
rect -1175 627 -1129 639
rect -1079 915 -1033 927
rect -1079 639 -1073 915
rect -1039 639 -1033 915
rect -1079 627 -1033 639
rect -983 915 -937 927
rect -983 639 -977 915
rect -943 639 -937 915
rect -983 627 -937 639
rect -887 915 -841 927
rect -887 639 -881 915
rect -847 639 -841 915
rect -887 627 -841 639
rect -791 915 -745 927
rect -791 639 -785 915
rect -751 639 -745 915
rect -791 627 -745 639
rect -695 915 -649 927
rect -695 639 -689 915
rect -655 639 -649 915
rect -695 627 -649 639
rect -599 915 -553 927
rect -599 639 -593 915
rect -559 639 -553 915
rect -599 627 -553 639
rect -503 915 -457 927
rect -503 639 -497 915
rect -463 639 -457 915
rect -503 627 -457 639
rect -407 915 -361 927
rect -407 639 -401 915
rect -367 639 -361 915
rect -407 627 -361 639
rect -311 915 -265 927
rect -311 639 -305 915
rect -271 639 -265 915
rect -311 627 -265 639
rect -215 915 -169 927
rect -215 639 -209 915
rect -175 639 -169 915
rect -215 627 -169 639
rect -119 915 -73 927
rect -119 639 -113 915
rect -79 639 -73 915
rect -119 627 -73 639
rect -23 915 23 927
rect -23 639 -17 915
rect 17 639 23 915
rect -23 627 23 639
rect 73 915 119 927
rect 73 639 79 915
rect 113 639 119 915
rect 73 627 119 639
rect 169 915 215 927
rect 169 639 175 915
rect 209 639 215 915
rect 169 627 215 639
rect 265 915 311 927
rect 265 639 271 915
rect 305 639 311 915
rect 265 627 311 639
rect 361 915 407 927
rect 361 639 367 915
rect 401 639 407 915
rect 361 627 407 639
rect 457 915 503 927
rect 457 639 463 915
rect 497 639 503 915
rect 457 627 503 639
rect 553 915 599 927
rect 553 639 559 915
rect 593 639 599 915
rect 553 627 599 639
rect 649 915 695 927
rect 649 639 655 915
rect 689 639 695 915
rect 649 627 695 639
rect 745 915 791 927
rect 745 639 751 915
rect 785 639 791 915
rect 745 627 791 639
rect 841 915 887 927
rect 841 639 847 915
rect 881 639 887 915
rect 841 627 887 639
rect 937 915 983 927
rect 937 639 943 915
rect 977 639 983 915
rect 937 627 983 639
rect 1033 915 1079 927
rect 1033 639 1039 915
rect 1073 639 1079 915
rect 1033 627 1079 639
rect 1129 915 1175 927
rect 1129 639 1135 915
rect 1169 639 1175 915
rect 1129 627 1175 639
rect 1225 915 1271 927
rect 1225 639 1231 915
rect 1265 639 1271 915
rect 1225 627 1271 639
rect 1321 915 1367 927
rect 1321 639 1327 915
rect 1361 639 1367 915
rect 1321 627 1367 639
rect 1417 915 1463 927
rect 1417 639 1423 915
rect 1457 639 1463 915
rect 1417 627 1463 639
rect 1513 915 1559 927
rect 1513 639 1519 915
rect 1553 639 1559 915
rect 1513 627 1559 639
rect 1609 915 1655 927
rect 1609 639 1615 915
rect 1649 639 1655 915
rect 1609 627 1655 639
rect 1705 915 1751 927
rect 1705 639 1711 915
rect 1745 639 1751 915
rect 1705 627 1751 639
rect 1801 915 1847 927
rect 1801 639 1807 915
rect 1841 639 1847 915
rect 1801 627 1847 639
rect 1897 915 1943 927
rect 1897 639 1903 915
rect 1937 639 1943 915
rect 1897 627 1943 639
rect 1993 915 2039 927
rect 1993 639 1999 915
rect 2033 639 2039 915
rect 1993 627 2039 639
rect 2089 915 2135 927
rect 2089 639 2095 915
rect 2129 639 2135 915
rect 2089 627 2135 639
rect 2185 915 2231 927
rect 2185 639 2191 915
rect 2225 639 2231 915
rect 2185 627 2231 639
rect 2281 915 2327 927
rect 2281 639 2287 915
rect 2321 639 2327 915
rect 2281 627 2327 639
rect 2377 915 2423 927
rect 2377 639 2383 915
rect 2417 639 2423 915
rect 2377 627 2423 639
rect 2473 915 2519 927
rect 2473 639 2479 915
rect 2513 639 2519 915
rect 2473 627 2519 639
rect 2569 915 2615 927
rect 2569 639 2575 915
rect 2609 639 2615 915
rect 2569 627 2615 639
rect 2665 915 2711 927
rect 2665 639 2671 915
rect 2705 639 2711 915
rect 2665 627 2711 639
rect 2761 915 2807 927
rect 2761 639 2767 915
rect 2801 639 2807 915
rect 2761 627 2807 639
rect 2857 915 2903 927
rect 2857 639 2863 915
rect 2897 639 2903 915
rect 2857 627 2903 639
rect 2953 915 2999 927
rect 2953 639 2959 915
rect 2993 639 2999 915
rect 2953 627 2999 639
rect 3049 915 3095 927
rect 3049 639 3055 915
rect 3089 639 3095 915
rect 3049 627 3095 639
rect 3145 915 3191 927
rect 3145 639 3151 915
rect 3185 639 3191 915
rect 3145 627 3191 639
rect 3241 915 3287 927
rect 3241 639 3247 915
rect 3281 639 3287 915
rect 3241 627 3287 639
rect 3337 915 3383 927
rect 3337 639 3343 915
rect 3377 639 3383 915
rect 3337 627 3383 639
rect 3433 915 3479 927
rect 3433 639 3439 915
rect 3473 639 3479 915
rect 3433 627 3479 639
rect 3529 915 3575 927
rect 3529 639 3535 915
rect 3569 639 3575 915
rect 3529 627 3575 639
rect 3625 915 3671 927
rect 3625 639 3631 915
rect 3665 639 3671 915
rect 3625 627 3671 639
rect 3721 915 3767 927
rect 3721 639 3727 915
rect 3761 639 3767 915
rect 3721 627 3767 639
rect 3817 915 3863 927
rect 3817 639 3823 915
rect 3857 639 3863 915
rect 3817 627 3863 639
rect 3913 915 3959 927
rect 3913 639 3919 915
rect 3953 639 3959 915
rect 3913 627 3959 639
rect 4009 915 4055 927
rect 4009 639 4015 915
rect 4049 639 4055 915
rect 4009 627 4055 639
rect 4105 915 4151 927
rect 4105 639 4111 915
rect 4145 639 4151 915
rect 4105 627 4151 639
rect 4201 915 4247 927
rect 4201 639 4207 915
rect 4241 639 4247 915
rect 4201 627 4247 639
rect 4297 915 4343 927
rect 4297 639 4303 915
rect 4337 639 4343 915
rect 4297 627 4343 639
rect 4393 915 4439 927
rect 4393 639 4399 915
rect 4433 639 4439 915
rect 4393 627 4439 639
rect 4489 915 4535 927
rect 4489 639 4495 915
rect 4529 639 4535 915
rect 4489 627 4535 639
rect 4585 915 4631 927
rect 4585 639 4591 915
rect 4625 639 4631 915
rect 4585 627 4631 639
rect 4681 915 4727 927
rect 4681 639 4687 915
rect 4721 639 4727 915
rect 4681 627 4727 639
rect 4777 915 4823 927
rect 4777 639 4783 915
rect 4817 639 4823 915
rect 4777 627 4823 639
rect -4685 589 -4627 595
rect -4685 555 -4673 589
rect -4639 555 -4627 589
rect -4685 549 -4627 555
rect -4493 589 -4435 595
rect -4493 555 -4481 589
rect -4447 555 -4435 589
rect -4493 549 -4435 555
rect -4301 589 -4243 595
rect -4301 555 -4289 589
rect -4255 555 -4243 589
rect -4301 549 -4243 555
rect -4109 589 -4051 595
rect -4109 555 -4097 589
rect -4063 555 -4051 589
rect -4109 549 -4051 555
rect -3917 589 -3859 595
rect -3917 555 -3905 589
rect -3871 555 -3859 589
rect -3917 549 -3859 555
rect -3725 589 -3667 595
rect -3725 555 -3713 589
rect -3679 555 -3667 589
rect -3725 549 -3667 555
rect -3533 589 -3475 595
rect -3533 555 -3521 589
rect -3487 555 -3475 589
rect -3533 549 -3475 555
rect -3341 589 -3283 595
rect -3341 555 -3329 589
rect -3295 555 -3283 589
rect -3341 549 -3283 555
rect -3149 589 -3091 595
rect -3149 555 -3137 589
rect -3103 555 -3091 589
rect -3149 549 -3091 555
rect -2957 589 -2899 595
rect -2957 555 -2945 589
rect -2911 555 -2899 589
rect -2957 549 -2899 555
rect -2765 589 -2707 595
rect -2765 555 -2753 589
rect -2719 555 -2707 589
rect -2765 549 -2707 555
rect -2573 589 -2515 595
rect -2573 555 -2561 589
rect -2527 555 -2515 589
rect -2573 549 -2515 555
rect -2381 589 -2323 595
rect -2381 555 -2369 589
rect -2335 555 -2323 589
rect -2381 549 -2323 555
rect -2189 589 -2131 595
rect -2189 555 -2177 589
rect -2143 555 -2131 589
rect -2189 549 -2131 555
rect -1997 589 -1939 595
rect -1997 555 -1985 589
rect -1951 555 -1939 589
rect -1997 549 -1939 555
rect -1805 589 -1747 595
rect -1805 555 -1793 589
rect -1759 555 -1747 589
rect -1805 549 -1747 555
rect -1613 589 -1555 595
rect -1613 555 -1601 589
rect -1567 555 -1555 589
rect -1613 549 -1555 555
rect -1421 589 -1363 595
rect -1421 555 -1409 589
rect -1375 555 -1363 589
rect -1421 549 -1363 555
rect -1229 589 -1171 595
rect -1229 555 -1217 589
rect -1183 555 -1171 589
rect -1229 549 -1171 555
rect -1037 589 -979 595
rect -1037 555 -1025 589
rect -991 555 -979 589
rect -1037 549 -979 555
rect -845 589 -787 595
rect -845 555 -833 589
rect -799 555 -787 589
rect -845 549 -787 555
rect -653 589 -595 595
rect -653 555 -641 589
rect -607 555 -595 589
rect -653 549 -595 555
rect -461 589 -403 595
rect -461 555 -449 589
rect -415 555 -403 589
rect -461 549 -403 555
rect -269 589 -211 595
rect -269 555 -257 589
rect -223 555 -211 589
rect -269 549 -211 555
rect -77 589 -19 595
rect -77 555 -65 589
rect -31 555 -19 589
rect -77 549 -19 555
rect 115 589 173 595
rect 115 555 127 589
rect 161 555 173 589
rect 115 549 173 555
rect 307 589 365 595
rect 307 555 319 589
rect 353 555 365 589
rect 307 549 365 555
rect 499 589 557 595
rect 499 555 511 589
rect 545 555 557 589
rect 499 549 557 555
rect 691 589 749 595
rect 691 555 703 589
rect 737 555 749 589
rect 691 549 749 555
rect 883 589 941 595
rect 883 555 895 589
rect 929 555 941 589
rect 883 549 941 555
rect 1075 589 1133 595
rect 1075 555 1087 589
rect 1121 555 1133 589
rect 1075 549 1133 555
rect 1267 589 1325 595
rect 1267 555 1279 589
rect 1313 555 1325 589
rect 1267 549 1325 555
rect 1459 589 1517 595
rect 1459 555 1471 589
rect 1505 555 1517 589
rect 1459 549 1517 555
rect 1651 589 1709 595
rect 1651 555 1663 589
rect 1697 555 1709 589
rect 1651 549 1709 555
rect 1843 589 1901 595
rect 1843 555 1855 589
rect 1889 555 1901 589
rect 1843 549 1901 555
rect 2035 589 2093 595
rect 2035 555 2047 589
rect 2081 555 2093 589
rect 2035 549 2093 555
rect 2227 589 2285 595
rect 2227 555 2239 589
rect 2273 555 2285 589
rect 2227 549 2285 555
rect 2419 589 2477 595
rect 2419 555 2431 589
rect 2465 555 2477 589
rect 2419 549 2477 555
rect 2611 589 2669 595
rect 2611 555 2623 589
rect 2657 555 2669 589
rect 2611 549 2669 555
rect 2803 589 2861 595
rect 2803 555 2815 589
rect 2849 555 2861 589
rect 2803 549 2861 555
rect 2995 589 3053 595
rect 2995 555 3007 589
rect 3041 555 3053 589
rect 2995 549 3053 555
rect 3187 589 3245 595
rect 3187 555 3199 589
rect 3233 555 3245 589
rect 3187 549 3245 555
rect 3379 589 3437 595
rect 3379 555 3391 589
rect 3425 555 3437 589
rect 3379 549 3437 555
rect 3571 589 3629 595
rect 3571 555 3583 589
rect 3617 555 3629 589
rect 3571 549 3629 555
rect 3763 589 3821 595
rect 3763 555 3775 589
rect 3809 555 3821 589
rect 3763 549 3821 555
rect 3955 589 4013 595
rect 3955 555 3967 589
rect 4001 555 4013 589
rect 3955 549 4013 555
rect 4147 589 4205 595
rect 4147 555 4159 589
rect 4193 555 4205 589
rect 4147 549 4205 555
rect 4339 589 4397 595
rect 4339 555 4351 589
rect 4385 555 4397 589
rect 4339 549 4397 555
rect 4531 589 4589 595
rect 4531 555 4543 589
rect 4577 555 4589 589
rect 4531 549 4589 555
rect 4723 589 4781 595
rect 4723 555 4735 589
rect 4769 555 4781 589
rect 4723 549 4781 555
rect -4685 481 -4627 487
rect -4685 447 -4673 481
rect -4639 447 -4627 481
rect -4685 441 -4627 447
rect -4493 481 -4435 487
rect -4493 447 -4481 481
rect -4447 447 -4435 481
rect -4493 441 -4435 447
rect -4301 481 -4243 487
rect -4301 447 -4289 481
rect -4255 447 -4243 481
rect -4301 441 -4243 447
rect -4109 481 -4051 487
rect -4109 447 -4097 481
rect -4063 447 -4051 481
rect -4109 441 -4051 447
rect -3917 481 -3859 487
rect -3917 447 -3905 481
rect -3871 447 -3859 481
rect -3917 441 -3859 447
rect -3725 481 -3667 487
rect -3725 447 -3713 481
rect -3679 447 -3667 481
rect -3725 441 -3667 447
rect -3533 481 -3475 487
rect -3533 447 -3521 481
rect -3487 447 -3475 481
rect -3533 441 -3475 447
rect -3341 481 -3283 487
rect -3341 447 -3329 481
rect -3295 447 -3283 481
rect -3341 441 -3283 447
rect -3149 481 -3091 487
rect -3149 447 -3137 481
rect -3103 447 -3091 481
rect -3149 441 -3091 447
rect -2957 481 -2899 487
rect -2957 447 -2945 481
rect -2911 447 -2899 481
rect -2957 441 -2899 447
rect -2765 481 -2707 487
rect -2765 447 -2753 481
rect -2719 447 -2707 481
rect -2765 441 -2707 447
rect -2573 481 -2515 487
rect -2573 447 -2561 481
rect -2527 447 -2515 481
rect -2573 441 -2515 447
rect -2381 481 -2323 487
rect -2381 447 -2369 481
rect -2335 447 -2323 481
rect -2381 441 -2323 447
rect -2189 481 -2131 487
rect -2189 447 -2177 481
rect -2143 447 -2131 481
rect -2189 441 -2131 447
rect -1997 481 -1939 487
rect -1997 447 -1985 481
rect -1951 447 -1939 481
rect -1997 441 -1939 447
rect -1805 481 -1747 487
rect -1805 447 -1793 481
rect -1759 447 -1747 481
rect -1805 441 -1747 447
rect -1613 481 -1555 487
rect -1613 447 -1601 481
rect -1567 447 -1555 481
rect -1613 441 -1555 447
rect -1421 481 -1363 487
rect -1421 447 -1409 481
rect -1375 447 -1363 481
rect -1421 441 -1363 447
rect -1229 481 -1171 487
rect -1229 447 -1217 481
rect -1183 447 -1171 481
rect -1229 441 -1171 447
rect -1037 481 -979 487
rect -1037 447 -1025 481
rect -991 447 -979 481
rect -1037 441 -979 447
rect -845 481 -787 487
rect -845 447 -833 481
rect -799 447 -787 481
rect -845 441 -787 447
rect -653 481 -595 487
rect -653 447 -641 481
rect -607 447 -595 481
rect -653 441 -595 447
rect -461 481 -403 487
rect -461 447 -449 481
rect -415 447 -403 481
rect -461 441 -403 447
rect -269 481 -211 487
rect -269 447 -257 481
rect -223 447 -211 481
rect -269 441 -211 447
rect -77 481 -19 487
rect -77 447 -65 481
rect -31 447 -19 481
rect -77 441 -19 447
rect 115 481 173 487
rect 115 447 127 481
rect 161 447 173 481
rect 115 441 173 447
rect 307 481 365 487
rect 307 447 319 481
rect 353 447 365 481
rect 307 441 365 447
rect 499 481 557 487
rect 499 447 511 481
rect 545 447 557 481
rect 499 441 557 447
rect 691 481 749 487
rect 691 447 703 481
rect 737 447 749 481
rect 691 441 749 447
rect 883 481 941 487
rect 883 447 895 481
rect 929 447 941 481
rect 883 441 941 447
rect 1075 481 1133 487
rect 1075 447 1087 481
rect 1121 447 1133 481
rect 1075 441 1133 447
rect 1267 481 1325 487
rect 1267 447 1279 481
rect 1313 447 1325 481
rect 1267 441 1325 447
rect 1459 481 1517 487
rect 1459 447 1471 481
rect 1505 447 1517 481
rect 1459 441 1517 447
rect 1651 481 1709 487
rect 1651 447 1663 481
rect 1697 447 1709 481
rect 1651 441 1709 447
rect 1843 481 1901 487
rect 1843 447 1855 481
rect 1889 447 1901 481
rect 1843 441 1901 447
rect 2035 481 2093 487
rect 2035 447 2047 481
rect 2081 447 2093 481
rect 2035 441 2093 447
rect 2227 481 2285 487
rect 2227 447 2239 481
rect 2273 447 2285 481
rect 2227 441 2285 447
rect 2419 481 2477 487
rect 2419 447 2431 481
rect 2465 447 2477 481
rect 2419 441 2477 447
rect 2611 481 2669 487
rect 2611 447 2623 481
rect 2657 447 2669 481
rect 2611 441 2669 447
rect 2803 481 2861 487
rect 2803 447 2815 481
rect 2849 447 2861 481
rect 2803 441 2861 447
rect 2995 481 3053 487
rect 2995 447 3007 481
rect 3041 447 3053 481
rect 2995 441 3053 447
rect 3187 481 3245 487
rect 3187 447 3199 481
rect 3233 447 3245 481
rect 3187 441 3245 447
rect 3379 481 3437 487
rect 3379 447 3391 481
rect 3425 447 3437 481
rect 3379 441 3437 447
rect 3571 481 3629 487
rect 3571 447 3583 481
rect 3617 447 3629 481
rect 3571 441 3629 447
rect 3763 481 3821 487
rect 3763 447 3775 481
rect 3809 447 3821 481
rect 3763 441 3821 447
rect 3955 481 4013 487
rect 3955 447 3967 481
rect 4001 447 4013 481
rect 3955 441 4013 447
rect 4147 481 4205 487
rect 4147 447 4159 481
rect 4193 447 4205 481
rect 4147 441 4205 447
rect 4339 481 4397 487
rect 4339 447 4351 481
rect 4385 447 4397 481
rect 4339 441 4397 447
rect 4531 481 4589 487
rect 4531 447 4543 481
rect 4577 447 4589 481
rect 4531 441 4589 447
rect 4723 481 4781 487
rect 4723 447 4735 481
rect 4769 447 4781 481
rect 4723 441 4781 447
rect -4823 397 -4777 409
rect -4823 121 -4817 397
rect -4783 121 -4777 397
rect -4823 109 -4777 121
rect -4727 397 -4681 409
rect -4727 121 -4721 397
rect -4687 121 -4681 397
rect -4727 109 -4681 121
rect -4631 397 -4585 409
rect -4631 121 -4625 397
rect -4591 121 -4585 397
rect -4631 109 -4585 121
rect -4535 397 -4489 409
rect -4535 121 -4529 397
rect -4495 121 -4489 397
rect -4535 109 -4489 121
rect -4439 397 -4393 409
rect -4439 121 -4433 397
rect -4399 121 -4393 397
rect -4439 109 -4393 121
rect -4343 397 -4297 409
rect -4343 121 -4337 397
rect -4303 121 -4297 397
rect -4343 109 -4297 121
rect -4247 397 -4201 409
rect -4247 121 -4241 397
rect -4207 121 -4201 397
rect -4247 109 -4201 121
rect -4151 397 -4105 409
rect -4151 121 -4145 397
rect -4111 121 -4105 397
rect -4151 109 -4105 121
rect -4055 397 -4009 409
rect -4055 121 -4049 397
rect -4015 121 -4009 397
rect -4055 109 -4009 121
rect -3959 397 -3913 409
rect -3959 121 -3953 397
rect -3919 121 -3913 397
rect -3959 109 -3913 121
rect -3863 397 -3817 409
rect -3863 121 -3857 397
rect -3823 121 -3817 397
rect -3863 109 -3817 121
rect -3767 397 -3721 409
rect -3767 121 -3761 397
rect -3727 121 -3721 397
rect -3767 109 -3721 121
rect -3671 397 -3625 409
rect -3671 121 -3665 397
rect -3631 121 -3625 397
rect -3671 109 -3625 121
rect -3575 397 -3529 409
rect -3575 121 -3569 397
rect -3535 121 -3529 397
rect -3575 109 -3529 121
rect -3479 397 -3433 409
rect -3479 121 -3473 397
rect -3439 121 -3433 397
rect -3479 109 -3433 121
rect -3383 397 -3337 409
rect -3383 121 -3377 397
rect -3343 121 -3337 397
rect -3383 109 -3337 121
rect -3287 397 -3241 409
rect -3287 121 -3281 397
rect -3247 121 -3241 397
rect -3287 109 -3241 121
rect -3191 397 -3145 409
rect -3191 121 -3185 397
rect -3151 121 -3145 397
rect -3191 109 -3145 121
rect -3095 397 -3049 409
rect -3095 121 -3089 397
rect -3055 121 -3049 397
rect -3095 109 -3049 121
rect -2999 397 -2953 409
rect -2999 121 -2993 397
rect -2959 121 -2953 397
rect -2999 109 -2953 121
rect -2903 397 -2857 409
rect -2903 121 -2897 397
rect -2863 121 -2857 397
rect -2903 109 -2857 121
rect -2807 397 -2761 409
rect -2807 121 -2801 397
rect -2767 121 -2761 397
rect -2807 109 -2761 121
rect -2711 397 -2665 409
rect -2711 121 -2705 397
rect -2671 121 -2665 397
rect -2711 109 -2665 121
rect -2615 397 -2569 409
rect -2615 121 -2609 397
rect -2575 121 -2569 397
rect -2615 109 -2569 121
rect -2519 397 -2473 409
rect -2519 121 -2513 397
rect -2479 121 -2473 397
rect -2519 109 -2473 121
rect -2423 397 -2377 409
rect -2423 121 -2417 397
rect -2383 121 -2377 397
rect -2423 109 -2377 121
rect -2327 397 -2281 409
rect -2327 121 -2321 397
rect -2287 121 -2281 397
rect -2327 109 -2281 121
rect -2231 397 -2185 409
rect -2231 121 -2225 397
rect -2191 121 -2185 397
rect -2231 109 -2185 121
rect -2135 397 -2089 409
rect -2135 121 -2129 397
rect -2095 121 -2089 397
rect -2135 109 -2089 121
rect -2039 397 -1993 409
rect -2039 121 -2033 397
rect -1999 121 -1993 397
rect -2039 109 -1993 121
rect -1943 397 -1897 409
rect -1943 121 -1937 397
rect -1903 121 -1897 397
rect -1943 109 -1897 121
rect -1847 397 -1801 409
rect -1847 121 -1841 397
rect -1807 121 -1801 397
rect -1847 109 -1801 121
rect -1751 397 -1705 409
rect -1751 121 -1745 397
rect -1711 121 -1705 397
rect -1751 109 -1705 121
rect -1655 397 -1609 409
rect -1655 121 -1649 397
rect -1615 121 -1609 397
rect -1655 109 -1609 121
rect -1559 397 -1513 409
rect -1559 121 -1553 397
rect -1519 121 -1513 397
rect -1559 109 -1513 121
rect -1463 397 -1417 409
rect -1463 121 -1457 397
rect -1423 121 -1417 397
rect -1463 109 -1417 121
rect -1367 397 -1321 409
rect -1367 121 -1361 397
rect -1327 121 -1321 397
rect -1367 109 -1321 121
rect -1271 397 -1225 409
rect -1271 121 -1265 397
rect -1231 121 -1225 397
rect -1271 109 -1225 121
rect -1175 397 -1129 409
rect -1175 121 -1169 397
rect -1135 121 -1129 397
rect -1175 109 -1129 121
rect -1079 397 -1033 409
rect -1079 121 -1073 397
rect -1039 121 -1033 397
rect -1079 109 -1033 121
rect -983 397 -937 409
rect -983 121 -977 397
rect -943 121 -937 397
rect -983 109 -937 121
rect -887 397 -841 409
rect -887 121 -881 397
rect -847 121 -841 397
rect -887 109 -841 121
rect -791 397 -745 409
rect -791 121 -785 397
rect -751 121 -745 397
rect -791 109 -745 121
rect -695 397 -649 409
rect -695 121 -689 397
rect -655 121 -649 397
rect -695 109 -649 121
rect -599 397 -553 409
rect -599 121 -593 397
rect -559 121 -553 397
rect -599 109 -553 121
rect -503 397 -457 409
rect -503 121 -497 397
rect -463 121 -457 397
rect -503 109 -457 121
rect -407 397 -361 409
rect -407 121 -401 397
rect -367 121 -361 397
rect -407 109 -361 121
rect -311 397 -265 409
rect -311 121 -305 397
rect -271 121 -265 397
rect -311 109 -265 121
rect -215 397 -169 409
rect -215 121 -209 397
rect -175 121 -169 397
rect -215 109 -169 121
rect -119 397 -73 409
rect -119 121 -113 397
rect -79 121 -73 397
rect -119 109 -73 121
rect -23 397 23 409
rect -23 121 -17 397
rect 17 121 23 397
rect -23 109 23 121
rect 73 397 119 409
rect 73 121 79 397
rect 113 121 119 397
rect 73 109 119 121
rect 169 397 215 409
rect 169 121 175 397
rect 209 121 215 397
rect 169 109 215 121
rect 265 397 311 409
rect 265 121 271 397
rect 305 121 311 397
rect 265 109 311 121
rect 361 397 407 409
rect 361 121 367 397
rect 401 121 407 397
rect 361 109 407 121
rect 457 397 503 409
rect 457 121 463 397
rect 497 121 503 397
rect 457 109 503 121
rect 553 397 599 409
rect 553 121 559 397
rect 593 121 599 397
rect 553 109 599 121
rect 649 397 695 409
rect 649 121 655 397
rect 689 121 695 397
rect 649 109 695 121
rect 745 397 791 409
rect 745 121 751 397
rect 785 121 791 397
rect 745 109 791 121
rect 841 397 887 409
rect 841 121 847 397
rect 881 121 887 397
rect 841 109 887 121
rect 937 397 983 409
rect 937 121 943 397
rect 977 121 983 397
rect 937 109 983 121
rect 1033 397 1079 409
rect 1033 121 1039 397
rect 1073 121 1079 397
rect 1033 109 1079 121
rect 1129 397 1175 409
rect 1129 121 1135 397
rect 1169 121 1175 397
rect 1129 109 1175 121
rect 1225 397 1271 409
rect 1225 121 1231 397
rect 1265 121 1271 397
rect 1225 109 1271 121
rect 1321 397 1367 409
rect 1321 121 1327 397
rect 1361 121 1367 397
rect 1321 109 1367 121
rect 1417 397 1463 409
rect 1417 121 1423 397
rect 1457 121 1463 397
rect 1417 109 1463 121
rect 1513 397 1559 409
rect 1513 121 1519 397
rect 1553 121 1559 397
rect 1513 109 1559 121
rect 1609 397 1655 409
rect 1609 121 1615 397
rect 1649 121 1655 397
rect 1609 109 1655 121
rect 1705 397 1751 409
rect 1705 121 1711 397
rect 1745 121 1751 397
rect 1705 109 1751 121
rect 1801 397 1847 409
rect 1801 121 1807 397
rect 1841 121 1847 397
rect 1801 109 1847 121
rect 1897 397 1943 409
rect 1897 121 1903 397
rect 1937 121 1943 397
rect 1897 109 1943 121
rect 1993 397 2039 409
rect 1993 121 1999 397
rect 2033 121 2039 397
rect 1993 109 2039 121
rect 2089 397 2135 409
rect 2089 121 2095 397
rect 2129 121 2135 397
rect 2089 109 2135 121
rect 2185 397 2231 409
rect 2185 121 2191 397
rect 2225 121 2231 397
rect 2185 109 2231 121
rect 2281 397 2327 409
rect 2281 121 2287 397
rect 2321 121 2327 397
rect 2281 109 2327 121
rect 2377 397 2423 409
rect 2377 121 2383 397
rect 2417 121 2423 397
rect 2377 109 2423 121
rect 2473 397 2519 409
rect 2473 121 2479 397
rect 2513 121 2519 397
rect 2473 109 2519 121
rect 2569 397 2615 409
rect 2569 121 2575 397
rect 2609 121 2615 397
rect 2569 109 2615 121
rect 2665 397 2711 409
rect 2665 121 2671 397
rect 2705 121 2711 397
rect 2665 109 2711 121
rect 2761 397 2807 409
rect 2761 121 2767 397
rect 2801 121 2807 397
rect 2761 109 2807 121
rect 2857 397 2903 409
rect 2857 121 2863 397
rect 2897 121 2903 397
rect 2857 109 2903 121
rect 2953 397 2999 409
rect 2953 121 2959 397
rect 2993 121 2999 397
rect 2953 109 2999 121
rect 3049 397 3095 409
rect 3049 121 3055 397
rect 3089 121 3095 397
rect 3049 109 3095 121
rect 3145 397 3191 409
rect 3145 121 3151 397
rect 3185 121 3191 397
rect 3145 109 3191 121
rect 3241 397 3287 409
rect 3241 121 3247 397
rect 3281 121 3287 397
rect 3241 109 3287 121
rect 3337 397 3383 409
rect 3337 121 3343 397
rect 3377 121 3383 397
rect 3337 109 3383 121
rect 3433 397 3479 409
rect 3433 121 3439 397
rect 3473 121 3479 397
rect 3433 109 3479 121
rect 3529 397 3575 409
rect 3529 121 3535 397
rect 3569 121 3575 397
rect 3529 109 3575 121
rect 3625 397 3671 409
rect 3625 121 3631 397
rect 3665 121 3671 397
rect 3625 109 3671 121
rect 3721 397 3767 409
rect 3721 121 3727 397
rect 3761 121 3767 397
rect 3721 109 3767 121
rect 3817 397 3863 409
rect 3817 121 3823 397
rect 3857 121 3863 397
rect 3817 109 3863 121
rect 3913 397 3959 409
rect 3913 121 3919 397
rect 3953 121 3959 397
rect 3913 109 3959 121
rect 4009 397 4055 409
rect 4009 121 4015 397
rect 4049 121 4055 397
rect 4009 109 4055 121
rect 4105 397 4151 409
rect 4105 121 4111 397
rect 4145 121 4151 397
rect 4105 109 4151 121
rect 4201 397 4247 409
rect 4201 121 4207 397
rect 4241 121 4247 397
rect 4201 109 4247 121
rect 4297 397 4343 409
rect 4297 121 4303 397
rect 4337 121 4343 397
rect 4297 109 4343 121
rect 4393 397 4439 409
rect 4393 121 4399 397
rect 4433 121 4439 397
rect 4393 109 4439 121
rect 4489 397 4535 409
rect 4489 121 4495 397
rect 4529 121 4535 397
rect 4489 109 4535 121
rect 4585 397 4631 409
rect 4585 121 4591 397
rect 4625 121 4631 397
rect 4585 109 4631 121
rect 4681 397 4727 409
rect 4681 121 4687 397
rect 4721 121 4727 397
rect 4681 109 4727 121
rect 4777 397 4823 409
rect 4777 121 4783 397
rect 4817 121 4823 397
rect 4777 109 4823 121
rect -4781 71 -4723 77
rect -4781 37 -4769 71
rect -4735 37 -4723 71
rect -4781 31 -4723 37
rect -4589 71 -4531 77
rect -4589 37 -4577 71
rect -4543 37 -4531 71
rect -4589 31 -4531 37
rect -4397 71 -4339 77
rect -4397 37 -4385 71
rect -4351 37 -4339 71
rect -4397 31 -4339 37
rect -4205 71 -4147 77
rect -4205 37 -4193 71
rect -4159 37 -4147 71
rect -4205 31 -4147 37
rect -4013 71 -3955 77
rect -4013 37 -4001 71
rect -3967 37 -3955 71
rect -4013 31 -3955 37
rect -3821 71 -3763 77
rect -3821 37 -3809 71
rect -3775 37 -3763 71
rect -3821 31 -3763 37
rect -3629 71 -3571 77
rect -3629 37 -3617 71
rect -3583 37 -3571 71
rect -3629 31 -3571 37
rect -3437 71 -3379 77
rect -3437 37 -3425 71
rect -3391 37 -3379 71
rect -3437 31 -3379 37
rect -3245 71 -3187 77
rect -3245 37 -3233 71
rect -3199 37 -3187 71
rect -3245 31 -3187 37
rect -3053 71 -2995 77
rect -3053 37 -3041 71
rect -3007 37 -2995 71
rect -3053 31 -2995 37
rect -2861 71 -2803 77
rect -2861 37 -2849 71
rect -2815 37 -2803 71
rect -2861 31 -2803 37
rect -2669 71 -2611 77
rect -2669 37 -2657 71
rect -2623 37 -2611 71
rect -2669 31 -2611 37
rect -2477 71 -2419 77
rect -2477 37 -2465 71
rect -2431 37 -2419 71
rect -2477 31 -2419 37
rect -2285 71 -2227 77
rect -2285 37 -2273 71
rect -2239 37 -2227 71
rect -2285 31 -2227 37
rect -2093 71 -2035 77
rect -2093 37 -2081 71
rect -2047 37 -2035 71
rect -2093 31 -2035 37
rect -1901 71 -1843 77
rect -1901 37 -1889 71
rect -1855 37 -1843 71
rect -1901 31 -1843 37
rect -1709 71 -1651 77
rect -1709 37 -1697 71
rect -1663 37 -1651 71
rect -1709 31 -1651 37
rect -1517 71 -1459 77
rect -1517 37 -1505 71
rect -1471 37 -1459 71
rect -1517 31 -1459 37
rect -1325 71 -1267 77
rect -1325 37 -1313 71
rect -1279 37 -1267 71
rect -1325 31 -1267 37
rect -1133 71 -1075 77
rect -1133 37 -1121 71
rect -1087 37 -1075 71
rect -1133 31 -1075 37
rect -941 71 -883 77
rect -941 37 -929 71
rect -895 37 -883 71
rect -941 31 -883 37
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect 979 71 1037 77
rect 979 37 991 71
rect 1025 37 1037 71
rect 979 31 1037 37
rect 1171 71 1229 77
rect 1171 37 1183 71
rect 1217 37 1229 71
rect 1171 31 1229 37
rect 1363 71 1421 77
rect 1363 37 1375 71
rect 1409 37 1421 71
rect 1363 31 1421 37
rect 1555 71 1613 77
rect 1555 37 1567 71
rect 1601 37 1613 71
rect 1555 31 1613 37
rect 1747 71 1805 77
rect 1747 37 1759 71
rect 1793 37 1805 71
rect 1747 31 1805 37
rect 1939 71 1997 77
rect 1939 37 1951 71
rect 1985 37 1997 71
rect 1939 31 1997 37
rect 2131 71 2189 77
rect 2131 37 2143 71
rect 2177 37 2189 71
rect 2131 31 2189 37
rect 2323 71 2381 77
rect 2323 37 2335 71
rect 2369 37 2381 71
rect 2323 31 2381 37
rect 2515 71 2573 77
rect 2515 37 2527 71
rect 2561 37 2573 71
rect 2515 31 2573 37
rect 2707 71 2765 77
rect 2707 37 2719 71
rect 2753 37 2765 71
rect 2707 31 2765 37
rect 2899 71 2957 77
rect 2899 37 2911 71
rect 2945 37 2957 71
rect 2899 31 2957 37
rect 3091 71 3149 77
rect 3091 37 3103 71
rect 3137 37 3149 71
rect 3091 31 3149 37
rect 3283 71 3341 77
rect 3283 37 3295 71
rect 3329 37 3341 71
rect 3283 31 3341 37
rect 3475 71 3533 77
rect 3475 37 3487 71
rect 3521 37 3533 71
rect 3475 31 3533 37
rect 3667 71 3725 77
rect 3667 37 3679 71
rect 3713 37 3725 71
rect 3667 31 3725 37
rect 3859 71 3917 77
rect 3859 37 3871 71
rect 3905 37 3917 71
rect 3859 31 3917 37
rect 4051 71 4109 77
rect 4051 37 4063 71
rect 4097 37 4109 71
rect 4051 31 4109 37
rect 4243 71 4301 77
rect 4243 37 4255 71
rect 4289 37 4301 71
rect 4243 31 4301 37
rect 4435 71 4493 77
rect 4435 37 4447 71
rect 4481 37 4493 71
rect 4435 31 4493 37
rect 4627 71 4685 77
rect 4627 37 4639 71
rect 4673 37 4685 71
rect 4627 31 4685 37
rect -4781 -37 -4723 -31
rect -4781 -71 -4769 -37
rect -4735 -71 -4723 -37
rect -4781 -77 -4723 -71
rect -4589 -37 -4531 -31
rect -4589 -71 -4577 -37
rect -4543 -71 -4531 -37
rect -4589 -77 -4531 -71
rect -4397 -37 -4339 -31
rect -4397 -71 -4385 -37
rect -4351 -71 -4339 -37
rect -4397 -77 -4339 -71
rect -4205 -37 -4147 -31
rect -4205 -71 -4193 -37
rect -4159 -71 -4147 -37
rect -4205 -77 -4147 -71
rect -4013 -37 -3955 -31
rect -4013 -71 -4001 -37
rect -3967 -71 -3955 -37
rect -4013 -77 -3955 -71
rect -3821 -37 -3763 -31
rect -3821 -71 -3809 -37
rect -3775 -71 -3763 -37
rect -3821 -77 -3763 -71
rect -3629 -37 -3571 -31
rect -3629 -71 -3617 -37
rect -3583 -71 -3571 -37
rect -3629 -77 -3571 -71
rect -3437 -37 -3379 -31
rect -3437 -71 -3425 -37
rect -3391 -71 -3379 -37
rect -3437 -77 -3379 -71
rect -3245 -37 -3187 -31
rect -3245 -71 -3233 -37
rect -3199 -71 -3187 -37
rect -3245 -77 -3187 -71
rect -3053 -37 -2995 -31
rect -3053 -71 -3041 -37
rect -3007 -71 -2995 -37
rect -3053 -77 -2995 -71
rect -2861 -37 -2803 -31
rect -2861 -71 -2849 -37
rect -2815 -71 -2803 -37
rect -2861 -77 -2803 -71
rect -2669 -37 -2611 -31
rect -2669 -71 -2657 -37
rect -2623 -71 -2611 -37
rect -2669 -77 -2611 -71
rect -2477 -37 -2419 -31
rect -2477 -71 -2465 -37
rect -2431 -71 -2419 -37
rect -2477 -77 -2419 -71
rect -2285 -37 -2227 -31
rect -2285 -71 -2273 -37
rect -2239 -71 -2227 -37
rect -2285 -77 -2227 -71
rect -2093 -37 -2035 -31
rect -2093 -71 -2081 -37
rect -2047 -71 -2035 -37
rect -2093 -77 -2035 -71
rect -1901 -37 -1843 -31
rect -1901 -71 -1889 -37
rect -1855 -71 -1843 -37
rect -1901 -77 -1843 -71
rect -1709 -37 -1651 -31
rect -1709 -71 -1697 -37
rect -1663 -71 -1651 -37
rect -1709 -77 -1651 -71
rect -1517 -37 -1459 -31
rect -1517 -71 -1505 -37
rect -1471 -71 -1459 -37
rect -1517 -77 -1459 -71
rect -1325 -37 -1267 -31
rect -1325 -71 -1313 -37
rect -1279 -71 -1267 -37
rect -1325 -77 -1267 -71
rect -1133 -37 -1075 -31
rect -1133 -71 -1121 -37
rect -1087 -71 -1075 -37
rect -1133 -77 -1075 -71
rect -941 -37 -883 -31
rect -941 -71 -929 -37
rect -895 -71 -883 -37
rect -941 -77 -883 -71
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect 979 -37 1037 -31
rect 979 -71 991 -37
rect 1025 -71 1037 -37
rect 979 -77 1037 -71
rect 1171 -37 1229 -31
rect 1171 -71 1183 -37
rect 1217 -71 1229 -37
rect 1171 -77 1229 -71
rect 1363 -37 1421 -31
rect 1363 -71 1375 -37
rect 1409 -71 1421 -37
rect 1363 -77 1421 -71
rect 1555 -37 1613 -31
rect 1555 -71 1567 -37
rect 1601 -71 1613 -37
rect 1555 -77 1613 -71
rect 1747 -37 1805 -31
rect 1747 -71 1759 -37
rect 1793 -71 1805 -37
rect 1747 -77 1805 -71
rect 1939 -37 1997 -31
rect 1939 -71 1951 -37
rect 1985 -71 1997 -37
rect 1939 -77 1997 -71
rect 2131 -37 2189 -31
rect 2131 -71 2143 -37
rect 2177 -71 2189 -37
rect 2131 -77 2189 -71
rect 2323 -37 2381 -31
rect 2323 -71 2335 -37
rect 2369 -71 2381 -37
rect 2323 -77 2381 -71
rect 2515 -37 2573 -31
rect 2515 -71 2527 -37
rect 2561 -71 2573 -37
rect 2515 -77 2573 -71
rect 2707 -37 2765 -31
rect 2707 -71 2719 -37
rect 2753 -71 2765 -37
rect 2707 -77 2765 -71
rect 2899 -37 2957 -31
rect 2899 -71 2911 -37
rect 2945 -71 2957 -37
rect 2899 -77 2957 -71
rect 3091 -37 3149 -31
rect 3091 -71 3103 -37
rect 3137 -71 3149 -37
rect 3091 -77 3149 -71
rect 3283 -37 3341 -31
rect 3283 -71 3295 -37
rect 3329 -71 3341 -37
rect 3283 -77 3341 -71
rect 3475 -37 3533 -31
rect 3475 -71 3487 -37
rect 3521 -71 3533 -37
rect 3475 -77 3533 -71
rect 3667 -37 3725 -31
rect 3667 -71 3679 -37
rect 3713 -71 3725 -37
rect 3667 -77 3725 -71
rect 3859 -37 3917 -31
rect 3859 -71 3871 -37
rect 3905 -71 3917 -37
rect 3859 -77 3917 -71
rect 4051 -37 4109 -31
rect 4051 -71 4063 -37
rect 4097 -71 4109 -37
rect 4051 -77 4109 -71
rect 4243 -37 4301 -31
rect 4243 -71 4255 -37
rect 4289 -71 4301 -37
rect 4243 -77 4301 -71
rect 4435 -37 4493 -31
rect 4435 -71 4447 -37
rect 4481 -71 4493 -37
rect 4435 -77 4493 -71
rect 4627 -37 4685 -31
rect 4627 -71 4639 -37
rect 4673 -71 4685 -37
rect 4627 -77 4685 -71
rect -4823 -121 -4777 -109
rect -4823 -397 -4817 -121
rect -4783 -397 -4777 -121
rect -4823 -409 -4777 -397
rect -4727 -121 -4681 -109
rect -4727 -397 -4721 -121
rect -4687 -397 -4681 -121
rect -4727 -409 -4681 -397
rect -4631 -121 -4585 -109
rect -4631 -397 -4625 -121
rect -4591 -397 -4585 -121
rect -4631 -409 -4585 -397
rect -4535 -121 -4489 -109
rect -4535 -397 -4529 -121
rect -4495 -397 -4489 -121
rect -4535 -409 -4489 -397
rect -4439 -121 -4393 -109
rect -4439 -397 -4433 -121
rect -4399 -397 -4393 -121
rect -4439 -409 -4393 -397
rect -4343 -121 -4297 -109
rect -4343 -397 -4337 -121
rect -4303 -397 -4297 -121
rect -4343 -409 -4297 -397
rect -4247 -121 -4201 -109
rect -4247 -397 -4241 -121
rect -4207 -397 -4201 -121
rect -4247 -409 -4201 -397
rect -4151 -121 -4105 -109
rect -4151 -397 -4145 -121
rect -4111 -397 -4105 -121
rect -4151 -409 -4105 -397
rect -4055 -121 -4009 -109
rect -4055 -397 -4049 -121
rect -4015 -397 -4009 -121
rect -4055 -409 -4009 -397
rect -3959 -121 -3913 -109
rect -3959 -397 -3953 -121
rect -3919 -397 -3913 -121
rect -3959 -409 -3913 -397
rect -3863 -121 -3817 -109
rect -3863 -397 -3857 -121
rect -3823 -397 -3817 -121
rect -3863 -409 -3817 -397
rect -3767 -121 -3721 -109
rect -3767 -397 -3761 -121
rect -3727 -397 -3721 -121
rect -3767 -409 -3721 -397
rect -3671 -121 -3625 -109
rect -3671 -397 -3665 -121
rect -3631 -397 -3625 -121
rect -3671 -409 -3625 -397
rect -3575 -121 -3529 -109
rect -3575 -397 -3569 -121
rect -3535 -397 -3529 -121
rect -3575 -409 -3529 -397
rect -3479 -121 -3433 -109
rect -3479 -397 -3473 -121
rect -3439 -397 -3433 -121
rect -3479 -409 -3433 -397
rect -3383 -121 -3337 -109
rect -3383 -397 -3377 -121
rect -3343 -397 -3337 -121
rect -3383 -409 -3337 -397
rect -3287 -121 -3241 -109
rect -3287 -397 -3281 -121
rect -3247 -397 -3241 -121
rect -3287 -409 -3241 -397
rect -3191 -121 -3145 -109
rect -3191 -397 -3185 -121
rect -3151 -397 -3145 -121
rect -3191 -409 -3145 -397
rect -3095 -121 -3049 -109
rect -3095 -397 -3089 -121
rect -3055 -397 -3049 -121
rect -3095 -409 -3049 -397
rect -2999 -121 -2953 -109
rect -2999 -397 -2993 -121
rect -2959 -397 -2953 -121
rect -2999 -409 -2953 -397
rect -2903 -121 -2857 -109
rect -2903 -397 -2897 -121
rect -2863 -397 -2857 -121
rect -2903 -409 -2857 -397
rect -2807 -121 -2761 -109
rect -2807 -397 -2801 -121
rect -2767 -397 -2761 -121
rect -2807 -409 -2761 -397
rect -2711 -121 -2665 -109
rect -2711 -397 -2705 -121
rect -2671 -397 -2665 -121
rect -2711 -409 -2665 -397
rect -2615 -121 -2569 -109
rect -2615 -397 -2609 -121
rect -2575 -397 -2569 -121
rect -2615 -409 -2569 -397
rect -2519 -121 -2473 -109
rect -2519 -397 -2513 -121
rect -2479 -397 -2473 -121
rect -2519 -409 -2473 -397
rect -2423 -121 -2377 -109
rect -2423 -397 -2417 -121
rect -2383 -397 -2377 -121
rect -2423 -409 -2377 -397
rect -2327 -121 -2281 -109
rect -2327 -397 -2321 -121
rect -2287 -397 -2281 -121
rect -2327 -409 -2281 -397
rect -2231 -121 -2185 -109
rect -2231 -397 -2225 -121
rect -2191 -397 -2185 -121
rect -2231 -409 -2185 -397
rect -2135 -121 -2089 -109
rect -2135 -397 -2129 -121
rect -2095 -397 -2089 -121
rect -2135 -409 -2089 -397
rect -2039 -121 -1993 -109
rect -2039 -397 -2033 -121
rect -1999 -397 -1993 -121
rect -2039 -409 -1993 -397
rect -1943 -121 -1897 -109
rect -1943 -397 -1937 -121
rect -1903 -397 -1897 -121
rect -1943 -409 -1897 -397
rect -1847 -121 -1801 -109
rect -1847 -397 -1841 -121
rect -1807 -397 -1801 -121
rect -1847 -409 -1801 -397
rect -1751 -121 -1705 -109
rect -1751 -397 -1745 -121
rect -1711 -397 -1705 -121
rect -1751 -409 -1705 -397
rect -1655 -121 -1609 -109
rect -1655 -397 -1649 -121
rect -1615 -397 -1609 -121
rect -1655 -409 -1609 -397
rect -1559 -121 -1513 -109
rect -1559 -397 -1553 -121
rect -1519 -397 -1513 -121
rect -1559 -409 -1513 -397
rect -1463 -121 -1417 -109
rect -1463 -397 -1457 -121
rect -1423 -397 -1417 -121
rect -1463 -409 -1417 -397
rect -1367 -121 -1321 -109
rect -1367 -397 -1361 -121
rect -1327 -397 -1321 -121
rect -1367 -409 -1321 -397
rect -1271 -121 -1225 -109
rect -1271 -397 -1265 -121
rect -1231 -397 -1225 -121
rect -1271 -409 -1225 -397
rect -1175 -121 -1129 -109
rect -1175 -397 -1169 -121
rect -1135 -397 -1129 -121
rect -1175 -409 -1129 -397
rect -1079 -121 -1033 -109
rect -1079 -397 -1073 -121
rect -1039 -397 -1033 -121
rect -1079 -409 -1033 -397
rect -983 -121 -937 -109
rect -983 -397 -977 -121
rect -943 -397 -937 -121
rect -983 -409 -937 -397
rect -887 -121 -841 -109
rect -887 -397 -881 -121
rect -847 -397 -841 -121
rect -887 -409 -841 -397
rect -791 -121 -745 -109
rect -791 -397 -785 -121
rect -751 -397 -745 -121
rect -791 -409 -745 -397
rect -695 -121 -649 -109
rect -695 -397 -689 -121
rect -655 -397 -649 -121
rect -695 -409 -649 -397
rect -599 -121 -553 -109
rect -599 -397 -593 -121
rect -559 -397 -553 -121
rect -599 -409 -553 -397
rect -503 -121 -457 -109
rect -503 -397 -497 -121
rect -463 -397 -457 -121
rect -503 -409 -457 -397
rect -407 -121 -361 -109
rect -407 -397 -401 -121
rect -367 -397 -361 -121
rect -407 -409 -361 -397
rect -311 -121 -265 -109
rect -311 -397 -305 -121
rect -271 -397 -265 -121
rect -311 -409 -265 -397
rect -215 -121 -169 -109
rect -215 -397 -209 -121
rect -175 -397 -169 -121
rect -215 -409 -169 -397
rect -119 -121 -73 -109
rect -119 -397 -113 -121
rect -79 -397 -73 -121
rect -119 -409 -73 -397
rect -23 -121 23 -109
rect -23 -397 -17 -121
rect 17 -397 23 -121
rect -23 -409 23 -397
rect 73 -121 119 -109
rect 73 -397 79 -121
rect 113 -397 119 -121
rect 73 -409 119 -397
rect 169 -121 215 -109
rect 169 -397 175 -121
rect 209 -397 215 -121
rect 169 -409 215 -397
rect 265 -121 311 -109
rect 265 -397 271 -121
rect 305 -397 311 -121
rect 265 -409 311 -397
rect 361 -121 407 -109
rect 361 -397 367 -121
rect 401 -397 407 -121
rect 361 -409 407 -397
rect 457 -121 503 -109
rect 457 -397 463 -121
rect 497 -397 503 -121
rect 457 -409 503 -397
rect 553 -121 599 -109
rect 553 -397 559 -121
rect 593 -397 599 -121
rect 553 -409 599 -397
rect 649 -121 695 -109
rect 649 -397 655 -121
rect 689 -397 695 -121
rect 649 -409 695 -397
rect 745 -121 791 -109
rect 745 -397 751 -121
rect 785 -397 791 -121
rect 745 -409 791 -397
rect 841 -121 887 -109
rect 841 -397 847 -121
rect 881 -397 887 -121
rect 841 -409 887 -397
rect 937 -121 983 -109
rect 937 -397 943 -121
rect 977 -397 983 -121
rect 937 -409 983 -397
rect 1033 -121 1079 -109
rect 1033 -397 1039 -121
rect 1073 -397 1079 -121
rect 1033 -409 1079 -397
rect 1129 -121 1175 -109
rect 1129 -397 1135 -121
rect 1169 -397 1175 -121
rect 1129 -409 1175 -397
rect 1225 -121 1271 -109
rect 1225 -397 1231 -121
rect 1265 -397 1271 -121
rect 1225 -409 1271 -397
rect 1321 -121 1367 -109
rect 1321 -397 1327 -121
rect 1361 -397 1367 -121
rect 1321 -409 1367 -397
rect 1417 -121 1463 -109
rect 1417 -397 1423 -121
rect 1457 -397 1463 -121
rect 1417 -409 1463 -397
rect 1513 -121 1559 -109
rect 1513 -397 1519 -121
rect 1553 -397 1559 -121
rect 1513 -409 1559 -397
rect 1609 -121 1655 -109
rect 1609 -397 1615 -121
rect 1649 -397 1655 -121
rect 1609 -409 1655 -397
rect 1705 -121 1751 -109
rect 1705 -397 1711 -121
rect 1745 -397 1751 -121
rect 1705 -409 1751 -397
rect 1801 -121 1847 -109
rect 1801 -397 1807 -121
rect 1841 -397 1847 -121
rect 1801 -409 1847 -397
rect 1897 -121 1943 -109
rect 1897 -397 1903 -121
rect 1937 -397 1943 -121
rect 1897 -409 1943 -397
rect 1993 -121 2039 -109
rect 1993 -397 1999 -121
rect 2033 -397 2039 -121
rect 1993 -409 2039 -397
rect 2089 -121 2135 -109
rect 2089 -397 2095 -121
rect 2129 -397 2135 -121
rect 2089 -409 2135 -397
rect 2185 -121 2231 -109
rect 2185 -397 2191 -121
rect 2225 -397 2231 -121
rect 2185 -409 2231 -397
rect 2281 -121 2327 -109
rect 2281 -397 2287 -121
rect 2321 -397 2327 -121
rect 2281 -409 2327 -397
rect 2377 -121 2423 -109
rect 2377 -397 2383 -121
rect 2417 -397 2423 -121
rect 2377 -409 2423 -397
rect 2473 -121 2519 -109
rect 2473 -397 2479 -121
rect 2513 -397 2519 -121
rect 2473 -409 2519 -397
rect 2569 -121 2615 -109
rect 2569 -397 2575 -121
rect 2609 -397 2615 -121
rect 2569 -409 2615 -397
rect 2665 -121 2711 -109
rect 2665 -397 2671 -121
rect 2705 -397 2711 -121
rect 2665 -409 2711 -397
rect 2761 -121 2807 -109
rect 2761 -397 2767 -121
rect 2801 -397 2807 -121
rect 2761 -409 2807 -397
rect 2857 -121 2903 -109
rect 2857 -397 2863 -121
rect 2897 -397 2903 -121
rect 2857 -409 2903 -397
rect 2953 -121 2999 -109
rect 2953 -397 2959 -121
rect 2993 -397 2999 -121
rect 2953 -409 2999 -397
rect 3049 -121 3095 -109
rect 3049 -397 3055 -121
rect 3089 -397 3095 -121
rect 3049 -409 3095 -397
rect 3145 -121 3191 -109
rect 3145 -397 3151 -121
rect 3185 -397 3191 -121
rect 3145 -409 3191 -397
rect 3241 -121 3287 -109
rect 3241 -397 3247 -121
rect 3281 -397 3287 -121
rect 3241 -409 3287 -397
rect 3337 -121 3383 -109
rect 3337 -397 3343 -121
rect 3377 -397 3383 -121
rect 3337 -409 3383 -397
rect 3433 -121 3479 -109
rect 3433 -397 3439 -121
rect 3473 -397 3479 -121
rect 3433 -409 3479 -397
rect 3529 -121 3575 -109
rect 3529 -397 3535 -121
rect 3569 -397 3575 -121
rect 3529 -409 3575 -397
rect 3625 -121 3671 -109
rect 3625 -397 3631 -121
rect 3665 -397 3671 -121
rect 3625 -409 3671 -397
rect 3721 -121 3767 -109
rect 3721 -397 3727 -121
rect 3761 -397 3767 -121
rect 3721 -409 3767 -397
rect 3817 -121 3863 -109
rect 3817 -397 3823 -121
rect 3857 -397 3863 -121
rect 3817 -409 3863 -397
rect 3913 -121 3959 -109
rect 3913 -397 3919 -121
rect 3953 -397 3959 -121
rect 3913 -409 3959 -397
rect 4009 -121 4055 -109
rect 4009 -397 4015 -121
rect 4049 -397 4055 -121
rect 4009 -409 4055 -397
rect 4105 -121 4151 -109
rect 4105 -397 4111 -121
rect 4145 -397 4151 -121
rect 4105 -409 4151 -397
rect 4201 -121 4247 -109
rect 4201 -397 4207 -121
rect 4241 -397 4247 -121
rect 4201 -409 4247 -397
rect 4297 -121 4343 -109
rect 4297 -397 4303 -121
rect 4337 -397 4343 -121
rect 4297 -409 4343 -397
rect 4393 -121 4439 -109
rect 4393 -397 4399 -121
rect 4433 -397 4439 -121
rect 4393 -409 4439 -397
rect 4489 -121 4535 -109
rect 4489 -397 4495 -121
rect 4529 -397 4535 -121
rect 4489 -409 4535 -397
rect 4585 -121 4631 -109
rect 4585 -397 4591 -121
rect 4625 -397 4631 -121
rect 4585 -409 4631 -397
rect 4681 -121 4727 -109
rect 4681 -397 4687 -121
rect 4721 -397 4727 -121
rect 4681 -409 4727 -397
rect 4777 -121 4823 -109
rect 4777 -397 4783 -121
rect 4817 -397 4823 -121
rect 4777 -409 4823 -397
rect -4685 -447 -4627 -441
rect -4685 -481 -4673 -447
rect -4639 -481 -4627 -447
rect -4685 -487 -4627 -481
rect -4493 -447 -4435 -441
rect -4493 -481 -4481 -447
rect -4447 -481 -4435 -447
rect -4493 -487 -4435 -481
rect -4301 -447 -4243 -441
rect -4301 -481 -4289 -447
rect -4255 -481 -4243 -447
rect -4301 -487 -4243 -481
rect -4109 -447 -4051 -441
rect -4109 -481 -4097 -447
rect -4063 -481 -4051 -447
rect -4109 -487 -4051 -481
rect -3917 -447 -3859 -441
rect -3917 -481 -3905 -447
rect -3871 -481 -3859 -447
rect -3917 -487 -3859 -481
rect -3725 -447 -3667 -441
rect -3725 -481 -3713 -447
rect -3679 -481 -3667 -447
rect -3725 -487 -3667 -481
rect -3533 -447 -3475 -441
rect -3533 -481 -3521 -447
rect -3487 -481 -3475 -447
rect -3533 -487 -3475 -481
rect -3341 -447 -3283 -441
rect -3341 -481 -3329 -447
rect -3295 -481 -3283 -447
rect -3341 -487 -3283 -481
rect -3149 -447 -3091 -441
rect -3149 -481 -3137 -447
rect -3103 -481 -3091 -447
rect -3149 -487 -3091 -481
rect -2957 -447 -2899 -441
rect -2957 -481 -2945 -447
rect -2911 -481 -2899 -447
rect -2957 -487 -2899 -481
rect -2765 -447 -2707 -441
rect -2765 -481 -2753 -447
rect -2719 -481 -2707 -447
rect -2765 -487 -2707 -481
rect -2573 -447 -2515 -441
rect -2573 -481 -2561 -447
rect -2527 -481 -2515 -447
rect -2573 -487 -2515 -481
rect -2381 -447 -2323 -441
rect -2381 -481 -2369 -447
rect -2335 -481 -2323 -447
rect -2381 -487 -2323 -481
rect -2189 -447 -2131 -441
rect -2189 -481 -2177 -447
rect -2143 -481 -2131 -447
rect -2189 -487 -2131 -481
rect -1997 -447 -1939 -441
rect -1997 -481 -1985 -447
rect -1951 -481 -1939 -447
rect -1997 -487 -1939 -481
rect -1805 -447 -1747 -441
rect -1805 -481 -1793 -447
rect -1759 -481 -1747 -447
rect -1805 -487 -1747 -481
rect -1613 -447 -1555 -441
rect -1613 -481 -1601 -447
rect -1567 -481 -1555 -447
rect -1613 -487 -1555 -481
rect -1421 -447 -1363 -441
rect -1421 -481 -1409 -447
rect -1375 -481 -1363 -447
rect -1421 -487 -1363 -481
rect -1229 -447 -1171 -441
rect -1229 -481 -1217 -447
rect -1183 -481 -1171 -447
rect -1229 -487 -1171 -481
rect -1037 -447 -979 -441
rect -1037 -481 -1025 -447
rect -991 -481 -979 -447
rect -1037 -487 -979 -481
rect -845 -447 -787 -441
rect -845 -481 -833 -447
rect -799 -481 -787 -447
rect -845 -487 -787 -481
rect -653 -447 -595 -441
rect -653 -481 -641 -447
rect -607 -481 -595 -447
rect -653 -487 -595 -481
rect -461 -447 -403 -441
rect -461 -481 -449 -447
rect -415 -481 -403 -447
rect -461 -487 -403 -481
rect -269 -447 -211 -441
rect -269 -481 -257 -447
rect -223 -481 -211 -447
rect -269 -487 -211 -481
rect -77 -447 -19 -441
rect -77 -481 -65 -447
rect -31 -481 -19 -447
rect -77 -487 -19 -481
rect 115 -447 173 -441
rect 115 -481 127 -447
rect 161 -481 173 -447
rect 115 -487 173 -481
rect 307 -447 365 -441
rect 307 -481 319 -447
rect 353 -481 365 -447
rect 307 -487 365 -481
rect 499 -447 557 -441
rect 499 -481 511 -447
rect 545 -481 557 -447
rect 499 -487 557 -481
rect 691 -447 749 -441
rect 691 -481 703 -447
rect 737 -481 749 -447
rect 691 -487 749 -481
rect 883 -447 941 -441
rect 883 -481 895 -447
rect 929 -481 941 -447
rect 883 -487 941 -481
rect 1075 -447 1133 -441
rect 1075 -481 1087 -447
rect 1121 -481 1133 -447
rect 1075 -487 1133 -481
rect 1267 -447 1325 -441
rect 1267 -481 1279 -447
rect 1313 -481 1325 -447
rect 1267 -487 1325 -481
rect 1459 -447 1517 -441
rect 1459 -481 1471 -447
rect 1505 -481 1517 -447
rect 1459 -487 1517 -481
rect 1651 -447 1709 -441
rect 1651 -481 1663 -447
rect 1697 -481 1709 -447
rect 1651 -487 1709 -481
rect 1843 -447 1901 -441
rect 1843 -481 1855 -447
rect 1889 -481 1901 -447
rect 1843 -487 1901 -481
rect 2035 -447 2093 -441
rect 2035 -481 2047 -447
rect 2081 -481 2093 -447
rect 2035 -487 2093 -481
rect 2227 -447 2285 -441
rect 2227 -481 2239 -447
rect 2273 -481 2285 -447
rect 2227 -487 2285 -481
rect 2419 -447 2477 -441
rect 2419 -481 2431 -447
rect 2465 -481 2477 -447
rect 2419 -487 2477 -481
rect 2611 -447 2669 -441
rect 2611 -481 2623 -447
rect 2657 -481 2669 -447
rect 2611 -487 2669 -481
rect 2803 -447 2861 -441
rect 2803 -481 2815 -447
rect 2849 -481 2861 -447
rect 2803 -487 2861 -481
rect 2995 -447 3053 -441
rect 2995 -481 3007 -447
rect 3041 -481 3053 -447
rect 2995 -487 3053 -481
rect 3187 -447 3245 -441
rect 3187 -481 3199 -447
rect 3233 -481 3245 -447
rect 3187 -487 3245 -481
rect 3379 -447 3437 -441
rect 3379 -481 3391 -447
rect 3425 -481 3437 -447
rect 3379 -487 3437 -481
rect 3571 -447 3629 -441
rect 3571 -481 3583 -447
rect 3617 -481 3629 -447
rect 3571 -487 3629 -481
rect 3763 -447 3821 -441
rect 3763 -481 3775 -447
rect 3809 -481 3821 -447
rect 3763 -487 3821 -481
rect 3955 -447 4013 -441
rect 3955 -481 3967 -447
rect 4001 -481 4013 -447
rect 3955 -487 4013 -481
rect 4147 -447 4205 -441
rect 4147 -481 4159 -447
rect 4193 -481 4205 -447
rect 4147 -487 4205 -481
rect 4339 -447 4397 -441
rect 4339 -481 4351 -447
rect 4385 -481 4397 -447
rect 4339 -487 4397 -481
rect 4531 -447 4589 -441
rect 4531 -481 4543 -447
rect 4577 -481 4589 -447
rect 4531 -487 4589 -481
rect 4723 -447 4781 -441
rect 4723 -481 4735 -447
rect 4769 -481 4781 -447
rect 4723 -487 4781 -481
rect -4685 -555 -4627 -549
rect -4685 -589 -4673 -555
rect -4639 -589 -4627 -555
rect -4685 -595 -4627 -589
rect -4493 -555 -4435 -549
rect -4493 -589 -4481 -555
rect -4447 -589 -4435 -555
rect -4493 -595 -4435 -589
rect -4301 -555 -4243 -549
rect -4301 -589 -4289 -555
rect -4255 -589 -4243 -555
rect -4301 -595 -4243 -589
rect -4109 -555 -4051 -549
rect -4109 -589 -4097 -555
rect -4063 -589 -4051 -555
rect -4109 -595 -4051 -589
rect -3917 -555 -3859 -549
rect -3917 -589 -3905 -555
rect -3871 -589 -3859 -555
rect -3917 -595 -3859 -589
rect -3725 -555 -3667 -549
rect -3725 -589 -3713 -555
rect -3679 -589 -3667 -555
rect -3725 -595 -3667 -589
rect -3533 -555 -3475 -549
rect -3533 -589 -3521 -555
rect -3487 -589 -3475 -555
rect -3533 -595 -3475 -589
rect -3341 -555 -3283 -549
rect -3341 -589 -3329 -555
rect -3295 -589 -3283 -555
rect -3341 -595 -3283 -589
rect -3149 -555 -3091 -549
rect -3149 -589 -3137 -555
rect -3103 -589 -3091 -555
rect -3149 -595 -3091 -589
rect -2957 -555 -2899 -549
rect -2957 -589 -2945 -555
rect -2911 -589 -2899 -555
rect -2957 -595 -2899 -589
rect -2765 -555 -2707 -549
rect -2765 -589 -2753 -555
rect -2719 -589 -2707 -555
rect -2765 -595 -2707 -589
rect -2573 -555 -2515 -549
rect -2573 -589 -2561 -555
rect -2527 -589 -2515 -555
rect -2573 -595 -2515 -589
rect -2381 -555 -2323 -549
rect -2381 -589 -2369 -555
rect -2335 -589 -2323 -555
rect -2381 -595 -2323 -589
rect -2189 -555 -2131 -549
rect -2189 -589 -2177 -555
rect -2143 -589 -2131 -555
rect -2189 -595 -2131 -589
rect -1997 -555 -1939 -549
rect -1997 -589 -1985 -555
rect -1951 -589 -1939 -555
rect -1997 -595 -1939 -589
rect -1805 -555 -1747 -549
rect -1805 -589 -1793 -555
rect -1759 -589 -1747 -555
rect -1805 -595 -1747 -589
rect -1613 -555 -1555 -549
rect -1613 -589 -1601 -555
rect -1567 -589 -1555 -555
rect -1613 -595 -1555 -589
rect -1421 -555 -1363 -549
rect -1421 -589 -1409 -555
rect -1375 -589 -1363 -555
rect -1421 -595 -1363 -589
rect -1229 -555 -1171 -549
rect -1229 -589 -1217 -555
rect -1183 -589 -1171 -555
rect -1229 -595 -1171 -589
rect -1037 -555 -979 -549
rect -1037 -589 -1025 -555
rect -991 -589 -979 -555
rect -1037 -595 -979 -589
rect -845 -555 -787 -549
rect -845 -589 -833 -555
rect -799 -589 -787 -555
rect -845 -595 -787 -589
rect -653 -555 -595 -549
rect -653 -589 -641 -555
rect -607 -589 -595 -555
rect -653 -595 -595 -589
rect -461 -555 -403 -549
rect -461 -589 -449 -555
rect -415 -589 -403 -555
rect -461 -595 -403 -589
rect -269 -555 -211 -549
rect -269 -589 -257 -555
rect -223 -589 -211 -555
rect -269 -595 -211 -589
rect -77 -555 -19 -549
rect -77 -589 -65 -555
rect -31 -589 -19 -555
rect -77 -595 -19 -589
rect 115 -555 173 -549
rect 115 -589 127 -555
rect 161 -589 173 -555
rect 115 -595 173 -589
rect 307 -555 365 -549
rect 307 -589 319 -555
rect 353 -589 365 -555
rect 307 -595 365 -589
rect 499 -555 557 -549
rect 499 -589 511 -555
rect 545 -589 557 -555
rect 499 -595 557 -589
rect 691 -555 749 -549
rect 691 -589 703 -555
rect 737 -589 749 -555
rect 691 -595 749 -589
rect 883 -555 941 -549
rect 883 -589 895 -555
rect 929 -589 941 -555
rect 883 -595 941 -589
rect 1075 -555 1133 -549
rect 1075 -589 1087 -555
rect 1121 -589 1133 -555
rect 1075 -595 1133 -589
rect 1267 -555 1325 -549
rect 1267 -589 1279 -555
rect 1313 -589 1325 -555
rect 1267 -595 1325 -589
rect 1459 -555 1517 -549
rect 1459 -589 1471 -555
rect 1505 -589 1517 -555
rect 1459 -595 1517 -589
rect 1651 -555 1709 -549
rect 1651 -589 1663 -555
rect 1697 -589 1709 -555
rect 1651 -595 1709 -589
rect 1843 -555 1901 -549
rect 1843 -589 1855 -555
rect 1889 -589 1901 -555
rect 1843 -595 1901 -589
rect 2035 -555 2093 -549
rect 2035 -589 2047 -555
rect 2081 -589 2093 -555
rect 2035 -595 2093 -589
rect 2227 -555 2285 -549
rect 2227 -589 2239 -555
rect 2273 -589 2285 -555
rect 2227 -595 2285 -589
rect 2419 -555 2477 -549
rect 2419 -589 2431 -555
rect 2465 -589 2477 -555
rect 2419 -595 2477 -589
rect 2611 -555 2669 -549
rect 2611 -589 2623 -555
rect 2657 -589 2669 -555
rect 2611 -595 2669 -589
rect 2803 -555 2861 -549
rect 2803 -589 2815 -555
rect 2849 -589 2861 -555
rect 2803 -595 2861 -589
rect 2995 -555 3053 -549
rect 2995 -589 3007 -555
rect 3041 -589 3053 -555
rect 2995 -595 3053 -589
rect 3187 -555 3245 -549
rect 3187 -589 3199 -555
rect 3233 -589 3245 -555
rect 3187 -595 3245 -589
rect 3379 -555 3437 -549
rect 3379 -589 3391 -555
rect 3425 -589 3437 -555
rect 3379 -595 3437 -589
rect 3571 -555 3629 -549
rect 3571 -589 3583 -555
rect 3617 -589 3629 -555
rect 3571 -595 3629 -589
rect 3763 -555 3821 -549
rect 3763 -589 3775 -555
rect 3809 -589 3821 -555
rect 3763 -595 3821 -589
rect 3955 -555 4013 -549
rect 3955 -589 3967 -555
rect 4001 -589 4013 -555
rect 3955 -595 4013 -589
rect 4147 -555 4205 -549
rect 4147 -589 4159 -555
rect 4193 -589 4205 -555
rect 4147 -595 4205 -589
rect 4339 -555 4397 -549
rect 4339 -589 4351 -555
rect 4385 -589 4397 -555
rect 4339 -595 4397 -589
rect 4531 -555 4589 -549
rect 4531 -589 4543 -555
rect 4577 -589 4589 -555
rect 4531 -595 4589 -589
rect 4723 -555 4781 -549
rect 4723 -589 4735 -555
rect 4769 -589 4781 -555
rect 4723 -595 4781 -589
rect -4823 -639 -4777 -627
rect -4823 -915 -4817 -639
rect -4783 -915 -4777 -639
rect -4823 -927 -4777 -915
rect -4727 -639 -4681 -627
rect -4727 -915 -4721 -639
rect -4687 -915 -4681 -639
rect -4727 -927 -4681 -915
rect -4631 -639 -4585 -627
rect -4631 -915 -4625 -639
rect -4591 -915 -4585 -639
rect -4631 -927 -4585 -915
rect -4535 -639 -4489 -627
rect -4535 -915 -4529 -639
rect -4495 -915 -4489 -639
rect -4535 -927 -4489 -915
rect -4439 -639 -4393 -627
rect -4439 -915 -4433 -639
rect -4399 -915 -4393 -639
rect -4439 -927 -4393 -915
rect -4343 -639 -4297 -627
rect -4343 -915 -4337 -639
rect -4303 -915 -4297 -639
rect -4343 -927 -4297 -915
rect -4247 -639 -4201 -627
rect -4247 -915 -4241 -639
rect -4207 -915 -4201 -639
rect -4247 -927 -4201 -915
rect -4151 -639 -4105 -627
rect -4151 -915 -4145 -639
rect -4111 -915 -4105 -639
rect -4151 -927 -4105 -915
rect -4055 -639 -4009 -627
rect -4055 -915 -4049 -639
rect -4015 -915 -4009 -639
rect -4055 -927 -4009 -915
rect -3959 -639 -3913 -627
rect -3959 -915 -3953 -639
rect -3919 -915 -3913 -639
rect -3959 -927 -3913 -915
rect -3863 -639 -3817 -627
rect -3863 -915 -3857 -639
rect -3823 -915 -3817 -639
rect -3863 -927 -3817 -915
rect -3767 -639 -3721 -627
rect -3767 -915 -3761 -639
rect -3727 -915 -3721 -639
rect -3767 -927 -3721 -915
rect -3671 -639 -3625 -627
rect -3671 -915 -3665 -639
rect -3631 -915 -3625 -639
rect -3671 -927 -3625 -915
rect -3575 -639 -3529 -627
rect -3575 -915 -3569 -639
rect -3535 -915 -3529 -639
rect -3575 -927 -3529 -915
rect -3479 -639 -3433 -627
rect -3479 -915 -3473 -639
rect -3439 -915 -3433 -639
rect -3479 -927 -3433 -915
rect -3383 -639 -3337 -627
rect -3383 -915 -3377 -639
rect -3343 -915 -3337 -639
rect -3383 -927 -3337 -915
rect -3287 -639 -3241 -627
rect -3287 -915 -3281 -639
rect -3247 -915 -3241 -639
rect -3287 -927 -3241 -915
rect -3191 -639 -3145 -627
rect -3191 -915 -3185 -639
rect -3151 -915 -3145 -639
rect -3191 -927 -3145 -915
rect -3095 -639 -3049 -627
rect -3095 -915 -3089 -639
rect -3055 -915 -3049 -639
rect -3095 -927 -3049 -915
rect -2999 -639 -2953 -627
rect -2999 -915 -2993 -639
rect -2959 -915 -2953 -639
rect -2999 -927 -2953 -915
rect -2903 -639 -2857 -627
rect -2903 -915 -2897 -639
rect -2863 -915 -2857 -639
rect -2903 -927 -2857 -915
rect -2807 -639 -2761 -627
rect -2807 -915 -2801 -639
rect -2767 -915 -2761 -639
rect -2807 -927 -2761 -915
rect -2711 -639 -2665 -627
rect -2711 -915 -2705 -639
rect -2671 -915 -2665 -639
rect -2711 -927 -2665 -915
rect -2615 -639 -2569 -627
rect -2615 -915 -2609 -639
rect -2575 -915 -2569 -639
rect -2615 -927 -2569 -915
rect -2519 -639 -2473 -627
rect -2519 -915 -2513 -639
rect -2479 -915 -2473 -639
rect -2519 -927 -2473 -915
rect -2423 -639 -2377 -627
rect -2423 -915 -2417 -639
rect -2383 -915 -2377 -639
rect -2423 -927 -2377 -915
rect -2327 -639 -2281 -627
rect -2327 -915 -2321 -639
rect -2287 -915 -2281 -639
rect -2327 -927 -2281 -915
rect -2231 -639 -2185 -627
rect -2231 -915 -2225 -639
rect -2191 -915 -2185 -639
rect -2231 -927 -2185 -915
rect -2135 -639 -2089 -627
rect -2135 -915 -2129 -639
rect -2095 -915 -2089 -639
rect -2135 -927 -2089 -915
rect -2039 -639 -1993 -627
rect -2039 -915 -2033 -639
rect -1999 -915 -1993 -639
rect -2039 -927 -1993 -915
rect -1943 -639 -1897 -627
rect -1943 -915 -1937 -639
rect -1903 -915 -1897 -639
rect -1943 -927 -1897 -915
rect -1847 -639 -1801 -627
rect -1847 -915 -1841 -639
rect -1807 -915 -1801 -639
rect -1847 -927 -1801 -915
rect -1751 -639 -1705 -627
rect -1751 -915 -1745 -639
rect -1711 -915 -1705 -639
rect -1751 -927 -1705 -915
rect -1655 -639 -1609 -627
rect -1655 -915 -1649 -639
rect -1615 -915 -1609 -639
rect -1655 -927 -1609 -915
rect -1559 -639 -1513 -627
rect -1559 -915 -1553 -639
rect -1519 -915 -1513 -639
rect -1559 -927 -1513 -915
rect -1463 -639 -1417 -627
rect -1463 -915 -1457 -639
rect -1423 -915 -1417 -639
rect -1463 -927 -1417 -915
rect -1367 -639 -1321 -627
rect -1367 -915 -1361 -639
rect -1327 -915 -1321 -639
rect -1367 -927 -1321 -915
rect -1271 -639 -1225 -627
rect -1271 -915 -1265 -639
rect -1231 -915 -1225 -639
rect -1271 -927 -1225 -915
rect -1175 -639 -1129 -627
rect -1175 -915 -1169 -639
rect -1135 -915 -1129 -639
rect -1175 -927 -1129 -915
rect -1079 -639 -1033 -627
rect -1079 -915 -1073 -639
rect -1039 -915 -1033 -639
rect -1079 -927 -1033 -915
rect -983 -639 -937 -627
rect -983 -915 -977 -639
rect -943 -915 -937 -639
rect -983 -927 -937 -915
rect -887 -639 -841 -627
rect -887 -915 -881 -639
rect -847 -915 -841 -639
rect -887 -927 -841 -915
rect -791 -639 -745 -627
rect -791 -915 -785 -639
rect -751 -915 -745 -639
rect -791 -927 -745 -915
rect -695 -639 -649 -627
rect -695 -915 -689 -639
rect -655 -915 -649 -639
rect -695 -927 -649 -915
rect -599 -639 -553 -627
rect -599 -915 -593 -639
rect -559 -915 -553 -639
rect -599 -927 -553 -915
rect -503 -639 -457 -627
rect -503 -915 -497 -639
rect -463 -915 -457 -639
rect -503 -927 -457 -915
rect -407 -639 -361 -627
rect -407 -915 -401 -639
rect -367 -915 -361 -639
rect -407 -927 -361 -915
rect -311 -639 -265 -627
rect -311 -915 -305 -639
rect -271 -915 -265 -639
rect -311 -927 -265 -915
rect -215 -639 -169 -627
rect -215 -915 -209 -639
rect -175 -915 -169 -639
rect -215 -927 -169 -915
rect -119 -639 -73 -627
rect -119 -915 -113 -639
rect -79 -915 -73 -639
rect -119 -927 -73 -915
rect -23 -639 23 -627
rect -23 -915 -17 -639
rect 17 -915 23 -639
rect -23 -927 23 -915
rect 73 -639 119 -627
rect 73 -915 79 -639
rect 113 -915 119 -639
rect 73 -927 119 -915
rect 169 -639 215 -627
rect 169 -915 175 -639
rect 209 -915 215 -639
rect 169 -927 215 -915
rect 265 -639 311 -627
rect 265 -915 271 -639
rect 305 -915 311 -639
rect 265 -927 311 -915
rect 361 -639 407 -627
rect 361 -915 367 -639
rect 401 -915 407 -639
rect 361 -927 407 -915
rect 457 -639 503 -627
rect 457 -915 463 -639
rect 497 -915 503 -639
rect 457 -927 503 -915
rect 553 -639 599 -627
rect 553 -915 559 -639
rect 593 -915 599 -639
rect 553 -927 599 -915
rect 649 -639 695 -627
rect 649 -915 655 -639
rect 689 -915 695 -639
rect 649 -927 695 -915
rect 745 -639 791 -627
rect 745 -915 751 -639
rect 785 -915 791 -639
rect 745 -927 791 -915
rect 841 -639 887 -627
rect 841 -915 847 -639
rect 881 -915 887 -639
rect 841 -927 887 -915
rect 937 -639 983 -627
rect 937 -915 943 -639
rect 977 -915 983 -639
rect 937 -927 983 -915
rect 1033 -639 1079 -627
rect 1033 -915 1039 -639
rect 1073 -915 1079 -639
rect 1033 -927 1079 -915
rect 1129 -639 1175 -627
rect 1129 -915 1135 -639
rect 1169 -915 1175 -639
rect 1129 -927 1175 -915
rect 1225 -639 1271 -627
rect 1225 -915 1231 -639
rect 1265 -915 1271 -639
rect 1225 -927 1271 -915
rect 1321 -639 1367 -627
rect 1321 -915 1327 -639
rect 1361 -915 1367 -639
rect 1321 -927 1367 -915
rect 1417 -639 1463 -627
rect 1417 -915 1423 -639
rect 1457 -915 1463 -639
rect 1417 -927 1463 -915
rect 1513 -639 1559 -627
rect 1513 -915 1519 -639
rect 1553 -915 1559 -639
rect 1513 -927 1559 -915
rect 1609 -639 1655 -627
rect 1609 -915 1615 -639
rect 1649 -915 1655 -639
rect 1609 -927 1655 -915
rect 1705 -639 1751 -627
rect 1705 -915 1711 -639
rect 1745 -915 1751 -639
rect 1705 -927 1751 -915
rect 1801 -639 1847 -627
rect 1801 -915 1807 -639
rect 1841 -915 1847 -639
rect 1801 -927 1847 -915
rect 1897 -639 1943 -627
rect 1897 -915 1903 -639
rect 1937 -915 1943 -639
rect 1897 -927 1943 -915
rect 1993 -639 2039 -627
rect 1993 -915 1999 -639
rect 2033 -915 2039 -639
rect 1993 -927 2039 -915
rect 2089 -639 2135 -627
rect 2089 -915 2095 -639
rect 2129 -915 2135 -639
rect 2089 -927 2135 -915
rect 2185 -639 2231 -627
rect 2185 -915 2191 -639
rect 2225 -915 2231 -639
rect 2185 -927 2231 -915
rect 2281 -639 2327 -627
rect 2281 -915 2287 -639
rect 2321 -915 2327 -639
rect 2281 -927 2327 -915
rect 2377 -639 2423 -627
rect 2377 -915 2383 -639
rect 2417 -915 2423 -639
rect 2377 -927 2423 -915
rect 2473 -639 2519 -627
rect 2473 -915 2479 -639
rect 2513 -915 2519 -639
rect 2473 -927 2519 -915
rect 2569 -639 2615 -627
rect 2569 -915 2575 -639
rect 2609 -915 2615 -639
rect 2569 -927 2615 -915
rect 2665 -639 2711 -627
rect 2665 -915 2671 -639
rect 2705 -915 2711 -639
rect 2665 -927 2711 -915
rect 2761 -639 2807 -627
rect 2761 -915 2767 -639
rect 2801 -915 2807 -639
rect 2761 -927 2807 -915
rect 2857 -639 2903 -627
rect 2857 -915 2863 -639
rect 2897 -915 2903 -639
rect 2857 -927 2903 -915
rect 2953 -639 2999 -627
rect 2953 -915 2959 -639
rect 2993 -915 2999 -639
rect 2953 -927 2999 -915
rect 3049 -639 3095 -627
rect 3049 -915 3055 -639
rect 3089 -915 3095 -639
rect 3049 -927 3095 -915
rect 3145 -639 3191 -627
rect 3145 -915 3151 -639
rect 3185 -915 3191 -639
rect 3145 -927 3191 -915
rect 3241 -639 3287 -627
rect 3241 -915 3247 -639
rect 3281 -915 3287 -639
rect 3241 -927 3287 -915
rect 3337 -639 3383 -627
rect 3337 -915 3343 -639
rect 3377 -915 3383 -639
rect 3337 -927 3383 -915
rect 3433 -639 3479 -627
rect 3433 -915 3439 -639
rect 3473 -915 3479 -639
rect 3433 -927 3479 -915
rect 3529 -639 3575 -627
rect 3529 -915 3535 -639
rect 3569 -915 3575 -639
rect 3529 -927 3575 -915
rect 3625 -639 3671 -627
rect 3625 -915 3631 -639
rect 3665 -915 3671 -639
rect 3625 -927 3671 -915
rect 3721 -639 3767 -627
rect 3721 -915 3727 -639
rect 3761 -915 3767 -639
rect 3721 -927 3767 -915
rect 3817 -639 3863 -627
rect 3817 -915 3823 -639
rect 3857 -915 3863 -639
rect 3817 -927 3863 -915
rect 3913 -639 3959 -627
rect 3913 -915 3919 -639
rect 3953 -915 3959 -639
rect 3913 -927 3959 -915
rect 4009 -639 4055 -627
rect 4009 -915 4015 -639
rect 4049 -915 4055 -639
rect 4009 -927 4055 -915
rect 4105 -639 4151 -627
rect 4105 -915 4111 -639
rect 4145 -915 4151 -639
rect 4105 -927 4151 -915
rect 4201 -639 4247 -627
rect 4201 -915 4207 -639
rect 4241 -915 4247 -639
rect 4201 -927 4247 -915
rect 4297 -639 4343 -627
rect 4297 -915 4303 -639
rect 4337 -915 4343 -639
rect 4297 -927 4343 -915
rect 4393 -639 4439 -627
rect 4393 -915 4399 -639
rect 4433 -915 4439 -639
rect 4393 -927 4439 -915
rect 4489 -639 4535 -627
rect 4489 -915 4495 -639
rect 4529 -915 4535 -639
rect 4489 -927 4535 -915
rect 4585 -639 4631 -627
rect 4585 -915 4591 -639
rect 4625 -915 4631 -639
rect 4585 -927 4631 -915
rect 4681 -639 4727 -627
rect 4681 -915 4687 -639
rect 4721 -915 4727 -639
rect 4681 -927 4727 -915
rect 4777 -639 4823 -627
rect 4777 -915 4783 -639
rect 4817 -915 4823 -639
rect 4777 -927 4823 -915
rect -4781 -965 -4723 -959
rect -4781 -999 -4769 -965
rect -4735 -999 -4723 -965
rect -4781 -1005 -4723 -999
rect -4589 -965 -4531 -959
rect -4589 -999 -4577 -965
rect -4543 -999 -4531 -965
rect -4589 -1005 -4531 -999
rect -4397 -965 -4339 -959
rect -4397 -999 -4385 -965
rect -4351 -999 -4339 -965
rect -4397 -1005 -4339 -999
rect -4205 -965 -4147 -959
rect -4205 -999 -4193 -965
rect -4159 -999 -4147 -965
rect -4205 -1005 -4147 -999
rect -4013 -965 -3955 -959
rect -4013 -999 -4001 -965
rect -3967 -999 -3955 -965
rect -4013 -1005 -3955 -999
rect -3821 -965 -3763 -959
rect -3821 -999 -3809 -965
rect -3775 -999 -3763 -965
rect -3821 -1005 -3763 -999
rect -3629 -965 -3571 -959
rect -3629 -999 -3617 -965
rect -3583 -999 -3571 -965
rect -3629 -1005 -3571 -999
rect -3437 -965 -3379 -959
rect -3437 -999 -3425 -965
rect -3391 -999 -3379 -965
rect -3437 -1005 -3379 -999
rect -3245 -965 -3187 -959
rect -3245 -999 -3233 -965
rect -3199 -999 -3187 -965
rect -3245 -1005 -3187 -999
rect -3053 -965 -2995 -959
rect -3053 -999 -3041 -965
rect -3007 -999 -2995 -965
rect -3053 -1005 -2995 -999
rect -2861 -965 -2803 -959
rect -2861 -999 -2849 -965
rect -2815 -999 -2803 -965
rect -2861 -1005 -2803 -999
rect -2669 -965 -2611 -959
rect -2669 -999 -2657 -965
rect -2623 -999 -2611 -965
rect -2669 -1005 -2611 -999
rect -2477 -965 -2419 -959
rect -2477 -999 -2465 -965
rect -2431 -999 -2419 -965
rect -2477 -1005 -2419 -999
rect -2285 -965 -2227 -959
rect -2285 -999 -2273 -965
rect -2239 -999 -2227 -965
rect -2285 -1005 -2227 -999
rect -2093 -965 -2035 -959
rect -2093 -999 -2081 -965
rect -2047 -999 -2035 -965
rect -2093 -1005 -2035 -999
rect -1901 -965 -1843 -959
rect -1901 -999 -1889 -965
rect -1855 -999 -1843 -965
rect -1901 -1005 -1843 -999
rect -1709 -965 -1651 -959
rect -1709 -999 -1697 -965
rect -1663 -999 -1651 -965
rect -1709 -1005 -1651 -999
rect -1517 -965 -1459 -959
rect -1517 -999 -1505 -965
rect -1471 -999 -1459 -965
rect -1517 -1005 -1459 -999
rect -1325 -965 -1267 -959
rect -1325 -999 -1313 -965
rect -1279 -999 -1267 -965
rect -1325 -1005 -1267 -999
rect -1133 -965 -1075 -959
rect -1133 -999 -1121 -965
rect -1087 -999 -1075 -965
rect -1133 -1005 -1075 -999
rect -941 -965 -883 -959
rect -941 -999 -929 -965
rect -895 -999 -883 -965
rect -941 -1005 -883 -999
rect -749 -965 -691 -959
rect -749 -999 -737 -965
rect -703 -999 -691 -965
rect -749 -1005 -691 -999
rect -557 -965 -499 -959
rect -557 -999 -545 -965
rect -511 -999 -499 -965
rect -557 -1005 -499 -999
rect -365 -965 -307 -959
rect -365 -999 -353 -965
rect -319 -999 -307 -965
rect -365 -1005 -307 -999
rect -173 -965 -115 -959
rect -173 -999 -161 -965
rect -127 -999 -115 -965
rect -173 -1005 -115 -999
rect 19 -965 77 -959
rect 19 -999 31 -965
rect 65 -999 77 -965
rect 19 -1005 77 -999
rect 211 -965 269 -959
rect 211 -999 223 -965
rect 257 -999 269 -965
rect 211 -1005 269 -999
rect 403 -965 461 -959
rect 403 -999 415 -965
rect 449 -999 461 -965
rect 403 -1005 461 -999
rect 595 -965 653 -959
rect 595 -999 607 -965
rect 641 -999 653 -965
rect 595 -1005 653 -999
rect 787 -965 845 -959
rect 787 -999 799 -965
rect 833 -999 845 -965
rect 787 -1005 845 -999
rect 979 -965 1037 -959
rect 979 -999 991 -965
rect 1025 -999 1037 -965
rect 979 -1005 1037 -999
rect 1171 -965 1229 -959
rect 1171 -999 1183 -965
rect 1217 -999 1229 -965
rect 1171 -1005 1229 -999
rect 1363 -965 1421 -959
rect 1363 -999 1375 -965
rect 1409 -999 1421 -965
rect 1363 -1005 1421 -999
rect 1555 -965 1613 -959
rect 1555 -999 1567 -965
rect 1601 -999 1613 -965
rect 1555 -1005 1613 -999
rect 1747 -965 1805 -959
rect 1747 -999 1759 -965
rect 1793 -999 1805 -965
rect 1747 -1005 1805 -999
rect 1939 -965 1997 -959
rect 1939 -999 1951 -965
rect 1985 -999 1997 -965
rect 1939 -1005 1997 -999
rect 2131 -965 2189 -959
rect 2131 -999 2143 -965
rect 2177 -999 2189 -965
rect 2131 -1005 2189 -999
rect 2323 -965 2381 -959
rect 2323 -999 2335 -965
rect 2369 -999 2381 -965
rect 2323 -1005 2381 -999
rect 2515 -965 2573 -959
rect 2515 -999 2527 -965
rect 2561 -999 2573 -965
rect 2515 -1005 2573 -999
rect 2707 -965 2765 -959
rect 2707 -999 2719 -965
rect 2753 -999 2765 -965
rect 2707 -1005 2765 -999
rect 2899 -965 2957 -959
rect 2899 -999 2911 -965
rect 2945 -999 2957 -965
rect 2899 -1005 2957 -999
rect 3091 -965 3149 -959
rect 3091 -999 3103 -965
rect 3137 -999 3149 -965
rect 3091 -1005 3149 -999
rect 3283 -965 3341 -959
rect 3283 -999 3295 -965
rect 3329 -999 3341 -965
rect 3283 -1005 3341 -999
rect 3475 -965 3533 -959
rect 3475 -999 3487 -965
rect 3521 -999 3533 -965
rect 3475 -1005 3533 -999
rect 3667 -965 3725 -959
rect 3667 -999 3679 -965
rect 3713 -999 3725 -965
rect 3667 -1005 3725 -999
rect 3859 -965 3917 -959
rect 3859 -999 3871 -965
rect 3905 -999 3917 -965
rect 3859 -1005 3917 -999
rect 4051 -965 4109 -959
rect 4051 -999 4063 -965
rect 4097 -999 4109 -965
rect 4051 -1005 4109 -999
rect 4243 -965 4301 -959
rect 4243 -999 4255 -965
rect 4289 -999 4301 -965
rect 4243 -1005 4301 -999
rect 4435 -965 4493 -959
rect 4435 -999 4447 -965
rect 4481 -999 4493 -965
rect 4435 -1005 4493 -999
rect 4627 -965 4685 -959
rect 4627 -999 4639 -965
rect 4673 -999 4685 -965
rect 4627 -1005 4685 -999
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -4914 -1084 4914 1084
string parameters w 1.5 l 0.15 m 4 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
