magic
tech sky130A
magscale 1 2
timestamp 1623959084
<< error_s >>
rect 9266 1136 9268 1158
rect 11726 569 11772 580
rect 1732 544 1751 546
rect 3393 493 3409 569
rect 3421 546 3446 548
rect 3421 520 3449 546
rect 5078 493 5096 569
rect 5106 545 5131 547
rect 5106 519 5134 545
rect 6762 493 6786 569
rect 6790 546 6815 548
rect 6790 520 6818 546
rect 8453 493 8474 568
rect 8481 540 8506 542
rect 8481 514 8509 540
rect 10140 493 10159 569
rect 11726 567 11744 569
rect 10168 542 10193 544
rect 10168 516 10196 542
rect 11727 510 11744 523
rect 9 141 21 168
rect -19 49 -7 77
rect 9 28 21 49
<< nwell >>
rect 10300 1147 10722 1823
rect 11303 1155 11816 1904
<< pwell >>
rect 10298 1904 10482 2452
rect 11528 1904 11816 2452
rect 10298 1877 10648 1904
rect 10318 1823 10648 1877
<< metal1 >>
rect 10332 2463 10476 2601
rect -54 2372 10476 2463
rect 11492 2452 11816 2601
rect -54 2280 -44 2372
rect 28 2326 10476 2372
rect 28 2280 38 2326
rect 9123 2320 10476 2326
rect -54 2186 4 2280
rect 10851 1913 10861 1976
rect 10949 1913 10959 1976
rect 11052 1794 11062 1877
rect 11150 1794 11160 1877
rect 547 1684 557 1756
rect 618 1684 628 1756
rect 1073 1684 1083 1756
rect 1144 1684 1154 1756
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 3495 1684 3505 1756
rect 3566 1684 3576 1756
rect 4021 1684 4031 1756
rect 4092 1684 4102 1756
rect 4969 1684 4979 1756
rect 5040 1684 5050 1756
rect 5495 1684 5505 1756
rect 5566 1684 5576 1756
rect 6443 1684 6453 1756
rect 6514 1684 6524 1756
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 7917 1684 7927 1756
rect 7988 1684 7998 1756
rect 8443 1684 8453 1756
rect 8514 1684 8524 1756
rect 9391 1684 9401 1756
rect 9462 1684 9472 1756
rect 9917 1684 9927 1756
rect 9988 1684 9998 1756
rect 328 1218 9266 1224
rect 0 1136 9266 1218
rect 10648 1136 11366 1190
rect 328 1130 9268 1136
rect -7 141 9 168
rect -7 49 3 141
rect 75 49 85 141
rect -7 28 9 49
<< via1 >>
rect -44 2280 28 2372
rect 10861 1913 10949 1976
rect 11062 1794 11150 1877
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
rect 3 49 75 141
<< metal2 >>
rect 62 2537 1547 2538
rect 62 2486 5975 2537
rect -44 2372 28 2382
rect -208 2280 -44 2365
rect -208 2278 28 2280
rect -208 124 -124 2278
rect -44 2270 28 2278
rect 15 1812 23 1838
rect 62 1826 114 2486
rect 1495 2485 5975 2486
rect 62 1812 79 1826
rect 1495 1811 1547 2485
rect 2972 2330 3043 2340
rect 2972 2246 3043 2256
rect 2981 1839 3033 2246
rect 2973 1813 3033 1839
rect 4451 1837 4503 2485
rect 2981 1812 3033 1813
rect 4436 1814 4503 1837
rect 5923 1817 5975 2485
rect 7396 2514 7467 2524
rect 7396 2420 7467 2430
rect 7404 1836 7456 2420
rect 4436 1811 4461 1814
rect 5923 1811 5948 1817
rect 7388 1813 7456 1836
rect 7388 1810 7413 1813
rect 8879 1810 8931 2443
rect 10861 1976 10949 1986
rect 10133 1970 10134 1973
rect 10087 1924 10861 1970
rect 10087 1804 10133 1924
rect 10861 1903 10949 1913
rect 11062 1877 11150 1887
rect 11062 1784 11150 1794
rect 557 1756 618 1766
rect 557 1674 618 1684
rect 1083 1756 1144 1766
rect 1083 1674 1144 1684
rect 2031 1756 2092 1766
rect 2031 1674 2092 1684
rect 2557 1756 2618 1766
rect 2557 1674 2618 1684
rect 3505 1756 3566 1766
rect 3505 1674 3566 1684
rect 4031 1756 4092 1766
rect 4031 1674 4092 1684
rect 4979 1756 5040 1766
rect 4979 1674 5040 1684
rect 5505 1756 5566 1766
rect 5505 1674 5566 1684
rect 6453 1756 6514 1766
rect 6453 1674 6514 1684
rect 6979 1756 7040 1766
rect 6979 1674 7040 1684
rect 7927 1756 7988 1766
rect 7927 1674 7988 1684
rect 8453 1756 8514 1766
rect 8453 1674 8514 1684
rect 9401 1756 9462 1766
rect 9401 1674 9462 1684
rect 9927 1756 9988 1766
rect 9927 1674 9988 1684
rect 11073 1409 11133 1784
rect 10952 1349 11133 1409
rect 10952 756 11012 1349
rect 10952 682 11012 692
rect 19 559 80 569
rect 19 493 80 503
rect 1671 559 1732 569
rect 3348 559 3409 569
rect 1732 518 1751 544
rect 1671 493 1732 503
rect 5035 559 5096 569
rect 3421 520 3446 546
rect 3348 493 3409 503
rect 6725 559 6786 569
rect 5106 519 5131 545
rect 5035 493 5096 503
rect 8413 559 8474 569
rect 6790 520 6815 546
rect 6725 493 6786 503
rect 10098 559 10159 569
rect 11744 567 11805 569
rect 8481 514 8506 540
rect 8413 493 8474 503
rect 11726 559 11805 567
rect 11726 552 11744 559
rect 10168 516 10193 542
rect 10098 493 10159 503
rect 11727 503 11744 510
rect 11727 495 11805 503
rect 11744 493 11805 495
rect 3 141 75 151
rect -208 49 3 124
rect -208 40 75 49
rect 3 39 75 40
<< via2 >>
rect 2972 2256 3043 2330
rect 7396 2430 7467 2514
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
rect 10952 692 11012 756
rect 19 503 80 559
rect 1671 503 1732 559
rect 3348 503 3409 559
rect 5035 503 5096 559
rect 6725 503 6786 559
rect 8413 503 8474 559
rect 10098 503 10159 559
rect 11744 503 11805 559
<< metal3 >>
rect 2981 2514 7477 2553
rect 2981 2493 7396 2514
rect 2981 2335 3041 2493
rect 7386 2430 7396 2493
rect 7467 2430 7477 2514
rect 7386 2425 7477 2430
rect 2962 2330 3053 2335
rect 2962 2256 2972 2330
rect 3043 2256 3053 2330
rect 2962 2251 3053 2256
rect 4497 2265 7957 2337
rect 1632 2014 3218 2086
rect 1632 1925 1704 2014
rect 1171 1853 1704 1925
rect 2753 1859 2903 1919
rect 2782 1848 2903 1859
rect 525 1756 628 1761
rect 525 1684 557 1756
rect 618 1684 628 1756
rect 525 1679 628 1684
rect 1054 1756 1154 1761
rect 1054 1684 1083 1756
rect 1144 1684 1154 1756
rect 1054 1679 1154 1684
rect 2021 1756 2102 1761
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2021 1679 2102 1684
rect 2547 1756 2628 1761
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 2547 1679 2628 1684
rect 525 1183 585 1679
rect 26 1123 585 1183
rect 1054 1173 1114 1679
rect 26 564 86 1123
rect 1054 1113 1725 1173
rect 1665 564 1725 1113
rect 2031 699 2091 1679
rect 2564 867 2624 1679
rect 2843 1536 2903 1848
rect 3146 1769 3218 2014
rect 4497 1925 4569 2265
rect 6173 2039 7718 2111
rect 6173 1925 6245 2039
rect 4119 1853 4569 1925
rect 5593 1853 6245 1925
rect 7067 1853 7366 1925
rect 3146 1761 3560 1769
rect 3146 1756 3576 1761
rect 3146 1697 3505 1756
rect 3495 1684 3505 1697
rect 3566 1684 3576 1756
rect 4021 1756 4102 1761
rect 4021 1734 4031 1756
rect 3495 1679 3576 1684
rect 4020 1684 4031 1734
rect 4092 1684 4102 1756
rect 4020 1679 4102 1684
rect 4969 1756 5050 1761
rect 4969 1684 4979 1756
rect 5040 1748 5050 1756
rect 5495 1756 5576 1761
rect 5040 1684 5060 1748
rect 4969 1679 5060 1684
rect 5495 1684 5505 1756
rect 5566 1743 5576 1756
rect 6443 1756 6524 1761
rect 5566 1684 5585 1743
rect 5495 1679 5585 1684
rect 6443 1684 6453 1756
rect 6514 1734 6524 1756
rect 6969 1756 7050 1761
rect 6514 1684 6525 1734
rect 6443 1679 6525 1684
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 6969 1679 7050 1684
rect 4020 1536 4080 1679
rect 2843 1476 4080 1536
rect 5000 1067 5060 1679
rect 5000 1007 5405 1067
rect 2564 807 5099 867
rect 2031 639 3414 699
rect 3354 564 3414 639
rect 5039 564 5099 807
rect 5345 809 5405 1007
rect 5525 950 5585 1679
rect 6465 1150 6525 1679
rect 6980 1335 7040 1679
rect 7294 1574 7366 1853
rect 7646 1774 7718 2039
rect 7885 2090 7957 2265
rect 7885 2018 9156 2090
rect 8541 1853 8845 1925
rect 7646 1761 7996 1774
rect 7646 1756 7998 1761
rect 7646 1702 7927 1756
rect 7917 1684 7927 1702
rect 7988 1684 7998 1756
rect 8443 1756 8524 1761
rect 8443 1742 8453 1756
rect 7917 1679 7998 1684
rect 8438 1684 8453 1742
rect 8514 1684 8524 1756
rect 8438 1679 8524 1684
rect 8438 1574 8510 1679
rect 7294 1502 8510 1574
rect 8773 1554 8845 1853
rect 9084 1769 9156 2018
rect 9084 1761 9446 1769
rect 9084 1756 9472 1761
rect 9084 1697 9401 1756
rect 9391 1684 9401 1697
rect 9462 1684 9472 1756
rect 9917 1756 9998 1761
rect 9917 1748 9927 1756
rect 9391 1679 9472 1684
rect 9902 1684 9927 1748
rect 9988 1684 9998 1756
rect 9902 1679 9998 1684
rect 9902 1554 9974 1679
rect 8773 1482 9974 1554
rect 6980 1275 10476 1335
rect 6465 1090 10166 1150
rect 5525 890 8474 950
rect 5345 749 6788 809
rect 6728 564 6788 749
rect 8414 564 8474 890
rect 10106 564 10166 1090
rect 10416 931 10476 1275
rect 10416 871 11810 931
rect 10942 756 11022 761
rect 10942 692 10952 756
rect 11012 692 11022 756
rect 10942 687 11022 692
rect 9 563 90 564
rect 9 559 145 563
rect 9 503 19 559
rect 80 503 145 559
rect 9 498 145 503
rect 1661 559 1742 564
rect 1661 503 1671 559
rect 1732 503 1742 559
rect 1661 498 1742 503
rect 3338 559 3419 564
rect 3338 503 3348 559
rect 3409 503 3419 559
rect 3338 498 3419 503
rect 5025 559 5106 564
rect 5025 503 5035 559
rect 5096 503 5106 559
rect 5025 498 5106 503
rect 6715 559 6796 564
rect 6715 503 6725 559
rect 6786 503 6796 559
rect 6715 498 6796 503
rect 8403 559 8484 564
rect 8403 503 8413 559
rect 8474 503 8484 559
rect 8403 498 8484 503
rect 10088 559 10169 564
rect 10088 503 10098 559
rect 10159 503 10169 559
rect 10088 498 10169 503
rect 85 112 145 498
rect 10952 112 11012 687
rect 11750 564 11810 871
rect 11734 559 11815 564
rect 11734 503 11744 559
rect 11805 503 11815 559
rect 11734 498 11815 503
rect 85 52 11012 112
use mux_2to1_logic  mux_2to1_logic_1
timestamp 1623959084
transform 1 0 1949 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_0
timestamp 1623959084
transform 1 0 475 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_0
timestamp 1623938174
transform 1 0 -10 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_1
timestamp 1623938174
transform 1 0 834 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_2
timestamp 1623959084
transform 1 0 3423 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_2
timestamp 1623938174
transform 1 0 1678 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_3
timestamp 1623938174
transform 1 0 2522 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_3
timestamp 1623959084
transform 1 0 4897 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_4
timestamp 1623938174
transform 1 0 3366 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_5
timestamp 1623938174
transform 1 0 4210 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_4
timestamp 1623959084
transform 1 0 6371 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_6
timestamp 1623938174
transform 1 0 5054 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_5
timestamp 1623959084
transform 1 0 7845 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_7
timestamp 1623938174
transform 1 0 5898 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_8
timestamp 1623938174
transform 1 0 6742 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_6
timestamp 1623959084
transform 1 0 9319 0 -1 1770
box -475 -633 999 607
use buffer_no_inv_x05  buffer_no_inv_x05_9
timestamp 1623938174
transform 1 0 7586 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_10
timestamp 1623938174
transform 1 0 8430 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_11
timestamp 1623938174
transform 1 0 9274 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_12
timestamp 1623938174
transform 1 0 10118 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_13
timestamp 1623938174
transform 1 0 10962 0 1 -10
box 10 10 854 1173
use nand_logic  nand_logic_0
timestamp 1623952422
transform 1 0 10695 0 -1 1870
box -219 -731 833 707
<< labels >>
rlabel via2 30 516 55 542 1 clk
rlabel metal2 8893 2121 8918 2147 1 reg0
rlabel metal3 6059 2508 6084 2534 1 reg1
rlabel space 11254 1972 11279 1998 1 clk_out
rlabel metal2 80 2501 105 2527 1 reg2
rlabel space 32 1216 57 1242 1 avdd1p8
rlabel space 146 2318 171 2344 1 avss1p8
<< end >>
