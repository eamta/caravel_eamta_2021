magic
tech sky130A
magscale 1 2
timestamp 1623250946
<< nwell >>
rect 574 13423 4975 13709
rect 605 9716 651 9807
<< pwell >>
rect 638 6873 5041 6937
rect 638 6866 668 6873
rect 723 6866 5041 6873
rect 638 -852 5041 6866
<< psubdiff >>
rect 2823 6860 2922 6861
rect 4971 6820 5005 6860
rect 675 3508 709 3546
rect 2823 3508 2857 3570
rect 4971 3507 5005 3584
rect 709 -836 733 -664
rect 4906 -836 4930 -664
<< nsubdiff >>
rect 670 13481 694 13653
rect 4867 13481 4891 13653
<< psubdiffcont >>
rect 675 3546 709 4712
rect 733 -836 4906 -664
<< nsubdiffcont >>
rect 694 13481 4867 13653
<< locali >>
rect 678 13481 694 13653
rect 4867 13481 4883 13653
rect 2823 6860 2922 6861
rect 4971 6820 5005 6860
rect 675 3508 709 3546
rect 2823 3508 2857 3570
rect 4971 3507 5005 3584
rect 717 -836 733 -664
rect 4906 -836 4922 -664
<< viali >>
rect 694 13481 4867 13653
rect 707 13389 4489 13423
rect 611 10224 645 13326
rect 4551 10224 4585 13326
rect 707 10127 3008 10161
rect 707 9767 2697 9801
rect 611 7502 645 9704
rect 2759 7589 2827 9704
rect 707 7405 2697 7439
rect 771 6827 2761 6861
rect 2919 6826 4909 6860
rect 675 4808 709 6764
rect 675 3546 709 4712
rect 4971 3608 5005 6764
rect 675 -456 709 3450
rect 4971 -456 5005 3450
rect 771 -552 2761 -518
rect 2919 -552 4909 -518
rect 733 -836 4906 -664
<< metal1 >>
rect 605 13653 4879 13659
rect 605 13481 694 13653
rect 4867 13481 4879 13653
rect 605 13423 4879 13481
rect 605 13389 707 13423
rect 4489 13389 4879 13423
rect 605 13383 4879 13389
rect 605 13326 651 13383
rect 605 10224 611 13326
rect 645 10224 651 13326
rect 704 10311 714 13319
rect 770 10311 780 13319
rect 847 13303 893 13383
rect 960 10311 970 13319
rect 1026 10311 1036 13319
rect 1103 13307 1149 13383
rect 1216 10311 1226 13319
rect 1282 10311 1292 13319
rect 1359 13308 1405 13383
rect 1472 10311 1482 13319
rect 1538 10311 1548 13319
rect 1615 13306 1661 13383
rect 1728 10311 1738 13319
rect 1794 10311 1804 13319
rect 1871 13307 1917 13383
rect 1984 10311 1994 13319
rect 2050 10311 2060 13319
rect 2127 13306 2173 13383
rect 2240 10311 2250 13319
rect 2306 10311 2316 13319
rect 2383 13307 2429 13383
rect 2496 10311 2506 13319
rect 2562 10311 2572 13319
rect 2639 13307 2685 13383
rect 2752 10311 2762 13319
rect 2818 10311 2828 13319
rect 2895 13307 2941 13383
rect 3008 10311 3018 13319
rect 3074 10311 3084 13319
rect 3151 13308 3197 13383
rect 3264 10311 3274 13319
rect 3330 10311 3340 13319
rect 3407 13308 3453 13383
rect 3520 10311 3530 13319
rect 3586 10311 3596 13319
rect 3663 13307 3709 13383
rect 3776 10311 3786 13319
rect 3842 10311 3852 13319
rect 3919 13310 3965 13383
rect 4032 10311 4042 13319
rect 4098 10311 4108 13319
rect 4175 13307 4221 13383
rect 4288 10311 4298 13319
rect 4354 10311 4364 13319
rect 4431 13306 4477 13383
rect 4545 13326 4591 13383
rect 605 10167 651 10224
rect 771 10219 4425 10275
rect 4545 10224 4551 13326
rect 4585 10224 4591 13326
rect 605 10161 3020 10167
rect 605 10127 707 10161
rect 3008 10127 3020 10161
rect 605 10121 3020 10127
rect 604 9801 2837 9807
rect 604 9767 707 9801
rect 2697 9767 2837 9801
rect 604 9761 2837 9767
rect 605 9704 651 9761
rect 605 7502 611 9704
rect 645 7502 651 9704
rect 2749 9704 2837 9761
rect 704 7585 714 9693
rect 770 7585 780 9693
rect 832 7585 842 9693
rect 898 7585 908 9693
rect 960 7585 970 9693
rect 1026 7585 1036 9693
rect 1088 7585 1098 9693
rect 1154 7585 1164 9693
rect 1216 7585 1226 9693
rect 1282 7585 1292 9693
rect 1344 7585 1354 9693
rect 1410 7585 1420 9693
rect 1472 7585 1482 9693
rect 1538 7585 1548 9693
rect 1600 7585 1610 9693
rect 1666 7585 1676 9693
rect 1728 7585 1738 9693
rect 1794 7585 1804 9693
rect 1856 7585 1866 9693
rect 1922 7585 1932 9693
rect 1984 7585 1994 9693
rect 2050 7585 2060 9693
rect 2112 7585 2122 9693
rect 2178 7585 2188 9693
rect 2240 7585 2250 9693
rect 2306 7585 2316 9693
rect 2368 7585 2378 9693
rect 2434 7585 2444 9693
rect 2496 7585 2506 9693
rect 2562 7585 2572 9693
rect 2624 7585 2634 9693
rect 2690 7585 2700 9693
rect 2749 7589 2759 9704
rect 2827 7589 2837 9704
rect 3563 9604 3844 10219
rect 4545 10212 4591 10224
rect 3553 9389 3563 9604
rect 3844 9389 3854 9604
rect 2931 8069 2941 8554
rect 3196 8069 3206 8554
rect 2753 7577 2833 7589
rect 2941 7548 3196 8069
rect 769 7502 3196 7548
rect 605 7445 651 7502
rect 605 7439 2709 7445
rect 605 7405 707 7439
rect 2697 7405 2709 7439
rect 605 7399 2709 7405
rect 605 7398 720 7399
rect 759 6866 5011 6867
rect 669 6861 5011 6866
rect 669 6827 771 6861
rect 2761 6860 5011 6861
rect 2761 6827 2919 6860
rect 669 6826 2919 6827
rect 4909 6826 5011 6860
rect 669 6821 5011 6826
rect 669 6772 716 6821
rect 2907 6820 5011 6821
rect 669 6764 715 6772
rect 669 4808 675 6764
rect 709 4808 715 6764
rect 2697 6725 3010 6790
rect 4965 6764 5011 6820
rect 764 4882 774 6690
rect 838 4882 848 6690
rect 669 4712 715 4808
rect 669 3546 675 4712
rect 709 3546 715 4712
rect 669 3450 715 3546
rect 879 4825 925 4894
rect 956 4882 966 6690
rect 1030 4882 1040 6690
rect 1071 4825 1117 4895
rect 1148 4882 1158 6690
rect 1222 4882 1232 6690
rect 1263 4825 1309 4893
rect 1340 4882 1350 6690
rect 1414 4882 1424 6690
rect 1455 4825 1501 4893
rect 1532 4882 1542 6690
rect 1606 4882 1616 6690
rect 1647 4825 1693 4894
rect 1724 4882 1734 6690
rect 1798 4882 1808 6690
rect 1839 4825 1885 4894
rect 1916 4882 1926 6690
rect 1990 4882 2000 6690
rect 2031 4825 2077 4894
rect 2108 4882 2118 6690
rect 2182 4882 2192 6690
rect 2223 4825 2269 4895
rect 2300 4882 2310 6690
rect 2374 4882 2384 6690
rect 2415 4825 2461 4894
rect 2492 4882 2502 6690
rect 2566 4882 2576 6690
rect 2607 4825 2653 4893
rect 2684 4882 2694 6690
rect 2758 4882 2768 6690
rect 879 3563 2653 4825
rect 2912 3682 2922 6690
rect 2986 3682 2996 6690
rect 3027 3623 3073 3693
rect 3104 3682 3114 6690
rect 3178 3682 3188 6690
rect 3219 3623 3265 3695
rect 3296 3681 3306 6689
rect 3370 3681 3380 6689
rect 3411 3623 3457 3701
rect 3488 3682 3498 6690
rect 3562 3682 3572 6690
rect 3603 3623 3649 3694
rect 3680 3682 3690 6690
rect 3754 3682 3764 6690
rect 3795 3623 3841 3697
rect 3872 3682 3882 6690
rect 3946 3682 3956 6690
rect 3987 3623 4033 3699
rect 4064 3682 4074 6690
rect 4138 3682 4148 6690
rect 4179 3623 4225 3700
rect 4256 3682 4266 6690
rect 4330 3682 4340 6690
rect 4371 3623 4417 3698
rect 4448 3682 4458 6690
rect 4522 3682 4532 6690
rect 4563 3623 4609 3698
rect 4640 3682 4650 6690
rect 4714 3682 4724 6690
rect 4755 3623 4801 3698
rect 4832 3682 4842 6690
rect 4906 3682 4916 6690
rect 879 3494 1360 3563
rect 1487 3494 2042 3563
rect 2169 3494 2653 3563
rect 3017 3536 3027 3623
rect 4801 3536 4811 3623
rect 4965 3608 4971 6764
rect 5005 3608 5011 6764
rect 879 3485 2653 3494
rect 879 3481 3036 3485
rect 879 3467 2653 3481
rect 879 3464 2075 3467
rect 947 3463 2075 3464
rect 947 3461 1062 3463
rect 1088 3461 2075 3463
rect 2085 3461 2653 3467
rect 669 -456 675 3450
rect 709 -456 715 3450
rect 879 3437 897 3461
rect 1002 3458 2653 3461
rect 1032 3453 2653 3458
rect 1061 3438 2653 3453
rect 879 3369 925 3437
rect 879 3364 923 3369
rect 1071 3365 1117 3438
rect 1263 3366 1309 3438
rect 1455 3367 1501 3438
rect 1647 3366 1693 3438
rect 1839 3363 1885 3438
rect 2031 3367 2077 3438
rect 2223 3368 2269 3438
rect 2415 3367 2461 3438
rect 2607 3367 2653 3438
rect 2665 3424 3036 3481
rect 4965 3450 5011 3608
rect 669 -459 715 -456
rect 783 -459 829 -365
rect 975 -459 1021 -367
rect 1167 -459 1213 -365
rect 1359 -459 1405 -366
rect 1551 -459 1597 -366
rect 1743 -459 1789 -363
rect 1935 -459 1981 -371
rect 2127 -459 2173 -366
rect 2319 -459 2365 -369
rect 2511 -459 2557 -373
rect 2703 -459 2749 -367
rect 2931 -459 2977 -366
rect 3008 -382 3018 3376
rect 3082 -382 3092 3376
rect 3123 -459 3169 -371
rect 3200 -382 3210 3376
rect 3274 -382 3284 3376
rect 3315 -459 3361 -368
rect 3392 -382 3402 3376
rect 3466 -382 3476 3376
rect 3507 -459 3553 -367
rect 3584 -382 3594 3376
rect 3658 -382 3668 3376
rect 3699 -459 3745 -367
rect 3776 -382 3786 3376
rect 3850 -382 3860 3376
rect 3891 -459 3937 -365
rect 3968 -382 3978 3376
rect 4042 -382 4052 3376
rect 4083 -459 4129 -363
rect 4160 -382 4170 3376
rect 4234 -382 4244 3376
rect 4275 -459 4321 -363
rect 4352 -382 4362 3376
rect 4426 -382 4436 3376
rect 4467 -459 4513 -363
rect 4544 -382 4554 3376
rect 4618 -382 4628 3376
rect 4659 -459 4705 -360
rect 4736 -382 4746 3376
rect 4810 -382 4820 3376
rect 4851 -459 4897 -366
rect 4965 -456 4971 3450
rect 5005 -456 5011 3450
rect 4965 -459 5011 -456
rect 669 -518 5011 -459
rect 669 -552 771 -518
rect 2761 -552 2919 -518
rect 4909 -552 5011 -518
rect 669 -664 5011 -552
rect 669 -836 733 -664
rect 4906 -836 5011 -664
rect 669 -842 5011 -836
<< via1 >>
rect 694 13481 4867 13653
rect 714 10311 770 13319
rect 970 10311 1026 13319
rect 1226 10311 1282 13319
rect 1482 10311 1538 13319
rect 1738 10311 1794 13319
rect 1994 10311 2050 13319
rect 2250 10311 2306 13319
rect 2506 10311 2562 13319
rect 2762 10311 2818 13319
rect 3018 10311 3074 13319
rect 3274 10311 3330 13319
rect 3530 10311 3586 13319
rect 3786 10311 3842 13319
rect 4042 10311 4098 13319
rect 4298 10311 4354 13319
rect 714 7585 770 9693
rect 842 7585 898 9693
rect 970 7585 1026 9693
rect 1098 7585 1154 9693
rect 1226 7585 1282 9693
rect 1354 7585 1410 9693
rect 1482 7585 1538 9693
rect 1610 7585 1666 9693
rect 1738 7585 1794 9693
rect 1866 7585 1922 9693
rect 1994 7585 2050 9693
rect 2122 7585 2178 9693
rect 2250 7585 2306 9693
rect 2378 7585 2434 9693
rect 2506 7585 2562 9693
rect 2634 7585 2690 9693
rect 2759 7589 2827 9704
rect 3563 9389 3844 9604
rect 2941 8069 3196 8554
rect 774 4882 838 6690
rect 966 4882 1030 6690
rect 1158 4882 1222 6690
rect 1350 4882 1414 6690
rect 1542 4882 1606 6690
rect 1734 4882 1798 6690
rect 1926 4882 1990 6690
rect 2118 4882 2182 6690
rect 2310 4882 2374 6690
rect 2502 4882 2566 6690
rect 2694 4882 2758 6690
rect 2922 3682 2986 6690
rect 3114 3682 3178 6690
rect 3306 3681 3370 6689
rect 3498 3682 3562 6690
rect 3690 3682 3754 6690
rect 3882 3682 3946 6690
rect 4074 3682 4138 6690
rect 4266 3682 4330 6690
rect 4458 3682 4522 6690
rect 4650 3682 4714 6690
rect 4842 3682 4906 6690
rect 3027 3536 4801 3623
rect 3018 -382 3082 3376
rect 3210 -382 3274 3376
rect 3402 -382 3466 3376
rect 3594 -382 3658 3376
rect 3786 -382 3850 3376
rect 3978 -382 4042 3376
rect 4170 -382 4234 3376
rect 4362 -382 4426 3376
rect 4554 -382 4618 3376
rect 4746 -382 4810 3376
rect 733 -836 4906 -664
<< metal2 >>
rect 694 13653 4867 13663
rect 694 13471 4867 13481
rect 714 13319 770 13329
rect 714 10118 770 10311
rect 970 13319 1026 13329
rect 970 10118 1026 10311
rect 1226 13319 1282 13329
rect 1226 10118 1282 10311
rect 1482 13319 1538 13329
rect 1482 10118 1538 10311
rect 1738 13319 1794 13329
rect 1738 10118 1794 10311
rect 1994 13319 2050 13329
rect 1994 10118 2050 10311
rect 2250 13319 2306 13329
rect 2250 10118 2306 10311
rect 2506 13319 2562 13329
rect 2506 10118 2562 10311
rect 2762 13319 2818 13329
rect 2762 10118 2818 10311
rect 3018 13319 3074 13329
rect 3018 10118 3074 10311
rect 3274 13319 3330 13329
rect 3274 10118 3330 10311
rect 3530 13319 3586 13329
rect 3530 10118 3586 10311
rect 3786 13319 3842 13329
rect 3786 10118 3842 10311
rect 4042 13319 4098 13329
rect 4042 10118 4098 10311
rect 4298 13319 4354 13329
rect 4298 10118 4354 10311
rect 714 9731 4354 10118
rect 714 9693 770 9731
rect 714 7575 770 7585
rect 842 9693 898 9703
rect 842 7393 898 7585
rect 970 9693 1026 9731
rect 970 7575 1026 7585
rect 1098 9693 1154 9703
rect 1098 7393 1154 7585
rect 1226 9693 1282 9731
rect 1226 7575 1282 7585
rect 1354 9693 1410 9703
rect 1354 7393 1410 7585
rect 1482 9693 1538 9731
rect 1482 7575 1538 7585
rect 1610 9693 1666 9703
rect 1610 7393 1666 7585
rect 1738 9693 1794 9731
rect 1738 7575 1794 7585
rect 1866 9693 1922 9703
rect 1866 7393 1922 7585
rect 1994 9693 2050 9731
rect 1994 7575 2050 7585
rect 2122 9693 2178 9703
rect 2122 7393 2178 7585
rect 2250 9693 2306 9731
rect 2250 7575 2306 7585
rect 2378 9693 2434 9703
rect 2378 7393 2434 7585
rect 2506 9693 2562 9731
rect 2759 9704 2827 9731
rect 2506 7575 2562 7585
rect 2634 9693 2690 9703
rect 2634 7393 2690 7585
rect 3563 9604 3844 9614
rect 3563 9379 3844 9389
rect 2941 8554 3196 8564
rect 2941 8059 3196 8069
rect 2759 7579 2827 7589
rect 774 7382 2690 7393
rect 774 7106 2689 7382
rect 774 6784 2690 7106
rect 3722 7087 4648 8053
rect 774 6726 2758 6784
rect 774 6725 900 6726
rect 774 6690 838 6725
rect 774 4872 838 4882
rect 966 6690 1030 6726
rect 966 4872 1030 4882
rect 1158 6690 1222 6726
rect 1158 4872 1222 4882
rect 1350 6690 1414 6726
rect 1350 4872 1414 4882
rect 1542 6690 1606 6726
rect 1542 4872 1606 4882
rect 1734 6690 1798 6726
rect 1734 4872 1798 4882
rect 1926 6690 1990 6726
rect 1926 4872 1990 4882
rect 2118 6690 2182 6726
rect 2118 4872 2182 4882
rect 2310 6690 2374 6726
rect 2310 4872 2374 4882
rect 2502 6690 2566 6726
rect 2683 6725 2758 6726
rect 2502 4872 2566 4882
rect 2694 6690 2758 6725
rect 2694 4872 2758 4882
rect 2922 6763 4906 7087
rect 2922 6690 2986 6763
rect 2922 3672 2986 3682
rect 3114 6690 3178 6763
rect 3114 3672 3178 3682
rect 3306 6689 3370 6763
rect 3306 3671 3370 3681
rect 3498 6690 3562 6763
rect 3498 3672 3562 3682
rect 3690 6690 3754 6763
rect 3690 3672 3754 3682
rect 3882 6690 3946 6763
rect 3882 3672 3946 3682
rect 4074 6690 4138 6763
rect 4074 3672 4138 3682
rect 4266 6690 4330 6763
rect 4266 3672 4330 3682
rect 4458 6690 4522 6763
rect 4458 3672 4522 3682
rect 4650 6690 4714 6763
rect 4650 3672 4714 3682
rect 4842 6690 4906 6763
rect 4842 3672 4906 3682
rect 3027 3623 4801 3633
rect 3018 3536 3027 3623
rect 4801 3536 4810 3623
rect 3018 3386 4810 3536
rect 3018 3376 3082 3386
rect 3018 -392 3082 -382
rect 3210 3376 3274 3386
rect 3210 -392 3274 -382
rect 3402 3376 3466 3386
rect 3402 -392 3466 -382
rect 3594 3376 3658 3386
rect 3594 -392 3658 -382
rect 3786 3376 3850 3386
rect 3786 -392 3850 -382
rect 3978 3376 4042 3386
rect 3978 -392 4042 -382
rect 4170 3376 4234 3386
rect 4170 -392 4234 -382
rect 4362 3376 4426 3386
rect 4362 -392 4426 -382
rect 4554 3376 4618 3386
rect 4554 -392 4618 -382
rect 4746 3376 4810 3386
rect 4746 -392 4810 -382
rect 733 -664 4906 -654
rect 733 -846 4906 -836
use sky130_fd_pr__nfet_01v8_lvt_SNTUMW  M1
timestamp 1623250946
transform 1 0 3914 0 1 5186
box -1127 -1710 1127 1710
use sky130_fd_pr__nfet_01v8_lvt_EU6LGP  M4
timestamp 1623250946
transform 1 0 1766 0 1 1497
box -1127 -2085 1127 2085
use sky130_fd_pr__nfet_01v8_lvt_5U6LBF  M2
timestamp 1623250946
transform 1 0 3914 0 1 1497
box -1127 -2085 1127 2085
use sky130_fd_pr__nfet_01v8_lvt_L5XAT6  M3
timestamp 1623248045
transform 1 0 1766 0 1 5786
box -1127 -1110 1127 1110
use sky130_fd_pr__pfet_01v8_lvt_QTSHDD  M5
timestamp 1623247083
transform 1 0 1702 0 1 8603
box -1127 -1234 1127 1234
use sky130_fd_pr__pfet_01v8_lvt_ND8574  M6
timestamp 1623247083
transform 1 0 2598 0 1 11775
box -2023 -1684 2023 1684
<< labels >>
rlabel via1 3563 9389 3844 9604 1 vbias_1
rlabel via1 2941 8069 3196 8554 1 vbias_2
rlabel metal2 3722 7557 4648 8053 1 ibias
rlabel nwell 694 13481 4867 13653 1 vdd
rlabel pwell 733 -836 4906 -664 1 vss
<< end >>
