magic
tech sky130A
magscale 1 2
timestamp 1623250946
<< pwell >>
rect -1127 -1710 1127 1710
<< nmoslvt >>
rect -927 -1500 -897 1500
rect -831 -1500 -801 1500
rect -735 -1500 -705 1500
rect -639 -1500 -609 1500
rect -543 -1500 -513 1500
rect -447 -1500 -417 1500
rect -351 -1500 -321 1500
rect -255 -1500 -225 1500
rect -159 -1500 -129 1500
rect -63 -1500 -33 1500
rect 33 -1500 63 1500
rect 129 -1500 159 1500
rect 225 -1500 255 1500
rect 321 -1500 351 1500
rect 417 -1500 447 1500
rect 513 -1500 543 1500
rect 609 -1500 639 1500
rect 705 -1500 735 1500
rect 801 -1500 831 1500
rect 897 -1500 927 1500
<< ndiff >>
rect -989 1488 -927 1500
rect -989 -1488 -977 1488
rect -943 -1488 -927 1488
rect -989 -1500 -927 -1488
rect -897 1488 -831 1500
rect -897 -1488 -881 1488
rect -847 -1488 -831 1488
rect -897 -1500 -831 -1488
rect -801 1488 -735 1500
rect -801 -1488 -785 1488
rect -751 -1488 -735 1488
rect -801 -1500 -735 -1488
rect -705 1488 -639 1500
rect -705 -1488 -689 1488
rect -655 -1488 -639 1488
rect -705 -1500 -639 -1488
rect -609 1488 -543 1500
rect -609 -1488 -593 1488
rect -559 -1488 -543 1488
rect -609 -1500 -543 -1488
rect -513 1488 -447 1500
rect -513 -1488 -497 1488
rect -463 -1488 -447 1488
rect -513 -1500 -447 -1488
rect -417 1488 -351 1500
rect -417 -1488 -401 1488
rect -367 -1488 -351 1488
rect -417 -1500 -351 -1488
rect -321 1488 -255 1500
rect -321 -1488 -305 1488
rect -271 -1488 -255 1488
rect -321 -1500 -255 -1488
rect -225 1488 -159 1500
rect -225 -1488 -209 1488
rect -175 -1488 -159 1488
rect -225 -1500 -159 -1488
rect -129 1488 -63 1500
rect -129 -1488 -113 1488
rect -79 -1488 -63 1488
rect -129 -1500 -63 -1488
rect -33 1488 33 1500
rect -33 -1488 -17 1488
rect 17 -1488 33 1488
rect -33 -1500 33 -1488
rect 63 1488 129 1500
rect 63 -1488 79 1488
rect 113 -1488 129 1488
rect 63 -1500 129 -1488
rect 159 1488 225 1500
rect 159 -1488 175 1488
rect 209 -1488 225 1488
rect 159 -1500 225 -1488
rect 255 1488 321 1500
rect 255 -1488 271 1488
rect 305 -1488 321 1488
rect 255 -1500 321 -1488
rect 351 1488 417 1500
rect 351 -1488 367 1488
rect 401 -1488 417 1488
rect 351 -1500 417 -1488
rect 447 1488 513 1500
rect 447 -1488 463 1488
rect 497 -1488 513 1488
rect 447 -1500 513 -1488
rect 543 1488 609 1500
rect 543 -1488 559 1488
rect 593 -1488 609 1488
rect 543 -1500 609 -1488
rect 639 1488 705 1500
rect 639 -1488 655 1488
rect 689 -1488 705 1488
rect 639 -1500 705 -1488
rect 735 1488 801 1500
rect 735 -1488 751 1488
rect 785 -1488 801 1488
rect 735 -1500 801 -1488
rect 831 1488 897 1500
rect 831 -1488 847 1488
rect 881 -1488 897 1488
rect 831 -1500 897 -1488
rect 927 1488 989 1500
rect 927 -1488 943 1488
rect 977 -1488 989 1488
rect 927 -1500 989 -1488
<< ndiffc >>
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
<< psubdiff >>
rect -1091 1640 -995 1674
rect 995 1640 1091 1674
rect -1091 -1640 -1057 1640
rect 1057 1578 1091 1640
rect 1057 -1640 1091 -1578
<< psubdiffcont >>
rect -995 1640 995 1674
rect 1057 -1578 1091 1578
<< poly >>
rect -927 1588 927 1611
rect -927 1554 -896 1588
rect 908 1554 927 1588
rect -927 1522 927 1554
rect -927 1500 -897 1522
rect -831 1500 -801 1522
rect -735 1500 -705 1522
rect -639 1500 -609 1522
rect -543 1500 -513 1522
rect -447 1500 -417 1522
rect -351 1500 -321 1522
rect -255 1500 -225 1522
rect -159 1500 -129 1522
rect -63 1500 -33 1522
rect 33 1500 63 1522
rect 129 1500 159 1522
rect 225 1500 255 1522
rect 321 1500 351 1522
rect 417 1500 447 1522
rect 513 1500 543 1522
rect 609 1500 639 1522
rect 705 1500 735 1522
rect 801 1500 831 1522
rect 897 1500 927 1522
rect -927 -1526 -897 -1500
rect -831 -1526 -801 -1500
rect -735 -1526 -705 -1500
rect -639 -1526 -609 -1500
rect -543 -1526 -513 -1500
rect -447 -1526 -417 -1500
rect -351 -1526 -321 -1500
rect -255 -1526 -225 -1500
rect -159 -1526 -129 -1500
rect -63 -1526 -33 -1500
rect 33 -1526 63 -1500
rect 129 -1526 159 -1500
rect 225 -1526 255 -1500
rect 321 -1526 351 -1500
rect 417 -1526 447 -1500
rect 513 -1526 543 -1500
rect 609 -1526 639 -1500
rect 705 -1526 735 -1500
rect 801 -1526 831 -1500
rect 897 -1526 927 -1500
<< polycont >>
rect -896 1554 908 1588
<< locali >>
rect -1091 1640 -995 1674
rect 995 1640 1091 1674
rect -1091 -1640 -1057 1640
rect -912 1591 924 1600
rect -912 1539 -899 1591
rect 917 1539 924 1591
rect -912 1538 924 1539
rect 1057 1578 1091 1640
rect -977 1488 -943 1504
rect -977 -1504 -943 -1488
rect -881 1488 -847 1504
rect -881 -1504 -847 -1488
rect -785 1488 -751 1504
rect -785 -1504 -751 -1488
rect -689 1488 -655 1504
rect -689 -1504 -655 -1488
rect -593 1488 -559 1504
rect -593 -1504 -559 -1488
rect -497 1488 -463 1504
rect -497 -1504 -463 -1488
rect -401 1488 -367 1504
rect -401 -1504 -367 -1488
rect -305 1488 -271 1504
rect -305 -1504 -271 -1488
rect -209 1488 -175 1504
rect -209 -1504 -175 -1488
rect -113 1488 -79 1504
rect -113 -1504 -79 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 79 1488 113 1504
rect 79 -1504 113 -1488
rect 175 1488 209 1504
rect 175 -1504 209 -1488
rect 271 1488 305 1504
rect 271 -1504 305 -1488
rect 367 1488 401 1504
rect 367 -1504 401 -1488
rect 463 1488 497 1504
rect 463 -1504 497 -1488
rect 559 1488 593 1504
rect 559 -1504 593 -1488
rect 655 1488 689 1504
rect 655 -1504 689 -1488
rect 751 1488 785 1504
rect 751 -1504 785 -1488
rect 847 1488 881 1504
rect 847 -1504 881 -1488
rect 943 1488 977 1504
rect 943 -1504 977 -1488
rect 1057 -1640 1091 -1578
<< viali >>
rect -899 1588 917 1591
rect -899 1554 -896 1588
rect -896 1554 908 1588
rect 908 1554 917 1588
rect -899 1539 917 1554
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
<< metal1 >>
rect -911 1591 929 1597
rect -911 1539 -899 1591
rect 917 1539 929 1591
rect -911 1533 929 1539
rect -983 1488 -937 1500
rect -983 -1488 -977 1488
rect -943 -1488 -937 1488
rect -983 -1500 -937 -1488
rect -887 1488 -841 1500
rect -887 -1488 -881 1488
rect -847 -1488 -841 1488
rect -887 -1500 -841 -1488
rect -791 1488 -745 1500
rect -791 -1488 -785 1488
rect -751 -1488 -745 1488
rect -791 -1500 -745 -1488
rect -695 1488 -649 1500
rect -695 -1488 -689 1488
rect -655 -1488 -649 1488
rect -695 -1500 -649 -1488
rect -599 1488 -553 1500
rect -599 -1488 -593 1488
rect -559 -1488 -553 1488
rect -599 -1500 -553 -1488
rect -503 1488 -457 1500
rect -503 -1488 -497 1488
rect -463 -1488 -457 1488
rect -503 -1500 -457 -1488
rect -407 1488 -361 1500
rect -407 -1488 -401 1488
rect -367 -1488 -361 1488
rect -407 -1500 -361 -1488
rect -311 1488 -265 1500
rect -311 -1488 -305 1488
rect -271 -1488 -265 1488
rect -311 -1500 -265 -1488
rect -215 1488 -169 1500
rect -215 -1488 -209 1488
rect -175 -1488 -169 1488
rect -215 -1500 -169 -1488
rect -119 1488 -73 1500
rect -119 -1488 -113 1488
rect -79 -1488 -73 1488
rect -119 -1500 -73 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 73 1488 119 1500
rect 73 -1488 79 1488
rect 113 -1488 119 1488
rect 73 -1500 119 -1488
rect 169 1488 215 1500
rect 169 -1488 175 1488
rect 209 -1488 215 1488
rect 169 -1500 215 -1488
rect 265 1488 311 1500
rect 265 -1488 271 1488
rect 305 -1488 311 1488
rect 265 -1500 311 -1488
rect 361 1488 407 1500
rect 361 -1488 367 1488
rect 401 -1488 407 1488
rect 361 -1500 407 -1488
rect 457 1488 503 1500
rect 457 -1488 463 1488
rect 497 -1488 503 1488
rect 457 -1500 503 -1488
rect 553 1488 599 1500
rect 553 -1488 559 1488
rect 593 -1488 599 1488
rect 553 -1500 599 -1488
rect 649 1488 695 1500
rect 649 -1488 655 1488
rect 689 -1488 695 1488
rect 649 -1500 695 -1488
rect 745 1488 791 1500
rect 745 -1488 751 1488
rect 785 -1488 791 1488
rect 745 -1500 791 -1488
rect 841 1488 887 1500
rect 841 -1488 847 1488
rect 881 -1488 887 1488
rect 841 -1500 887 -1488
rect 937 1488 983 1500
rect 937 -1488 943 1488
rect 977 -1488 983 1488
rect 937 -1500 983 -1488
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1074 -1657 1074 1657
string parameters w 15 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
