magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 298 1077 333 1111
rect 299 1058 333 1077
rect 129 1009 187 1015
rect 129 975 141 1009
rect 129 969 187 975
rect 318 821 333 1058
rect 352 1024 387 1058
rect 667 1024 702 1058
rect 352 821 386 1024
rect 668 1005 702 1024
rect 498 956 556 962
rect 498 922 510 956
rect 498 916 556 922
rect 466 821 500 872
rect 554 821 588 872
rect -53 547 647 821
rect 316 494 647 547
rect 687 530 702 1005
rect 721 971 756 1005
rect 1036 971 1071 1005
rect 721 530 755 971
rect 1037 952 1071 971
rect 1423 952 1476 953
rect 867 903 925 909
rect 867 869 879 903
rect 867 863 925 869
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1056 477 1071 952
rect 1090 918 1125 952
rect 1405 918 1476 952
rect 1090 477 1124 918
rect 1406 917 1476 918
rect 1423 883 1494 917
rect 1774 883 1809 917
rect 1236 850 1294 856
rect 1236 816 1248 850
rect 1236 810 1294 816
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1423 424 1493 883
rect 1775 864 1809 883
rect 1605 815 1663 821
rect 1605 781 1617 815
rect 1605 775 1663 781
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1794 371 1809 864
rect 1828 830 1863 864
rect 2143 830 2178 864
rect 1828 371 1862 830
rect 2144 811 2178 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 811
rect 2197 777 2232 811
rect 2512 777 2547 811
rect 2197 318 2231 777
rect 2513 758 2547 777
rect 2343 709 2401 715
rect 2343 675 2355 709
rect 2343 669 2401 675
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2532 265 2547 758
rect 2566 724 2601 758
rect 2881 724 2916 758
rect 2566 265 2600 724
rect 2882 705 2916 724
rect 2712 656 2770 662
rect 2712 622 2724 656
rect 2712 616 2770 622
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 2901 212 2916 705
rect 2935 671 2970 705
rect 3250 671 3285 705
rect 2935 212 2969 671
rect 3251 652 3285 671
rect 3081 603 3139 609
rect 3081 569 3093 603
rect 3081 563 3139 569
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3270 159 3285 652
rect 3304 618 3339 652
rect 3304 159 3338 618
rect 3450 550 3508 556
rect 3450 516 3462 550
rect 3620 527 3654 545
rect 3450 510 3508 516
rect 3620 491 3690 527
rect 3637 457 3708 491
rect 3988 457 4023 491
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3637 106 3707 457
rect 3989 438 4023 457
rect 3819 389 3877 395
rect 3819 355 3831 389
rect 3819 349 3877 355
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3637 70 3690 106
rect 4008 53 4023 438
rect 4042 404 4077 438
rect 4042 53 4076 404
rect 4188 336 4246 342
rect 4188 302 4200 336
rect 4188 296 4246 302
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 24 0 101 21
rect 131 0 200 21
rect 4042 19 4057 53
rect 24 -28 101 -7
rect 131 -28 228 -7
<< nwell >>
rect -354 820 647 821
rect -355 384 647 820
rect -355 381 -354 384
rect -342 381 647 384
<< psubdiff >>
rect -269 -117 -245 -83
rect 555 -117 579 -83
<< nsubdiff >>
rect -273 751 43 785
rect 353 751 576 785
<< psubdiffcont >>
rect -245 -117 555 -83
<< nsubdiffcont >>
rect 43 751 353 785
<< poly >>
rect 43 691 352 721
rect -260 428 -230 649
rect -60 428 -30 649
rect -260 398 -30 428
rect -260 384 -230 398
rect -295 368 -230 384
rect -295 334 -285 368
rect -251 334 -230 368
rect -295 318 -230 334
rect -260 -39 -230 318
rect -66 318 -12 333
rect 43 318 73 691
rect 146 363 176 649
rect 234 375 264 649
rect 322 417 352 691
rect 522 375 552 649
rect -66 317 73 318
rect -66 283 -56 317
rect -22 288 73 317
rect 138 347 192 363
rect 138 313 148 347
rect 182 313 192 347
rect 234 345 552 375
rect 138 297 192 313
rect -22 283 -12 288
rect -66 267 -12 283
rect -54 23 -24 267
rect 146 5 176 297
rect 522 276 552 345
rect 522 260 624 276
rect 234 -39 264 237
rect 322 5 352 237
rect 522 226 580 260
rect 614 226 624 260
rect 522 210 624 226
rect 522 5 552 210
rect 322 -25 552 5
rect -260 -69 264 -39
<< polycont >>
rect -285 334 -251 368
rect -56 283 -22 317
rect 148 313 182 347
rect 580 226 614 260
<< locali >>
rect -295 368 -241 384
rect -295 334 -285 368
rect -251 334 -241 368
rect -295 318 -241 334
rect 138 347 192 363
rect -66 317 -12 333
rect -66 283 -56 317
rect -22 283 -12 317
rect 138 313 148 347
rect 182 313 192 347
rect 138 297 192 313
rect -66 267 -12 283
rect 570 260 624 276
rect 570 226 580 260
rect 614 226 624 260
rect 570 210 624 226
<< viali >>
rect -273 751 43 785
rect 43 751 353 785
rect 353 751 576 785
rect -285 334 -251 368
rect -56 283 -22 317
rect 148 313 182 347
rect 580 226 614 260
rect -270 -117 -245 -83
rect -245 -117 555 -83
rect 555 -117 580 -83
rect -270 -118 580 -117
<< metal1 >>
rect -354 785 647 821
rect -354 751 -273 785
rect 576 751 647 785
rect -354 745 647 751
rect -301 638 -270 745
rect -309 559 -270 638
rect -109 624 -69 745
rect -109 611 -68 624
rect -309 452 -271 559
rect -220 452 -180 611
rect -108 459 -68 611
rect -21 587 19 617
rect 99 587 139 619
rect -21 483 139 587
rect -21 475 24 483
rect 95 475 139 483
rect 187 481 227 621
rect 362 617 402 745
rect -21 452 19 475
rect 99 454 139 475
rect 184 456 227 481
rect 361 608 402 617
rect -223 446 -180 452
rect -223 445 -195 446
rect -223 443 -189 445
rect 184 443 224 456
rect 361 452 401 608
rect 471 485 511 622
rect 567 616 598 745
rect 471 457 512 485
rect -342 368 -241 384
rect -342 334 -285 368
rect -251 334 -241 368
rect -342 318 -241 334
rect -212 316 -184 443
rect 182 433 224 443
rect 472 437 512 457
rect 564 451 604 616
rect 182 415 210 433
rect 56 387 210 415
rect 56 355 84 387
rect -66 317 -12 333
rect -66 316 -56 317
rect -212 287 -56 316
rect -310 46 -274 135
rect -212 133 -184 287
rect -66 283 -56 287
rect -22 283 -12 317
rect 31 303 41 355
rect 93 303 103 355
rect 138 347 192 359
rect 138 313 148 347
rect 182 327 192 347
rect 476 327 507 437
rect 182 313 507 327
rect -66 267 -12 283
rect 56 269 84 303
rect 138 299 507 313
rect 138 297 192 299
rect 56 239 210 269
rect -217 132 -186 133
rect -310 -76 -279 46
rect -222 45 -186 132
rect -107 77 -61 227
rect 182 217 210 239
rect 182 211 231 217
rect 89 200 137 202
rect 183 200 231 211
rect 0 157 231 200
rect -103 -76 -63 77
rect -6 42 231 157
rect -6 0 200 42
rect 270 25 318 200
rect 358 32 406 207
rect 476 154 507 299
rect 570 260 625 276
rect 570 226 580 260
rect 614 226 625 260
rect 570 210 625 226
rect 473 33 513 154
rect -6 -7 24 0
rect 101 -7 131 0
rect 278 -7 308 25
rect -6 -35 308 -7
rect 362 -76 402 32
rect 561 30 601 113
rect 565 -76 596 30
rect -355 -83 647 -76
rect -355 -118 -270 -83
rect 580 -118 647 -83
rect -355 -124 647 -118
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
<< via1 >>
rect 41 303 93 355
<< metal2 >>
rect 31 355 103 365
rect 31 303 41 355
rect 93 303 103 355
rect 31 293 103 303
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615150785
transform 1 0 -245 0 1 88
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_0
timestamp 1615077590
transform 1 0 -39 0 1 139
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_1
timestamp 1615077590
transform 1 0 161 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_3
timestamp 1615077590
transform 1 0 337 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_2
timestamp 1615077590
transform 1 0 249 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_1
timestamp 1615150785
transform 1 0 537 0 1 76
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_XSLFBL  XM7
timestamp 1624053917
transform 1 0 2372 0 1 538
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM6
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 1634 0 1 644
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM9
timestamp 1624053917
transform 1 0 3110 0 1 432
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM8
timestamp 1624053917
transform 1 0 2741 0 1 485
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM12
timestamp 1624053917
transform 1 0 4217 0 1 219
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM11
timestamp 1624053917
transform 1 0 3848 0 1 272
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM10
timestamp 1624053917
transform 1 0 3479 0 1 379
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_0
timestamp 1614978561
transform 1 0 -45 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_4
timestamp 1614978561
transform 1 0 -245 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_1
timestamp 1614978561
transform 1 0 161 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_2
timestamp 1614978561
transform 1 0 249 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_3
timestamp 1614978561
transform 1 0 337 0 1 533
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_L9ESED  XM2
timestamp 1624053917
transform 1 0 527 0 1 794
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM1
timestamp 1624053917
transform 1 0 158 0 1 847
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_5
timestamp 1614978561
transform 1 0 537 0 1 533
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_L9ESED  XM4
timestamp 1624053917
transform 1 0 1265 0 1 688
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM3
timestamp 1624053917
transform 1 0 896 0 1 741
box -211 -300 211 300
<< labels >>
rlabel metal1 -354 -124 646 -76 1 vss
rlabel nwell -354 745 646 821 1 vdd
rlabel metal2 31 293 103 365 1 out
rlabel metal1 570 210 625 276 1 in1
rlabel metal1 -342 318 -241 384 1 in2
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 in1
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 in2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 out
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
<< end >>
