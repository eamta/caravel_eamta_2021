magic
tech sky130A
magscale 1 2
timestamp 1622937437
<< error_p >>
rect -1085 1572 -1027 1578
rect -893 1572 -835 1578
rect -701 1572 -643 1578
rect -509 1572 -451 1578
rect -317 1572 -259 1578
rect -125 1572 -67 1578
rect 67 1572 125 1578
rect 259 1572 317 1578
rect 451 1572 509 1578
rect 643 1572 701 1578
rect 835 1572 893 1578
rect 1027 1572 1085 1578
rect -1085 1538 -1073 1572
rect -893 1538 -881 1572
rect -701 1538 -689 1572
rect -509 1538 -497 1572
rect -317 1538 -305 1572
rect -125 1538 -113 1572
rect 67 1538 79 1572
rect 259 1538 271 1572
rect 451 1538 463 1572
rect 643 1538 655 1572
rect 835 1538 847 1572
rect 1027 1538 1039 1572
rect -1085 1532 -1027 1538
rect -893 1532 -835 1538
rect -701 1532 -643 1538
rect -509 1532 -451 1538
rect -317 1532 -259 1538
rect -125 1532 -67 1538
rect 67 1532 125 1538
rect 259 1532 317 1538
rect 451 1532 509 1538
rect 643 1532 701 1538
rect 835 1532 893 1538
rect 1027 1532 1085 1538
rect -1181 -1538 -1123 -1532
rect -989 -1538 -931 -1532
rect -797 -1538 -739 -1532
rect -605 -1538 -547 -1532
rect -413 -1538 -355 -1532
rect -221 -1538 -163 -1532
rect -29 -1538 29 -1532
rect 163 -1538 221 -1532
rect 355 -1538 413 -1532
rect 547 -1538 605 -1532
rect 739 -1538 797 -1532
rect 931 -1538 989 -1532
rect 1123 -1538 1181 -1532
rect -1181 -1572 -1169 -1538
rect -989 -1572 -977 -1538
rect -797 -1572 -785 -1538
rect -605 -1572 -593 -1538
rect -413 -1572 -401 -1538
rect -221 -1572 -209 -1538
rect -29 -1572 -17 -1538
rect 163 -1572 175 -1538
rect 355 -1572 367 -1538
rect 547 -1572 559 -1538
rect 739 -1572 751 -1538
rect 931 -1572 943 -1538
rect 1123 -1572 1135 -1538
rect -1181 -1578 -1123 -1572
rect -989 -1578 -931 -1572
rect -797 -1578 -739 -1572
rect -605 -1578 -547 -1572
rect -413 -1578 -355 -1572
rect -221 -1578 -163 -1572
rect -29 -1578 29 -1572
rect 163 -1578 221 -1572
rect 355 -1578 413 -1572
rect 547 -1578 605 -1572
rect 739 -1578 797 -1572
rect 931 -1578 989 -1572
rect 1123 -1578 1181 -1572
<< pwell >>
rect -1367 -1710 1367 1710
<< nmoslvt >>
rect -1167 -1500 -1137 1500
rect -1071 -1500 -1041 1500
rect -975 -1500 -945 1500
rect -879 -1500 -849 1500
rect -783 -1500 -753 1500
rect -687 -1500 -657 1500
rect -591 -1500 -561 1500
rect -495 -1500 -465 1500
rect -399 -1500 -369 1500
rect -303 -1500 -273 1500
rect -207 -1500 -177 1500
rect -111 -1500 -81 1500
rect -15 -1500 15 1500
rect 81 -1500 111 1500
rect 177 -1500 207 1500
rect 273 -1500 303 1500
rect 369 -1500 399 1500
rect 465 -1500 495 1500
rect 561 -1500 591 1500
rect 657 -1500 687 1500
rect 753 -1500 783 1500
rect 849 -1500 879 1500
rect 945 -1500 975 1500
rect 1041 -1500 1071 1500
rect 1137 -1500 1167 1500
<< ndiff >>
rect -1229 1488 -1167 1500
rect -1229 -1488 -1217 1488
rect -1183 -1488 -1167 1488
rect -1229 -1500 -1167 -1488
rect -1137 1488 -1071 1500
rect -1137 -1488 -1121 1488
rect -1087 -1488 -1071 1488
rect -1137 -1500 -1071 -1488
rect -1041 1488 -975 1500
rect -1041 -1488 -1025 1488
rect -991 -1488 -975 1488
rect -1041 -1500 -975 -1488
rect -945 1488 -879 1500
rect -945 -1488 -929 1488
rect -895 -1488 -879 1488
rect -945 -1500 -879 -1488
rect -849 1488 -783 1500
rect -849 -1488 -833 1488
rect -799 -1488 -783 1488
rect -849 -1500 -783 -1488
rect -753 1488 -687 1500
rect -753 -1488 -737 1488
rect -703 -1488 -687 1488
rect -753 -1500 -687 -1488
rect -657 1488 -591 1500
rect -657 -1488 -641 1488
rect -607 -1488 -591 1488
rect -657 -1500 -591 -1488
rect -561 1488 -495 1500
rect -561 -1488 -545 1488
rect -511 -1488 -495 1488
rect -561 -1500 -495 -1488
rect -465 1488 -399 1500
rect -465 -1488 -449 1488
rect -415 -1488 -399 1488
rect -465 -1500 -399 -1488
rect -369 1488 -303 1500
rect -369 -1488 -353 1488
rect -319 -1488 -303 1488
rect -369 -1500 -303 -1488
rect -273 1488 -207 1500
rect -273 -1488 -257 1488
rect -223 -1488 -207 1488
rect -273 -1500 -207 -1488
rect -177 1488 -111 1500
rect -177 -1488 -161 1488
rect -127 -1488 -111 1488
rect -177 -1500 -111 -1488
rect -81 1488 -15 1500
rect -81 -1488 -65 1488
rect -31 -1488 -15 1488
rect -81 -1500 -15 -1488
rect 15 1488 81 1500
rect 15 -1488 31 1488
rect 65 -1488 81 1488
rect 15 -1500 81 -1488
rect 111 1488 177 1500
rect 111 -1488 127 1488
rect 161 -1488 177 1488
rect 111 -1500 177 -1488
rect 207 1488 273 1500
rect 207 -1488 223 1488
rect 257 -1488 273 1488
rect 207 -1500 273 -1488
rect 303 1488 369 1500
rect 303 -1488 319 1488
rect 353 -1488 369 1488
rect 303 -1500 369 -1488
rect 399 1488 465 1500
rect 399 -1488 415 1488
rect 449 -1488 465 1488
rect 399 -1500 465 -1488
rect 495 1488 561 1500
rect 495 -1488 511 1488
rect 545 -1488 561 1488
rect 495 -1500 561 -1488
rect 591 1488 657 1500
rect 591 -1488 607 1488
rect 641 -1488 657 1488
rect 591 -1500 657 -1488
rect 687 1488 753 1500
rect 687 -1488 703 1488
rect 737 -1488 753 1488
rect 687 -1500 753 -1488
rect 783 1488 849 1500
rect 783 -1488 799 1488
rect 833 -1488 849 1488
rect 783 -1500 849 -1488
rect 879 1488 945 1500
rect 879 -1488 895 1488
rect 929 -1488 945 1488
rect 879 -1500 945 -1488
rect 975 1488 1041 1500
rect 975 -1488 991 1488
rect 1025 -1488 1041 1488
rect 975 -1500 1041 -1488
rect 1071 1488 1137 1500
rect 1071 -1488 1087 1488
rect 1121 -1488 1137 1488
rect 1071 -1500 1137 -1488
rect 1167 1488 1229 1500
rect 1167 -1488 1183 1488
rect 1217 -1488 1229 1488
rect 1167 -1500 1229 -1488
<< ndiffc >>
rect -1217 -1488 -1183 1488
rect -1121 -1488 -1087 1488
rect -1025 -1488 -991 1488
rect -929 -1488 -895 1488
rect -833 -1488 -799 1488
rect -737 -1488 -703 1488
rect -641 -1488 -607 1488
rect -545 -1488 -511 1488
rect -449 -1488 -415 1488
rect -353 -1488 -319 1488
rect -257 -1488 -223 1488
rect -161 -1488 -127 1488
rect -65 -1488 -31 1488
rect 31 -1488 65 1488
rect 127 -1488 161 1488
rect 223 -1488 257 1488
rect 319 -1488 353 1488
rect 415 -1488 449 1488
rect 511 -1488 545 1488
rect 607 -1488 641 1488
rect 703 -1488 737 1488
rect 799 -1488 833 1488
rect 895 -1488 929 1488
rect 991 -1488 1025 1488
rect 1087 -1488 1121 1488
rect 1183 -1488 1217 1488
<< psubdiff >>
rect -1331 1640 -1235 1674
rect 1235 1640 1331 1674
rect -1331 1578 -1297 1640
rect 1297 1578 1331 1640
rect -1331 -1640 -1297 -1578
rect 1297 -1640 1331 -1578
rect -1331 -1674 -1235 -1640
rect 1235 -1674 1331 -1640
<< psubdiffcont >>
rect -1235 1640 1235 1674
rect -1331 -1578 -1297 1578
rect 1297 -1578 1331 1578
rect -1235 -1674 1235 -1640
<< poly >>
rect -1089 1572 -1023 1588
rect -1089 1538 -1073 1572
rect -1039 1538 -1023 1572
rect -1167 1500 -1137 1526
rect -1089 1522 -1023 1538
rect -897 1572 -831 1588
rect -897 1538 -881 1572
rect -847 1538 -831 1572
rect -1071 1500 -1041 1522
rect -975 1500 -945 1526
rect -897 1522 -831 1538
rect -705 1572 -639 1588
rect -705 1538 -689 1572
rect -655 1538 -639 1572
rect -879 1500 -849 1522
rect -783 1500 -753 1526
rect -705 1522 -639 1538
rect -513 1572 -447 1588
rect -513 1538 -497 1572
rect -463 1538 -447 1572
rect -687 1500 -657 1522
rect -591 1500 -561 1526
rect -513 1522 -447 1538
rect -321 1572 -255 1588
rect -321 1538 -305 1572
rect -271 1538 -255 1572
rect -495 1500 -465 1522
rect -399 1500 -369 1526
rect -321 1522 -255 1538
rect -129 1572 -63 1588
rect -129 1538 -113 1572
rect -79 1538 -63 1572
rect -303 1500 -273 1522
rect -207 1500 -177 1526
rect -129 1522 -63 1538
rect 63 1572 129 1588
rect 63 1538 79 1572
rect 113 1538 129 1572
rect -111 1500 -81 1522
rect -15 1500 15 1526
rect 63 1522 129 1538
rect 255 1572 321 1588
rect 255 1538 271 1572
rect 305 1538 321 1572
rect 81 1500 111 1522
rect 177 1500 207 1526
rect 255 1522 321 1538
rect 447 1572 513 1588
rect 447 1538 463 1572
rect 497 1538 513 1572
rect 273 1500 303 1522
rect 369 1500 399 1526
rect 447 1522 513 1538
rect 639 1572 705 1588
rect 639 1538 655 1572
rect 689 1538 705 1572
rect 465 1500 495 1522
rect 561 1500 591 1526
rect 639 1522 705 1538
rect 831 1572 897 1588
rect 831 1538 847 1572
rect 881 1538 897 1572
rect 657 1500 687 1522
rect 753 1500 783 1526
rect 831 1522 897 1538
rect 1023 1572 1089 1588
rect 1023 1538 1039 1572
rect 1073 1538 1089 1572
rect 849 1500 879 1522
rect 945 1500 975 1526
rect 1023 1522 1089 1538
rect 1041 1500 1071 1522
rect 1137 1500 1167 1526
rect -1167 -1522 -1137 -1500
rect -1185 -1538 -1119 -1522
rect -1071 -1526 -1041 -1500
rect -975 -1522 -945 -1500
rect -1185 -1572 -1169 -1538
rect -1135 -1572 -1119 -1538
rect -1185 -1588 -1119 -1572
rect -993 -1538 -927 -1522
rect -879 -1526 -849 -1500
rect -783 -1522 -753 -1500
rect -993 -1572 -977 -1538
rect -943 -1572 -927 -1538
rect -993 -1588 -927 -1572
rect -801 -1538 -735 -1522
rect -687 -1526 -657 -1500
rect -591 -1522 -561 -1500
rect -801 -1572 -785 -1538
rect -751 -1572 -735 -1538
rect -801 -1588 -735 -1572
rect -609 -1538 -543 -1522
rect -495 -1526 -465 -1500
rect -399 -1522 -369 -1500
rect -609 -1572 -593 -1538
rect -559 -1572 -543 -1538
rect -609 -1588 -543 -1572
rect -417 -1538 -351 -1522
rect -303 -1526 -273 -1500
rect -207 -1522 -177 -1500
rect -417 -1572 -401 -1538
rect -367 -1572 -351 -1538
rect -417 -1588 -351 -1572
rect -225 -1538 -159 -1522
rect -111 -1526 -81 -1500
rect -15 -1522 15 -1500
rect -225 -1572 -209 -1538
rect -175 -1572 -159 -1538
rect -225 -1588 -159 -1572
rect -33 -1538 33 -1522
rect 81 -1526 111 -1500
rect 177 -1522 207 -1500
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect -33 -1588 33 -1572
rect 159 -1538 225 -1522
rect 273 -1526 303 -1500
rect 369 -1522 399 -1500
rect 159 -1572 175 -1538
rect 209 -1572 225 -1538
rect 159 -1588 225 -1572
rect 351 -1538 417 -1522
rect 465 -1526 495 -1500
rect 561 -1522 591 -1500
rect 351 -1572 367 -1538
rect 401 -1572 417 -1538
rect 351 -1588 417 -1572
rect 543 -1538 609 -1522
rect 657 -1526 687 -1500
rect 753 -1522 783 -1500
rect 543 -1572 559 -1538
rect 593 -1572 609 -1538
rect 543 -1588 609 -1572
rect 735 -1538 801 -1522
rect 849 -1526 879 -1500
rect 945 -1522 975 -1500
rect 735 -1572 751 -1538
rect 785 -1572 801 -1538
rect 735 -1588 801 -1572
rect 927 -1538 993 -1522
rect 1041 -1526 1071 -1500
rect 1137 -1522 1167 -1500
rect 927 -1572 943 -1538
rect 977 -1572 993 -1538
rect 927 -1588 993 -1572
rect 1119 -1538 1185 -1522
rect 1119 -1572 1135 -1538
rect 1169 -1572 1185 -1538
rect 1119 -1588 1185 -1572
<< polycont >>
rect -1073 1538 -1039 1572
rect -881 1538 -847 1572
rect -689 1538 -655 1572
rect -497 1538 -463 1572
rect -305 1538 -271 1572
rect -113 1538 -79 1572
rect 79 1538 113 1572
rect 271 1538 305 1572
rect 463 1538 497 1572
rect 655 1538 689 1572
rect 847 1538 881 1572
rect 1039 1538 1073 1572
rect -1169 -1572 -1135 -1538
rect -977 -1572 -943 -1538
rect -785 -1572 -751 -1538
rect -593 -1572 -559 -1538
rect -401 -1572 -367 -1538
rect -209 -1572 -175 -1538
rect -17 -1572 17 -1538
rect 175 -1572 209 -1538
rect 367 -1572 401 -1538
rect 559 -1572 593 -1538
rect 751 -1572 785 -1538
rect 943 -1572 977 -1538
rect 1135 -1572 1169 -1538
<< locali >>
rect -1331 1640 -1235 1674
rect 1235 1640 1331 1674
rect -1331 1578 -1297 1640
rect 1297 1578 1331 1640
rect -1089 1538 -1073 1572
rect -1039 1538 -1023 1572
rect -897 1538 -881 1572
rect -847 1538 -831 1572
rect -705 1538 -689 1572
rect -655 1538 -639 1572
rect -513 1538 -497 1572
rect -463 1538 -447 1572
rect -321 1538 -305 1572
rect -271 1538 -255 1572
rect -129 1538 -113 1572
rect -79 1538 -63 1572
rect 63 1538 79 1572
rect 113 1538 129 1572
rect 255 1538 271 1572
rect 305 1538 321 1572
rect 447 1538 463 1572
rect 497 1538 513 1572
rect 639 1538 655 1572
rect 689 1538 705 1572
rect 831 1538 847 1572
rect 881 1538 897 1572
rect 1023 1538 1039 1572
rect 1073 1538 1089 1572
rect -1217 1488 -1183 1504
rect -1217 -1504 -1183 -1488
rect -1121 1488 -1087 1504
rect -1121 -1504 -1087 -1488
rect -1025 1488 -991 1504
rect -1025 -1504 -991 -1488
rect -929 1488 -895 1504
rect -929 -1504 -895 -1488
rect -833 1488 -799 1504
rect -833 -1504 -799 -1488
rect -737 1488 -703 1504
rect -737 -1504 -703 -1488
rect -641 1488 -607 1504
rect -641 -1504 -607 -1488
rect -545 1488 -511 1504
rect -545 -1504 -511 -1488
rect -449 1488 -415 1504
rect -449 -1504 -415 -1488
rect -353 1488 -319 1504
rect -353 -1504 -319 -1488
rect -257 1488 -223 1504
rect -257 -1504 -223 -1488
rect -161 1488 -127 1504
rect -161 -1504 -127 -1488
rect -65 1488 -31 1504
rect -65 -1504 -31 -1488
rect 31 1488 65 1504
rect 31 -1504 65 -1488
rect 127 1488 161 1504
rect 127 -1504 161 -1488
rect 223 1488 257 1504
rect 223 -1504 257 -1488
rect 319 1488 353 1504
rect 319 -1504 353 -1488
rect 415 1488 449 1504
rect 415 -1504 449 -1488
rect 511 1488 545 1504
rect 511 -1504 545 -1488
rect 607 1488 641 1504
rect 607 -1504 641 -1488
rect 703 1488 737 1504
rect 703 -1504 737 -1488
rect 799 1488 833 1504
rect 799 -1504 833 -1488
rect 895 1488 929 1504
rect 895 -1504 929 -1488
rect 991 1488 1025 1504
rect 991 -1504 1025 -1488
rect 1087 1488 1121 1504
rect 1087 -1504 1121 -1488
rect 1183 1488 1217 1504
rect 1183 -1504 1217 -1488
rect -1185 -1572 -1169 -1538
rect -1135 -1572 -1119 -1538
rect -993 -1572 -977 -1538
rect -943 -1572 -927 -1538
rect -801 -1572 -785 -1538
rect -751 -1572 -735 -1538
rect -609 -1572 -593 -1538
rect -559 -1572 -543 -1538
rect -417 -1572 -401 -1538
rect -367 -1572 -351 -1538
rect -225 -1572 -209 -1538
rect -175 -1572 -159 -1538
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect 159 -1572 175 -1538
rect 209 -1572 225 -1538
rect 351 -1572 367 -1538
rect 401 -1572 417 -1538
rect 543 -1572 559 -1538
rect 593 -1572 609 -1538
rect 735 -1572 751 -1538
rect 785 -1572 801 -1538
rect 927 -1572 943 -1538
rect 977 -1572 993 -1538
rect 1119 -1572 1135 -1538
rect 1169 -1572 1185 -1538
rect -1331 -1640 -1297 -1578
rect 1297 -1640 1331 -1578
rect -1331 -1674 -1235 -1640
rect 1235 -1674 1331 -1640
<< viali >>
rect -1073 1538 -1039 1572
rect -881 1538 -847 1572
rect -689 1538 -655 1572
rect -497 1538 -463 1572
rect -305 1538 -271 1572
rect -113 1538 -79 1572
rect 79 1538 113 1572
rect 271 1538 305 1572
rect 463 1538 497 1572
rect 655 1538 689 1572
rect 847 1538 881 1572
rect 1039 1538 1073 1572
rect -1217 -1488 -1183 1488
rect -1121 -1488 -1087 1488
rect -1025 -1488 -991 1488
rect -929 -1488 -895 1488
rect -833 -1488 -799 1488
rect -737 -1488 -703 1488
rect -641 -1488 -607 1488
rect -545 -1488 -511 1488
rect -449 -1488 -415 1488
rect -353 -1488 -319 1488
rect -257 -1488 -223 1488
rect -161 -1488 -127 1488
rect -65 -1488 -31 1488
rect 31 -1488 65 1488
rect 127 -1488 161 1488
rect 223 -1488 257 1488
rect 319 -1488 353 1488
rect 415 -1488 449 1488
rect 511 -1488 545 1488
rect 607 -1488 641 1488
rect 703 -1488 737 1488
rect 799 -1488 833 1488
rect 895 -1488 929 1488
rect 991 -1488 1025 1488
rect 1087 -1488 1121 1488
rect 1183 -1488 1217 1488
rect -1169 -1572 -1135 -1538
rect -977 -1572 -943 -1538
rect -785 -1572 -751 -1538
rect -593 -1572 -559 -1538
rect -401 -1572 -367 -1538
rect -209 -1572 -175 -1538
rect -17 -1572 17 -1538
rect 175 -1572 209 -1538
rect 367 -1572 401 -1538
rect 559 -1572 593 -1538
rect 751 -1572 785 -1538
rect 943 -1572 977 -1538
rect 1135 -1572 1169 -1538
<< metal1 >>
rect -1085 1572 -1027 1578
rect -1085 1538 -1073 1572
rect -1039 1538 -1027 1572
rect -1085 1532 -1027 1538
rect -893 1572 -835 1578
rect -893 1538 -881 1572
rect -847 1538 -835 1572
rect -893 1532 -835 1538
rect -701 1572 -643 1578
rect -701 1538 -689 1572
rect -655 1538 -643 1572
rect -701 1532 -643 1538
rect -509 1572 -451 1578
rect -509 1538 -497 1572
rect -463 1538 -451 1572
rect -509 1532 -451 1538
rect -317 1572 -259 1578
rect -317 1538 -305 1572
rect -271 1538 -259 1572
rect -317 1532 -259 1538
rect -125 1572 -67 1578
rect -125 1538 -113 1572
rect -79 1538 -67 1572
rect -125 1532 -67 1538
rect 67 1572 125 1578
rect 67 1538 79 1572
rect 113 1538 125 1572
rect 67 1532 125 1538
rect 259 1572 317 1578
rect 259 1538 271 1572
rect 305 1538 317 1572
rect 259 1532 317 1538
rect 451 1572 509 1578
rect 451 1538 463 1572
rect 497 1538 509 1572
rect 451 1532 509 1538
rect 643 1572 701 1578
rect 643 1538 655 1572
rect 689 1538 701 1572
rect 643 1532 701 1538
rect 835 1572 893 1578
rect 835 1538 847 1572
rect 881 1538 893 1572
rect 835 1532 893 1538
rect 1027 1572 1085 1578
rect 1027 1538 1039 1572
rect 1073 1538 1085 1572
rect 1027 1532 1085 1538
rect -1223 1488 -1177 1500
rect -1223 -1488 -1217 1488
rect -1183 -1488 -1177 1488
rect -1223 -1500 -1177 -1488
rect -1127 1488 -1081 1500
rect -1127 -1488 -1121 1488
rect -1087 -1488 -1081 1488
rect -1127 -1500 -1081 -1488
rect -1031 1488 -985 1500
rect -1031 -1488 -1025 1488
rect -991 -1488 -985 1488
rect -1031 -1500 -985 -1488
rect -935 1488 -889 1500
rect -935 -1488 -929 1488
rect -895 -1488 -889 1488
rect -935 -1500 -889 -1488
rect -839 1488 -793 1500
rect -839 -1488 -833 1488
rect -799 -1488 -793 1488
rect -839 -1500 -793 -1488
rect -743 1488 -697 1500
rect -743 -1488 -737 1488
rect -703 -1488 -697 1488
rect -743 -1500 -697 -1488
rect -647 1488 -601 1500
rect -647 -1488 -641 1488
rect -607 -1488 -601 1488
rect -647 -1500 -601 -1488
rect -551 1488 -505 1500
rect -551 -1488 -545 1488
rect -511 -1488 -505 1488
rect -551 -1500 -505 -1488
rect -455 1488 -409 1500
rect -455 -1488 -449 1488
rect -415 -1488 -409 1488
rect -455 -1500 -409 -1488
rect -359 1488 -313 1500
rect -359 -1488 -353 1488
rect -319 -1488 -313 1488
rect -359 -1500 -313 -1488
rect -263 1488 -217 1500
rect -263 -1488 -257 1488
rect -223 -1488 -217 1488
rect -263 -1500 -217 -1488
rect -167 1488 -121 1500
rect -167 -1488 -161 1488
rect -127 -1488 -121 1488
rect -167 -1500 -121 -1488
rect -71 1488 -25 1500
rect -71 -1488 -65 1488
rect -31 -1488 -25 1488
rect -71 -1500 -25 -1488
rect 25 1488 71 1500
rect 25 -1488 31 1488
rect 65 -1488 71 1488
rect 25 -1500 71 -1488
rect 121 1488 167 1500
rect 121 -1488 127 1488
rect 161 -1488 167 1488
rect 121 -1500 167 -1488
rect 217 1488 263 1500
rect 217 -1488 223 1488
rect 257 -1488 263 1488
rect 217 -1500 263 -1488
rect 313 1488 359 1500
rect 313 -1488 319 1488
rect 353 -1488 359 1488
rect 313 -1500 359 -1488
rect 409 1488 455 1500
rect 409 -1488 415 1488
rect 449 -1488 455 1488
rect 409 -1500 455 -1488
rect 505 1488 551 1500
rect 505 -1488 511 1488
rect 545 -1488 551 1488
rect 505 -1500 551 -1488
rect 601 1488 647 1500
rect 601 -1488 607 1488
rect 641 -1488 647 1488
rect 601 -1500 647 -1488
rect 697 1488 743 1500
rect 697 -1488 703 1488
rect 737 -1488 743 1488
rect 697 -1500 743 -1488
rect 793 1488 839 1500
rect 793 -1488 799 1488
rect 833 -1488 839 1488
rect 793 -1500 839 -1488
rect 889 1488 935 1500
rect 889 -1488 895 1488
rect 929 -1488 935 1488
rect 889 -1500 935 -1488
rect 985 1488 1031 1500
rect 985 -1488 991 1488
rect 1025 -1488 1031 1488
rect 985 -1500 1031 -1488
rect 1081 1488 1127 1500
rect 1081 -1488 1087 1488
rect 1121 -1488 1127 1488
rect 1081 -1500 1127 -1488
rect 1177 1488 1223 1500
rect 1177 -1488 1183 1488
rect 1217 -1488 1223 1488
rect 1177 -1500 1223 -1488
rect -1181 -1538 -1123 -1532
rect -1181 -1572 -1169 -1538
rect -1135 -1572 -1123 -1538
rect -1181 -1578 -1123 -1572
rect -989 -1538 -931 -1532
rect -989 -1572 -977 -1538
rect -943 -1572 -931 -1538
rect -989 -1578 -931 -1572
rect -797 -1538 -739 -1532
rect -797 -1572 -785 -1538
rect -751 -1572 -739 -1538
rect -797 -1578 -739 -1572
rect -605 -1538 -547 -1532
rect -605 -1572 -593 -1538
rect -559 -1572 -547 -1538
rect -605 -1578 -547 -1572
rect -413 -1538 -355 -1532
rect -413 -1572 -401 -1538
rect -367 -1572 -355 -1538
rect -413 -1578 -355 -1572
rect -221 -1538 -163 -1532
rect -221 -1572 -209 -1538
rect -175 -1572 -163 -1538
rect -221 -1578 -163 -1572
rect -29 -1538 29 -1532
rect -29 -1572 -17 -1538
rect 17 -1572 29 -1538
rect -29 -1578 29 -1572
rect 163 -1538 221 -1532
rect 163 -1572 175 -1538
rect 209 -1572 221 -1538
rect 163 -1578 221 -1572
rect 355 -1538 413 -1532
rect 355 -1572 367 -1538
rect 401 -1572 413 -1538
rect 355 -1578 413 -1572
rect 547 -1538 605 -1532
rect 547 -1572 559 -1538
rect 593 -1572 605 -1538
rect 547 -1578 605 -1572
rect 739 -1538 797 -1532
rect 739 -1572 751 -1538
rect 785 -1572 797 -1538
rect 739 -1578 797 -1572
rect 931 -1538 989 -1532
rect 931 -1572 943 -1538
rect 977 -1572 989 -1538
rect 931 -1578 989 -1572
rect 1123 -1538 1181 -1532
rect 1123 -1572 1135 -1538
rect 1169 -1572 1181 -1538
rect 1123 -1578 1181 -1572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1314 -1657 1314 1657
string parameters w 15 l 0.15 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
