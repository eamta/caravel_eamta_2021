magic
tech sky130A
magscale 1 2
timestamp 1615909117
<< error_p >>
rect -14720 -311 -14662 -305
rect -14602 -311 -14544 -305
rect -14484 -311 -14426 -305
rect -14366 -311 -14308 -305
rect -14248 -311 -14190 -305
rect -14130 -311 -14072 -305
rect -14012 -311 -13954 -305
rect -13894 -311 -13836 -305
rect -13776 -311 -13718 -305
rect -13658 -311 -13600 -305
rect -13540 -311 -13482 -305
rect -13422 -311 -13364 -305
rect -13304 -311 -13246 -305
rect -13186 -311 -13128 -305
rect -13068 -311 -13010 -305
rect -12950 -311 -12892 -305
rect -12832 -311 -12774 -305
rect -12714 -311 -12656 -305
rect -12596 -311 -12538 -305
rect -12478 -311 -12420 -305
rect -12360 -311 -12302 -305
rect -12242 -311 -12184 -305
rect -12124 -311 -12066 -305
rect -12006 -311 -11948 -305
rect -11888 -311 -11830 -305
rect -11770 -311 -11712 -305
rect -11652 -311 -11594 -305
rect -11534 -311 -11476 -305
rect -11416 -311 -11358 -305
rect -11298 -311 -11240 -305
rect -11180 -311 -11122 -305
rect -11062 -311 -11004 -305
rect -10944 -311 -10886 -305
rect -10826 -311 -10768 -305
rect -10708 -311 -10650 -305
rect -10590 -311 -10532 -305
rect -10472 -311 -10414 -305
rect -10354 -311 -10296 -305
rect -10236 -311 -10178 -305
rect -10118 -311 -10060 -305
rect -10000 -311 -9942 -305
rect -9882 -311 -9824 -305
rect -9764 -311 -9706 -305
rect -9646 -311 -9588 -305
rect -9528 -311 -9470 -305
rect -9410 -311 -9352 -305
rect -9292 -311 -9234 -305
rect -9174 -311 -9116 -305
rect -9056 -311 -8998 -305
rect -8938 -311 -8880 -305
rect -8820 -311 -8762 -305
rect -8702 -311 -8644 -305
rect -8584 -311 -8526 -305
rect -8466 -311 -8408 -305
rect -8348 -311 -8290 -305
rect -8230 -311 -8172 -305
rect -8112 -311 -8054 -305
rect -7994 -311 -7936 -305
rect -7876 -311 -7818 -305
rect -7758 -311 -7700 -305
rect -7640 -311 -7582 -305
rect -7522 -311 -7464 -305
rect -7404 -311 -7346 -305
rect -7286 -311 -7228 -305
rect -7168 -311 -7110 -305
rect -7050 -311 -6992 -305
rect -6932 -311 -6874 -305
rect -6814 -311 -6756 -305
rect -6696 -311 -6638 -305
rect -6578 -311 -6520 -305
rect -6460 -311 -6402 -305
rect -6342 -311 -6284 -305
rect -6224 -311 -6166 -305
rect -6106 -311 -6048 -305
rect -5988 -311 -5930 -305
rect -5870 -311 -5812 -305
rect -5752 -311 -5694 -305
rect -5634 -311 -5576 -305
rect -5516 -311 -5458 -305
rect -5398 -311 -5340 -305
rect -5280 -311 -5222 -305
rect -5162 -311 -5104 -305
rect -5044 -311 -4986 -305
rect -4926 -311 -4868 -305
rect -4808 -311 -4750 -305
rect -4690 -311 -4632 -305
rect -4572 -311 -4514 -305
rect -4454 -311 -4396 -305
rect -4336 -311 -4278 -305
rect -4218 -311 -4160 -305
rect -4100 -311 -4042 -305
rect -3982 -311 -3924 -305
rect -3864 -311 -3806 -305
rect -3746 -311 -3688 -305
rect -3628 -311 -3570 -305
rect -3510 -311 -3452 -305
rect -3392 -311 -3334 -305
rect -3274 -311 -3216 -305
rect -3156 -311 -3098 -305
rect -3038 -311 -2980 -305
rect -2920 -311 -2862 -305
rect -2802 -311 -2744 -305
rect -2684 -311 -2626 -305
rect -2566 -311 -2508 -305
rect -2448 -311 -2390 -305
rect -2330 -311 -2272 -305
rect -2212 -311 -2154 -305
rect -2094 -311 -2036 -305
rect -1976 -311 -1918 -305
rect -1858 -311 -1800 -305
rect -1740 -311 -1682 -305
rect -1622 -311 -1564 -305
rect -1504 -311 -1446 -305
rect -1386 -311 -1328 -305
rect -1268 -311 -1210 -305
rect -1150 -311 -1092 -305
rect -1032 -311 -974 -305
rect -914 -311 -856 -305
rect -796 -311 -738 -305
rect -678 -311 -620 -305
rect -560 -311 -502 -305
rect -442 -311 -384 -305
rect -324 -311 -266 -305
rect -206 -311 -148 -305
rect -88 -311 -30 -305
rect 30 -311 88 -305
rect 148 -311 206 -305
rect 266 -311 324 -305
rect 384 -311 442 -305
rect 502 -311 560 -305
rect 620 -311 678 -305
rect 738 -311 796 -305
rect 856 -311 914 -305
rect 974 -311 1032 -305
rect 1092 -311 1150 -305
rect 1210 -311 1268 -305
rect 1328 -311 1386 -305
rect 1446 -311 1504 -305
rect 1564 -311 1622 -305
rect 1682 -311 1740 -305
rect 1800 -311 1858 -305
rect 1918 -311 1976 -305
rect 2036 -311 2094 -305
rect 2154 -311 2212 -305
rect 2272 -311 2330 -305
rect 2390 -311 2448 -305
rect 2508 -311 2566 -305
rect 2626 -311 2684 -305
rect 2744 -311 2802 -305
rect 2862 -311 2920 -305
rect 2980 -311 3038 -305
rect 3098 -311 3156 -305
rect 3216 -311 3274 -305
rect 3334 -311 3392 -305
rect 3452 -311 3510 -305
rect 3570 -311 3628 -305
rect 3688 -311 3746 -305
rect 3806 -311 3864 -305
rect 3924 -311 3982 -305
rect 4042 -311 4100 -305
rect 4160 -311 4218 -305
rect 4278 -311 4336 -305
rect 4396 -311 4454 -305
rect 4514 -311 4572 -305
rect 4632 -311 4690 -305
rect 4750 -311 4808 -305
rect 4868 -311 4926 -305
rect 4986 -311 5044 -305
rect 5104 -311 5162 -305
rect 5222 -311 5280 -305
rect 5340 -311 5398 -305
rect 5458 -311 5516 -305
rect 5576 -311 5634 -305
rect 5694 -311 5752 -305
rect 5812 -311 5870 -305
rect 5930 -311 5988 -305
rect 6048 -311 6106 -305
rect 6166 -311 6224 -305
rect 6284 -311 6342 -305
rect 6402 -311 6460 -305
rect 6520 -311 6578 -305
rect 6638 -311 6696 -305
rect 6756 -311 6814 -305
rect 6874 -311 6932 -305
rect 6992 -311 7050 -305
rect 7110 -311 7168 -305
rect 7228 -311 7286 -305
rect 7346 -311 7404 -305
rect 7464 -311 7522 -305
rect 7582 -311 7640 -305
rect 7700 -311 7758 -305
rect 7818 -311 7876 -305
rect 7936 -311 7994 -305
rect 8054 -311 8112 -305
rect 8172 -311 8230 -305
rect 8290 -311 8348 -305
rect 8408 -311 8466 -305
rect 8526 -311 8584 -305
rect 8644 -311 8702 -305
rect 8762 -311 8820 -305
rect 8880 -311 8938 -305
rect 8998 -311 9056 -305
rect 9116 -311 9174 -305
rect 9234 -311 9292 -305
rect 9352 -311 9410 -305
rect 9470 -311 9528 -305
rect 9588 -311 9646 -305
rect 9706 -311 9764 -305
rect 9824 -311 9882 -305
rect 9942 -311 10000 -305
rect 10060 -311 10118 -305
rect 10178 -311 10236 -305
rect 10296 -311 10354 -305
rect 10414 -311 10472 -305
rect 10532 -311 10590 -305
rect 10650 -311 10708 -305
rect 10768 -311 10826 -305
rect 10886 -311 10944 -305
rect 11004 -311 11062 -305
rect 11122 -311 11180 -305
rect 11240 -311 11298 -305
rect 11358 -311 11416 -305
rect 11476 -311 11534 -305
rect 11594 -311 11652 -305
rect 11712 -311 11770 -305
rect 11830 -311 11888 -305
rect 11948 -311 12006 -305
rect 12066 -311 12124 -305
rect 12184 -311 12242 -305
rect 12302 -311 12360 -305
rect 12420 -311 12478 -305
rect 12538 -311 12596 -305
rect 12656 -311 12714 -305
rect 12774 -311 12832 -305
rect 12892 -311 12950 -305
rect 13010 -311 13068 -305
rect 13128 -311 13186 -305
rect 13246 -311 13304 -305
rect 13364 -311 13422 -305
rect 13482 -311 13540 -305
rect 13600 -311 13658 -305
rect 13718 -311 13776 -305
rect 13836 -311 13894 -305
rect 13954 -311 14012 -305
rect 14072 -311 14130 -305
rect 14190 -311 14248 -305
rect 14308 -311 14366 -305
rect 14426 -311 14484 -305
rect 14544 -311 14602 -305
rect 14662 -311 14720 -305
rect -14720 -345 -14708 -311
rect -14602 -345 -14590 -311
rect -14484 -345 -14472 -311
rect -14366 -345 -14354 -311
rect -14248 -345 -14236 -311
rect -14130 -345 -14118 -311
rect -14012 -345 -14000 -311
rect -13894 -345 -13882 -311
rect -13776 -345 -13764 -311
rect -13658 -345 -13646 -311
rect -13540 -345 -13528 -311
rect -13422 -345 -13410 -311
rect -13304 -345 -13292 -311
rect -13186 -345 -13174 -311
rect -13068 -345 -13056 -311
rect -12950 -345 -12938 -311
rect -12832 -345 -12820 -311
rect -12714 -345 -12702 -311
rect -12596 -345 -12584 -311
rect -12478 -345 -12466 -311
rect -12360 -345 -12348 -311
rect -12242 -345 -12230 -311
rect -12124 -345 -12112 -311
rect -12006 -345 -11994 -311
rect -11888 -345 -11876 -311
rect -11770 -345 -11758 -311
rect -11652 -345 -11640 -311
rect -11534 -345 -11522 -311
rect -11416 -345 -11404 -311
rect -11298 -345 -11286 -311
rect -11180 -345 -11168 -311
rect -11062 -345 -11050 -311
rect -10944 -345 -10932 -311
rect -10826 -345 -10814 -311
rect -10708 -345 -10696 -311
rect -10590 -345 -10578 -311
rect -10472 -345 -10460 -311
rect -10354 -345 -10342 -311
rect -10236 -345 -10224 -311
rect -10118 -345 -10106 -311
rect -10000 -345 -9988 -311
rect -9882 -345 -9870 -311
rect -9764 -345 -9752 -311
rect -9646 -345 -9634 -311
rect -9528 -345 -9516 -311
rect -9410 -345 -9398 -311
rect -9292 -345 -9280 -311
rect -9174 -345 -9162 -311
rect -9056 -345 -9044 -311
rect -8938 -345 -8926 -311
rect -8820 -345 -8808 -311
rect -8702 -345 -8690 -311
rect -8584 -345 -8572 -311
rect -8466 -345 -8454 -311
rect -8348 -345 -8336 -311
rect -8230 -345 -8218 -311
rect -8112 -345 -8100 -311
rect -7994 -345 -7982 -311
rect -7876 -345 -7864 -311
rect -7758 -345 -7746 -311
rect -7640 -345 -7628 -311
rect -7522 -345 -7510 -311
rect -7404 -345 -7392 -311
rect -7286 -345 -7274 -311
rect -7168 -345 -7156 -311
rect -7050 -345 -7038 -311
rect -6932 -345 -6920 -311
rect -6814 -345 -6802 -311
rect -6696 -345 -6684 -311
rect -6578 -345 -6566 -311
rect -6460 -345 -6448 -311
rect -6342 -345 -6330 -311
rect -6224 -345 -6212 -311
rect -6106 -345 -6094 -311
rect -5988 -345 -5976 -311
rect -5870 -345 -5858 -311
rect -5752 -345 -5740 -311
rect -5634 -345 -5622 -311
rect -5516 -345 -5504 -311
rect -5398 -345 -5386 -311
rect -5280 -345 -5268 -311
rect -5162 -345 -5150 -311
rect -5044 -345 -5032 -311
rect -4926 -345 -4914 -311
rect -4808 -345 -4796 -311
rect -4690 -345 -4678 -311
rect -4572 -345 -4560 -311
rect -4454 -345 -4442 -311
rect -4336 -345 -4324 -311
rect -4218 -345 -4206 -311
rect -4100 -345 -4088 -311
rect -3982 -345 -3970 -311
rect -3864 -345 -3852 -311
rect -3746 -345 -3734 -311
rect -3628 -345 -3616 -311
rect -3510 -345 -3498 -311
rect -3392 -345 -3380 -311
rect -3274 -345 -3262 -311
rect -3156 -345 -3144 -311
rect -3038 -345 -3026 -311
rect -2920 -345 -2908 -311
rect -2802 -345 -2790 -311
rect -2684 -345 -2672 -311
rect -2566 -345 -2554 -311
rect -2448 -345 -2436 -311
rect -2330 -345 -2318 -311
rect -2212 -345 -2200 -311
rect -2094 -345 -2082 -311
rect -1976 -345 -1964 -311
rect -1858 -345 -1846 -311
rect -1740 -345 -1728 -311
rect -1622 -345 -1610 -311
rect -1504 -345 -1492 -311
rect -1386 -345 -1374 -311
rect -1268 -345 -1256 -311
rect -1150 -345 -1138 -311
rect -1032 -345 -1020 -311
rect -914 -345 -902 -311
rect -796 -345 -784 -311
rect -678 -345 -666 -311
rect -560 -345 -548 -311
rect -442 -345 -430 -311
rect -324 -345 -312 -311
rect -206 -345 -194 -311
rect -88 -345 -76 -311
rect 30 -345 42 -311
rect 148 -345 160 -311
rect 266 -345 278 -311
rect 384 -345 396 -311
rect 502 -345 514 -311
rect 620 -345 632 -311
rect 738 -345 750 -311
rect 856 -345 868 -311
rect 974 -345 986 -311
rect 1092 -345 1104 -311
rect 1210 -345 1222 -311
rect 1328 -345 1340 -311
rect 1446 -345 1458 -311
rect 1564 -345 1576 -311
rect 1682 -345 1694 -311
rect 1800 -345 1812 -311
rect 1918 -345 1930 -311
rect 2036 -345 2048 -311
rect 2154 -345 2166 -311
rect 2272 -345 2284 -311
rect 2390 -345 2402 -311
rect 2508 -345 2520 -311
rect 2626 -345 2638 -311
rect 2744 -345 2756 -311
rect 2862 -345 2874 -311
rect 2980 -345 2992 -311
rect 3098 -345 3110 -311
rect 3216 -345 3228 -311
rect 3334 -345 3346 -311
rect 3452 -345 3464 -311
rect 3570 -345 3582 -311
rect 3688 -345 3700 -311
rect 3806 -345 3818 -311
rect 3924 -345 3936 -311
rect 4042 -345 4054 -311
rect 4160 -345 4172 -311
rect 4278 -345 4290 -311
rect 4396 -345 4408 -311
rect 4514 -345 4526 -311
rect 4632 -345 4644 -311
rect 4750 -345 4762 -311
rect 4868 -345 4880 -311
rect 4986 -345 4998 -311
rect 5104 -345 5116 -311
rect 5222 -345 5234 -311
rect 5340 -345 5352 -311
rect 5458 -345 5470 -311
rect 5576 -345 5588 -311
rect 5694 -345 5706 -311
rect 5812 -345 5824 -311
rect 5930 -345 5942 -311
rect 6048 -345 6060 -311
rect 6166 -345 6178 -311
rect 6284 -345 6296 -311
rect 6402 -345 6414 -311
rect 6520 -345 6532 -311
rect 6638 -345 6650 -311
rect 6756 -345 6768 -311
rect 6874 -345 6886 -311
rect 6992 -345 7004 -311
rect 7110 -345 7122 -311
rect 7228 -345 7240 -311
rect 7346 -345 7358 -311
rect 7464 -345 7476 -311
rect 7582 -345 7594 -311
rect 7700 -345 7712 -311
rect 7818 -345 7830 -311
rect 7936 -345 7948 -311
rect 8054 -345 8066 -311
rect 8172 -345 8184 -311
rect 8290 -345 8302 -311
rect 8408 -345 8420 -311
rect 8526 -345 8538 -311
rect 8644 -345 8656 -311
rect 8762 -345 8774 -311
rect 8880 -345 8892 -311
rect 8998 -345 9010 -311
rect 9116 -345 9128 -311
rect 9234 -345 9246 -311
rect 9352 -345 9364 -311
rect 9470 -345 9482 -311
rect 9588 -345 9600 -311
rect 9706 -345 9718 -311
rect 9824 -345 9836 -311
rect 9942 -345 9954 -311
rect 10060 -345 10072 -311
rect 10178 -345 10190 -311
rect 10296 -345 10308 -311
rect 10414 -345 10426 -311
rect 10532 -345 10544 -311
rect 10650 -345 10662 -311
rect 10768 -345 10780 -311
rect 10886 -345 10898 -311
rect 11004 -345 11016 -311
rect 11122 -345 11134 -311
rect 11240 -345 11252 -311
rect 11358 -345 11370 -311
rect 11476 -345 11488 -311
rect 11594 -345 11606 -311
rect 11712 -345 11724 -311
rect 11830 -345 11842 -311
rect 11948 -345 11960 -311
rect 12066 -345 12078 -311
rect 12184 -345 12196 -311
rect 12302 -345 12314 -311
rect 12420 -345 12432 -311
rect 12538 -345 12550 -311
rect 12656 -345 12668 -311
rect 12774 -345 12786 -311
rect 12892 -345 12904 -311
rect 13010 -345 13022 -311
rect 13128 -345 13140 -311
rect 13246 -345 13258 -311
rect 13364 -345 13376 -311
rect 13482 -345 13494 -311
rect 13600 -345 13612 -311
rect 13718 -345 13730 -311
rect 13836 -345 13848 -311
rect 13954 -345 13966 -311
rect 14072 -345 14084 -311
rect 14190 -345 14202 -311
rect 14308 -345 14320 -311
rect 14426 -345 14438 -311
rect 14544 -345 14556 -311
rect 14662 -345 14674 -311
rect -14720 -351 -14662 -345
rect -14602 -351 -14544 -345
rect -14484 -351 -14426 -345
rect -14366 -351 -14308 -345
rect -14248 -351 -14190 -345
rect -14130 -351 -14072 -345
rect -14012 -351 -13954 -345
rect -13894 -351 -13836 -345
rect -13776 -351 -13718 -345
rect -13658 -351 -13600 -345
rect -13540 -351 -13482 -345
rect -13422 -351 -13364 -345
rect -13304 -351 -13246 -345
rect -13186 -351 -13128 -345
rect -13068 -351 -13010 -345
rect -12950 -351 -12892 -345
rect -12832 -351 -12774 -345
rect -12714 -351 -12656 -345
rect -12596 -351 -12538 -345
rect -12478 -351 -12420 -345
rect -12360 -351 -12302 -345
rect -12242 -351 -12184 -345
rect -12124 -351 -12066 -345
rect -12006 -351 -11948 -345
rect -11888 -351 -11830 -345
rect -11770 -351 -11712 -345
rect -11652 -351 -11594 -345
rect -11534 -351 -11476 -345
rect -11416 -351 -11358 -345
rect -11298 -351 -11240 -345
rect -11180 -351 -11122 -345
rect -11062 -351 -11004 -345
rect -10944 -351 -10886 -345
rect -10826 -351 -10768 -345
rect -10708 -351 -10650 -345
rect -10590 -351 -10532 -345
rect -10472 -351 -10414 -345
rect -10354 -351 -10296 -345
rect -10236 -351 -10178 -345
rect -10118 -351 -10060 -345
rect -10000 -351 -9942 -345
rect -9882 -351 -9824 -345
rect -9764 -351 -9706 -345
rect -9646 -351 -9588 -345
rect -9528 -351 -9470 -345
rect -9410 -351 -9352 -345
rect -9292 -351 -9234 -345
rect -9174 -351 -9116 -345
rect -9056 -351 -8998 -345
rect -8938 -351 -8880 -345
rect -8820 -351 -8762 -345
rect -8702 -351 -8644 -345
rect -8584 -351 -8526 -345
rect -8466 -351 -8408 -345
rect -8348 -351 -8290 -345
rect -8230 -351 -8172 -345
rect -8112 -351 -8054 -345
rect -7994 -351 -7936 -345
rect -7876 -351 -7818 -345
rect -7758 -351 -7700 -345
rect -7640 -351 -7582 -345
rect -7522 -351 -7464 -345
rect -7404 -351 -7346 -345
rect -7286 -351 -7228 -345
rect -7168 -351 -7110 -345
rect -7050 -351 -6992 -345
rect -6932 -351 -6874 -345
rect -6814 -351 -6756 -345
rect -6696 -351 -6638 -345
rect -6578 -351 -6520 -345
rect -6460 -351 -6402 -345
rect -6342 -351 -6284 -345
rect -6224 -351 -6166 -345
rect -6106 -351 -6048 -345
rect -5988 -351 -5930 -345
rect -5870 -351 -5812 -345
rect -5752 -351 -5694 -345
rect -5634 -351 -5576 -345
rect -5516 -351 -5458 -345
rect -5398 -351 -5340 -345
rect -5280 -351 -5222 -345
rect -5162 -351 -5104 -345
rect -5044 -351 -4986 -345
rect -4926 -351 -4868 -345
rect -4808 -351 -4750 -345
rect -4690 -351 -4632 -345
rect -4572 -351 -4514 -345
rect -4454 -351 -4396 -345
rect -4336 -351 -4278 -345
rect -4218 -351 -4160 -345
rect -4100 -351 -4042 -345
rect -3982 -351 -3924 -345
rect -3864 -351 -3806 -345
rect -3746 -351 -3688 -345
rect -3628 -351 -3570 -345
rect -3510 -351 -3452 -345
rect -3392 -351 -3334 -345
rect -3274 -351 -3216 -345
rect -3156 -351 -3098 -345
rect -3038 -351 -2980 -345
rect -2920 -351 -2862 -345
rect -2802 -351 -2744 -345
rect -2684 -351 -2626 -345
rect -2566 -351 -2508 -345
rect -2448 -351 -2390 -345
rect -2330 -351 -2272 -345
rect -2212 -351 -2154 -345
rect -2094 -351 -2036 -345
rect -1976 -351 -1918 -345
rect -1858 -351 -1800 -345
rect -1740 -351 -1682 -345
rect -1622 -351 -1564 -345
rect -1504 -351 -1446 -345
rect -1386 -351 -1328 -345
rect -1268 -351 -1210 -345
rect -1150 -351 -1092 -345
rect -1032 -351 -974 -345
rect -914 -351 -856 -345
rect -796 -351 -738 -345
rect -678 -351 -620 -345
rect -560 -351 -502 -345
rect -442 -351 -384 -345
rect -324 -351 -266 -345
rect -206 -351 -148 -345
rect -88 -351 -30 -345
rect 30 -351 88 -345
rect 148 -351 206 -345
rect 266 -351 324 -345
rect 384 -351 442 -345
rect 502 -351 560 -345
rect 620 -351 678 -345
rect 738 -351 796 -345
rect 856 -351 914 -345
rect 974 -351 1032 -345
rect 1092 -351 1150 -345
rect 1210 -351 1268 -345
rect 1328 -351 1386 -345
rect 1446 -351 1504 -345
rect 1564 -351 1622 -345
rect 1682 -351 1740 -345
rect 1800 -351 1858 -345
rect 1918 -351 1976 -345
rect 2036 -351 2094 -345
rect 2154 -351 2212 -345
rect 2272 -351 2330 -345
rect 2390 -351 2448 -345
rect 2508 -351 2566 -345
rect 2626 -351 2684 -345
rect 2744 -351 2802 -345
rect 2862 -351 2920 -345
rect 2980 -351 3038 -345
rect 3098 -351 3156 -345
rect 3216 -351 3274 -345
rect 3334 -351 3392 -345
rect 3452 -351 3510 -345
rect 3570 -351 3628 -345
rect 3688 -351 3746 -345
rect 3806 -351 3864 -345
rect 3924 -351 3982 -345
rect 4042 -351 4100 -345
rect 4160 -351 4218 -345
rect 4278 -351 4336 -345
rect 4396 -351 4454 -345
rect 4514 -351 4572 -345
rect 4632 -351 4690 -345
rect 4750 -351 4808 -345
rect 4868 -351 4926 -345
rect 4986 -351 5044 -345
rect 5104 -351 5162 -345
rect 5222 -351 5280 -345
rect 5340 -351 5398 -345
rect 5458 -351 5516 -345
rect 5576 -351 5634 -345
rect 5694 -351 5752 -345
rect 5812 -351 5870 -345
rect 5930 -351 5988 -345
rect 6048 -351 6106 -345
rect 6166 -351 6224 -345
rect 6284 -351 6342 -345
rect 6402 -351 6460 -345
rect 6520 -351 6578 -345
rect 6638 -351 6696 -345
rect 6756 -351 6814 -345
rect 6874 -351 6932 -345
rect 6992 -351 7050 -345
rect 7110 -351 7168 -345
rect 7228 -351 7286 -345
rect 7346 -351 7404 -345
rect 7464 -351 7522 -345
rect 7582 -351 7640 -345
rect 7700 -351 7758 -345
rect 7818 -351 7876 -345
rect 7936 -351 7994 -345
rect 8054 -351 8112 -345
rect 8172 -351 8230 -345
rect 8290 -351 8348 -345
rect 8408 -351 8466 -345
rect 8526 -351 8584 -345
rect 8644 -351 8702 -345
rect 8762 -351 8820 -345
rect 8880 -351 8938 -345
rect 8998 -351 9056 -345
rect 9116 -351 9174 -345
rect 9234 -351 9292 -345
rect 9352 -351 9410 -345
rect 9470 -351 9528 -345
rect 9588 -351 9646 -345
rect 9706 -351 9764 -345
rect 9824 -351 9882 -345
rect 9942 -351 10000 -345
rect 10060 -351 10118 -345
rect 10178 -351 10236 -345
rect 10296 -351 10354 -345
rect 10414 -351 10472 -345
rect 10532 -351 10590 -345
rect 10650 -351 10708 -345
rect 10768 -351 10826 -345
rect 10886 -351 10944 -345
rect 11004 -351 11062 -345
rect 11122 -351 11180 -345
rect 11240 -351 11298 -345
rect 11358 -351 11416 -345
rect 11476 -351 11534 -345
rect 11594 -351 11652 -345
rect 11712 -351 11770 -345
rect 11830 -351 11888 -345
rect 11948 -351 12006 -345
rect 12066 -351 12124 -345
rect 12184 -351 12242 -345
rect 12302 -351 12360 -345
rect 12420 -351 12478 -345
rect 12538 -351 12596 -345
rect 12656 -351 12714 -345
rect 12774 -351 12832 -345
rect 12892 -351 12950 -345
rect 13010 -351 13068 -345
rect 13128 -351 13186 -345
rect 13246 -351 13304 -345
rect 13364 -351 13422 -345
rect 13482 -351 13540 -345
rect 13600 -351 13658 -345
rect 13718 -351 13776 -345
rect 13836 -351 13894 -345
rect 13954 -351 14012 -345
rect 14072 -351 14130 -345
rect 14190 -351 14248 -345
rect 14308 -351 14366 -345
rect 14426 -351 14484 -345
rect 14544 -351 14602 -345
rect 14662 -351 14720 -345
<< nwell >>
rect -14917 -484 14917 484
<< pmos >>
rect -14721 -264 -14661 336
rect -14603 -264 -14543 336
rect -14485 -264 -14425 336
rect -14367 -264 -14307 336
rect -14249 -264 -14189 336
rect -14131 -264 -14071 336
rect -14013 -264 -13953 336
rect -13895 -264 -13835 336
rect -13777 -264 -13717 336
rect -13659 -264 -13599 336
rect -13541 -264 -13481 336
rect -13423 -264 -13363 336
rect -13305 -264 -13245 336
rect -13187 -264 -13127 336
rect -13069 -264 -13009 336
rect -12951 -264 -12891 336
rect -12833 -264 -12773 336
rect -12715 -264 -12655 336
rect -12597 -264 -12537 336
rect -12479 -264 -12419 336
rect -12361 -264 -12301 336
rect -12243 -264 -12183 336
rect -12125 -264 -12065 336
rect -12007 -264 -11947 336
rect -11889 -264 -11829 336
rect -11771 -264 -11711 336
rect -11653 -264 -11593 336
rect -11535 -264 -11475 336
rect -11417 -264 -11357 336
rect -11299 -264 -11239 336
rect -11181 -264 -11121 336
rect -11063 -264 -11003 336
rect -10945 -264 -10885 336
rect -10827 -264 -10767 336
rect -10709 -264 -10649 336
rect -10591 -264 -10531 336
rect -10473 -264 -10413 336
rect -10355 -264 -10295 336
rect -10237 -264 -10177 336
rect -10119 -264 -10059 336
rect -10001 -264 -9941 336
rect -9883 -264 -9823 336
rect -9765 -264 -9705 336
rect -9647 -264 -9587 336
rect -9529 -264 -9469 336
rect -9411 -264 -9351 336
rect -9293 -264 -9233 336
rect -9175 -264 -9115 336
rect -9057 -264 -8997 336
rect -8939 -264 -8879 336
rect -8821 -264 -8761 336
rect -8703 -264 -8643 336
rect -8585 -264 -8525 336
rect -8467 -264 -8407 336
rect -8349 -264 -8289 336
rect -8231 -264 -8171 336
rect -8113 -264 -8053 336
rect -7995 -264 -7935 336
rect -7877 -264 -7817 336
rect -7759 -264 -7699 336
rect -7641 -264 -7581 336
rect -7523 -264 -7463 336
rect -7405 -264 -7345 336
rect -7287 -264 -7227 336
rect -7169 -264 -7109 336
rect -7051 -264 -6991 336
rect -6933 -264 -6873 336
rect -6815 -264 -6755 336
rect -6697 -264 -6637 336
rect -6579 -264 -6519 336
rect -6461 -264 -6401 336
rect -6343 -264 -6283 336
rect -6225 -264 -6165 336
rect -6107 -264 -6047 336
rect -5989 -264 -5929 336
rect -5871 -264 -5811 336
rect -5753 -264 -5693 336
rect -5635 -264 -5575 336
rect -5517 -264 -5457 336
rect -5399 -264 -5339 336
rect -5281 -264 -5221 336
rect -5163 -264 -5103 336
rect -5045 -264 -4985 336
rect -4927 -264 -4867 336
rect -4809 -264 -4749 336
rect -4691 -264 -4631 336
rect -4573 -264 -4513 336
rect -4455 -264 -4395 336
rect -4337 -264 -4277 336
rect -4219 -264 -4159 336
rect -4101 -264 -4041 336
rect -3983 -264 -3923 336
rect -3865 -264 -3805 336
rect -3747 -264 -3687 336
rect -3629 -264 -3569 336
rect -3511 -264 -3451 336
rect -3393 -264 -3333 336
rect -3275 -264 -3215 336
rect -3157 -264 -3097 336
rect -3039 -264 -2979 336
rect -2921 -264 -2861 336
rect -2803 -264 -2743 336
rect -2685 -264 -2625 336
rect -2567 -264 -2507 336
rect -2449 -264 -2389 336
rect -2331 -264 -2271 336
rect -2213 -264 -2153 336
rect -2095 -264 -2035 336
rect -1977 -264 -1917 336
rect -1859 -264 -1799 336
rect -1741 -264 -1681 336
rect -1623 -264 -1563 336
rect -1505 -264 -1445 336
rect -1387 -264 -1327 336
rect -1269 -264 -1209 336
rect -1151 -264 -1091 336
rect -1033 -264 -973 336
rect -915 -264 -855 336
rect -797 -264 -737 336
rect -679 -264 -619 336
rect -561 -264 -501 336
rect -443 -264 -383 336
rect -325 -264 -265 336
rect -207 -264 -147 336
rect -89 -264 -29 336
rect 29 -264 89 336
rect 147 -264 207 336
rect 265 -264 325 336
rect 383 -264 443 336
rect 501 -264 561 336
rect 619 -264 679 336
rect 737 -264 797 336
rect 855 -264 915 336
rect 973 -264 1033 336
rect 1091 -264 1151 336
rect 1209 -264 1269 336
rect 1327 -264 1387 336
rect 1445 -264 1505 336
rect 1563 -264 1623 336
rect 1681 -264 1741 336
rect 1799 -264 1859 336
rect 1917 -264 1977 336
rect 2035 -264 2095 336
rect 2153 -264 2213 336
rect 2271 -264 2331 336
rect 2389 -264 2449 336
rect 2507 -264 2567 336
rect 2625 -264 2685 336
rect 2743 -264 2803 336
rect 2861 -264 2921 336
rect 2979 -264 3039 336
rect 3097 -264 3157 336
rect 3215 -264 3275 336
rect 3333 -264 3393 336
rect 3451 -264 3511 336
rect 3569 -264 3629 336
rect 3687 -264 3747 336
rect 3805 -264 3865 336
rect 3923 -264 3983 336
rect 4041 -264 4101 336
rect 4159 -264 4219 336
rect 4277 -264 4337 336
rect 4395 -264 4455 336
rect 4513 -264 4573 336
rect 4631 -264 4691 336
rect 4749 -264 4809 336
rect 4867 -264 4927 336
rect 4985 -264 5045 336
rect 5103 -264 5163 336
rect 5221 -264 5281 336
rect 5339 -264 5399 336
rect 5457 -264 5517 336
rect 5575 -264 5635 336
rect 5693 -264 5753 336
rect 5811 -264 5871 336
rect 5929 -264 5989 336
rect 6047 -264 6107 336
rect 6165 -264 6225 336
rect 6283 -264 6343 336
rect 6401 -264 6461 336
rect 6519 -264 6579 336
rect 6637 -264 6697 336
rect 6755 -264 6815 336
rect 6873 -264 6933 336
rect 6991 -264 7051 336
rect 7109 -264 7169 336
rect 7227 -264 7287 336
rect 7345 -264 7405 336
rect 7463 -264 7523 336
rect 7581 -264 7641 336
rect 7699 -264 7759 336
rect 7817 -264 7877 336
rect 7935 -264 7995 336
rect 8053 -264 8113 336
rect 8171 -264 8231 336
rect 8289 -264 8349 336
rect 8407 -264 8467 336
rect 8525 -264 8585 336
rect 8643 -264 8703 336
rect 8761 -264 8821 336
rect 8879 -264 8939 336
rect 8997 -264 9057 336
rect 9115 -264 9175 336
rect 9233 -264 9293 336
rect 9351 -264 9411 336
rect 9469 -264 9529 336
rect 9587 -264 9647 336
rect 9705 -264 9765 336
rect 9823 -264 9883 336
rect 9941 -264 10001 336
rect 10059 -264 10119 336
rect 10177 -264 10237 336
rect 10295 -264 10355 336
rect 10413 -264 10473 336
rect 10531 -264 10591 336
rect 10649 -264 10709 336
rect 10767 -264 10827 336
rect 10885 -264 10945 336
rect 11003 -264 11063 336
rect 11121 -264 11181 336
rect 11239 -264 11299 336
rect 11357 -264 11417 336
rect 11475 -264 11535 336
rect 11593 -264 11653 336
rect 11711 -264 11771 336
rect 11829 -264 11889 336
rect 11947 -264 12007 336
rect 12065 -264 12125 336
rect 12183 -264 12243 336
rect 12301 -264 12361 336
rect 12419 -264 12479 336
rect 12537 -264 12597 336
rect 12655 -264 12715 336
rect 12773 -264 12833 336
rect 12891 -264 12951 336
rect 13009 -264 13069 336
rect 13127 -264 13187 336
rect 13245 -264 13305 336
rect 13363 -264 13423 336
rect 13481 -264 13541 336
rect 13599 -264 13659 336
rect 13717 -264 13777 336
rect 13835 -264 13895 336
rect 13953 -264 14013 336
rect 14071 -264 14131 336
rect 14189 -264 14249 336
rect 14307 -264 14367 336
rect 14425 -264 14485 336
rect 14543 -264 14603 336
rect 14661 -264 14721 336
<< pdiff >>
rect -14779 324 -14721 336
rect -14779 -252 -14767 324
rect -14733 -252 -14721 324
rect -14779 -264 -14721 -252
rect -14661 324 -14603 336
rect -14661 -252 -14649 324
rect -14615 -252 -14603 324
rect -14661 -264 -14603 -252
rect -14543 324 -14485 336
rect -14543 -252 -14531 324
rect -14497 -252 -14485 324
rect -14543 -264 -14485 -252
rect -14425 324 -14367 336
rect -14425 -252 -14413 324
rect -14379 -252 -14367 324
rect -14425 -264 -14367 -252
rect -14307 324 -14249 336
rect -14307 -252 -14295 324
rect -14261 -252 -14249 324
rect -14307 -264 -14249 -252
rect -14189 324 -14131 336
rect -14189 -252 -14177 324
rect -14143 -252 -14131 324
rect -14189 -264 -14131 -252
rect -14071 324 -14013 336
rect -14071 -252 -14059 324
rect -14025 -252 -14013 324
rect -14071 -264 -14013 -252
rect -13953 324 -13895 336
rect -13953 -252 -13941 324
rect -13907 -252 -13895 324
rect -13953 -264 -13895 -252
rect -13835 324 -13777 336
rect -13835 -252 -13823 324
rect -13789 -252 -13777 324
rect -13835 -264 -13777 -252
rect -13717 324 -13659 336
rect -13717 -252 -13705 324
rect -13671 -252 -13659 324
rect -13717 -264 -13659 -252
rect -13599 324 -13541 336
rect -13599 -252 -13587 324
rect -13553 -252 -13541 324
rect -13599 -264 -13541 -252
rect -13481 324 -13423 336
rect -13481 -252 -13469 324
rect -13435 -252 -13423 324
rect -13481 -264 -13423 -252
rect -13363 324 -13305 336
rect -13363 -252 -13351 324
rect -13317 -252 -13305 324
rect -13363 -264 -13305 -252
rect -13245 324 -13187 336
rect -13245 -252 -13233 324
rect -13199 -252 -13187 324
rect -13245 -264 -13187 -252
rect -13127 324 -13069 336
rect -13127 -252 -13115 324
rect -13081 -252 -13069 324
rect -13127 -264 -13069 -252
rect -13009 324 -12951 336
rect -13009 -252 -12997 324
rect -12963 -252 -12951 324
rect -13009 -264 -12951 -252
rect -12891 324 -12833 336
rect -12891 -252 -12879 324
rect -12845 -252 -12833 324
rect -12891 -264 -12833 -252
rect -12773 324 -12715 336
rect -12773 -252 -12761 324
rect -12727 -252 -12715 324
rect -12773 -264 -12715 -252
rect -12655 324 -12597 336
rect -12655 -252 -12643 324
rect -12609 -252 -12597 324
rect -12655 -264 -12597 -252
rect -12537 324 -12479 336
rect -12537 -252 -12525 324
rect -12491 -252 -12479 324
rect -12537 -264 -12479 -252
rect -12419 324 -12361 336
rect -12419 -252 -12407 324
rect -12373 -252 -12361 324
rect -12419 -264 -12361 -252
rect -12301 324 -12243 336
rect -12301 -252 -12289 324
rect -12255 -252 -12243 324
rect -12301 -264 -12243 -252
rect -12183 324 -12125 336
rect -12183 -252 -12171 324
rect -12137 -252 -12125 324
rect -12183 -264 -12125 -252
rect -12065 324 -12007 336
rect -12065 -252 -12053 324
rect -12019 -252 -12007 324
rect -12065 -264 -12007 -252
rect -11947 324 -11889 336
rect -11947 -252 -11935 324
rect -11901 -252 -11889 324
rect -11947 -264 -11889 -252
rect -11829 324 -11771 336
rect -11829 -252 -11817 324
rect -11783 -252 -11771 324
rect -11829 -264 -11771 -252
rect -11711 324 -11653 336
rect -11711 -252 -11699 324
rect -11665 -252 -11653 324
rect -11711 -264 -11653 -252
rect -11593 324 -11535 336
rect -11593 -252 -11581 324
rect -11547 -252 -11535 324
rect -11593 -264 -11535 -252
rect -11475 324 -11417 336
rect -11475 -252 -11463 324
rect -11429 -252 -11417 324
rect -11475 -264 -11417 -252
rect -11357 324 -11299 336
rect -11357 -252 -11345 324
rect -11311 -252 -11299 324
rect -11357 -264 -11299 -252
rect -11239 324 -11181 336
rect -11239 -252 -11227 324
rect -11193 -252 -11181 324
rect -11239 -264 -11181 -252
rect -11121 324 -11063 336
rect -11121 -252 -11109 324
rect -11075 -252 -11063 324
rect -11121 -264 -11063 -252
rect -11003 324 -10945 336
rect -11003 -252 -10991 324
rect -10957 -252 -10945 324
rect -11003 -264 -10945 -252
rect -10885 324 -10827 336
rect -10885 -252 -10873 324
rect -10839 -252 -10827 324
rect -10885 -264 -10827 -252
rect -10767 324 -10709 336
rect -10767 -252 -10755 324
rect -10721 -252 -10709 324
rect -10767 -264 -10709 -252
rect -10649 324 -10591 336
rect -10649 -252 -10637 324
rect -10603 -252 -10591 324
rect -10649 -264 -10591 -252
rect -10531 324 -10473 336
rect -10531 -252 -10519 324
rect -10485 -252 -10473 324
rect -10531 -264 -10473 -252
rect -10413 324 -10355 336
rect -10413 -252 -10401 324
rect -10367 -252 -10355 324
rect -10413 -264 -10355 -252
rect -10295 324 -10237 336
rect -10295 -252 -10283 324
rect -10249 -252 -10237 324
rect -10295 -264 -10237 -252
rect -10177 324 -10119 336
rect -10177 -252 -10165 324
rect -10131 -252 -10119 324
rect -10177 -264 -10119 -252
rect -10059 324 -10001 336
rect -10059 -252 -10047 324
rect -10013 -252 -10001 324
rect -10059 -264 -10001 -252
rect -9941 324 -9883 336
rect -9941 -252 -9929 324
rect -9895 -252 -9883 324
rect -9941 -264 -9883 -252
rect -9823 324 -9765 336
rect -9823 -252 -9811 324
rect -9777 -252 -9765 324
rect -9823 -264 -9765 -252
rect -9705 324 -9647 336
rect -9705 -252 -9693 324
rect -9659 -252 -9647 324
rect -9705 -264 -9647 -252
rect -9587 324 -9529 336
rect -9587 -252 -9575 324
rect -9541 -252 -9529 324
rect -9587 -264 -9529 -252
rect -9469 324 -9411 336
rect -9469 -252 -9457 324
rect -9423 -252 -9411 324
rect -9469 -264 -9411 -252
rect -9351 324 -9293 336
rect -9351 -252 -9339 324
rect -9305 -252 -9293 324
rect -9351 -264 -9293 -252
rect -9233 324 -9175 336
rect -9233 -252 -9221 324
rect -9187 -252 -9175 324
rect -9233 -264 -9175 -252
rect -9115 324 -9057 336
rect -9115 -252 -9103 324
rect -9069 -252 -9057 324
rect -9115 -264 -9057 -252
rect -8997 324 -8939 336
rect -8997 -252 -8985 324
rect -8951 -252 -8939 324
rect -8997 -264 -8939 -252
rect -8879 324 -8821 336
rect -8879 -252 -8867 324
rect -8833 -252 -8821 324
rect -8879 -264 -8821 -252
rect -8761 324 -8703 336
rect -8761 -252 -8749 324
rect -8715 -252 -8703 324
rect -8761 -264 -8703 -252
rect -8643 324 -8585 336
rect -8643 -252 -8631 324
rect -8597 -252 -8585 324
rect -8643 -264 -8585 -252
rect -8525 324 -8467 336
rect -8525 -252 -8513 324
rect -8479 -252 -8467 324
rect -8525 -264 -8467 -252
rect -8407 324 -8349 336
rect -8407 -252 -8395 324
rect -8361 -252 -8349 324
rect -8407 -264 -8349 -252
rect -8289 324 -8231 336
rect -8289 -252 -8277 324
rect -8243 -252 -8231 324
rect -8289 -264 -8231 -252
rect -8171 324 -8113 336
rect -8171 -252 -8159 324
rect -8125 -252 -8113 324
rect -8171 -264 -8113 -252
rect -8053 324 -7995 336
rect -8053 -252 -8041 324
rect -8007 -252 -7995 324
rect -8053 -264 -7995 -252
rect -7935 324 -7877 336
rect -7935 -252 -7923 324
rect -7889 -252 -7877 324
rect -7935 -264 -7877 -252
rect -7817 324 -7759 336
rect -7817 -252 -7805 324
rect -7771 -252 -7759 324
rect -7817 -264 -7759 -252
rect -7699 324 -7641 336
rect -7699 -252 -7687 324
rect -7653 -252 -7641 324
rect -7699 -264 -7641 -252
rect -7581 324 -7523 336
rect -7581 -252 -7569 324
rect -7535 -252 -7523 324
rect -7581 -264 -7523 -252
rect -7463 324 -7405 336
rect -7463 -252 -7451 324
rect -7417 -252 -7405 324
rect -7463 -264 -7405 -252
rect -7345 324 -7287 336
rect -7345 -252 -7333 324
rect -7299 -252 -7287 324
rect -7345 -264 -7287 -252
rect -7227 324 -7169 336
rect -7227 -252 -7215 324
rect -7181 -252 -7169 324
rect -7227 -264 -7169 -252
rect -7109 324 -7051 336
rect -7109 -252 -7097 324
rect -7063 -252 -7051 324
rect -7109 -264 -7051 -252
rect -6991 324 -6933 336
rect -6991 -252 -6979 324
rect -6945 -252 -6933 324
rect -6991 -264 -6933 -252
rect -6873 324 -6815 336
rect -6873 -252 -6861 324
rect -6827 -252 -6815 324
rect -6873 -264 -6815 -252
rect -6755 324 -6697 336
rect -6755 -252 -6743 324
rect -6709 -252 -6697 324
rect -6755 -264 -6697 -252
rect -6637 324 -6579 336
rect -6637 -252 -6625 324
rect -6591 -252 -6579 324
rect -6637 -264 -6579 -252
rect -6519 324 -6461 336
rect -6519 -252 -6507 324
rect -6473 -252 -6461 324
rect -6519 -264 -6461 -252
rect -6401 324 -6343 336
rect -6401 -252 -6389 324
rect -6355 -252 -6343 324
rect -6401 -264 -6343 -252
rect -6283 324 -6225 336
rect -6283 -252 -6271 324
rect -6237 -252 -6225 324
rect -6283 -264 -6225 -252
rect -6165 324 -6107 336
rect -6165 -252 -6153 324
rect -6119 -252 -6107 324
rect -6165 -264 -6107 -252
rect -6047 324 -5989 336
rect -6047 -252 -6035 324
rect -6001 -252 -5989 324
rect -6047 -264 -5989 -252
rect -5929 324 -5871 336
rect -5929 -252 -5917 324
rect -5883 -252 -5871 324
rect -5929 -264 -5871 -252
rect -5811 324 -5753 336
rect -5811 -252 -5799 324
rect -5765 -252 -5753 324
rect -5811 -264 -5753 -252
rect -5693 324 -5635 336
rect -5693 -252 -5681 324
rect -5647 -252 -5635 324
rect -5693 -264 -5635 -252
rect -5575 324 -5517 336
rect -5575 -252 -5563 324
rect -5529 -252 -5517 324
rect -5575 -264 -5517 -252
rect -5457 324 -5399 336
rect -5457 -252 -5445 324
rect -5411 -252 -5399 324
rect -5457 -264 -5399 -252
rect -5339 324 -5281 336
rect -5339 -252 -5327 324
rect -5293 -252 -5281 324
rect -5339 -264 -5281 -252
rect -5221 324 -5163 336
rect -5221 -252 -5209 324
rect -5175 -252 -5163 324
rect -5221 -264 -5163 -252
rect -5103 324 -5045 336
rect -5103 -252 -5091 324
rect -5057 -252 -5045 324
rect -5103 -264 -5045 -252
rect -4985 324 -4927 336
rect -4985 -252 -4973 324
rect -4939 -252 -4927 324
rect -4985 -264 -4927 -252
rect -4867 324 -4809 336
rect -4867 -252 -4855 324
rect -4821 -252 -4809 324
rect -4867 -264 -4809 -252
rect -4749 324 -4691 336
rect -4749 -252 -4737 324
rect -4703 -252 -4691 324
rect -4749 -264 -4691 -252
rect -4631 324 -4573 336
rect -4631 -252 -4619 324
rect -4585 -252 -4573 324
rect -4631 -264 -4573 -252
rect -4513 324 -4455 336
rect -4513 -252 -4501 324
rect -4467 -252 -4455 324
rect -4513 -264 -4455 -252
rect -4395 324 -4337 336
rect -4395 -252 -4383 324
rect -4349 -252 -4337 324
rect -4395 -264 -4337 -252
rect -4277 324 -4219 336
rect -4277 -252 -4265 324
rect -4231 -252 -4219 324
rect -4277 -264 -4219 -252
rect -4159 324 -4101 336
rect -4159 -252 -4147 324
rect -4113 -252 -4101 324
rect -4159 -264 -4101 -252
rect -4041 324 -3983 336
rect -4041 -252 -4029 324
rect -3995 -252 -3983 324
rect -4041 -264 -3983 -252
rect -3923 324 -3865 336
rect -3923 -252 -3911 324
rect -3877 -252 -3865 324
rect -3923 -264 -3865 -252
rect -3805 324 -3747 336
rect -3805 -252 -3793 324
rect -3759 -252 -3747 324
rect -3805 -264 -3747 -252
rect -3687 324 -3629 336
rect -3687 -252 -3675 324
rect -3641 -252 -3629 324
rect -3687 -264 -3629 -252
rect -3569 324 -3511 336
rect -3569 -252 -3557 324
rect -3523 -252 -3511 324
rect -3569 -264 -3511 -252
rect -3451 324 -3393 336
rect -3451 -252 -3439 324
rect -3405 -252 -3393 324
rect -3451 -264 -3393 -252
rect -3333 324 -3275 336
rect -3333 -252 -3321 324
rect -3287 -252 -3275 324
rect -3333 -264 -3275 -252
rect -3215 324 -3157 336
rect -3215 -252 -3203 324
rect -3169 -252 -3157 324
rect -3215 -264 -3157 -252
rect -3097 324 -3039 336
rect -3097 -252 -3085 324
rect -3051 -252 -3039 324
rect -3097 -264 -3039 -252
rect -2979 324 -2921 336
rect -2979 -252 -2967 324
rect -2933 -252 -2921 324
rect -2979 -264 -2921 -252
rect -2861 324 -2803 336
rect -2861 -252 -2849 324
rect -2815 -252 -2803 324
rect -2861 -264 -2803 -252
rect -2743 324 -2685 336
rect -2743 -252 -2731 324
rect -2697 -252 -2685 324
rect -2743 -264 -2685 -252
rect -2625 324 -2567 336
rect -2625 -252 -2613 324
rect -2579 -252 -2567 324
rect -2625 -264 -2567 -252
rect -2507 324 -2449 336
rect -2507 -252 -2495 324
rect -2461 -252 -2449 324
rect -2507 -264 -2449 -252
rect -2389 324 -2331 336
rect -2389 -252 -2377 324
rect -2343 -252 -2331 324
rect -2389 -264 -2331 -252
rect -2271 324 -2213 336
rect -2271 -252 -2259 324
rect -2225 -252 -2213 324
rect -2271 -264 -2213 -252
rect -2153 324 -2095 336
rect -2153 -252 -2141 324
rect -2107 -252 -2095 324
rect -2153 -264 -2095 -252
rect -2035 324 -1977 336
rect -2035 -252 -2023 324
rect -1989 -252 -1977 324
rect -2035 -264 -1977 -252
rect -1917 324 -1859 336
rect -1917 -252 -1905 324
rect -1871 -252 -1859 324
rect -1917 -264 -1859 -252
rect -1799 324 -1741 336
rect -1799 -252 -1787 324
rect -1753 -252 -1741 324
rect -1799 -264 -1741 -252
rect -1681 324 -1623 336
rect -1681 -252 -1669 324
rect -1635 -252 -1623 324
rect -1681 -264 -1623 -252
rect -1563 324 -1505 336
rect -1563 -252 -1551 324
rect -1517 -252 -1505 324
rect -1563 -264 -1505 -252
rect -1445 324 -1387 336
rect -1445 -252 -1433 324
rect -1399 -252 -1387 324
rect -1445 -264 -1387 -252
rect -1327 324 -1269 336
rect -1327 -252 -1315 324
rect -1281 -252 -1269 324
rect -1327 -264 -1269 -252
rect -1209 324 -1151 336
rect -1209 -252 -1197 324
rect -1163 -252 -1151 324
rect -1209 -264 -1151 -252
rect -1091 324 -1033 336
rect -1091 -252 -1079 324
rect -1045 -252 -1033 324
rect -1091 -264 -1033 -252
rect -973 324 -915 336
rect -973 -252 -961 324
rect -927 -252 -915 324
rect -973 -264 -915 -252
rect -855 324 -797 336
rect -855 -252 -843 324
rect -809 -252 -797 324
rect -855 -264 -797 -252
rect -737 324 -679 336
rect -737 -252 -725 324
rect -691 -252 -679 324
rect -737 -264 -679 -252
rect -619 324 -561 336
rect -619 -252 -607 324
rect -573 -252 -561 324
rect -619 -264 -561 -252
rect -501 324 -443 336
rect -501 -252 -489 324
rect -455 -252 -443 324
rect -501 -264 -443 -252
rect -383 324 -325 336
rect -383 -252 -371 324
rect -337 -252 -325 324
rect -383 -264 -325 -252
rect -265 324 -207 336
rect -265 -252 -253 324
rect -219 -252 -207 324
rect -265 -264 -207 -252
rect -147 324 -89 336
rect -147 -252 -135 324
rect -101 -252 -89 324
rect -147 -264 -89 -252
rect -29 324 29 336
rect -29 -252 -17 324
rect 17 -252 29 324
rect -29 -264 29 -252
rect 89 324 147 336
rect 89 -252 101 324
rect 135 -252 147 324
rect 89 -264 147 -252
rect 207 324 265 336
rect 207 -252 219 324
rect 253 -252 265 324
rect 207 -264 265 -252
rect 325 324 383 336
rect 325 -252 337 324
rect 371 -252 383 324
rect 325 -264 383 -252
rect 443 324 501 336
rect 443 -252 455 324
rect 489 -252 501 324
rect 443 -264 501 -252
rect 561 324 619 336
rect 561 -252 573 324
rect 607 -252 619 324
rect 561 -264 619 -252
rect 679 324 737 336
rect 679 -252 691 324
rect 725 -252 737 324
rect 679 -264 737 -252
rect 797 324 855 336
rect 797 -252 809 324
rect 843 -252 855 324
rect 797 -264 855 -252
rect 915 324 973 336
rect 915 -252 927 324
rect 961 -252 973 324
rect 915 -264 973 -252
rect 1033 324 1091 336
rect 1033 -252 1045 324
rect 1079 -252 1091 324
rect 1033 -264 1091 -252
rect 1151 324 1209 336
rect 1151 -252 1163 324
rect 1197 -252 1209 324
rect 1151 -264 1209 -252
rect 1269 324 1327 336
rect 1269 -252 1281 324
rect 1315 -252 1327 324
rect 1269 -264 1327 -252
rect 1387 324 1445 336
rect 1387 -252 1399 324
rect 1433 -252 1445 324
rect 1387 -264 1445 -252
rect 1505 324 1563 336
rect 1505 -252 1517 324
rect 1551 -252 1563 324
rect 1505 -264 1563 -252
rect 1623 324 1681 336
rect 1623 -252 1635 324
rect 1669 -252 1681 324
rect 1623 -264 1681 -252
rect 1741 324 1799 336
rect 1741 -252 1753 324
rect 1787 -252 1799 324
rect 1741 -264 1799 -252
rect 1859 324 1917 336
rect 1859 -252 1871 324
rect 1905 -252 1917 324
rect 1859 -264 1917 -252
rect 1977 324 2035 336
rect 1977 -252 1989 324
rect 2023 -252 2035 324
rect 1977 -264 2035 -252
rect 2095 324 2153 336
rect 2095 -252 2107 324
rect 2141 -252 2153 324
rect 2095 -264 2153 -252
rect 2213 324 2271 336
rect 2213 -252 2225 324
rect 2259 -252 2271 324
rect 2213 -264 2271 -252
rect 2331 324 2389 336
rect 2331 -252 2343 324
rect 2377 -252 2389 324
rect 2331 -264 2389 -252
rect 2449 324 2507 336
rect 2449 -252 2461 324
rect 2495 -252 2507 324
rect 2449 -264 2507 -252
rect 2567 324 2625 336
rect 2567 -252 2579 324
rect 2613 -252 2625 324
rect 2567 -264 2625 -252
rect 2685 324 2743 336
rect 2685 -252 2697 324
rect 2731 -252 2743 324
rect 2685 -264 2743 -252
rect 2803 324 2861 336
rect 2803 -252 2815 324
rect 2849 -252 2861 324
rect 2803 -264 2861 -252
rect 2921 324 2979 336
rect 2921 -252 2933 324
rect 2967 -252 2979 324
rect 2921 -264 2979 -252
rect 3039 324 3097 336
rect 3039 -252 3051 324
rect 3085 -252 3097 324
rect 3039 -264 3097 -252
rect 3157 324 3215 336
rect 3157 -252 3169 324
rect 3203 -252 3215 324
rect 3157 -264 3215 -252
rect 3275 324 3333 336
rect 3275 -252 3287 324
rect 3321 -252 3333 324
rect 3275 -264 3333 -252
rect 3393 324 3451 336
rect 3393 -252 3405 324
rect 3439 -252 3451 324
rect 3393 -264 3451 -252
rect 3511 324 3569 336
rect 3511 -252 3523 324
rect 3557 -252 3569 324
rect 3511 -264 3569 -252
rect 3629 324 3687 336
rect 3629 -252 3641 324
rect 3675 -252 3687 324
rect 3629 -264 3687 -252
rect 3747 324 3805 336
rect 3747 -252 3759 324
rect 3793 -252 3805 324
rect 3747 -264 3805 -252
rect 3865 324 3923 336
rect 3865 -252 3877 324
rect 3911 -252 3923 324
rect 3865 -264 3923 -252
rect 3983 324 4041 336
rect 3983 -252 3995 324
rect 4029 -252 4041 324
rect 3983 -264 4041 -252
rect 4101 324 4159 336
rect 4101 -252 4113 324
rect 4147 -252 4159 324
rect 4101 -264 4159 -252
rect 4219 324 4277 336
rect 4219 -252 4231 324
rect 4265 -252 4277 324
rect 4219 -264 4277 -252
rect 4337 324 4395 336
rect 4337 -252 4349 324
rect 4383 -252 4395 324
rect 4337 -264 4395 -252
rect 4455 324 4513 336
rect 4455 -252 4467 324
rect 4501 -252 4513 324
rect 4455 -264 4513 -252
rect 4573 324 4631 336
rect 4573 -252 4585 324
rect 4619 -252 4631 324
rect 4573 -264 4631 -252
rect 4691 324 4749 336
rect 4691 -252 4703 324
rect 4737 -252 4749 324
rect 4691 -264 4749 -252
rect 4809 324 4867 336
rect 4809 -252 4821 324
rect 4855 -252 4867 324
rect 4809 -264 4867 -252
rect 4927 324 4985 336
rect 4927 -252 4939 324
rect 4973 -252 4985 324
rect 4927 -264 4985 -252
rect 5045 324 5103 336
rect 5045 -252 5057 324
rect 5091 -252 5103 324
rect 5045 -264 5103 -252
rect 5163 324 5221 336
rect 5163 -252 5175 324
rect 5209 -252 5221 324
rect 5163 -264 5221 -252
rect 5281 324 5339 336
rect 5281 -252 5293 324
rect 5327 -252 5339 324
rect 5281 -264 5339 -252
rect 5399 324 5457 336
rect 5399 -252 5411 324
rect 5445 -252 5457 324
rect 5399 -264 5457 -252
rect 5517 324 5575 336
rect 5517 -252 5529 324
rect 5563 -252 5575 324
rect 5517 -264 5575 -252
rect 5635 324 5693 336
rect 5635 -252 5647 324
rect 5681 -252 5693 324
rect 5635 -264 5693 -252
rect 5753 324 5811 336
rect 5753 -252 5765 324
rect 5799 -252 5811 324
rect 5753 -264 5811 -252
rect 5871 324 5929 336
rect 5871 -252 5883 324
rect 5917 -252 5929 324
rect 5871 -264 5929 -252
rect 5989 324 6047 336
rect 5989 -252 6001 324
rect 6035 -252 6047 324
rect 5989 -264 6047 -252
rect 6107 324 6165 336
rect 6107 -252 6119 324
rect 6153 -252 6165 324
rect 6107 -264 6165 -252
rect 6225 324 6283 336
rect 6225 -252 6237 324
rect 6271 -252 6283 324
rect 6225 -264 6283 -252
rect 6343 324 6401 336
rect 6343 -252 6355 324
rect 6389 -252 6401 324
rect 6343 -264 6401 -252
rect 6461 324 6519 336
rect 6461 -252 6473 324
rect 6507 -252 6519 324
rect 6461 -264 6519 -252
rect 6579 324 6637 336
rect 6579 -252 6591 324
rect 6625 -252 6637 324
rect 6579 -264 6637 -252
rect 6697 324 6755 336
rect 6697 -252 6709 324
rect 6743 -252 6755 324
rect 6697 -264 6755 -252
rect 6815 324 6873 336
rect 6815 -252 6827 324
rect 6861 -252 6873 324
rect 6815 -264 6873 -252
rect 6933 324 6991 336
rect 6933 -252 6945 324
rect 6979 -252 6991 324
rect 6933 -264 6991 -252
rect 7051 324 7109 336
rect 7051 -252 7063 324
rect 7097 -252 7109 324
rect 7051 -264 7109 -252
rect 7169 324 7227 336
rect 7169 -252 7181 324
rect 7215 -252 7227 324
rect 7169 -264 7227 -252
rect 7287 324 7345 336
rect 7287 -252 7299 324
rect 7333 -252 7345 324
rect 7287 -264 7345 -252
rect 7405 324 7463 336
rect 7405 -252 7417 324
rect 7451 -252 7463 324
rect 7405 -264 7463 -252
rect 7523 324 7581 336
rect 7523 -252 7535 324
rect 7569 -252 7581 324
rect 7523 -264 7581 -252
rect 7641 324 7699 336
rect 7641 -252 7653 324
rect 7687 -252 7699 324
rect 7641 -264 7699 -252
rect 7759 324 7817 336
rect 7759 -252 7771 324
rect 7805 -252 7817 324
rect 7759 -264 7817 -252
rect 7877 324 7935 336
rect 7877 -252 7889 324
rect 7923 -252 7935 324
rect 7877 -264 7935 -252
rect 7995 324 8053 336
rect 7995 -252 8007 324
rect 8041 -252 8053 324
rect 7995 -264 8053 -252
rect 8113 324 8171 336
rect 8113 -252 8125 324
rect 8159 -252 8171 324
rect 8113 -264 8171 -252
rect 8231 324 8289 336
rect 8231 -252 8243 324
rect 8277 -252 8289 324
rect 8231 -264 8289 -252
rect 8349 324 8407 336
rect 8349 -252 8361 324
rect 8395 -252 8407 324
rect 8349 -264 8407 -252
rect 8467 324 8525 336
rect 8467 -252 8479 324
rect 8513 -252 8525 324
rect 8467 -264 8525 -252
rect 8585 324 8643 336
rect 8585 -252 8597 324
rect 8631 -252 8643 324
rect 8585 -264 8643 -252
rect 8703 324 8761 336
rect 8703 -252 8715 324
rect 8749 -252 8761 324
rect 8703 -264 8761 -252
rect 8821 324 8879 336
rect 8821 -252 8833 324
rect 8867 -252 8879 324
rect 8821 -264 8879 -252
rect 8939 324 8997 336
rect 8939 -252 8951 324
rect 8985 -252 8997 324
rect 8939 -264 8997 -252
rect 9057 324 9115 336
rect 9057 -252 9069 324
rect 9103 -252 9115 324
rect 9057 -264 9115 -252
rect 9175 324 9233 336
rect 9175 -252 9187 324
rect 9221 -252 9233 324
rect 9175 -264 9233 -252
rect 9293 324 9351 336
rect 9293 -252 9305 324
rect 9339 -252 9351 324
rect 9293 -264 9351 -252
rect 9411 324 9469 336
rect 9411 -252 9423 324
rect 9457 -252 9469 324
rect 9411 -264 9469 -252
rect 9529 324 9587 336
rect 9529 -252 9541 324
rect 9575 -252 9587 324
rect 9529 -264 9587 -252
rect 9647 324 9705 336
rect 9647 -252 9659 324
rect 9693 -252 9705 324
rect 9647 -264 9705 -252
rect 9765 324 9823 336
rect 9765 -252 9777 324
rect 9811 -252 9823 324
rect 9765 -264 9823 -252
rect 9883 324 9941 336
rect 9883 -252 9895 324
rect 9929 -252 9941 324
rect 9883 -264 9941 -252
rect 10001 324 10059 336
rect 10001 -252 10013 324
rect 10047 -252 10059 324
rect 10001 -264 10059 -252
rect 10119 324 10177 336
rect 10119 -252 10131 324
rect 10165 -252 10177 324
rect 10119 -264 10177 -252
rect 10237 324 10295 336
rect 10237 -252 10249 324
rect 10283 -252 10295 324
rect 10237 -264 10295 -252
rect 10355 324 10413 336
rect 10355 -252 10367 324
rect 10401 -252 10413 324
rect 10355 -264 10413 -252
rect 10473 324 10531 336
rect 10473 -252 10485 324
rect 10519 -252 10531 324
rect 10473 -264 10531 -252
rect 10591 324 10649 336
rect 10591 -252 10603 324
rect 10637 -252 10649 324
rect 10591 -264 10649 -252
rect 10709 324 10767 336
rect 10709 -252 10721 324
rect 10755 -252 10767 324
rect 10709 -264 10767 -252
rect 10827 324 10885 336
rect 10827 -252 10839 324
rect 10873 -252 10885 324
rect 10827 -264 10885 -252
rect 10945 324 11003 336
rect 10945 -252 10957 324
rect 10991 -252 11003 324
rect 10945 -264 11003 -252
rect 11063 324 11121 336
rect 11063 -252 11075 324
rect 11109 -252 11121 324
rect 11063 -264 11121 -252
rect 11181 324 11239 336
rect 11181 -252 11193 324
rect 11227 -252 11239 324
rect 11181 -264 11239 -252
rect 11299 324 11357 336
rect 11299 -252 11311 324
rect 11345 -252 11357 324
rect 11299 -264 11357 -252
rect 11417 324 11475 336
rect 11417 -252 11429 324
rect 11463 -252 11475 324
rect 11417 -264 11475 -252
rect 11535 324 11593 336
rect 11535 -252 11547 324
rect 11581 -252 11593 324
rect 11535 -264 11593 -252
rect 11653 324 11711 336
rect 11653 -252 11665 324
rect 11699 -252 11711 324
rect 11653 -264 11711 -252
rect 11771 324 11829 336
rect 11771 -252 11783 324
rect 11817 -252 11829 324
rect 11771 -264 11829 -252
rect 11889 324 11947 336
rect 11889 -252 11901 324
rect 11935 -252 11947 324
rect 11889 -264 11947 -252
rect 12007 324 12065 336
rect 12007 -252 12019 324
rect 12053 -252 12065 324
rect 12007 -264 12065 -252
rect 12125 324 12183 336
rect 12125 -252 12137 324
rect 12171 -252 12183 324
rect 12125 -264 12183 -252
rect 12243 324 12301 336
rect 12243 -252 12255 324
rect 12289 -252 12301 324
rect 12243 -264 12301 -252
rect 12361 324 12419 336
rect 12361 -252 12373 324
rect 12407 -252 12419 324
rect 12361 -264 12419 -252
rect 12479 324 12537 336
rect 12479 -252 12491 324
rect 12525 -252 12537 324
rect 12479 -264 12537 -252
rect 12597 324 12655 336
rect 12597 -252 12609 324
rect 12643 -252 12655 324
rect 12597 -264 12655 -252
rect 12715 324 12773 336
rect 12715 -252 12727 324
rect 12761 -252 12773 324
rect 12715 -264 12773 -252
rect 12833 324 12891 336
rect 12833 -252 12845 324
rect 12879 -252 12891 324
rect 12833 -264 12891 -252
rect 12951 324 13009 336
rect 12951 -252 12963 324
rect 12997 -252 13009 324
rect 12951 -264 13009 -252
rect 13069 324 13127 336
rect 13069 -252 13081 324
rect 13115 -252 13127 324
rect 13069 -264 13127 -252
rect 13187 324 13245 336
rect 13187 -252 13199 324
rect 13233 -252 13245 324
rect 13187 -264 13245 -252
rect 13305 324 13363 336
rect 13305 -252 13317 324
rect 13351 -252 13363 324
rect 13305 -264 13363 -252
rect 13423 324 13481 336
rect 13423 -252 13435 324
rect 13469 -252 13481 324
rect 13423 -264 13481 -252
rect 13541 324 13599 336
rect 13541 -252 13553 324
rect 13587 -252 13599 324
rect 13541 -264 13599 -252
rect 13659 324 13717 336
rect 13659 -252 13671 324
rect 13705 -252 13717 324
rect 13659 -264 13717 -252
rect 13777 324 13835 336
rect 13777 -252 13789 324
rect 13823 -252 13835 324
rect 13777 -264 13835 -252
rect 13895 324 13953 336
rect 13895 -252 13907 324
rect 13941 -252 13953 324
rect 13895 -264 13953 -252
rect 14013 324 14071 336
rect 14013 -252 14025 324
rect 14059 -252 14071 324
rect 14013 -264 14071 -252
rect 14131 324 14189 336
rect 14131 -252 14143 324
rect 14177 -252 14189 324
rect 14131 -264 14189 -252
rect 14249 324 14307 336
rect 14249 -252 14261 324
rect 14295 -252 14307 324
rect 14249 -264 14307 -252
rect 14367 324 14425 336
rect 14367 -252 14379 324
rect 14413 -252 14425 324
rect 14367 -264 14425 -252
rect 14485 324 14543 336
rect 14485 -252 14497 324
rect 14531 -252 14543 324
rect 14485 -264 14543 -252
rect 14603 324 14661 336
rect 14603 -252 14615 324
rect 14649 -252 14661 324
rect 14603 -264 14661 -252
rect 14721 324 14779 336
rect 14721 -252 14733 324
rect 14767 -252 14779 324
rect 14721 -264 14779 -252
<< pdiffc >>
rect -14767 -252 -14733 324
rect -14649 -252 -14615 324
rect -14531 -252 -14497 324
rect -14413 -252 -14379 324
rect -14295 -252 -14261 324
rect -14177 -252 -14143 324
rect -14059 -252 -14025 324
rect -13941 -252 -13907 324
rect -13823 -252 -13789 324
rect -13705 -252 -13671 324
rect -13587 -252 -13553 324
rect -13469 -252 -13435 324
rect -13351 -252 -13317 324
rect -13233 -252 -13199 324
rect -13115 -252 -13081 324
rect -12997 -252 -12963 324
rect -12879 -252 -12845 324
rect -12761 -252 -12727 324
rect -12643 -252 -12609 324
rect -12525 -252 -12491 324
rect -12407 -252 -12373 324
rect -12289 -252 -12255 324
rect -12171 -252 -12137 324
rect -12053 -252 -12019 324
rect -11935 -252 -11901 324
rect -11817 -252 -11783 324
rect -11699 -252 -11665 324
rect -11581 -252 -11547 324
rect -11463 -252 -11429 324
rect -11345 -252 -11311 324
rect -11227 -252 -11193 324
rect -11109 -252 -11075 324
rect -10991 -252 -10957 324
rect -10873 -252 -10839 324
rect -10755 -252 -10721 324
rect -10637 -252 -10603 324
rect -10519 -252 -10485 324
rect -10401 -252 -10367 324
rect -10283 -252 -10249 324
rect -10165 -252 -10131 324
rect -10047 -252 -10013 324
rect -9929 -252 -9895 324
rect -9811 -252 -9777 324
rect -9693 -252 -9659 324
rect -9575 -252 -9541 324
rect -9457 -252 -9423 324
rect -9339 -252 -9305 324
rect -9221 -252 -9187 324
rect -9103 -252 -9069 324
rect -8985 -252 -8951 324
rect -8867 -252 -8833 324
rect -8749 -252 -8715 324
rect -8631 -252 -8597 324
rect -8513 -252 -8479 324
rect -8395 -252 -8361 324
rect -8277 -252 -8243 324
rect -8159 -252 -8125 324
rect -8041 -252 -8007 324
rect -7923 -252 -7889 324
rect -7805 -252 -7771 324
rect -7687 -252 -7653 324
rect -7569 -252 -7535 324
rect -7451 -252 -7417 324
rect -7333 -252 -7299 324
rect -7215 -252 -7181 324
rect -7097 -252 -7063 324
rect -6979 -252 -6945 324
rect -6861 -252 -6827 324
rect -6743 -252 -6709 324
rect -6625 -252 -6591 324
rect -6507 -252 -6473 324
rect -6389 -252 -6355 324
rect -6271 -252 -6237 324
rect -6153 -252 -6119 324
rect -6035 -252 -6001 324
rect -5917 -252 -5883 324
rect -5799 -252 -5765 324
rect -5681 -252 -5647 324
rect -5563 -252 -5529 324
rect -5445 -252 -5411 324
rect -5327 -252 -5293 324
rect -5209 -252 -5175 324
rect -5091 -252 -5057 324
rect -4973 -252 -4939 324
rect -4855 -252 -4821 324
rect -4737 -252 -4703 324
rect -4619 -252 -4585 324
rect -4501 -252 -4467 324
rect -4383 -252 -4349 324
rect -4265 -252 -4231 324
rect -4147 -252 -4113 324
rect -4029 -252 -3995 324
rect -3911 -252 -3877 324
rect -3793 -252 -3759 324
rect -3675 -252 -3641 324
rect -3557 -252 -3523 324
rect -3439 -252 -3405 324
rect -3321 -252 -3287 324
rect -3203 -252 -3169 324
rect -3085 -252 -3051 324
rect -2967 -252 -2933 324
rect -2849 -252 -2815 324
rect -2731 -252 -2697 324
rect -2613 -252 -2579 324
rect -2495 -252 -2461 324
rect -2377 -252 -2343 324
rect -2259 -252 -2225 324
rect -2141 -252 -2107 324
rect -2023 -252 -1989 324
rect -1905 -252 -1871 324
rect -1787 -252 -1753 324
rect -1669 -252 -1635 324
rect -1551 -252 -1517 324
rect -1433 -252 -1399 324
rect -1315 -252 -1281 324
rect -1197 -252 -1163 324
rect -1079 -252 -1045 324
rect -961 -252 -927 324
rect -843 -252 -809 324
rect -725 -252 -691 324
rect -607 -252 -573 324
rect -489 -252 -455 324
rect -371 -252 -337 324
rect -253 -252 -219 324
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
rect 219 -252 253 324
rect 337 -252 371 324
rect 455 -252 489 324
rect 573 -252 607 324
rect 691 -252 725 324
rect 809 -252 843 324
rect 927 -252 961 324
rect 1045 -252 1079 324
rect 1163 -252 1197 324
rect 1281 -252 1315 324
rect 1399 -252 1433 324
rect 1517 -252 1551 324
rect 1635 -252 1669 324
rect 1753 -252 1787 324
rect 1871 -252 1905 324
rect 1989 -252 2023 324
rect 2107 -252 2141 324
rect 2225 -252 2259 324
rect 2343 -252 2377 324
rect 2461 -252 2495 324
rect 2579 -252 2613 324
rect 2697 -252 2731 324
rect 2815 -252 2849 324
rect 2933 -252 2967 324
rect 3051 -252 3085 324
rect 3169 -252 3203 324
rect 3287 -252 3321 324
rect 3405 -252 3439 324
rect 3523 -252 3557 324
rect 3641 -252 3675 324
rect 3759 -252 3793 324
rect 3877 -252 3911 324
rect 3995 -252 4029 324
rect 4113 -252 4147 324
rect 4231 -252 4265 324
rect 4349 -252 4383 324
rect 4467 -252 4501 324
rect 4585 -252 4619 324
rect 4703 -252 4737 324
rect 4821 -252 4855 324
rect 4939 -252 4973 324
rect 5057 -252 5091 324
rect 5175 -252 5209 324
rect 5293 -252 5327 324
rect 5411 -252 5445 324
rect 5529 -252 5563 324
rect 5647 -252 5681 324
rect 5765 -252 5799 324
rect 5883 -252 5917 324
rect 6001 -252 6035 324
rect 6119 -252 6153 324
rect 6237 -252 6271 324
rect 6355 -252 6389 324
rect 6473 -252 6507 324
rect 6591 -252 6625 324
rect 6709 -252 6743 324
rect 6827 -252 6861 324
rect 6945 -252 6979 324
rect 7063 -252 7097 324
rect 7181 -252 7215 324
rect 7299 -252 7333 324
rect 7417 -252 7451 324
rect 7535 -252 7569 324
rect 7653 -252 7687 324
rect 7771 -252 7805 324
rect 7889 -252 7923 324
rect 8007 -252 8041 324
rect 8125 -252 8159 324
rect 8243 -252 8277 324
rect 8361 -252 8395 324
rect 8479 -252 8513 324
rect 8597 -252 8631 324
rect 8715 -252 8749 324
rect 8833 -252 8867 324
rect 8951 -252 8985 324
rect 9069 -252 9103 324
rect 9187 -252 9221 324
rect 9305 -252 9339 324
rect 9423 -252 9457 324
rect 9541 -252 9575 324
rect 9659 -252 9693 324
rect 9777 -252 9811 324
rect 9895 -252 9929 324
rect 10013 -252 10047 324
rect 10131 -252 10165 324
rect 10249 -252 10283 324
rect 10367 -252 10401 324
rect 10485 -252 10519 324
rect 10603 -252 10637 324
rect 10721 -252 10755 324
rect 10839 -252 10873 324
rect 10957 -252 10991 324
rect 11075 -252 11109 324
rect 11193 -252 11227 324
rect 11311 -252 11345 324
rect 11429 -252 11463 324
rect 11547 -252 11581 324
rect 11665 -252 11699 324
rect 11783 -252 11817 324
rect 11901 -252 11935 324
rect 12019 -252 12053 324
rect 12137 -252 12171 324
rect 12255 -252 12289 324
rect 12373 -252 12407 324
rect 12491 -252 12525 324
rect 12609 -252 12643 324
rect 12727 -252 12761 324
rect 12845 -252 12879 324
rect 12963 -252 12997 324
rect 13081 -252 13115 324
rect 13199 -252 13233 324
rect 13317 -252 13351 324
rect 13435 -252 13469 324
rect 13553 -252 13587 324
rect 13671 -252 13705 324
rect 13789 -252 13823 324
rect 13907 -252 13941 324
rect 14025 -252 14059 324
rect 14143 -252 14177 324
rect 14261 -252 14295 324
rect 14379 -252 14413 324
rect 14497 -252 14531 324
rect 14615 -252 14649 324
rect 14733 -252 14767 324
<< nsubdiff >>
rect -14881 414 -14785 448
rect 14785 414 14881 448
rect -14881 351 -14847 414
rect 14847 351 14881 414
rect -14881 -414 -14847 -351
rect 14847 -414 14881 -351
rect -14881 -448 -14785 -414
rect 14785 -448 14881 -414
<< nsubdiffcont >>
rect -14785 414 14785 448
rect -14881 -351 -14847 351
rect 14847 -351 14881 351
rect -14785 -448 14785 -414
<< poly >>
rect -14721 336 -14661 362
rect -14603 336 -14543 362
rect -14485 336 -14425 362
rect -14367 336 -14307 362
rect -14249 336 -14189 362
rect -14131 336 -14071 362
rect -14013 336 -13953 362
rect -13895 336 -13835 362
rect -13777 336 -13717 362
rect -13659 336 -13599 362
rect -13541 336 -13481 362
rect -13423 336 -13363 362
rect -13305 336 -13245 362
rect -13187 336 -13127 362
rect -13069 336 -13009 362
rect -12951 336 -12891 362
rect -12833 336 -12773 362
rect -12715 336 -12655 362
rect -12597 336 -12537 362
rect -12479 336 -12419 362
rect -12361 336 -12301 362
rect -12243 336 -12183 362
rect -12125 336 -12065 362
rect -12007 336 -11947 362
rect -11889 336 -11829 362
rect -11771 336 -11711 362
rect -11653 336 -11593 362
rect -11535 336 -11475 362
rect -11417 336 -11357 362
rect -11299 336 -11239 362
rect -11181 336 -11121 362
rect -11063 336 -11003 362
rect -10945 336 -10885 362
rect -10827 336 -10767 362
rect -10709 336 -10649 362
rect -10591 336 -10531 362
rect -10473 336 -10413 362
rect -10355 336 -10295 362
rect -10237 336 -10177 362
rect -10119 336 -10059 362
rect -10001 336 -9941 362
rect -9883 336 -9823 362
rect -9765 336 -9705 362
rect -9647 336 -9587 362
rect -9529 336 -9469 362
rect -9411 336 -9351 362
rect -9293 336 -9233 362
rect -9175 336 -9115 362
rect -9057 336 -8997 362
rect -8939 336 -8879 362
rect -8821 336 -8761 362
rect -8703 336 -8643 362
rect -8585 336 -8525 362
rect -8467 336 -8407 362
rect -8349 336 -8289 362
rect -8231 336 -8171 362
rect -8113 336 -8053 362
rect -7995 336 -7935 362
rect -7877 336 -7817 362
rect -7759 336 -7699 362
rect -7641 336 -7581 362
rect -7523 336 -7463 362
rect -7405 336 -7345 362
rect -7287 336 -7227 362
rect -7169 336 -7109 362
rect -7051 336 -6991 362
rect -6933 336 -6873 362
rect -6815 336 -6755 362
rect -6697 336 -6637 362
rect -6579 336 -6519 362
rect -6461 336 -6401 362
rect -6343 336 -6283 362
rect -6225 336 -6165 362
rect -6107 336 -6047 362
rect -5989 336 -5929 362
rect -5871 336 -5811 362
rect -5753 336 -5693 362
rect -5635 336 -5575 362
rect -5517 336 -5457 362
rect -5399 336 -5339 362
rect -5281 336 -5221 362
rect -5163 336 -5103 362
rect -5045 336 -4985 362
rect -4927 336 -4867 362
rect -4809 336 -4749 362
rect -4691 336 -4631 362
rect -4573 336 -4513 362
rect -4455 336 -4395 362
rect -4337 336 -4277 362
rect -4219 336 -4159 362
rect -4101 336 -4041 362
rect -3983 336 -3923 362
rect -3865 336 -3805 362
rect -3747 336 -3687 362
rect -3629 336 -3569 362
rect -3511 336 -3451 362
rect -3393 336 -3333 362
rect -3275 336 -3215 362
rect -3157 336 -3097 362
rect -3039 336 -2979 362
rect -2921 336 -2861 362
rect -2803 336 -2743 362
rect -2685 336 -2625 362
rect -2567 336 -2507 362
rect -2449 336 -2389 362
rect -2331 336 -2271 362
rect -2213 336 -2153 362
rect -2095 336 -2035 362
rect -1977 336 -1917 362
rect -1859 336 -1799 362
rect -1741 336 -1681 362
rect -1623 336 -1563 362
rect -1505 336 -1445 362
rect -1387 336 -1327 362
rect -1269 336 -1209 362
rect -1151 336 -1091 362
rect -1033 336 -973 362
rect -915 336 -855 362
rect -797 336 -737 362
rect -679 336 -619 362
rect -561 336 -501 362
rect -443 336 -383 362
rect -325 336 -265 362
rect -207 336 -147 362
rect -89 336 -29 362
rect 29 336 89 362
rect 147 336 207 362
rect 265 336 325 362
rect 383 336 443 362
rect 501 336 561 362
rect 619 336 679 362
rect 737 336 797 362
rect 855 336 915 362
rect 973 336 1033 362
rect 1091 336 1151 362
rect 1209 336 1269 362
rect 1327 336 1387 362
rect 1445 336 1505 362
rect 1563 336 1623 362
rect 1681 336 1741 362
rect 1799 336 1859 362
rect 1917 336 1977 362
rect 2035 336 2095 362
rect 2153 336 2213 362
rect 2271 336 2331 362
rect 2389 336 2449 362
rect 2507 336 2567 362
rect 2625 336 2685 362
rect 2743 336 2803 362
rect 2861 336 2921 362
rect 2979 336 3039 362
rect 3097 336 3157 362
rect 3215 336 3275 362
rect 3333 336 3393 362
rect 3451 336 3511 362
rect 3569 336 3629 362
rect 3687 336 3747 362
rect 3805 336 3865 362
rect 3923 336 3983 362
rect 4041 336 4101 362
rect 4159 336 4219 362
rect 4277 336 4337 362
rect 4395 336 4455 362
rect 4513 336 4573 362
rect 4631 336 4691 362
rect 4749 336 4809 362
rect 4867 336 4927 362
rect 4985 336 5045 362
rect 5103 336 5163 362
rect 5221 336 5281 362
rect 5339 336 5399 362
rect 5457 336 5517 362
rect 5575 336 5635 362
rect 5693 336 5753 362
rect 5811 336 5871 362
rect 5929 336 5989 362
rect 6047 336 6107 362
rect 6165 336 6225 362
rect 6283 336 6343 362
rect 6401 336 6461 362
rect 6519 336 6579 362
rect 6637 336 6697 362
rect 6755 336 6815 362
rect 6873 336 6933 362
rect 6991 336 7051 362
rect 7109 336 7169 362
rect 7227 336 7287 362
rect 7345 336 7405 362
rect 7463 336 7523 362
rect 7581 336 7641 362
rect 7699 336 7759 362
rect 7817 336 7877 362
rect 7935 336 7995 362
rect 8053 336 8113 362
rect 8171 336 8231 362
rect 8289 336 8349 362
rect 8407 336 8467 362
rect 8525 336 8585 362
rect 8643 336 8703 362
rect 8761 336 8821 362
rect 8879 336 8939 362
rect 8997 336 9057 362
rect 9115 336 9175 362
rect 9233 336 9293 362
rect 9351 336 9411 362
rect 9469 336 9529 362
rect 9587 336 9647 362
rect 9705 336 9765 362
rect 9823 336 9883 362
rect 9941 336 10001 362
rect 10059 336 10119 362
rect 10177 336 10237 362
rect 10295 336 10355 362
rect 10413 336 10473 362
rect 10531 336 10591 362
rect 10649 336 10709 362
rect 10767 336 10827 362
rect 10885 336 10945 362
rect 11003 336 11063 362
rect 11121 336 11181 362
rect 11239 336 11299 362
rect 11357 336 11417 362
rect 11475 336 11535 362
rect 11593 336 11653 362
rect 11711 336 11771 362
rect 11829 336 11889 362
rect 11947 336 12007 362
rect 12065 336 12125 362
rect 12183 336 12243 362
rect 12301 336 12361 362
rect 12419 336 12479 362
rect 12537 336 12597 362
rect 12655 336 12715 362
rect 12773 336 12833 362
rect 12891 336 12951 362
rect 13009 336 13069 362
rect 13127 336 13187 362
rect 13245 336 13305 362
rect 13363 336 13423 362
rect 13481 336 13541 362
rect 13599 336 13659 362
rect 13717 336 13777 362
rect 13835 336 13895 362
rect 13953 336 14013 362
rect 14071 336 14131 362
rect 14189 336 14249 362
rect 14307 336 14367 362
rect 14425 336 14485 362
rect 14543 336 14603 362
rect 14661 336 14721 362
rect -14721 -295 -14661 -264
rect -14603 -295 -14543 -264
rect -14485 -295 -14425 -264
rect -14367 -295 -14307 -264
rect -14249 -295 -14189 -264
rect -14131 -295 -14071 -264
rect -14013 -295 -13953 -264
rect -13895 -295 -13835 -264
rect -13777 -295 -13717 -264
rect -13659 -295 -13599 -264
rect -13541 -295 -13481 -264
rect -13423 -295 -13363 -264
rect -13305 -295 -13245 -264
rect -13187 -295 -13127 -264
rect -13069 -295 -13009 -264
rect -12951 -295 -12891 -264
rect -12833 -295 -12773 -264
rect -12715 -295 -12655 -264
rect -12597 -295 -12537 -264
rect -12479 -295 -12419 -264
rect -12361 -295 -12301 -264
rect -12243 -295 -12183 -264
rect -12125 -295 -12065 -264
rect -12007 -295 -11947 -264
rect -11889 -295 -11829 -264
rect -11771 -295 -11711 -264
rect -11653 -295 -11593 -264
rect -11535 -295 -11475 -264
rect -11417 -295 -11357 -264
rect -11299 -295 -11239 -264
rect -11181 -295 -11121 -264
rect -11063 -295 -11003 -264
rect -10945 -295 -10885 -264
rect -10827 -295 -10767 -264
rect -10709 -295 -10649 -264
rect -10591 -295 -10531 -264
rect -10473 -295 -10413 -264
rect -10355 -295 -10295 -264
rect -10237 -295 -10177 -264
rect -10119 -295 -10059 -264
rect -10001 -295 -9941 -264
rect -9883 -295 -9823 -264
rect -9765 -295 -9705 -264
rect -9647 -295 -9587 -264
rect -9529 -295 -9469 -264
rect -9411 -295 -9351 -264
rect -9293 -295 -9233 -264
rect -9175 -295 -9115 -264
rect -9057 -295 -8997 -264
rect -8939 -295 -8879 -264
rect -8821 -295 -8761 -264
rect -8703 -295 -8643 -264
rect -8585 -295 -8525 -264
rect -8467 -295 -8407 -264
rect -8349 -295 -8289 -264
rect -8231 -295 -8171 -264
rect -8113 -295 -8053 -264
rect -7995 -295 -7935 -264
rect -7877 -295 -7817 -264
rect -7759 -295 -7699 -264
rect -7641 -295 -7581 -264
rect -7523 -295 -7463 -264
rect -7405 -295 -7345 -264
rect -7287 -295 -7227 -264
rect -7169 -295 -7109 -264
rect -7051 -295 -6991 -264
rect -6933 -295 -6873 -264
rect -6815 -295 -6755 -264
rect -6697 -295 -6637 -264
rect -6579 -295 -6519 -264
rect -6461 -295 -6401 -264
rect -6343 -295 -6283 -264
rect -6225 -295 -6165 -264
rect -6107 -295 -6047 -264
rect -5989 -295 -5929 -264
rect -5871 -295 -5811 -264
rect -5753 -295 -5693 -264
rect -5635 -295 -5575 -264
rect -5517 -295 -5457 -264
rect -5399 -295 -5339 -264
rect -5281 -295 -5221 -264
rect -5163 -295 -5103 -264
rect -5045 -295 -4985 -264
rect -4927 -295 -4867 -264
rect -4809 -295 -4749 -264
rect -4691 -295 -4631 -264
rect -4573 -295 -4513 -264
rect -4455 -295 -4395 -264
rect -4337 -295 -4277 -264
rect -4219 -295 -4159 -264
rect -4101 -295 -4041 -264
rect -3983 -295 -3923 -264
rect -3865 -295 -3805 -264
rect -3747 -295 -3687 -264
rect -3629 -295 -3569 -264
rect -3511 -295 -3451 -264
rect -3393 -295 -3333 -264
rect -3275 -295 -3215 -264
rect -3157 -295 -3097 -264
rect -3039 -295 -2979 -264
rect -2921 -295 -2861 -264
rect -2803 -295 -2743 -264
rect -2685 -295 -2625 -264
rect -2567 -295 -2507 -264
rect -2449 -295 -2389 -264
rect -2331 -295 -2271 -264
rect -2213 -295 -2153 -264
rect -2095 -295 -2035 -264
rect -1977 -295 -1917 -264
rect -1859 -295 -1799 -264
rect -1741 -295 -1681 -264
rect -1623 -295 -1563 -264
rect -1505 -295 -1445 -264
rect -1387 -295 -1327 -264
rect -1269 -295 -1209 -264
rect -1151 -295 -1091 -264
rect -1033 -295 -973 -264
rect -915 -295 -855 -264
rect -797 -295 -737 -264
rect -679 -295 -619 -264
rect -561 -295 -501 -264
rect -443 -295 -383 -264
rect -325 -295 -265 -264
rect -207 -295 -147 -264
rect -89 -295 -29 -264
rect 29 -295 89 -264
rect 147 -295 207 -264
rect 265 -295 325 -264
rect 383 -295 443 -264
rect 501 -295 561 -264
rect 619 -295 679 -264
rect 737 -295 797 -264
rect 855 -295 915 -264
rect 973 -295 1033 -264
rect 1091 -295 1151 -264
rect 1209 -295 1269 -264
rect 1327 -295 1387 -264
rect 1445 -295 1505 -264
rect 1563 -295 1623 -264
rect 1681 -295 1741 -264
rect 1799 -295 1859 -264
rect 1917 -295 1977 -264
rect 2035 -295 2095 -264
rect 2153 -295 2213 -264
rect 2271 -295 2331 -264
rect 2389 -295 2449 -264
rect 2507 -295 2567 -264
rect 2625 -295 2685 -264
rect 2743 -295 2803 -264
rect 2861 -295 2921 -264
rect 2979 -295 3039 -264
rect 3097 -295 3157 -264
rect 3215 -295 3275 -264
rect 3333 -295 3393 -264
rect 3451 -295 3511 -264
rect 3569 -295 3629 -264
rect 3687 -295 3747 -264
rect 3805 -295 3865 -264
rect 3923 -295 3983 -264
rect 4041 -295 4101 -264
rect 4159 -295 4219 -264
rect 4277 -295 4337 -264
rect 4395 -295 4455 -264
rect 4513 -295 4573 -264
rect 4631 -295 4691 -264
rect 4749 -295 4809 -264
rect 4867 -295 4927 -264
rect 4985 -295 5045 -264
rect 5103 -295 5163 -264
rect 5221 -295 5281 -264
rect 5339 -295 5399 -264
rect 5457 -295 5517 -264
rect 5575 -295 5635 -264
rect 5693 -295 5753 -264
rect 5811 -295 5871 -264
rect 5929 -295 5989 -264
rect 6047 -295 6107 -264
rect 6165 -295 6225 -264
rect 6283 -295 6343 -264
rect 6401 -295 6461 -264
rect 6519 -295 6579 -264
rect 6637 -295 6697 -264
rect 6755 -295 6815 -264
rect 6873 -295 6933 -264
rect 6991 -295 7051 -264
rect 7109 -295 7169 -264
rect 7227 -295 7287 -264
rect 7345 -295 7405 -264
rect 7463 -295 7523 -264
rect 7581 -295 7641 -264
rect 7699 -295 7759 -264
rect 7817 -295 7877 -264
rect 7935 -295 7995 -264
rect 8053 -295 8113 -264
rect 8171 -295 8231 -264
rect 8289 -295 8349 -264
rect 8407 -295 8467 -264
rect 8525 -295 8585 -264
rect 8643 -295 8703 -264
rect 8761 -295 8821 -264
rect 8879 -295 8939 -264
rect 8997 -295 9057 -264
rect 9115 -295 9175 -264
rect 9233 -295 9293 -264
rect 9351 -295 9411 -264
rect 9469 -295 9529 -264
rect 9587 -295 9647 -264
rect 9705 -295 9765 -264
rect 9823 -295 9883 -264
rect 9941 -295 10001 -264
rect 10059 -295 10119 -264
rect 10177 -295 10237 -264
rect 10295 -295 10355 -264
rect 10413 -295 10473 -264
rect 10531 -295 10591 -264
rect 10649 -295 10709 -264
rect 10767 -295 10827 -264
rect 10885 -295 10945 -264
rect 11003 -295 11063 -264
rect 11121 -295 11181 -264
rect 11239 -295 11299 -264
rect 11357 -295 11417 -264
rect 11475 -295 11535 -264
rect 11593 -295 11653 -264
rect 11711 -295 11771 -264
rect 11829 -295 11889 -264
rect 11947 -295 12007 -264
rect 12065 -295 12125 -264
rect 12183 -295 12243 -264
rect 12301 -295 12361 -264
rect 12419 -295 12479 -264
rect 12537 -295 12597 -264
rect 12655 -295 12715 -264
rect 12773 -295 12833 -264
rect 12891 -295 12951 -264
rect 13009 -295 13069 -264
rect 13127 -295 13187 -264
rect 13245 -295 13305 -264
rect 13363 -295 13423 -264
rect 13481 -295 13541 -264
rect 13599 -295 13659 -264
rect 13717 -295 13777 -264
rect 13835 -295 13895 -264
rect 13953 -295 14013 -264
rect 14071 -295 14131 -264
rect 14189 -295 14249 -264
rect 14307 -295 14367 -264
rect 14425 -295 14485 -264
rect 14543 -295 14603 -264
rect 14661 -295 14721 -264
rect -14724 -311 -14658 -295
rect -14724 -345 -14708 -311
rect -14674 -345 -14658 -311
rect -14724 -361 -14658 -345
rect -14606 -311 -14540 -295
rect -14606 -345 -14590 -311
rect -14556 -345 -14540 -311
rect -14606 -361 -14540 -345
rect -14488 -311 -14422 -295
rect -14488 -345 -14472 -311
rect -14438 -345 -14422 -311
rect -14488 -361 -14422 -345
rect -14370 -311 -14304 -295
rect -14370 -345 -14354 -311
rect -14320 -345 -14304 -311
rect -14370 -361 -14304 -345
rect -14252 -311 -14186 -295
rect -14252 -345 -14236 -311
rect -14202 -345 -14186 -311
rect -14252 -361 -14186 -345
rect -14134 -311 -14068 -295
rect -14134 -345 -14118 -311
rect -14084 -345 -14068 -311
rect -14134 -361 -14068 -345
rect -14016 -311 -13950 -295
rect -14016 -345 -14000 -311
rect -13966 -345 -13950 -311
rect -14016 -361 -13950 -345
rect -13898 -311 -13832 -295
rect -13898 -345 -13882 -311
rect -13848 -345 -13832 -311
rect -13898 -361 -13832 -345
rect -13780 -311 -13714 -295
rect -13780 -345 -13764 -311
rect -13730 -345 -13714 -311
rect -13780 -361 -13714 -345
rect -13662 -311 -13596 -295
rect -13662 -345 -13646 -311
rect -13612 -345 -13596 -311
rect -13662 -361 -13596 -345
rect -13544 -311 -13478 -295
rect -13544 -345 -13528 -311
rect -13494 -345 -13478 -311
rect -13544 -361 -13478 -345
rect -13426 -311 -13360 -295
rect -13426 -345 -13410 -311
rect -13376 -345 -13360 -311
rect -13426 -361 -13360 -345
rect -13308 -311 -13242 -295
rect -13308 -345 -13292 -311
rect -13258 -345 -13242 -311
rect -13308 -361 -13242 -345
rect -13190 -311 -13124 -295
rect -13190 -345 -13174 -311
rect -13140 -345 -13124 -311
rect -13190 -361 -13124 -345
rect -13072 -311 -13006 -295
rect -13072 -345 -13056 -311
rect -13022 -345 -13006 -311
rect -13072 -361 -13006 -345
rect -12954 -311 -12888 -295
rect -12954 -345 -12938 -311
rect -12904 -345 -12888 -311
rect -12954 -361 -12888 -345
rect -12836 -311 -12770 -295
rect -12836 -345 -12820 -311
rect -12786 -345 -12770 -311
rect -12836 -361 -12770 -345
rect -12718 -311 -12652 -295
rect -12718 -345 -12702 -311
rect -12668 -345 -12652 -311
rect -12718 -361 -12652 -345
rect -12600 -311 -12534 -295
rect -12600 -345 -12584 -311
rect -12550 -345 -12534 -311
rect -12600 -361 -12534 -345
rect -12482 -311 -12416 -295
rect -12482 -345 -12466 -311
rect -12432 -345 -12416 -311
rect -12482 -361 -12416 -345
rect -12364 -311 -12298 -295
rect -12364 -345 -12348 -311
rect -12314 -345 -12298 -311
rect -12364 -361 -12298 -345
rect -12246 -311 -12180 -295
rect -12246 -345 -12230 -311
rect -12196 -345 -12180 -311
rect -12246 -361 -12180 -345
rect -12128 -311 -12062 -295
rect -12128 -345 -12112 -311
rect -12078 -345 -12062 -311
rect -12128 -361 -12062 -345
rect -12010 -311 -11944 -295
rect -12010 -345 -11994 -311
rect -11960 -345 -11944 -311
rect -12010 -361 -11944 -345
rect -11892 -311 -11826 -295
rect -11892 -345 -11876 -311
rect -11842 -345 -11826 -311
rect -11892 -361 -11826 -345
rect -11774 -311 -11708 -295
rect -11774 -345 -11758 -311
rect -11724 -345 -11708 -311
rect -11774 -361 -11708 -345
rect -11656 -311 -11590 -295
rect -11656 -345 -11640 -311
rect -11606 -345 -11590 -311
rect -11656 -361 -11590 -345
rect -11538 -311 -11472 -295
rect -11538 -345 -11522 -311
rect -11488 -345 -11472 -311
rect -11538 -361 -11472 -345
rect -11420 -311 -11354 -295
rect -11420 -345 -11404 -311
rect -11370 -345 -11354 -311
rect -11420 -361 -11354 -345
rect -11302 -311 -11236 -295
rect -11302 -345 -11286 -311
rect -11252 -345 -11236 -311
rect -11302 -361 -11236 -345
rect -11184 -311 -11118 -295
rect -11184 -345 -11168 -311
rect -11134 -345 -11118 -311
rect -11184 -361 -11118 -345
rect -11066 -311 -11000 -295
rect -11066 -345 -11050 -311
rect -11016 -345 -11000 -311
rect -11066 -361 -11000 -345
rect -10948 -311 -10882 -295
rect -10948 -345 -10932 -311
rect -10898 -345 -10882 -311
rect -10948 -361 -10882 -345
rect -10830 -311 -10764 -295
rect -10830 -345 -10814 -311
rect -10780 -345 -10764 -311
rect -10830 -361 -10764 -345
rect -10712 -311 -10646 -295
rect -10712 -345 -10696 -311
rect -10662 -345 -10646 -311
rect -10712 -361 -10646 -345
rect -10594 -311 -10528 -295
rect -10594 -345 -10578 -311
rect -10544 -345 -10528 -311
rect -10594 -361 -10528 -345
rect -10476 -311 -10410 -295
rect -10476 -345 -10460 -311
rect -10426 -345 -10410 -311
rect -10476 -361 -10410 -345
rect -10358 -311 -10292 -295
rect -10358 -345 -10342 -311
rect -10308 -345 -10292 -311
rect -10358 -361 -10292 -345
rect -10240 -311 -10174 -295
rect -10240 -345 -10224 -311
rect -10190 -345 -10174 -311
rect -10240 -361 -10174 -345
rect -10122 -311 -10056 -295
rect -10122 -345 -10106 -311
rect -10072 -345 -10056 -311
rect -10122 -361 -10056 -345
rect -10004 -311 -9938 -295
rect -10004 -345 -9988 -311
rect -9954 -345 -9938 -311
rect -10004 -361 -9938 -345
rect -9886 -311 -9820 -295
rect -9886 -345 -9870 -311
rect -9836 -345 -9820 -311
rect -9886 -361 -9820 -345
rect -9768 -311 -9702 -295
rect -9768 -345 -9752 -311
rect -9718 -345 -9702 -311
rect -9768 -361 -9702 -345
rect -9650 -311 -9584 -295
rect -9650 -345 -9634 -311
rect -9600 -345 -9584 -311
rect -9650 -361 -9584 -345
rect -9532 -311 -9466 -295
rect -9532 -345 -9516 -311
rect -9482 -345 -9466 -311
rect -9532 -361 -9466 -345
rect -9414 -311 -9348 -295
rect -9414 -345 -9398 -311
rect -9364 -345 -9348 -311
rect -9414 -361 -9348 -345
rect -9296 -311 -9230 -295
rect -9296 -345 -9280 -311
rect -9246 -345 -9230 -311
rect -9296 -361 -9230 -345
rect -9178 -311 -9112 -295
rect -9178 -345 -9162 -311
rect -9128 -345 -9112 -311
rect -9178 -361 -9112 -345
rect -9060 -311 -8994 -295
rect -9060 -345 -9044 -311
rect -9010 -345 -8994 -311
rect -9060 -361 -8994 -345
rect -8942 -311 -8876 -295
rect -8942 -345 -8926 -311
rect -8892 -345 -8876 -311
rect -8942 -361 -8876 -345
rect -8824 -311 -8758 -295
rect -8824 -345 -8808 -311
rect -8774 -345 -8758 -311
rect -8824 -361 -8758 -345
rect -8706 -311 -8640 -295
rect -8706 -345 -8690 -311
rect -8656 -345 -8640 -311
rect -8706 -361 -8640 -345
rect -8588 -311 -8522 -295
rect -8588 -345 -8572 -311
rect -8538 -345 -8522 -311
rect -8588 -361 -8522 -345
rect -8470 -311 -8404 -295
rect -8470 -345 -8454 -311
rect -8420 -345 -8404 -311
rect -8470 -361 -8404 -345
rect -8352 -311 -8286 -295
rect -8352 -345 -8336 -311
rect -8302 -345 -8286 -311
rect -8352 -361 -8286 -345
rect -8234 -311 -8168 -295
rect -8234 -345 -8218 -311
rect -8184 -345 -8168 -311
rect -8234 -361 -8168 -345
rect -8116 -311 -8050 -295
rect -8116 -345 -8100 -311
rect -8066 -345 -8050 -311
rect -8116 -361 -8050 -345
rect -7998 -311 -7932 -295
rect -7998 -345 -7982 -311
rect -7948 -345 -7932 -311
rect -7998 -361 -7932 -345
rect -7880 -311 -7814 -295
rect -7880 -345 -7864 -311
rect -7830 -345 -7814 -311
rect -7880 -361 -7814 -345
rect -7762 -311 -7696 -295
rect -7762 -345 -7746 -311
rect -7712 -345 -7696 -311
rect -7762 -361 -7696 -345
rect -7644 -311 -7578 -295
rect -7644 -345 -7628 -311
rect -7594 -345 -7578 -311
rect -7644 -361 -7578 -345
rect -7526 -311 -7460 -295
rect -7526 -345 -7510 -311
rect -7476 -345 -7460 -311
rect -7526 -361 -7460 -345
rect -7408 -311 -7342 -295
rect -7408 -345 -7392 -311
rect -7358 -345 -7342 -311
rect -7408 -361 -7342 -345
rect -7290 -311 -7224 -295
rect -7290 -345 -7274 -311
rect -7240 -345 -7224 -311
rect -7290 -361 -7224 -345
rect -7172 -311 -7106 -295
rect -7172 -345 -7156 -311
rect -7122 -345 -7106 -311
rect -7172 -361 -7106 -345
rect -7054 -311 -6988 -295
rect -7054 -345 -7038 -311
rect -7004 -345 -6988 -311
rect -7054 -361 -6988 -345
rect -6936 -311 -6870 -295
rect -6936 -345 -6920 -311
rect -6886 -345 -6870 -311
rect -6936 -361 -6870 -345
rect -6818 -311 -6752 -295
rect -6818 -345 -6802 -311
rect -6768 -345 -6752 -311
rect -6818 -361 -6752 -345
rect -6700 -311 -6634 -295
rect -6700 -345 -6684 -311
rect -6650 -345 -6634 -311
rect -6700 -361 -6634 -345
rect -6582 -311 -6516 -295
rect -6582 -345 -6566 -311
rect -6532 -345 -6516 -311
rect -6582 -361 -6516 -345
rect -6464 -311 -6398 -295
rect -6464 -345 -6448 -311
rect -6414 -345 -6398 -311
rect -6464 -361 -6398 -345
rect -6346 -311 -6280 -295
rect -6346 -345 -6330 -311
rect -6296 -345 -6280 -311
rect -6346 -361 -6280 -345
rect -6228 -311 -6162 -295
rect -6228 -345 -6212 -311
rect -6178 -345 -6162 -311
rect -6228 -361 -6162 -345
rect -6110 -311 -6044 -295
rect -6110 -345 -6094 -311
rect -6060 -345 -6044 -311
rect -6110 -361 -6044 -345
rect -5992 -311 -5926 -295
rect -5992 -345 -5976 -311
rect -5942 -345 -5926 -311
rect -5992 -361 -5926 -345
rect -5874 -311 -5808 -295
rect -5874 -345 -5858 -311
rect -5824 -345 -5808 -311
rect -5874 -361 -5808 -345
rect -5756 -311 -5690 -295
rect -5756 -345 -5740 -311
rect -5706 -345 -5690 -311
rect -5756 -361 -5690 -345
rect -5638 -311 -5572 -295
rect -5638 -345 -5622 -311
rect -5588 -345 -5572 -311
rect -5638 -361 -5572 -345
rect -5520 -311 -5454 -295
rect -5520 -345 -5504 -311
rect -5470 -345 -5454 -311
rect -5520 -361 -5454 -345
rect -5402 -311 -5336 -295
rect -5402 -345 -5386 -311
rect -5352 -345 -5336 -311
rect -5402 -361 -5336 -345
rect -5284 -311 -5218 -295
rect -5284 -345 -5268 -311
rect -5234 -345 -5218 -311
rect -5284 -361 -5218 -345
rect -5166 -311 -5100 -295
rect -5166 -345 -5150 -311
rect -5116 -345 -5100 -311
rect -5166 -361 -5100 -345
rect -5048 -311 -4982 -295
rect -5048 -345 -5032 -311
rect -4998 -345 -4982 -311
rect -5048 -361 -4982 -345
rect -4930 -311 -4864 -295
rect -4930 -345 -4914 -311
rect -4880 -345 -4864 -311
rect -4930 -361 -4864 -345
rect -4812 -311 -4746 -295
rect -4812 -345 -4796 -311
rect -4762 -345 -4746 -311
rect -4812 -361 -4746 -345
rect -4694 -311 -4628 -295
rect -4694 -345 -4678 -311
rect -4644 -345 -4628 -311
rect -4694 -361 -4628 -345
rect -4576 -311 -4510 -295
rect -4576 -345 -4560 -311
rect -4526 -345 -4510 -311
rect -4576 -361 -4510 -345
rect -4458 -311 -4392 -295
rect -4458 -345 -4442 -311
rect -4408 -345 -4392 -311
rect -4458 -361 -4392 -345
rect -4340 -311 -4274 -295
rect -4340 -345 -4324 -311
rect -4290 -345 -4274 -311
rect -4340 -361 -4274 -345
rect -4222 -311 -4156 -295
rect -4222 -345 -4206 -311
rect -4172 -345 -4156 -311
rect -4222 -361 -4156 -345
rect -4104 -311 -4038 -295
rect -4104 -345 -4088 -311
rect -4054 -345 -4038 -311
rect -4104 -361 -4038 -345
rect -3986 -311 -3920 -295
rect -3986 -345 -3970 -311
rect -3936 -345 -3920 -311
rect -3986 -361 -3920 -345
rect -3868 -311 -3802 -295
rect -3868 -345 -3852 -311
rect -3818 -345 -3802 -311
rect -3868 -361 -3802 -345
rect -3750 -311 -3684 -295
rect -3750 -345 -3734 -311
rect -3700 -345 -3684 -311
rect -3750 -361 -3684 -345
rect -3632 -311 -3566 -295
rect -3632 -345 -3616 -311
rect -3582 -345 -3566 -311
rect -3632 -361 -3566 -345
rect -3514 -311 -3448 -295
rect -3514 -345 -3498 -311
rect -3464 -345 -3448 -311
rect -3514 -361 -3448 -345
rect -3396 -311 -3330 -295
rect -3396 -345 -3380 -311
rect -3346 -345 -3330 -311
rect -3396 -361 -3330 -345
rect -3278 -311 -3212 -295
rect -3278 -345 -3262 -311
rect -3228 -345 -3212 -311
rect -3278 -361 -3212 -345
rect -3160 -311 -3094 -295
rect -3160 -345 -3144 -311
rect -3110 -345 -3094 -311
rect -3160 -361 -3094 -345
rect -3042 -311 -2976 -295
rect -3042 -345 -3026 -311
rect -2992 -345 -2976 -311
rect -3042 -361 -2976 -345
rect -2924 -311 -2858 -295
rect -2924 -345 -2908 -311
rect -2874 -345 -2858 -311
rect -2924 -361 -2858 -345
rect -2806 -311 -2740 -295
rect -2806 -345 -2790 -311
rect -2756 -345 -2740 -311
rect -2806 -361 -2740 -345
rect -2688 -311 -2622 -295
rect -2688 -345 -2672 -311
rect -2638 -345 -2622 -311
rect -2688 -361 -2622 -345
rect -2570 -311 -2504 -295
rect -2570 -345 -2554 -311
rect -2520 -345 -2504 -311
rect -2570 -361 -2504 -345
rect -2452 -311 -2386 -295
rect -2452 -345 -2436 -311
rect -2402 -345 -2386 -311
rect -2452 -361 -2386 -345
rect -2334 -311 -2268 -295
rect -2334 -345 -2318 -311
rect -2284 -345 -2268 -311
rect -2334 -361 -2268 -345
rect -2216 -311 -2150 -295
rect -2216 -345 -2200 -311
rect -2166 -345 -2150 -311
rect -2216 -361 -2150 -345
rect -2098 -311 -2032 -295
rect -2098 -345 -2082 -311
rect -2048 -345 -2032 -311
rect -2098 -361 -2032 -345
rect -1980 -311 -1914 -295
rect -1980 -345 -1964 -311
rect -1930 -345 -1914 -311
rect -1980 -361 -1914 -345
rect -1862 -311 -1796 -295
rect -1862 -345 -1846 -311
rect -1812 -345 -1796 -311
rect -1862 -361 -1796 -345
rect -1744 -311 -1678 -295
rect -1744 -345 -1728 -311
rect -1694 -345 -1678 -311
rect -1744 -361 -1678 -345
rect -1626 -311 -1560 -295
rect -1626 -345 -1610 -311
rect -1576 -345 -1560 -311
rect -1626 -361 -1560 -345
rect -1508 -311 -1442 -295
rect -1508 -345 -1492 -311
rect -1458 -345 -1442 -311
rect -1508 -361 -1442 -345
rect -1390 -311 -1324 -295
rect -1390 -345 -1374 -311
rect -1340 -345 -1324 -311
rect -1390 -361 -1324 -345
rect -1272 -311 -1206 -295
rect -1272 -345 -1256 -311
rect -1222 -345 -1206 -311
rect -1272 -361 -1206 -345
rect -1154 -311 -1088 -295
rect -1154 -345 -1138 -311
rect -1104 -345 -1088 -311
rect -1154 -361 -1088 -345
rect -1036 -311 -970 -295
rect -1036 -345 -1020 -311
rect -986 -345 -970 -311
rect -1036 -361 -970 -345
rect -918 -311 -852 -295
rect -918 -345 -902 -311
rect -868 -345 -852 -311
rect -918 -361 -852 -345
rect -800 -311 -734 -295
rect -800 -345 -784 -311
rect -750 -345 -734 -311
rect -800 -361 -734 -345
rect -682 -311 -616 -295
rect -682 -345 -666 -311
rect -632 -345 -616 -311
rect -682 -361 -616 -345
rect -564 -311 -498 -295
rect -564 -345 -548 -311
rect -514 -345 -498 -311
rect -564 -361 -498 -345
rect -446 -311 -380 -295
rect -446 -345 -430 -311
rect -396 -345 -380 -311
rect -446 -361 -380 -345
rect -328 -311 -262 -295
rect -328 -345 -312 -311
rect -278 -345 -262 -311
rect -328 -361 -262 -345
rect -210 -311 -144 -295
rect -210 -345 -194 -311
rect -160 -345 -144 -311
rect -210 -361 -144 -345
rect -92 -311 -26 -295
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect -92 -361 -26 -345
rect 26 -311 92 -295
rect 26 -345 42 -311
rect 76 -345 92 -311
rect 26 -361 92 -345
rect 144 -311 210 -295
rect 144 -345 160 -311
rect 194 -345 210 -311
rect 144 -361 210 -345
rect 262 -311 328 -295
rect 262 -345 278 -311
rect 312 -345 328 -311
rect 262 -361 328 -345
rect 380 -311 446 -295
rect 380 -345 396 -311
rect 430 -345 446 -311
rect 380 -361 446 -345
rect 498 -311 564 -295
rect 498 -345 514 -311
rect 548 -345 564 -311
rect 498 -361 564 -345
rect 616 -311 682 -295
rect 616 -345 632 -311
rect 666 -345 682 -311
rect 616 -361 682 -345
rect 734 -311 800 -295
rect 734 -345 750 -311
rect 784 -345 800 -311
rect 734 -361 800 -345
rect 852 -311 918 -295
rect 852 -345 868 -311
rect 902 -345 918 -311
rect 852 -361 918 -345
rect 970 -311 1036 -295
rect 970 -345 986 -311
rect 1020 -345 1036 -311
rect 970 -361 1036 -345
rect 1088 -311 1154 -295
rect 1088 -345 1104 -311
rect 1138 -345 1154 -311
rect 1088 -361 1154 -345
rect 1206 -311 1272 -295
rect 1206 -345 1222 -311
rect 1256 -345 1272 -311
rect 1206 -361 1272 -345
rect 1324 -311 1390 -295
rect 1324 -345 1340 -311
rect 1374 -345 1390 -311
rect 1324 -361 1390 -345
rect 1442 -311 1508 -295
rect 1442 -345 1458 -311
rect 1492 -345 1508 -311
rect 1442 -361 1508 -345
rect 1560 -311 1626 -295
rect 1560 -345 1576 -311
rect 1610 -345 1626 -311
rect 1560 -361 1626 -345
rect 1678 -311 1744 -295
rect 1678 -345 1694 -311
rect 1728 -345 1744 -311
rect 1678 -361 1744 -345
rect 1796 -311 1862 -295
rect 1796 -345 1812 -311
rect 1846 -345 1862 -311
rect 1796 -361 1862 -345
rect 1914 -311 1980 -295
rect 1914 -345 1930 -311
rect 1964 -345 1980 -311
rect 1914 -361 1980 -345
rect 2032 -311 2098 -295
rect 2032 -345 2048 -311
rect 2082 -345 2098 -311
rect 2032 -361 2098 -345
rect 2150 -311 2216 -295
rect 2150 -345 2166 -311
rect 2200 -345 2216 -311
rect 2150 -361 2216 -345
rect 2268 -311 2334 -295
rect 2268 -345 2284 -311
rect 2318 -345 2334 -311
rect 2268 -361 2334 -345
rect 2386 -311 2452 -295
rect 2386 -345 2402 -311
rect 2436 -345 2452 -311
rect 2386 -361 2452 -345
rect 2504 -311 2570 -295
rect 2504 -345 2520 -311
rect 2554 -345 2570 -311
rect 2504 -361 2570 -345
rect 2622 -311 2688 -295
rect 2622 -345 2638 -311
rect 2672 -345 2688 -311
rect 2622 -361 2688 -345
rect 2740 -311 2806 -295
rect 2740 -345 2756 -311
rect 2790 -345 2806 -311
rect 2740 -361 2806 -345
rect 2858 -311 2924 -295
rect 2858 -345 2874 -311
rect 2908 -345 2924 -311
rect 2858 -361 2924 -345
rect 2976 -311 3042 -295
rect 2976 -345 2992 -311
rect 3026 -345 3042 -311
rect 2976 -361 3042 -345
rect 3094 -311 3160 -295
rect 3094 -345 3110 -311
rect 3144 -345 3160 -311
rect 3094 -361 3160 -345
rect 3212 -311 3278 -295
rect 3212 -345 3228 -311
rect 3262 -345 3278 -311
rect 3212 -361 3278 -345
rect 3330 -311 3396 -295
rect 3330 -345 3346 -311
rect 3380 -345 3396 -311
rect 3330 -361 3396 -345
rect 3448 -311 3514 -295
rect 3448 -345 3464 -311
rect 3498 -345 3514 -311
rect 3448 -361 3514 -345
rect 3566 -311 3632 -295
rect 3566 -345 3582 -311
rect 3616 -345 3632 -311
rect 3566 -361 3632 -345
rect 3684 -311 3750 -295
rect 3684 -345 3700 -311
rect 3734 -345 3750 -311
rect 3684 -361 3750 -345
rect 3802 -311 3868 -295
rect 3802 -345 3818 -311
rect 3852 -345 3868 -311
rect 3802 -361 3868 -345
rect 3920 -311 3986 -295
rect 3920 -345 3936 -311
rect 3970 -345 3986 -311
rect 3920 -361 3986 -345
rect 4038 -311 4104 -295
rect 4038 -345 4054 -311
rect 4088 -345 4104 -311
rect 4038 -361 4104 -345
rect 4156 -311 4222 -295
rect 4156 -345 4172 -311
rect 4206 -345 4222 -311
rect 4156 -361 4222 -345
rect 4274 -311 4340 -295
rect 4274 -345 4290 -311
rect 4324 -345 4340 -311
rect 4274 -361 4340 -345
rect 4392 -311 4458 -295
rect 4392 -345 4408 -311
rect 4442 -345 4458 -311
rect 4392 -361 4458 -345
rect 4510 -311 4576 -295
rect 4510 -345 4526 -311
rect 4560 -345 4576 -311
rect 4510 -361 4576 -345
rect 4628 -311 4694 -295
rect 4628 -345 4644 -311
rect 4678 -345 4694 -311
rect 4628 -361 4694 -345
rect 4746 -311 4812 -295
rect 4746 -345 4762 -311
rect 4796 -345 4812 -311
rect 4746 -361 4812 -345
rect 4864 -311 4930 -295
rect 4864 -345 4880 -311
rect 4914 -345 4930 -311
rect 4864 -361 4930 -345
rect 4982 -311 5048 -295
rect 4982 -345 4998 -311
rect 5032 -345 5048 -311
rect 4982 -361 5048 -345
rect 5100 -311 5166 -295
rect 5100 -345 5116 -311
rect 5150 -345 5166 -311
rect 5100 -361 5166 -345
rect 5218 -311 5284 -295
rect 5218 -345 5234 -311
rect 5268 -345 5284 -311
rect 5218 -361 5284 -345
rect 5336 -311 5402 -295
rect 5336 -345 5352 -311
rect 5386 -345 5402 -311
rect 5336 -361 5402 -345
rect 5454 -311 5520 -295
rect 5454 -345 5470 -311
rect 5504 -345 5520 -311
rect 5454 -361 5520 -345
rect 5572 -311 5638 -295
rect 5572 -345 5588 -311
rect 5622 -345 5638 -311
rect 5572 -361 5638 -345
rect 5690 -311 5756 -295
rect 5690 -345 5706 -311
rect 5740 -345 5756 -311
rect 5690 -361 5756 -345
rect 5808 -311 5874 -295
rect 5808 -345 5824 -311
rect 5858 -345 5874 -311
rect 5808 -361 5874 -345
rect 5926 -311 5992 -295
rect 5926 -345 5942 -311
rect 5976 -345 5992 -311
rect 5926 -361 5992 -345
rect 6044 -311 6110 -295
rect 6044 -345 6060 -311
rect 6094 -345 6110 -311
rect 6044 -361 6110 -345
rect 6162 -311 6228 -295
rect 6162 -345 6178 -311
rect 6212 -345 6228 -311
rect 6162 -361 6228 -345
rect 6280 -311 6346 -295
rect 6280 -345 6296 -311
rect 6330 -345 6346 -311
rect 6280 -361 6346 -345
rect 6398 -311 6464 -295
rect 6398 -345 6414 -311
rect 6448 -345 6464 -311
rect 6398 -361 6464 -345
rect 6516 -311 6582 -295
rect 6516 -345 6532 -311
rect 6566 -345 6582 -311
rect 6516 -361 6582 -345
rect 6634 -311 6700 -295
rect 6634 -345 6650 -311
rect 6684 -345 6700 -311
rect 6634 -361 6700 -345
rect 6752 -311 6818 -295
rect 6752 -345 6768 -311
rect 6802 -345 6818 -311
rect 6752 -361 6818 -345
rect 6870 -311 6936 -295
rect 6870 -345 6886 -311
rect 6920 -345 6936 -311
rect 6870 -361 6936 -345
rect 6988 -311 7054 -295
rect 6988 -345 7004 -311
rect 7038 -345 7054 -311
rect 6988 -361 7054 -345
rect 7106 -311 7172 -295
rect 7106 -345 7122 -311
rect 7156 -345 7172 -311
rect 7106 -361 7172 -345
rect 7224 -311 7290 -295
rect 7224 -345 7240 -311
rect 7274 -345 7290 -311
rect 7224 -361 7290 -345
rect 7342 -311 7408 -295
rect 7342 -345 7358 -311
rect 7392 -345 7408 -311
rect 7342 -361 7408 -345
rect 7460 -311 7526 -295
rect 7460 -345 7476 -311
rect 7510 -345 7526 -311
rect 7460 -361 7526 -345
rect 7578 -311 7644 -295
rect 7578 -345 7594 -311
rect 7628 -345 7644 -311
rect 7578 -361 7644 -345
rect 7696 -311 7762 -295
rect 7696 -345 7712 -311
rect 7746 -345 7762 -311
rect 7696 -361 7762 -345
rect 7814 -311 7880 -295
rect 7814 -345 7830 -311
rect 7864 -345 7880 -311
rect 7814 -361 7880 -345
rect 7932 -311 7998 -295
rect 7932 -345 7948 -311
rect 7982 -345 7998 -311
rect 7932 -361 7998 -345
rect 8050 -311 8116 -295
rect 8050 -345 8066 -311
rect 8100 -345 8116 -311
rect 8050 -361 8116 -345
rect 8168 -311 8234 -295
rect 8168 -345 8184 -311
rect 8218 -345 8234 -311
rect 8168 -361 8234 -345
rect 8286 -311 8352 -295
rect 8286 -345 8302 -311
rect 8336 -345 8352 -311
rect 8286 -361 8352 -345
rect 8404 -311 8470 -295
rect 8404 -345 8420 -311
rect 8454 -345 8470 -311
rect 8404 -361 8470 -345
rect 8522 -311 8588 -295
rect 8522 -345 8538 -311
rect 8572 -345 8588 -311
rect 8522 -361 8588 -345
rect 8640 -311 8706 -295
rect 8640 -345 8656 -311
rect 8690 -345 8706 -311
rect 8640 -361 8706 -345
rect 8758 -311 8824 -295
rect 8758 -345 8774 -311
rect 8808 -345 8824 -311
rect 8758 -361 8824 -345
rect 8876 -311 8942 -295
rect 8876 -345 8892 -311
rect 8926 -345 8942 -311
rect 8876 -361 8942 -345
rect 8994 -311 9060 -295
rect 8994 -345 9010 -311
rect 9044 -345 9060 -311
rect 8994 -361 9060 -345
rect 9112 -311 9178 -295
rect 9112 -345 9128 -311
rect 9162 -345 9178 -311
rect 9112 -361 9178 -345
rect 9230 -311 9296 -295
rect 9230 -345 9246 -311
rect 9280 -345 9296 -311
rect 9230 -361 9296 -345
rect 9348 -311 9414 -295
rect 9348 -345 9364 -311
rect 9398 -345 9414 -311
rect 9348 -361 9414 -345
rect 9466 -311 9532 -295
rect 9466 -345 9482 -311
rect 9516 -345 9532 -311
rect 9466 -361 9532 -345
rect 9584 -311 9650 -295
rect 9584 -345 9600 -311
rect 9634 -345 9650 -311
rect 9584 -361 9650 -345
rect 9702 -311 9768 -295
rect 9702 -345 9718 -311
rect 9752 -345 9768 -311
rect 9702 -361 9768 -345
rect 9820 -311 9886 -295
rect 9820 -345 9836 -311
rect 9870 -345 9886 -311
rect 9820 -361 9886 -345
rect 9938 -311 10004 -295
rect 9938 -345 9954 -311
rect 9988 -345 10004 -311
rect 9938 -361 10004 -345
rect 10056 -311 10122 -295
rect 10056 -345 10072 -311
rect 10106 -345 10122 -311
rect 10056 -361 10122 -345
rect 10174 -311 10240 -295
rect 10174 -345 10190 -311
rect 10224 -345 10240 -311
rect 10174 -361 10240 -345
rect 10292 -311 10358 -295
rect 10292 -345 10308 -311
rect 10342 -345 10358 -311
rect 10292 -361 10358 -345
rect 10410 -311 10476 -295
rect 10410 -345 10426 -311
rect 10460 -345 10476 -311
rect 10410 -361 10476 -345
rect 10528 -311 10594 -295
rect 10528 -345 10544 -311
rect 10578 -345 10594 -311
rect 10528 -361 10594 -345
rect 10646 -311 10712 -295
rect 10646 -345 10662 -311
rect 10696 -345 10712 -311
rect 10646 -361 10712 -345
rect 10764 -311 10830 -295
rect 10764 -345 10780 -311
rect 10814 -345 10830 -311
rect 10764 -361 10830 -345
rect 10882 -311 10948 -295
rect 10882 -345 10898 -311
rect 10932 -345 10948 -311
rect 10882 -361 10948 -345
rect 11000 -311 11066 -295
rect 11000 -345 11016 -311
rect 11050 -345 11066 -311
rect 11000 -361 11066 -345
rect 11118 -311 11184 -295
rect 11118 -345 11134 -311
rect 11168 -345 11184 -311
rect 11118 -361 11184 -345
rect 11236 -311 11302 -295
rect 11236 -345 11252 -311
rect 11286 -345 11302 -311
rect 11236 -361 11302 -345
rect 11354 -311 11420 -295
rect 11354 -345 11370 -311
rect 11404 -345 11420 -311
rect 11354 -361 11420 -345
rect 11472 -311 11538 -295
rect 11472 -345 11488 -311
rect 11522 -345 11538 -311
rect 11472 -361 11538 -345
rect 11590 -311 11656 -295
rect 11590 -345 11606 -311
rect 11640 -345 11656 -311
rect 11590 -361 11656 -345
rect 11708 -311 11774 -295
rect 11708 -345 11724 -311
rect 11758 -345 11774 -311
rect 11708 -361 11774 -345
rect 11826 -311 11892 -295
rect 11826 -345 11842 -311
rect 11876 -345 11892 -311
rect 11826 -361 11892 -345
rect 11944 -311 12010 -295
rect 11944 -345 11960 -311
rect 11994 -345 12010 -311
rect 11944 -361 12010 -345
rect 12062 -311 12128 -295
rect 12062 -345 12078 -311
rect 12112 -345 12128 -311
rect 12062 -361 12128 -345
rect 12180 -311 12246 -295
rect 12180 -345 12196 -311
rect 12230 -345 12246 -311
rect 12180 -361 12246 -345
rect 12298 -311 12364 -295
rect 12298 -345 12314 -311
rect 12348 -345 12364 -311
rect 12298 -361 12364 -345
rect 12416 -311 12482 -295
rect 12416 -345 12432 -311
rect 12466 -345 12482 -311
rect 12416 -361 12482 -345
rect 12534 -311 12600 -295
rect 12534 -345 12550 -311
rect 12584 -345 12600 -311
rect 12534 -361 12600 -345
rect 12652 -311 12718 -295
rect 12652 -345 12668 -311
rect 12702 -345 12718 -311
rect 12652 -361 12718 -345
rect 12770 -311 12836 -295
rect 12770 -345 12786 -311
rect 12820 -345 12836 -311
rect 12770 -361 12836 -345
rect 12888 -311 12954 -295
rect 12888 -345 12904 -311
rect 12938 -345 12954 -311
rect 12888 -361 12954 -345
rect 13006 -311 13072 -295
rect 13006 -345 13022 -311
rect 13056 -345 13072 -311
rect 13006 -361 13072 -345
rect 13124 -311 13190 -295
rect 13124 -345 13140 -311
rect 13174 -345 13190 -311
rect 13124 -361 13190 -345
rect 13242 -311 13308 -295
rect 13242 -345 13258 -311
rect 13292 -345 13308 -311
rect 13242 -361 13308 -345
rect 13360 -311 13426 -295
rect 13360 -345 13376 -311
rect 13410 -345 13426 -311
rect 13360 -361 13426 -345
rect 13478 -311 13544 -295
rect 13478 -345 13494 -311
rect 13528 -345 13544 -311
rect 13478 -361 13544 -345
rect 13596 -311 13662 -295
rect 13596 -345 13612 -311
rect 13646 -345 13662 -311
rect 13596 -361 13662 -345
rect 13714 -311 13780 -295
rect 13714 -345 13730 -311
rect 13764 -345 13780 -311
rect 13714 -361 13780 -345
rect 13832 -311 13898 -295
rect 13832 -345 13848 -311
rect 13882 -345 13898 -311
rect 13832 -361 13898 -345
rect 13950 -311 14016 -295
rect 13950 -345 13966 -311
rect 14000 -345 14016 -311
rect 13950 -361 14016 -345
rect 14068 -311 14134 -295
rect 14068 -345 14084 -311
rect 14118 -345 14134 -311
rect 14068 -361 14134 -345
rect 14186 -311 14252 -295
rect 14186 -345 14202 -311
rect 14236 -345 14252 -311
rect 14186 -361 14252 -345
rect 14304 -311 14370 -295
rect 14304 -345 14320 -311
rect 14354 -345 14370 -311
rect 14304 -361 14370 -345
rect 14422 -311 14488 -295
rect 14422 -345 14438 -311
rect 14472 -345 14488 -311
rect 14422 -361 14488 -345
rect 14540 -311 14606 -295
rect 14540 -345 14556 -311
rect 14590 -345 14606 -311
rect 14540 -361 14606 -345
rect 14658 -311 14724 -295
rect 14658 -345 14674 -311
rect 14708 -345 14724 -311
rect 14658 -361 14724 -345
<< polycont >>
rect -14708 -345 -14674 -311
rect -14590 -345 -14556 -311
rect -14472 -345 -14438 -311
rect -14354 -345 -14320 -311
rect -14236 -345 -14202 -311
rect -14118 -345 -14084 -311
rect -14000 -345 -13966 -311
rect -13882 -345 -13848 -311
rect -13764 -345 -13730 -311
rect -13646 -345 -13612 -311
rect -13528 -345 -13494 -311
rect -13410 -345 -13376 -311
rect -13292 -345 -13258 -311
rect -13174 -345 -13140 -311
rect -13056 -345 -13022 -311
rect -12938 -345 -12904 -311
rect -12820 -345 -12786 -311
rect -12702 -345 -12668 -311
rect -12584 -345 -12550 -311
rect -12466 -345 -12432 -311
rect -12348 -345 -12314 -311
rect -12230 -345 -12196 -311
rect -12112 -345 -12078 -311
rect -11994 -345 -11960 -311
rect -11876 -345 -11842 -311
rect -11758 -345 -11724 -311
rect -11640 -345 -11606 -311
rect -11522 -345 -11488 -311
rect -11404 -345 -11370 -311
rect -11286 -345 -11252 -311
rect -11168 -345 -11134 -311
rect -11050 -345 -11016 -311
rect -10932 -345 -10898 -311
rect -10814 -345 -10780 -311
rect -10696 -345 -10662 -311
rect -10578 -345 -10544 -311
rect -10460 -345 -10426 -311
rect -10342 -345 -10308 -311
rect -10224 -345 -10190 -311
rect -10106 -345 -10072 -311
rect -9988 -345 -9954 -311
rect -9870 -345 -9836 -311
rect -9752 -345 -9718 -311
rect -9634 -345 -9600 -311
rect -9516 -345 -9482 -311
rect -9398 -345 -9364 -311
rect -9280 -345 -9246 -311
rect -9162 -345 -9128 -311
rect -9044 -345 -9010 -311
rect -8926 -345 -8892 -311
rect -8808 -345 -8774 -311
rect -8690 -345 -8656 -311
rect -8572 -345 -8538 -311
rect -8454 -345 -8420 -311
rect -8336 -345 -8302 -311
rect -8218 -345 -8184 -311
rect -8100 -345 -8066 -311
rect -7982 -345 -7948 -311
rect -7864 -345 -7830 -311
rect -7746 -345 -7712 -311
rect -7628 -345 -7594 -311
rect -7510 -345 -7476 -311
rect -7392 -345 -7358 -311
rect -7274 -345 -7240 -311
rect -7156 -345 -7122 -311
rect -7038 -345 -7004 -311
rect -6920 -345 -6886 -311
rect -6802 -345 -6768 -311
rect -6684 -345 -6650 -311
rect -6566 -345 -6532 -311
rect -6448 -345 -6414 -311
rect -6330 -345 -6296 -311
rect -6212 -345 -6178 -311
rect -6094 -345 -6060 -311
rect -5976 -345 -5942 -311
rect -5858 -345 -5824 -311
rect -5740 -345 -5706 -311
rect -5622 -345 -5588 -311
rect -5504 -345 -5470 -311
rect -5386 -345 -5352 -311
rect -5268 -345 -5234 -311
rect -5150 -345 -5116 -311
rect -5032 -345 -4998 -311
rect -4914 -345 -4880 -311
rect -4796 -345 -4762 -311
rect -4678 -345 -4644 -311
rect -4560 -345 -4526 -311
rect -4442 -345 -4408 -311
rect -4324 -345 -4290 -311
rect -4206 -345 -4172 -311
rect -4088 -345 -4054 -311
rect -3970 -345 -3936 -311
rect -3852 -345 -3818 -311
rect -3734 -345 -3700 -311
rect -3616 -345 -3582 -311
rect -3498 -345 -3464 -311
rect -3380 -345 -3346 -311
rect -3262 -345 -3228 -311
rect -3144 -345 -3110 -311
rect -3026 -345 -2992 -311
rect -2908 -345 -2874 -311
rect -2790 -345 -2756 -311
rect -2672 -345 -2638 -311
rect -2554 -345 -2520 -311
rect -2436 -345 -2402 -311
rect -2318 -345 -2284 -311
rect -2200 -345 -2166 -311
rect -2082 -345 -2048 -311
rect -1964 -345 -1930 -311
rect -1846 -345 -1812 -311
rect -1728 -345 -1694 -311
rect -1610 -345 -1576 -311
rect -1492 -345 -1458 -311
rect -1374 -345 -1340 -311
rect -1256 -345 -1222 -311
rect -1138 -345 -1104 -311
rect -1020 -345 -986 -311
rect -902 -345 -868 -311
rect -784 -345 -750 -311
rect -666 -345 -632 -311
rect -548 -345 -514 -311
rect -430 -345 -396 -311
rect -312 -345 -278 -311
rect -194 -345 -160 -311
rect -76 -345 -42 -311
rect 42 -345 76 -311
rect 160 -345 194 -311
rect 278 -345 312 -311
rect 396 -345 430 -311
rect 514 -345 548 -311
rect 632 -345 666 -311
rect 750 -345 784 -311
rect 868 -345 902 -311
rect 986 -345 1020 -311
rect 1104 -345 1138 -311
rect 1222 -345 1256 -311
rect 1340 -345 1374 -311
rect 1458 -345 1492 -311
rect 1576 -345 1610 -311
rect 1694 -345 1728 -311
rect 1812 -345 1846 -311
rect 1930 -345 1964 -311
rect 2048 -345 2082 -311
rect 2166 -345 2200 -311
rect 2284 -345 2318 -311
rect 2402 -345 2436 -311
rect 2520 -345 2554 -311
rect 2638 -345 2672 -311
rect 2756 -345 2790 -311
rect 2874 -345 2908 -311
rect 2992 -345 3026 -311
rect 3110 -345 3144 -311
rect 3228 -345 3262 -311
rect 3346 -345 3380 -311
rect 3464 -345 3498 -311
rect 3582 -345 3616 -311
rect 3700 -345 3734 -311
rect 3818 -345 3852 -311
rect 3936 -345 3970 -311
rect 4054 -345 4088 -311
rect 4172 -345 4206 -311
rect 4290 -345 4324 -311
rect 4408 -345 4442 -311
rect 4526 -345 4560 -311
rect 4644 -345 4678 -311
rect 4762 -345 4796 -311
rect 4880 -345 4914 -311
rect 4998 -345 5032 -311
rect 5116 -345 5150 -311
rect 5234 -345 5268 -311
rect 5352 -345 5386 -311
rect 5470 -345 5504 -311
rect 5588 -345 5622 -311
rect 5706 -345 5740 -311
rect 5824 -345 5858 -311
rect 5942 -345 5976 -311
rect 6060 -345 6094 -311
rect 6178 -345 6212 -311
rect 6296 -345 6330 -311
rect 6414 -345 6448 -311
rect 6532 -345 6566 -311
rect 6650 -345 6684 -311
rect 6768 -345 6802 -311
rect 6886 -345 6920 -311
rect 7004 -345 7038 -311
rect 7122 -345 7156 -311
rect 7240 -345 7274 -311
rect 7358 -345 7392 -311
rect 7476 -345 7510 -311
rect 7594 -345 7628 -311
rect 7712 -345 7746 -311
rect 7830 -345 7864 -311
rect 7948 -345 7982 -311
rect 8066 -345 8100 -311
rect 8184 -345 8218 -311
rect 8302 -345 8336 -311
rect 8420 -345 8454 -311
rect 8538 -345 8572 -311
rect 8656 -345 8690 -311
rect 8774 -345 8808 -311
rect 8892 -345 8926 -311
rect 9010 -345 9044 -311
rect 9128 -345 9162 -311
rect 9246 -345 9280 -311
rect 9364 -345 9398 -311
rect 9482 -345 9516 -311
rect 9600 -345 9634 -311
rect 9718 -345 9752 -311
rect 9836 -345 9870 -311
rect 9954 -345 9988 -311
rect 10072 -345 10106 -311
rect 10190 -345 10224 -311
rect 10308 -345 10342 -311
rect 10426 -345 10460 -311
rect 10544 -345 10578 -311
rect 10662 -345 10696 -311
rect 10780 -345 10814 -311
rect 10898 -345 10932 -311
rect 11016 -345 11050 -311
rect 11134 -345 11168 -311
rect 11252 -345 11286 -311
rect 11370 -345 11404 -311
rect 11488 -345 11522 -311
rect 11606 -345 11640 -311
rect 11724 -345 11758 -311
rect 11842 -345 11876 -311
rect 11960 -345 11994 -311
rect 12078 -345 12112 -311
rect 12196 -345 12230 -311
rect 12314 -345 12348 -311
rect 12432 -345 12466 -311
rect 12550 -345 12584 -311
rect 12668 -345 12702 -311
rect 12786 -345 12820 -311
rect 12904 -345 12938 -311
rect 13022 -345 13056 -311
rect 13140 -345 13174 -311
rect 13258 -345 13292 -311
rect 13376 -345 13410 -311
rect 13494 -345 13528 -311
rect 13612 -345 13646 -311
rect 13730 -345 13764 -311
rect 13848 -345 13882 -311
rect 13966 -345 14000 -311
rect 14084 -345 14118 -311
rect 14202 -345 14236 -311
rect 14320 -345 14354 -311
rect 14438 -345 14472 -311
rect 14556 -345 14590 -311
rect 14674 -345 14708 -311
<< locali >>
rect -14881 414 -14785 448
rect 14785 414 14881 448
rect -14881 351 -14847 414
rect 14847 351 14881 414
rect -14767 324 -14733 340
rect -14767 -268 -14733 -252
rect -14649 324 -14615 340
rect -14649 -268 -14615 -252
rect -14531 324 -14497 340
rect -14531 -268 -14497 -252
rect -14413 324 -14379 340
rect -14413 -268 -14379 -252
rect -14295 324 -14261 340
rect -14295 -268 -14261 -252
rect -14177 324 -14143 340
rect -14177 -268 -14143 -252
rect -14059 324 -14025 340
rect -14059 -268 -14025 -252
rect -13941 324 -13907 340
rect -13941 -268 -13907 -252
rect -13823 324 -13789 340
rect -13823 -268 -13789 -252
rect -13705 324 -13671 340
rect -13705 -268 -13671 -252
rect -13587 324 -13553 340
rect -13587 -268 -13553 -252
rect -13469 324 -13435 340
rect -13469 -268 -13435 -252
rect -13351 324 -13317 340
rect -13351 -268 -13317 -252
rect -13233 324 -13199 340
rect -13233 -268 -13199 -252
rect -13115 324 -13081 340
rect -13115 -268 -13081 -252
rect -12997 324 -12963 340
rect -12997 -268 -12963 -252
rect -12879 324 -12845 340
rect -12879 -268 -12845 -252
rect -12761 324 -12727 340
rect -12761 -268 -12727 -252
rect -12643 324 -12609 340
rect -12643 -268 -12609 -252
rect -12525 324 -12491 340
rect -12525 -268 -12491 -252
rect -12407 324 -12373 340
rect -12407 -268 -12373 -252
rect -12289 324 -12255 340
rect -12289 -268 -12255 -252
rect -12171 324 -12137 340
rect -12171 -268 -12137 -252
rect -12053 324 -12019 340
rect -12053 -268 -12019 -252
rect -11935 324 -11901 340
rect -11935 -268 -11901 -252
rect -11817 324 -11783 340
rect -11817 -268 -11783 -252
rect -11699 324 -11665 340
rect -11699 -268 -11665 -252
rect -11581 324 -11547 340
rect -11581 -268 -11547 -252
rect -11463 324 -11429 340
rect -11463 -268 -11429 -252
rect -11345 324 -11311 340
rect -11345 -268 -11311 -252
rect -11227 324 -11193 340
rect -11227 -268 -11193 -252
rect -11109 324 -11075 340
rect -11109 -268 -11075 -252
rect -10991 324 -10957 340
rect -10991 -268 -10957 -252
rect -10873 324 -10839 340
rect -10873 -268 -10839 -252
rect -10755 324 -10721 340
rect -10755 -268 -10721 -252
rect -10637 324 -10603 340
rect -10637 -268 -10603 -252
rect -10519 324 -10485 340
rect -10519 -268 -10485 -252
rect -10401 324 -10367 340
rect -10401 -268 -10367 -252
rect -10283 324 -10249 340
rect -10283 -268 -10249 -252
rect -10165 324 -10131 340
rect -10165 -268 -10131 -252
rect -10047 324 -10013 340
rect -10047 -268 -10013 -252
rect -9929 324 -9895 340
rect -9929 -268 -9895 -252
rect -9811 324 -9777 340
rect -9811 -268 -9777 -252
rect -9693 324 -9659 340
rect -9693 -268 -9659 -252
rect -9575 324 -9541 340
rect -9575 -268 -9541 -252
rect -9457 324 -9423 340
rect -9457 -268 -9423 -252
rect -9339 324 -9305 340
rect -9339 -268 -9305 -252
rect -9221 324 -9187 340
rect -9221 -268 -9187 -252
rect -9103 324 -9069 340
rect -9103 -268 -9069 -252
rect -8985 324 -8951 340
rect -8985 -268 -8951 -252
rect -8867 324 -8833 340
rect -8867 -268 -8833 -252
rect -8749 324 -8715 340
rect -8749 -268 -8715 -252
rect -8631 324 -8597 340
rect -8631 -268 -8597 -252
rect -8513 324 -8479 340
rect -8513 -268 -8479 -252
rect -8395 324 -8361 340
rect -8395 -268 -8361 -252
rect -8277 324 -8243 340
rect -8277 -268 -8243 -252
rect -8159 324 -8125 340
rect -8159 -268 -8125 -252
rect -8041 324 -8007 340
rect -8041 -268 -8007 -252
rect -7923 324 -7889 340
rect -7923 -268 -7889 -252
rect -7805 324 -7771 340
rect -7805 -268 -7771 -252
rect -7687 324 -7653 340
rect -7687 -268 -7653 -252
rect -7569 324 -7535 340
rect -7569 -268 -7535 -252
rect -7451 324 -7417 340
rect -7451 -268 -7417 -252
rect -7333 324 -7299 340
rect -7333 -268 -7299 -252
rect -7215 324 -7181 340
rect -7215 -268 -7181 -252
rect -7097 324 -7063 340
rect -7097 -268 -7063 -252
rect -6979 324 -6945 340
rect -6979 -268 -6945 -252
rect -6861 324 -6827 340
rect -6861 -268 -6827 -252
rect -6743 324 -6709 340
rect -6743 -268 -6709 -252
rect -6625 324 -6591 340
rect -6625 -268 -6591 -252
rect -6507 324 -6473 340
rect -6507 -268 -6473 -252
rect -6389 324 -6355 340
rect -6389 -268 -6355 -252
rect -6271 324 -6237 340
rect -6271 -268 -6237 -252
rect -6153 324 -6119 340
rect -6153 -268 -6119 -252
rect -6035 324 -6001 340
rect -6035 -268 -6001 -252
rect -5917 324 -5883 340
rect -5917 -268 -5883 -252
rect -5799 324 -5765 340
rect -5799 -268 -5765 -252
rect -5681 324 -5647 340
rect -5681 -268 -5647 -252
rect -5563 324 -5529 340
rect -5563 -268 -5529 -252
rect -5445 324 -5411 340
rect -5445 -268 -5411 -252
rect -5327 324 -5293 340
rect -5327 -268 -5293 -252
rect -5209 324 -5175 340
rect -5209 -268 -5175 -252
rect -5091 324 -5057 340
rect -5091 -268 -5057 -252
rect -4973 324 -4939 340
rect -4973 -268 -4939 -252
rect -4855 324 -4821 340
rect -4855 -268 -4821 -252
rect -4737 324 -4703 340
rect -4737 -268 -4703 -252
rect -4619 324 -4585 340
rect -4619 -268 -4585 -252
rect -4501 324 -4467 340
rect -4501 -268 -4467 -252
rect -4383 324 -4349 340
rect -4383 -268 -4349 -252
rect -4265 324 -4231 340
rect -4265 -268 -4231 -252
rect -4147 324 -4113 340
rect -4147 -268 -4113 -252
rect -4029 324 -3995 340
rect -4029 -268 -3995 -252
rect -3911 324 -3877 340
rect -3911 -268 -3877 -252
rect -3793 324 -3759 340
rect -3793 -268 -3759 -252
rect -3675 324 -3641 340
rect -3675 -268 -3641 -252
rect -3557 324 -3523 340
rect -3557 -268 -3523 -252
rect -3439 324 -3405 340
rect -3439 -268 -3405 -252
rect -3321 324 -3287 340
rect -3321 -268 -3287 -252
rect -3203 324 -3169 340
rect -3203 -268 -3169 -252
rect -3085 324 -3051 340
rect -3085 -268 -3051 -252
rect -2967 324 -2933 340
rect -2967 -268 -2933 -252
rect -2849 324 -2815 340
rect -2849 -268 -2815 -252
rect -2731 324 -2697 340
rect -2731 -268 -2697 -252
rect -2613 324 -2579 340
rect -2613 -268 -2579 -252
rect -2495 324 -2461 340
rect -2495 -268 -2461 -252
rect -2377 324 -2343 340
rect -2377 -268 -2343 -252
rect -2259 324 -2225 340
rect -2259 -268 -2225 -252
rect -2141 324 -2107 340
rect -2141 -268 -2107 -252
rect -2023 324 -1989 340
rect -2023 -268 -1989 -252
rect -1905 324 -1871 340
rect -1905 -268 -1871 -252
rect -1787 324 -1753 340
rect -1787 -268 -1753 -252
rect -1669 324 -1635 340
rect -1669 -268 -1635 -252
rect -1551 324 -1517 340
rect -1551 -268 -1517 -252
rect -1433 324 -1399 340
rect -1433 -268 -1399 -252
rect -1315 324 -1281 340
rect -1315 -268 -1281 -252
rect -1197 324 -1163 340
rect -1197 -268 -1163 -252
rect -1079 324 -1045 340
rect -1079 -268 -1045 -252
rect -961 324 -927 340
rect -961 -268 -927 -252
rect -843 324 -809 340
rect -843 -268 -809 -252
rect -725 324 -691 340
rect -725 -268 -691 -252
rect -607 324 -573 340
rect -607 -268 -573 -252
rect -489 324 -455 340
rect -489 -268 -455 -252
rect -371 324 -337 340
rect -371 -268 -337 -252
rect -253 324 -219 340
rect -253 -268 -219 -252
rect -135 324 -101 340
rect -135 -268 -101 -252
rect -17 324 17 340
rect -17 -268 17 -252
rect 101 324 135 340
rect 101 -268 135 -252
rect 219 324 253 340
rect 219 -268 253 -252
rect 337 324 371 340
rect 337 -268 371 -252
rect 455 324 489 340
rect 455 -268 489 -252
rect 573 324 607 340
rect 573 -268 607 -252
rect 691 324 725 340
rect 691 -268 725 -252
rect 809 324 843 340
rect 809 -268 843 -252
rect 927 324 961 340
rect 927 -268 961 -252
rect 1045 324 1079 340
rect 1045 -268 1079 -252
rect 1163 324 1197 340
rect 1163 -268 1197 -252
rect 1281 324 1315 340
rect 1281 -268 1315 -252
rect 1399 324 1433 340
rect 1399 -268 1433 -252
rect 1517 324 1551 340
rect 1517 -268 1551 -252
rect 1635 324 1669 340
rect 1635 -268 1669 -252
rect 1753 324 1787 340
rect 1753 -268 1787 -252
rect 1871 324 1905 340
rect 1871 -268 1905 -252
rect 1989 324 2023 340
rect 1989 -268 2023 -252
rect 2107 324 2141 340
rect 2107 -268 2141 -252
rect 2225 324 2259 340
rect 2225 -268 2259 -252
rect 2343 324 2377 340
rect 2343 -268 2377 -252
rect 2461 324 2495 340
rect 2461 -268 2495 -252
rect 2579 324 2613 340
rect 2579 -268 2613 -252
rect 2697 324 2731 340
rect 2697 -268 2731 -252
rect 2815 324 2849 340
rect 2815 -268 2849 -252
rect 2933 324 2967 340
rect 2933 -268 2967 -252
rect 3051 324 3085 340
rect 3051 -268 3085 -252
rect 3169 324 3203 340
rect 3169 -268 3203 -252
rect 3287 324 3321 340
rect 3287 -268 3321 -252
rect 3405 324 3439 340
rect 3405 -268 3439 -252
rect 3523 324 3557 340
rect 3523 -268 3557 -252
rect 3641 324 3675 340
rect 3641 -268 3675 -252
rect 3759 324 3793 340
rect 3759 -268 3793 -252
rect 3877 324 3911 340
rect 3877 -268 3911 -252
rect 3995 324 4029 340
rect 3995 -268 4029 -252
rect 4113 324 4147 340
rect 4113 -268 4147 -252
rect 4231 324 4265 340
rect 4231 -268 4265 -252
rect 4349 324 4383 340
rect 4349 -268 4383 -252
rect 4467 324 4501 340
rect 4467 -268 4501 -252
rect 4585 324 4619 340
rect 4585 -268 4619 -252
rect 4703 324 4737 340
rect 4703 -268 4737 -252
rect 4821 324 4855 340
rect 4821 -268 4855 -252
rect 4939 324 4973 340
rect 4939 -268 4973 -252
rect 5057 324 5091 340
rect 5057 -268 5091 -252
rect 5175 324 5209 340
rect 5175 -268 5209 -252
rect 5293 324 5327 340
rect 5293 -268 5327 -252
rect 5411 324 5445 340
rect 5411 -268 5445 -252
rect 5529 324 5563 340
rect 5529 -268 5563 -252
rect 5647 324 5681 340
rect 5647 -268 5681 -252
rect 5765 324 5799 340
rect 5765 -268 5799 -252
rect 5883 324 5917 340
rect 5883 -268 5917 -252
rect 6001 324 6035 340
rect 6001 -268 6035 -252
rect 6119 324 6153 340
rect 6119 -268 6153 -252
rect 6237 324 6271 340
rect 6237 -268 6271 -252
rect 6355 324 6389 340
rect 6355 -268 6389 -252
rect 6473 324 6507 340
rect 6473 -268 6507 -252
rect 6591 324 6625 340
rect 6591 -268 6625 -252
rect 6709 324 6743 340
rect 6709 -268 6743 -252
rect 6827 324 6861 340
rect 6827 -268 6861 -252
rect 6945 324 6979 340
rect 6945 -268 6979 -252
rect 7063 324 7097 340
rect 7063 -268 7097 -252
rect 7181 324 7215 340
rect 7181 -268 7215 -252
rect 7299 324 7333 340
rect 7299 -268 7333 -252
rect 7417 324 7451 340
rect 7417 -268 7451 -252
rect 7535 324 7569 340
rect 7535 -268 7569 -252
rect 7653 324 7687 340
rect 7653 -268 7687 -252
rect 7771 324 7805 340
rect 7771 -268 7805 -252
rect 7889 324 7923 340
rect 7889 -268 7923 -252
rect 8007 324 8041 340
rect 8007 -268 8041 -252
rect 8125 324 8159 340
rect 8125 -268 8159 -252
rect 8243 324 8277 340
rect 8243 -268 8277 -252
rect 8361 324 8395 340
rect 8361 -268 8395 -252
rect 8479 324 8513 340
rect 8479 -268 8513 -252
rect 8597 324 8631 340
rect 8597 -268 8631 -252
rect 8715 324 8749 340
rect 8715 -268 8749 -252
rect 8833 324 8867 340
rect 8833 -268 8867 -252
rect 8951 324 8985 340
rect 8951 -268 8985 -252
rect 9069 324 9103 340
rect 9069 -268 9103 -252
rect 9187 324 9221 340
rect 9187 -268 9221 -252
rect 9305 324 9339 340
rect 9305 -268 9339 -252
rect 9423 324 9457 340
rect 9423 -268 9457 -252
rect 9541 324 9575 340
rect 9541 -268 9575 -252
rect 9659 324 9693 340
rect 9659 -268 9693 -252
rect 9777 324 9811 340
rect 9777 -268 9811 -252
rect 9895 324 9929 340
rect 9895 -268 9929 -252
rect 10013 324 10047 340
rect 10013 -268 10047 -252
rect 10131 324 10165 340
rect 10131 -268 10165 -252
rect 10249 324 10283 340
rect 10249 -268 10283 -252
rect 10367 324 10401 340
rect 10367 -268 10401 -252
rect 10485 324 10519 340
rect 10485 -268 10519 -252
rect 10603 324 10637 340
rect 10603 -268 10637 -252
rect 10721 324 10755 340
rect 10721 -268 10755 -252
rect 10839 324 10873 340
rect 10839 -268 10873 -252
rect 10957 324 10991 340
rect 10957 -268 10991 -252
rect 11075 324 11109 340
rect 11075 -268 11109 -252
rect 11193 324 11227 340
rect 11193 -268 11227 -252
rect 11311 324 11345 340
rect 11311 -268 11345 -252
rect 11429 324 11463 340
rect 11429 -268 11463 -252
rect 11547 324 11581 340
rect 11547 -268 11581 -252
rect 11665 324 11699 340
rect 11665 -268 11699 -252
rect 11783 324 11817 340
rect 11783 -268 11817 -252
rect 11901 324 11935 340
rect 11901 -268 11935 -252
rect 12019 324 12053 340
rect 12019 -268 12053 -252
rect 12137 324 12171 340
rect 12137 -268 12171 -252
rect 12255 324 12289 340
rect 12255 -268 12289 -252
rect 12373 324 12407 340
rect 12373 -268 12407 -252
rect 12491 324 12525 340
rect 12491 -268 12525 -252
rect 12609 324 12643 340
rect 12609 -268 12643 -252
rect 12727 324 12761 340
rect 12727 -268 12761 -252
rect 12845 324 12879 340
rect 12845 -268 12879 -252
rect 12963 324 12997 340
rect 12963 -268 12997 -252
rect 13081 324 13115 340
rect 13081 -268 13115 -252
rect 13199 324 13233 340
rect 13199 -268 13233 -252
rect 13317 324 13351 340
rect 13317 -268 13351 -252
rect 13435 324 13469 340
rect 13435 -268 13469 -252
rect 13553 324 13587 340
rect 13553 -268 13587 -252
rect 13671 324 13705 340
rect 13671 -268 13705 -252
rect 13789 324 13823 340
rect 13789 -268 13823 -252
rect 13907 324 13941 340
rect 13907 -268 13941 -252
rect 14025 324 14059 340
rect 14025 -268 14059 -252
rect 14143 324 14177 340
rect 14143 -268 14177 -252
rect 14261 324 14295 340
rect 14261 -268 14295 -252
rect 14379 324 14413 340
rect 14379 -268 14413 -252
rect 14497 324 14531 340
rect 14497 -268 14531 -252
rect 14615 324 14649 340
rect 14615 -268 14649 -252
rect 14733 324 14767 340
rect 14733 -268 14767 -252
rect -14724 -345 -14708 -311
rect -14674 -345 -14658 -311
rect -14606 -345 -14590 -311
rect -14556 -345 -14540 -311
rect -14488 -345 -14472 -311
rect -14438 -345 -14422 -311
rect -14370 -345 -14354 -311
rect -14320 -345 -14304 -311
rect -14252 -345 -14236 -311
rect -14202 -345 -14186 -311
rect -14134 -345 -14118 -311
rect -14084 -345 -14068 -311
rect -14016 -345 -14000 -311
rect -13966 -345 -13950 -311
rect -13898 -345 -13882 -311
rect -13848 -345 -13832 -311
rect -13780 -345 -13764 -311
rect -13730 -345 -13714 -311
rect -13662 -345 -13646 -311
rect -13612 -345 -13596 -311
rect -13544 -345 -13528 -311
rect -13494 -345 -13478 -311
rect -13426 -345 -13410 -311
rect -13376 -345 -13360 -311
rect -13308 -345 -13292 -311
rect -13258 -345 -13242 -311
rect -13190 -345 -13174 -311
rect -13140 -345 -13124 -311
rect -13072 -345 -13056 -311
rect -13022 -345 -13006 -311
rect -12954 -345 -12938 -311
rect -12904 -345 -12888 -311
rect -12836 -345 -12820 -311
rect -12786 -345 -12770 -311
rect -12718 -345 -12702 -311
rect -12668 -345 -12652 -311
rect -12600 -345 -12584 -311
rect -12550 -345 -12534 -311
rect -12482 -345 -12466 -311
rect -12432 -345 -12416 -311
rect -12364 -345 -12348 -311
rect -12314 -345 -12298 -311
rect -12246 -345 -12230 -311
rect -12196 -345 -12180 -311
rect -12128 -345 -12112 -311
rect -12078 -345 -12062 -311
rect -12010 -345 -11994 -311
rect -11960 -345 -11944 -311
rect -11892 -345 -11876 -311
rect -11842 -345 -11826 -311
rect -11774 -345 -11758 -311
rect -11724 -345 -11708 -311
rect -11656 -345 -11640 -311
rect -11606 -345 -11590 -311
rect -11538 -345 -11522 -311
rect -11488 -345 -11472 -311
rect -11420 -345 -11404 -311
rect -11370 -345 -11354 -311
rect -11302 -345 -11286 -311
rect -11252 -345 -11236 -311
rect -11184 -345 -11168 -311
rect -11134 -345 -11118 -311
rect -11066 -345 -11050 -311
rect -11016 -345 -11000 -311
rect -10948 -345 -10932 -311
rect -10898 -345 -10882 -311
rect -10830 -345 -10814 -311
rect -10780 -345 -10764 -311
rect -10712 -345 -10696 -311
rect -10662 -345 -10646 -311
rect -10594 -345 -10578 -311
rect -10544 -345 -10528 -311
rect -10476 -345 -10460 -311
rect -10426 -345 -10410 -311
rect -10358 -345 -10342 -311
rect -10308 -345 -10292 -311
rect -10240 -345 -10224 -311
rect -10190 -345 -10174 -311
rect -10122 -345 -10106 -311
rect -10072 -345 -10056 -311
rect -10004 -345 -9988 -311
rect -9954 -345 -9938 -311
rect -9886 -345 -9870 -311
rect -9836 -345 -9820 -311
rect -9768 -345 -9752 -311
rect -9718 -345 -9702 -311
rect -9650 -345 -9634 -311
rect -9600 -345 -9584 -311
rect -9532 -345 -9516 -311
rect -9482 -345 -9466 -311
rect -9414 -345 -9398 -311
rect -9364 -345 -9348 -311
rect -9296 -345 -9280 -311
rect -9246 -345 -9230 -311
rect -9178 -345 -9162 -311
rect -9128 -345 -9112 -311
rect -9060 -345 -9044 -311
rect -9010 -345 -8994 -311
rect -8942 -345 -8926 -311
rect -8892 -345 -8876 -311
rect -8824 -345 -8808 -311
rect -8774 -345 -8758 -311
rect -8706 -345 -8690 -311
rect -8656 -345 -8640 -311
rect -8588 -345 -8572 -311
rect -8538 -345 -8522 -311
rect -8470 -345 -8454 -311
rect -8420 -345 -8404 -311
rect -8352 -345 -8336 -311
rect -8302 -345 -8286 -311
rect -8234 -345 -8218 -311
rect -8184 -345 -8168 -311
rect -8116 -345 -8100 -311
rect -8066 -345 -8050 -311
rect -7998 -345 -7982 -311
rect -7948 -345 -7932 -311
rect -7880 -345 -7864 -311
rect -7830 -345 -7814 -311
rect -7762 -345 -7746 -311
rect -7712 -345 -7696 -311
rect -7644 -345 -7628 -311
rect -7594 -345 -7578 -311
rect -7526 -345 -7510 -311
rect -7476 -345 -7460 -311
rect -7408 -345 -7392 -311
rect -7358 -345 -7342 -311
rect -7290 -345 -7274 -311
rect -7240 -345 -7224 -311
rect -7172 -345 -7156 -311
rect -7122 -345 -7106 -311
rect -7054 -345 -7038 -311
rect -7004 -345 -6988 -311
rect -6936 -345 -6920 -311
rect -6886 -345 -6870 -311
rect -6818 -345 -6802 -311
rect -6768 -345 -6752 -311
rect -6700 -345 -6684 -311
rect -6650 -345 -6634 -311
rect -6582 -345 -6566 -311
rect -6532 -345 -6516 -311
rect -6464 -345 -6448 -311
rect -6414 -345 -6398 -311
rect -6346 -345 -6330 -311
rect -6296 -345 -6280 -311
rect -6228 -345 -6212 -311
rect -6178 -345 -6162 -311
rect -6110 -345 -6094 -311
rect -6060 -345 -6044 -311
rect -5992 -345 -5976 -311
rect -5942 -345 -5926 -311
rect -5874 -345 -5858 -311
rect -5824 -345 -5808 -311
rect -5756 -345 -5740 -311
rect -5706 -345 -5690 -311
rect -5638 -345 -5622 -311
rect -5588 -345 -5572 -311
rect -5520 -345 -5504 -311
rect -5470 -345 -5454 -311
rect -5402 -345 -5386 -311
rect -5352 -345 -5336 -311
rect -5284 -345 -5268 -311
rect -5234 -345 -5218 -311
rect -5166 -345 -5150 -311
rect -5116 -345 -5100 -311
rect -5048 -345 -5032 -311
rect -4998 -345 -4982 -311
rect -4930 -345 -4914 -311
rect -4880 -345 -4864 -311
rect -4812 -345 -4796 -311
rect -4762 -345 -4746 -311
rect -4694 -345 -4678 -311
rect -4644 -345 -4628 -311
rect -4576 -345 -4560 -311
rect -4526 -345 -4510 -311
rect -4458 -345 -4442 -311
rect -4408 -345 -4392 -311
rect -4340 -345 -4324 -311
rect -4290 -345 -4274 -311
rect -4222 -345 -4206 -311
rect -4172 -345 -4156 -311
rect -4104 -345 -4088 -311
rect -4054 -345 -4038 -311
rect -3986 -345 -3970 -311
rect -3936 -345 -3920 -311
rect -3868 -345 -3852 -311
rect -3818 -345 -3802 -311
rect -3750 -345 -3734 -311
rect -3700 -345 -3684 -311
rect -3632 -345 -3616 -311
rect -3582 -345 -3566 -311
rect -3514 -345 -3498 -311
rect -3464 -345 -3448 -311
rect -3396 -345 -3380 -311
rect -3346 -345 -3330 -311
rect -3278 -345 -3262 -311
rect -3228 -345 -3212 -311
rect -3160 -345 -3144 -311
rect -3110 -345 -3094 -311
rect -3042 -345 -3026 -311
rect -2992 -345 -2976 -311
rect -2924 -345 -2908 -311
rect -2874 -345 -2858 -311
rect -2806 -345 -2790 -311
rect -2756 -345 -2740 -311
rect -2688 -345 -2672 -311
rect -2638 -345 -2622 -311
rect -2570 -345 -2554 -311
rect -2520 -345 -2504 -311
rect -2452 -345 -2436 -311
rect -2402 -345 -2386 -311
rect -2334 -345 -2318 -311
rect -2284 -345 -2268 -311
rect -2216 -345 -2200 -311
rect -2166 -345 -2150 -311
rect -2098 -345 -2082 -311
rect -2048 -345 -2032 -311
rect -1980 -345 -1964 -311
rect -1930 -345 -1914 -311
rect -1862 -345 -1846 -311
rect -1812 -345 -1796 -311
rect -1744 -345 -1728 -311
rect -1694 -345 -1678 -311
rect -1626 -345 -1610 -311
rect -1576 -345 -1560 -311
rect -1508 -345 -1492 -311
rect -1458 -345 -1442 -311
rect -1390 -345 -1374 -311
rect -1340 -345 -1324 -311
rect -1272 -345 -1256 -311
rect -1222 -345 -1206 -311
rect -1154 -345 -1138 -311
rect -1104 -345 -1088 -311
rect -1036 -345 -1020 -311
rect -986 -345 -970 -311
rect -918 -345 -902 -311
rect -868 -345 -852 -311
rect -800 -345 -784 -311
rect -750 -345 -734 -311
rect -682 -345 -666 -311
rect -632 -345 -616 -311
rect -564 -345 -548 -311
rect -514 -345 -498 -311
rect -446 -345 -430 -311
rect -396 -345 -380 -311
rect -328 -345 -312 -311
rect -278 -345 -262 -311
rect -210 -345 -194 -311
rect -160 -345 -144 -311
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect 26 -345 42 -311
rect 76 -345 92 -311
rect 144 -345 160 -311
rect 194 -345 210 -311
rect 262 -345 278 -311
rect 312 -345 328 -311
rect 380 -345 396 -311
rect 430 -345 446 -311
rect 498 -345 514 -311
rect 548 -345 564 -311
rect 616 -345 632 -311
rect 666 -345 682 -311
rect 734 -345 750 -311
rect 784 -345 800 -311
rect 852 -345 868 -311
rect 902 -345 918 -311
rect 970 -345 986 -311
rect 1020 -345 1036 -311
rect 1088 -345 1104 -311
rect 1138 -345 1154 -311
rect 1206 -345 1222 -311
rect 1256 -345 1272 -311
rect 1324 -345 1340 -311
rect 1374 -345 1390 -311
rect 1442 -345 1458 -311
rect 1492 -345 1508 -311
rect 1560 -345 1576 -311
rect 1610 -345 1626 -311
rect 1678 -345 1694 -311
rect 1728 -345 1744 -311
rect 1796 -345 1812 -311
rect 1846 -345 1862 -311
rect 1914 -345 1930 -311
rect 1964 -345 1980 -311
rect 2032 -345 2048 -311
rect 2082 -345 2098 -311
rect 2150 -345 2166 -311
rect 2200 -345 2216 -311
rect 2268 -345 2284 -311
rect 2318 -345 2334 -311
rect 2386 -345 2402 -311
rect 2436 -345 2452 -311
rect 2504 -345 2520 -311
rect 2554 -345 2570 -311
rect 2622 -345 2638 -311
rect 2672 -345 2688 -311
rect 2740 -345 2756 -311
rect 2790 -345 2806 -311
rect 2858 -345 2874 -311
rect 2908 -345 2924 -311
rect 2976 -345 2992 -311
rect 3026 -345 3042 -311
rect 3094 -345 3110 -311
rect 3144 -345 3160 -311
rect 3212 -345 3228 -311
rect 3262 -345 3278 -311
rect 3330 -345 3346 -311
rect 3380 -345 3396 -311
rect 3448 -345 3464 -311
rect 3498 -345 3514 -311
rect 3566 -345 3582 -311
rect 3616 -345 3632 -311
rect 3684 -345 3700 -311
rect 3734 -345 3750 -311
rect 3802 -345 3818 -311
rect 3852 -345 3868 -311
rect 3920 -345 3936 -311
rect 3970 -345 3986 -311
rect 4038 -345 4054 -311
rect 4088 -345 4104 -311
rect 4156 -345 4172 -311
rect 4206 -345 4222 -311
rect 4274 -345 4290 -311
rect 4324 -345 4340 -311
rect 4392 -345 4408 -311
rect 4442 -345 4458 -311
rect 4510 -345 4526 -311
rect 4560 -345 4576 -311
rect 4628 -345 4644 -311
rect 4678 -345 4694 -311
rect 4746 -345 4762 -311
rect 4796 -345 4812 -311
rect 4864 -345 4880 -311
rect 4914 -345 4930 -311
rect 4982 -345 4998 -311
rect 5032 -345 5048 -311
rect 5100 -345 5116 -311
rect 5150 -345 5166 -311
rect 5218 -345 5234 -311
rect 5268 -345 5284 -311
rect 5336 -345 5352 -311
rect 5386 -345 5402 -311
rect 5454 -345 5470 -311
rect 5504 -345 5520 -311
rect 5572 -345 5588 -311
rect 5622 -345 5638 -311
rect 5690 -345 5706 -311
rect 5740 -345 5756 -311
rect 5808 -345 5824 -311
rect 5858 -345 5874 -311
rect 5926 -345 5942 -311
rect 5976 -345 5992 -311
rect 6044 -345 6060 -311
rect 6094 -345 6110 -311
rect 6162 -345 6178 -311
rect 6212 -345 6228 -311
rect 6280 -345 6296 -311
rect 6330 -345 6346 -311
rect 6398 -345 6414 -311
rect 6448 -345 6464 -311
rect 6516 -345 6532 -311
rect 6566 -345 6582 -311
rect 6634 -345 6650 -311
rect 6684 -345 6700 -311
rect 6752 -345 6768 -311
rect 6802 -345 6818 -311
rect 6870 -345 6886 -311
rect 6920 -345 6936 -311
rect 6988 -345 7004 -311
rect 7038 -345 7054 -311
rect 7106 -345 7122 -311
rect 7156 -345 7172 -311
rect 7224 -345 7240 -311
rect 7274 -345 7290 -311
rect 7342 -345 7358 -311
rect 7392 -345 7408 -311
rect 7460 -345 7476 -311
rect 7510 -345 7526 -311
rect 7578 -345 7594 -311
rect 7628 -345 7644 -311
rect 7696 -345 7712 -311
rect 7746 -345 7762 -311
rect 7814 -345 7830 -311
rect 7864 -345 7880 -311
rect 7932 -345 7948 -311
rect 7982 -345 7998 -311
rect 8050 -345 8066 -311
rect 8100 -345 8116 -311
rect 8168 -345 8184 -311
rect 8218 -345 8234 -311
rect 8286 -345 8302 -311
rect 8336 -345 8352 -311
rect 8404 -345 8420 -311
rect 8454 -345 8470 -311
rect 8522 -345 8538 -311
rect 8572 -345 8588 -311
rect 8640 -345 8656 -311
rect 8690 -345 8706 -311
rect 8758 -345 8774 -311
rect 8808 -345 8824 -311
rect 8876 -345 8892 -311
rect 8926 -345 8942 -311
rect 8994 -345 9010 -311
rect 9044 -345 9060 -311
rect 9112 -345 9128 -311
rect 9162 -345 9178 -311
rect 9230 -345 9246 -311
rect 9280 -345 9296 -311
rect 9348 -345 9364 -311
rect 9398 -345 9414 -311
rect 9466 -345 9482 -311
rect 9516 -345 9532 -311
rect 9584 -345 9600 -311
rect 9634 -345 9650 -311
rect 9702 -345 9718 -311
rect 9752 -345 9768 -311
rect 9820 -345 9836 -311
rect 9870 -345 9886 -311
rect 9938 -345 9954 -311
rect 9988 -345 10004 -311
rect 10056 -345 10072 -311
rect 10106 -345 10122 -311
rect 10174 -345 10190 -311
rect 10224 -345 10240 -311
rect 10292 -345 10308 -311
rect 10342 -345 10358 -311
rect 10410 -345 10426 -311
rect 10460 -345 10476 -311
rect 10528 -345 10544 -311
rect 10578 -345 10594 -311
rect 10646 -345 10662 -311
rect 10696 -345 10712 -311
rect 10764 -345 10780 -311
rect 10814 -345 10830 -311
rect 10882 -345 10898 -311
rect 10932 -345 10948 -311
rect 11000 -345 11016 -311
rect 11050 -345 11066 -311
rect 11118 -345 11134 -311
rect 11168 -345 11184 -311
rect 11236 -345 11252 -311
rect 11286 -345 11302 -311
rect 11354 -345 11370 -311
rect 11404 -345 11420 -311
rect 11472 -345 11488 -311
rect 11522 -345 11538 -311
rect 11590 -345 11606 -311
rect 11640 -345 11656 -311
rect 11708 -345 11724 -311
rect 11758 -345 11774 -311
rect 11826 -345 11842 -311
rect 11876 -345 11892 -311
rect 11944 -345 11960 -311
rect 11994 -345 12010 -311
rect 12062 -345 12078 -311
rect 12112 -345 12128 -311
rect 12180 -345 12196 -311
rect 12230 -345 12246 -311
rect 12298 -345 12314 -311
rect 12348 -345 12364 -311
rect 12416 -345 12432 -311
rect 12466 -345 12482 -311
rect 12534 -345 12550 -311
rect 12584 -345 12600 -311
rect 12652 -345 12668 -311
rect 12702 -345 12718 -311
rect 12770 -345 12786 -311
rect 12820 -345 12836 -311
rect 12888 -345 12904 -311
rect 12938 -345 12954 -311
rect 13006 -345 13022 -311
rect 13056 -345 13072 -311
rect 13124 -345 13140 -311
rect 13174 -345 13190 -311
rect 13242 -345 13258 -311
rect 13292 -345 13308 -311
rect 13360 -345 13376 -311
rect 13410 -345 13426 -311
rect 13478 -345 13494 -311
rect 13528 -345 13544 -311
rect 13596 -345 13612 -311
rect 13646 -345 13662 -311
rect 13714 -345 13730 -311
rect 13764 -345 13780 -311
rect 13832 -345 13848 -311
rect 13882 -345 13898 -311
rect 13950 -345 13966 -311
rect 14000 -345 14016 -311
rect 14068 -345 14084 -311
rect 14118 -345 14134 -311
rect 14186 -345 14202 -311
rect 14236 -345 14252 -311
rect 14304 -345 14320 -311
rect 14354 -345 14370 -311
rect 14422 -345 14438 -311
rect 14472 -345 14488 -311
rect 14540 -345 14556 -311
rect 14590 -345 14606 -311
rect 14658 -345 14674 -311
rect 14708 -345 14724 -311
rect -14881 -414 -14847 -351
rect 14847 -414 14881 -351
rect -14881 -448 -14785 -414
rect 14785 -448 14881 -414
<< viali >>
rect -14767 -252 -14733 324
rect -14649 -252 -14615 324
rect -14531 -252 -14497 324
rect -14413 -252 -14379 324
rect -14295 -252 -14261 324
rect -14177 -252 -14143 324
rect -14059 -252 -14025 324
rect -13941 -252 -13907 324
rect -13823 -252 -13789 324
rect -13705 -252 -13671 324
rect -13587 -252 -13553 324
rect -13469 -252 -13435 324
rect -13351 -252 -13317 324
rect -13233 -252 -13199 324
rect -13115 -252 -13081 324
rect -12997 -252 -12963 324
rect -12879 -252 -12845 324
rect -12761 -252 -12727 324
rect -12643 -252 -12609 324
rect -12525 -252 -12491 324
rect -12407 -252 -12373 324
rect -12289 -252 -12255 324
rect -12171 -252 -12137 324
rect -12053 -252 -12019 324
rect -11935 -252 -11901 324
rect -11817 -252 -11783 324
rect -11699 -252 -11665 324
rect -11581 -252 -11547 324
rect -11463 -252 -11429 324
rect -11345 -252 -11311 324
rect -11227 -252 -11193 324
rect -11109 -252 -11075 324
rect -10991 -252 -10957 324
rect -10873 -252 -10839 324
rect -10755 -252 -10721 324
rect -10637 -252 -10603 324
rect -10519 -252 -10485 324
rect -10401 -252 -10367 324
rect -10283 -252 -10249 324
rect -10165 -252 -10131 324
rect -10047 -252 -10013 324
rect -9929 -252 -9895 324
rect -9811 -252 -9777 324
rect -9693 -252 -9659 324
rect -9575 -252 -9541 324
rect -9457 -252 -9423 324
rect -9339 -252 -9305 324
rect -9221 -252 -9187 324
rect -9103 -252 -9069 324
rect -8985 -252 -8951 324
rect -8867 -252 -8833 324
rect -8749 -252 -8715 324
rect -8631 -252 -8597 324
rect -8513 -252 -8479 324
rect -8395 -252 -8361 324
rect -8277 -252 -8243 324
rect -8159 -252 -8125 324
rect -8041 -252 -8007 324
rect -7923 -252 -7889 324
rect -7805 -252 -7771 324
rect -7687 -252 -7653 324
rect -7569 -252 -7535 324
rect -7451 -252 -7417 324
rect -7333 -252 -7299 324
rect -7215 -252 -7181 324
rect -7097 -252 -7063 324
rect -6979 -252 -6945 324
rect -6861 -252 -6827 324
rect -6743 -252 -6709 324
rect -6625 -252 -6591 324
rect -6507 -252 -6473 324
rect -6389 -252 -6355 324
rect -6271 -252 -6237 324
rect -6153 -252 -6119 324
rect -6035 -252 -6001 324
rect -5917 -252 -5883 324
rect -5799 -252 -5765 324
rect -5681 -252 -5647 324
rect -5563 -252 -5529 324
rect -5445 -252 -5411 324
rect -5327 -252 -5293 324
rect -5209 -252 -5175 324
rect -5091 -252 -5057 324
rect -4973 -252 -4939 324
rect -4855 -252 -4821 324
rect -4737 -252 -4703 324
rect -4619 -252 -4585 324
rect -4501 -252 -4467 324
rect -4383 -252 -4349 324
rect -4265 -252 -4231 324
rect -4147 -252 -4113 324
rect -4029 -252 -3995 324
rect -3911 -252 -3877 324
rect -3793 -252 -3759 324
rect -3675 -252 -3641 324
rect -3557 -252 -3523 324
rect -3439 -252 -3405 324
rect -3321 -252 -3287 324
rect -3203 -252 -3169 324
rect -3085 -252 -3051 324
rect -2967 -252 -2933 324
rect -2849 -252 -2815 324
rect -2731 -252 -2697 324
rect -2613 -252 -2579 324
rect -2495 -252 -2461 324
rect -2377 -252 -2343 324
rect -2259 -252 -2225 324
rect -2141 -252 -2107 324
rect -2023 -252 -1989 324
rect -1905 -252 -1871 324
rect -1787 -252 -1753 324
rect -1669 -252 -1635 324
rect -1551 -252 -1517 324
rect -1433 -252 -1399 324
rect -1315 -252 -1281 324
rect -1197 -252 -1163 324
rect -1079 -252 -1045 324
rect -961 -252 -927 324
rect -843 -252 -809 324
rect -725 -252 -691 324
rect -607 -252 -573 324
rect -489 -252 -455 324
rect -371 -252 -337 324
rect -253 -252 -219 324
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
rect 219 -252 253 324
rect 337 -252 371 324
rect 455 -252 489 324
rect 573 -252 607 324
rect 691 -252 725 324
rect 809 -252 843 324
rect 927 -252 961 324
rect 1045 -252 1079 324
rect 1163 -252 1197 324
rect 1281 -252 1315 324
rect 1399 -252 1433 324
rect 1517 -252 1551 324
rect 1635 -252 1669 324
rect 1753 -252 1787 324
rect 1871 -252 1905 324
rect 1989 -252 2023 324
rect 2107 -252 2141 324
rect 2225 -252 2259 324
rect 2343 -252 2377 324
rect 2461 -252 2495 324
rect 2579 -252 2613 324
rect 2697 -252 2731 324
rect 2815 -252 2849 324
rect 2933 -252 2967 324
rect 3051 -252 3085 324
rect 3169 -252 3203 324
rect 3287 -252 3321 324
rect 3405 -252 3439 324
rect 3523 -252 3557 324
rect 3641 -252 3675 324
rect 3759 -252 3793 324
rect 3877 -252 3911 324
rect 3995 -252 4029 324
rect 4113 -252 4147 324
rect 4231 -252 4265 324
rect 4349 -252 4383 324
rect 4467 -252 4501 324
rect 4585 -252 4619 324
rect 4703 -252 4737 324
rect 4821 -252 4855 324
rect 4939 -252 4973 324
rect 5057 -252 5091 324
rect 5175 -252 5209 324
rect 5293 -252 5327 324
rect 5411 -252 5445 324
rect 5529 -252 5563 324
rect 5647 -252 5681 324
rect 5765 -252 5799 324
rect 5883 -252 5917 324
rect 6001 -252 6035 324
rect 6119 -252 6153 324
rect 6237 -252 6271 324
rect 6355 -252 6389 324
rect 6473 -252 6507 324
rect 6591 -252 6625 324
rect 6709 -252 6743 324
rect 6827 -252 6861 324
rect 6945 -252 6979 324
rect 7063 -252 7097 324
rect 7181 -252 7215 324
rect 7299 -252 7333 324
rect 7417 -252 7451 324
rect 7535 -252 7569 324
rect 7653 -252 7687 324
rect 7771 -252 7805 324
rect 7889 -252 7923 324
rect 8007 -252 8041 324
rect 8125 -252 8159 324
rect 8243 -252 8277 324
rect 8361 -252 8395 324
rect 8479 -252 8513 324
rect 8597 -252 8631 324
rect 8715 -252 8749 324
rect 8833 -252 8867 324
rect 8951 -252 8985 324
rect 9069 -252 9103 324
rect 9187 -252 9221 324
rect 9305 -252 9339 324
rect 9423 -252 9457 324
rect 9541 -252 9575 324
rect 9659 -252 9693 324
rect 9777 -252 9811 324
rect 9895 -252 9929 324
rect 10013 -252 10047 324
rect 10131 -252 10165 324
rect 10249 -252 10283 324
rect 10367 -252 10401 324
rect 10485 -252 10519 324
rect 10603 -252 10637 324
rect 10721 -252 10755 324
rect 10839 -252 10873 324
rect 10957 -252 10991 324
rect 11075 -252 11109 324
rect 11193 -252 11227 324
rect 11311 -252 11345 324
rect 11429 -252 11463 324
rect 11547 -252 11581 324
rect 11665 -252 11699 324
rect 11783 -252 11817 324
rect 11901 -252 11935 324
rect 12019 -252 12053 324
rect 12137 -252 12171 324
rect 12255 -252 12289 324
rect 12373 -252 12407 324
rect 12491 -252 12525 324
rect 12609 -252 12643 324
rect 12727 -252 12761 324
rect 12845 -252 12879 324
rect 12963 -252 12997 324
rect 13081 -252 13115 324
rect 13199 -252 13233 324
rect 13317 -252 13351 324
rect 13435 -252 13469 324
rect 13553 -252 13587 324
rect 13671 -252 13705 324
rect 13789 -252 13823 324
rect 13907 -252 13941 324
rect 14025 -252 14059 324
rect 14143 -252 14177 324
rect 14261 -252 14295 324
rect 14379 -252 14413 324
rect 14497 -252 14531 324
rect 14615 -252 14649 324
rect 14733 -252 14767 324
rect -14708 -345 -14674 -311
rect -14590 -345 -14556 -311
rect -14472 -345 -14438 -311
rect -14354 -345 -14320 -311
rect -14236 -345 -14202 -311
rect -14118 -345 -14084 -311
rect -14000 -345 -13966 -311
rect -13882 -345 -13848 -311
rect -13764 -345 -13730 -311
rect -13646 -345 -13612 -311
rect -13528 -345 -13494 -311
rect -13410 -345 -13376 -311
rect -13292 -345 -13258 -311
rect -13174 -345 -13140 -311
rect -13056 -345 -13022 -311
rect -12938 -345 -12904 -311
rect -12820 -345 -12786 -311
rect -12702 -345 -12668 -311
rect -12584 -345 -12550 -311
rect -12466 -345 -12432 -311
rect -12348 -345 -12314 -311
rect -12230 -345 -12196 -311
rect -12112 -345 -12078 -311
rect -11994 -345 -11960 -311
rect -11876 -345 -11842 -311
rect -11758 -345 -11724 -311
rect -11640 -345 -11606 -311
rect -11522 -345 -11488 -311
rect -11404 -345 -11370 -311
rect -11286 -345 -11252 -311
rect -11168 -345 -11134 -311
rect -11050 -345 -11016 -311
rect -10932 -345 -10898 -311
rect -10814 -345 -10780 -311
rect -10696 -345 -10662 -311
rect -10578 -345 -10544 -311
rect -10460 -345 -10426 -311
rect -10342 -345 -10308 -311
rect -10224 -345 -10190 -311
rect -10106 -345 -10072 -311
rect -9988 -345 -9954 -311
rect -9870 -345 -9836 -311
rect -9752 -345 -9718 -311
rect -9634 -345 -9600 -311
rect -9516 -345 -9482 -311
rect -9398 -345 -9364 -311
rect -9280 -345 -9246 -311
rect -9162 -345 -9128 -311
rect -9044 -345 -9010 -311
rect -8926 -345 -8892 -311
rect -8808 -345 -8774 -311
rect -8690 -345 -8656 -311
rect -8572 -345 -8538 -311
rect -8454 -345 -8420 -311
rect -8336 -345 -8302 -311
rect -8218 -345 -8184 -311
rect -8100 -345 -8066 -311
rect -7982 -345 -7948 -311
rect -7864 -345 -7830 -311
rect -7746 -345 -7712 -311
rect -7628 -345 -7594 -311
rect -7510 -345 -7476 -311
rect -7392 -345 -7358 -311
rect -7274 -345 -7240 -311
rect -7156 -345 -7122 -311
rect -7038 -345 -7004 -311
rect -6920 -345 -6886 -311
rect -6802 -345 -6768 -311
rect -6684 -345 -6650 -311
rect -6566 -345 -6532 -311
rect -6448 -345 -6414 -311
rect -6330 -345 -6296 -311
rect -6212 -345 -6178 -311
rect -6094 -345 -6060 -311
rect -5976 -345 -5942 -311
rect -5858 -345 -5824 -311
rect -5740 -345 -5706 -311
rect -5622 -345 -5588 -311
rect -5504 -345 -5470 -311
rect -5386 -345 -5352 -311
rect -5268 -345 -5234 -311
rect -5150 -345 -5116 -311
rect -5032 -345 -4998 -311
rect -4914 -345 -4880 -311
rect -4796 -345 -4762 -311
rect -4678 -345 -4644 -311
rect -4560 -345 -4526 -311
rect -4442 -345 -4408 -311
rect -4324 -345 -4290 -311
rect -4206 -345 -4172 -311
rect -4088 -345 -4054 -311
rect -3970 -345 -3936 -311
rect -3852 -345 -3818 -311
rect -3734 -345 -3700 -311
rect -3616 -345 -3582 -311
rect -3498 -345 -3464 -311
rect -3380 -345 -3346 -311
rect -3262 -345 -3228 -311
rect -3144 -345 -3110 -311
rect -3026 -345 -2992 -311
rect -2908 -345 -2874 -311
rect -2790 -345 -2756 -311
rect -2672 -345 -2638 -311
rect -2554 -345 -2520 -311
rect -2436 -345 -2402 -311
rect -2318 -345 -2284 -311
rect -2200 -345 -2166 -311
rect -2082 -345 -2048 -311
rect -1964 -345 -1930 -311
rect -1846 -345 -1812 -311
rect -1728 -345 -1694 -311
rect -1610 -345 -1576 -311
rect -1492 -345 -1458 -311
rect -1374 -345 -1340 -311
rect -1256 -345 -1222 -311
rect -1138 -345 -1104 -311
rect -1020 -345 -986 -311
rect -902 -345 -868 -311
rect -784 -345 -750 -311
rect -666 -345 -632 -311
rect -548 -345 -514 -311
rect -430 -345 -396 -311
rect -312 -345 -278 -311
rect -194 -345 -160 -311
rect -76 -345 -42 -311
rect 42 -345 76 -311
rect 160 -345 194 -311
rect 278 -345 312 -311
rect 396 -345 430 -311
rect 514 -345 548 -311
rect 632 -345 666 -311
rect 750 -345 784 -311
rect 868 -345 902 -311
rect 986 -345 1020 -311
rect 1104 -345 1138 -311
rect 1222 -345 1256 -311
rect 1340 -345 1374 -311
rect 1458 -345 1492 -311
rect 1576 -345 1610 -311
rect 1694 -345 1728 -311
rect 1812 -345 1846 -311
rect 1930 -345 1964 -311
rect 2048 -345 2082 -311
rect 2166 -345 2200 -311
rect 2284 -345 2318 -311
rect 2402 -345 2436 -311
rect 2520 -345 2554 -311
rect 2638 -345 2672 -311
rect 2756 -345 2790 -311
rect 2874 -345 2908 -311
rect 2992 -345 3026 -311
rect 3110 -345 3144 -311
rect 3228 -345 3262 -311
rect 3346 -345 3380 -311
rect 3464 -345 3498 -311
rect 3582 -345 3616 -311
rect 3700 -345 3734 -311
rect 3818 -345 3852 -311
rect 3936 -345 3970 -311
rect 4054 -345 4088 -311
rect 4172 -345 4206 -311
rect 4290 -345 4324 -311
rect 4408 -345 4442 -311
rect 4526 -345 4560 -311
rect 4644 -345 4678 -311
rect 4762 -345 4796 -311
rect 4880 -345 4914 -311
rect 4998 -345 5032 -311
rect 5116 -345 5150 -311
rect 5234 -345 5268 -311
rect 5352 -345 5386 -311
rect 5470 -345 5504 -311
rect 5588 -345 5622 -311
rect 5706 -345 5740 -311
rect 5824 -345 5858 -311
rect 5942 -345 5976 -311
rect 6060 -345 6094 -311
rect 6178 -345 6212 -311
rect 6296 -345 6330 -311
rect 6414 -345 6448 -311
rect 6532 -345 6566 -311
rect 6650 -345 6684 -311
rect 6768 -345 6802 -311
rect 6886 -345 6920 -311
rect 7004 -345 7038 -311
rect 7122 -345 7156 -311
rect 7240 -345 7274 -311
rect 7358 -345 7392 -311
rect 7476 -345 7510 -311
rect 7594 -345 7628 -311
rect 7712 -345 7746 -311
rect 7830 -345 7864 -311
rect 7948 -345 7982 -311
rect 8066 -345 8100 -311
rect 8184 -345 8218 -311
rect 8302 -345 8336 -311
rect 8420 -345 8454 -311
rect 8538 -345 8572 -311
rect 8656 -345 8690 -311
rect 8774 -345 8808 -311
rect 8892 -345 8926 -311
rect 9010 -345 9044 -311
rect 9128 -345 9162 -311
rect 9246 -345 9280 -311
rect 9364 -345 9398 -311
rect 9482 -345 9516 -311
rect 9600 -345 9634 -311
rect 9718 -345 9752 -311
rect 9836 -345 9870 -311
rect 9954 -345 9988 -311
rect 10072 -345 10106 -311
rect 10190 -345 10224 -311
rect 10308 -345 10342 -311
rect 10426 -345 10460 -311
rect 10544 -345 10578 -311
rect 10662 -345 10696 -311
rect 10780 -345 10814 -311
rect 10898 -345 10932 -311
rect 11016 -345 11050 -311
rect 11134 -345 11168 -311
rect 11252 -345 11286 -311
rect 11370 -345 11404 -311
rect 11488 -345 11522 -311
rect 11606 -345 11640 -311
rect 11724 -345 11758 -311
rect 11842 -345 11876 -311
rect 11960 -345 11994 -311
rect 12078 -345 12112 -311
rect 12196 -345 12230 -311
rect 12314 -345 12348 -311
rect 12432 -345 12466 -311
rect 12550 -345 12584 -311
rect 12668 -345 12702 -311
rect 12786 -345 12820 -311
rect 12904 -345 12938 -311
rect 13022 -345 13056 -311
rect 13140 -345 13174 -311
rect 13258 -345 13292 -311
rect 13376 -345 13410 -311
rect 13494 -345 13528 -311
rect 13612 -345 13646 -311
rect 13730 -345 13764 -311
rect 13848 -345 13882 -311
rect 13966 -345 14000 -311
rect 14084 -345 14118 -311
rect 14202 -345 14236 -311
rect 14320 -345 14354 -311
rect 14438 -345 14472 -311
rect 14556 -345 14590 -311
rect 14674 -345 14708 -311
<< metal1 >>
rect -14773 324 -14727 336
rect -14773 -252 -14767 324
rect -14733 -252 -14727 324
rect -14773 -264 -14727 -252
rect -14655 324 -14609 336
rect -14655 -252 -14649 324
rect -14615 -252 -14609 324
rect -14655 -264 -14609 -252
rect -14537 324 -14491 336
rect -14537 -252 -14531 324
rect -14497 -252 -14491 324
rect -14537 -264 -14491 -252
rect -14419 324 -14373 336
rect -14419 -252 -14413 324
rect -14379 -252 -14373 324
rect -14419 -264 -14373 -252
rect -14301 324 -14255 336
rect -14301 -252 -14295 324
rect -14261 -252 -14255 324
rect -14301 -264 -14255 -252
rect -14183 324 -14137 336
rect -14183 -252 -14177 324
rect -14143 -252 -14137 324
rect -14183 -264 -14137 -252
rect -14065 324 -14019 336
rect -14065 -252 -14059 324
rect -14025 -252 -14019 324
rect -14065 -264 -14019 -252
rect -13947 324 -13901 336
rect -13947 -252 -13941 324
rect -13907 -252 -13901 324
rect -13947 -264 -13901 -252
rect -13829 324 -13783 336
rect -13829 -252 -13823 324
rect -13789 -252 -13783 324
rect -13829 -264 -13783 -252
rect -13711 324 -13665 336
rect -13711 -252 -13705 324
rect -13671 -252 -13665 324
rect -13711 -264 -13665 -252
rect -13593 324 -13547 336
rect -13593 -252 -13587 324
rect -13553 -252 -13547 324
rect -13593 -264 -13547 -252
rect -13475 324 -13429 336
rect -13475 -252 -13469 324
rect -13435 -252 -13429 324
rect -13475 -264 -13429 -252
rect -13357 324 -13311 336
rect -13357 -252 -13351 324
rect -13317 -252 -13311 324
rect -13357 -264 -13311 -252
rect -13239 324 -13193 336
rect -13239 -252 -13233 324
rect -13199 -252 -13193 324
rect -13239 -264 -13193 -252
rect -13121 324 -13075 336
rect -13121 -252 -13115 324
rect -13081 -252 -13075 324
rect -13121 -264 -13075 -252
rect -13003 324 -12957 336
rect -13003 -252 -12997 324
rect -12963 -252 -12957 324
rect -13003 -264 -12957 -252
rect -12885 324 -12839 336
rect -12885 -252 -12879 324
rect -12845 -252 -12839 324
rect -12885 -264 -12839 -252
rect -12767 324 -12721 336
rect -12767 -252 -12761 324
rect -12727 -252 -12721 324
rect -12767 -264 -12721 -252
rect -12649 324 -12603 336
rect -12649 -252 -12643 324
rect -12609 -252 -12603 324
rect -12649 -264 -12603 -252
rect -12531 324 -12485 336
rect -12531 -252 -12525 324
rect -12491 -252 -12485 324
rect -12531 -264 -12485 -252
rect -12413 324 -12367 336
rect -12413 -252 -12407 324
rect -12373 -252 -12367 324
rect -12413 -264 -12367 -252
rect -12295 324 -12249 336
rect -12295 -252 -12289 324
rect -12255 -252 -12249 324
rect -12295 -264 -12249 -252
rect -12177 324 -12131 336
rect -12177 -252 -12171 324
rect -12137 -252 -12131 324
rect -12177 -264 -12131 -252
rect -12059 324 -12013 336
rect -12059 -252 -12053 324
rect -12019 -252 -12013 324
rect -12059 -264 -12013 -252
rect -11941 324 -11895 336
rect -11941 -252 -11935 324
rect -11901 -252 -11895 324
rect -11941 -264 -11895 -252
rect -11823 324 -11777 336
rect -11823 -252 -11817 324
rect -11783 -252 -11777 324
rect -11823 -264 -11777 -252
rect -11705 324 -11659 336
rect -11705 -252 -11699 324
rect -11665 -252 -11659 324
rect -11705 -264 -11659 -252
rect -11587 324 -11541 336
rect -11587 -252 -11581 324
rect -11547 -252 -11541 324
rect -11587 -264 -11541 -252
rect -11469 324 -11423 336
rect -11469 -252 -11463 324
rect -11429 -252 -11423 324
rect -11469 -264 -11423 -252
rect -11351 324 -11305 336
rect -11351 -252 -11345 324
rect -11311 -252 -11305 324
rect -11351 -264 -11305 -252
rect -11233 324 -11187 336
rect -11233 -252 -11227 324
rect -11193 -252 -11187 324
rect -11233 -264 -11187 -252
rect -11115 324 -11069 336
rect -11115 -252 -11109 324
rect -11075 -252 -11069 324
rect -11115 -264 -11069 -252
rect -10997 324 -10951 336
rect -10997 -252 -10991 324
rect -10957 -252 -10951 324
rect -10997 -264 -10951 -252
rect -10879 324 -10833 336
rect -10879 -252 -10873 324
rect -10839 -252 -10833 324
rect -10879 -264 -10833 -252
rect -10761 324 -10715 336
rect -10761 -252 -10755 324
rect -10721 -252 -10715 324
rect -10761 -264 -10715 -252
rect -10643 324 -10597 336
rect -10643 -252 -10637 324
rect -10603 -252 -10597 324
rect -10643 -264 -10597 -252
rect -10525 324 -10479 336
rect -10525 -252 -10519 324
rect -10485 -252 -10479 324
rect -10525 -264 -10479 -252
rect -10407 324 -10361 336
rect -10407 -252 -10401 324
rect -10367 -252 -10361 324
rect -10407 -264 -10361 -252
rect -10289 324 -10243 336
rect -10289 -252 -10283 324
rect -10249 -252 -10243 324
rect -10289 -264 -10243 -252
rect -10171 324 -10125 336
rect -10171 -252 -10165 324
rect -10131 -252 -10125 324
rect -10171 -264 -10125 -252
rect -10053 324 -10007 336
rect -10053 -252 -10047 324
rect -10013 -252 -10007 324
rect -10053 -264 -10007 -252
rect -9935 324 -9889 336
rect -9935 -252 -9929 324
rect -9895 -252 -9889 324
rect -9935 -264 -9889 -252
rect -9817 324 -9771 336
rect -9817 -252 -9811 324
rect -9777 -252 -9771 324
rect -9817 -264 -9771 -252
rect -9699 324 -9653 336
rect -9699 -252 -9693 324
rect -9659 -252 -9653 324
rect -9699 -264 -9653 -252
rect -9581 324 -9535 336
rect -9581 -252 -9575 324
rect -9541 -252 -9535 324
rect -9581 -264 -9535 -252
rect -9463 324 -9417 336
rect -9463 -252 -9457 324
rect -9423 -252 -9417 324
rect -9463 -264 -9417 -252
rect -9345 324 -9299 336
rect -9345 -252 -9339 324
rect -9305 -252 -9299 324
rect -9345 -264 -9299 -252
rect -9227 324 -9181 336
rect -9227 -252 -9221 324
rect -9187 -252 -9181 324
rect -9227 -264 -9181 -252
rect -9109 324 -9063 336
rect -9109 -252 -9103 324
rect -9069 -252 -9063 324
rect -9109 -264 -9063 -252
rect -8991 324 -8945 336
rect -8991 -252 -8985 324
rect -8951 -252 -8945 324
rect -8991 -264 -8945 -252
rect -8873 324 -8827 336
rect -8873 -252 -8867 324
rect -8833 -252 -8827 324
rect -8873 -264 -8827 -252
rect -8755 324 -8709 336
rect -8755 -252 -8749 324
rect -8715 -252 -8709 324
rect -8755 -264 -8709 -252
rect -8637 324 -8591 336
rect -8637 -252 -8631 324
rect -8597 -252 -8591 324
rect -8637 -264 -8591 -252
rect -8519 324 -8473 336
rect -8519 -252 -8513 324
rect -8479 -252 -8473 324
rect -8519 -264 -8473 -252
rect -8401 324 -8355 336
rect -8401 -252 -8395 324
rect -8361 -252 -8355 324
rect -8401 -264 -8355 -252
rect -8283 324 -8237 336
rect -8283 -252 -8277 324
rect -8243 -252 -8237 324
rect -8283 -264 -8237 -252
rect -8165 324 -8119 336
rect -8165 -252 -8159 324
rect -8125 -252 -8119 324
rect -8165 -264 -8119 -252
rect -8047 324 -8001 336
rect -8047 -252 -8041 324
rect -8007 -252 -8001 324
rect -8047 -264 -8001 -252
rect -7929 324 -7883 336
rect -7929 -252 -7923 324
rect -7889 -252 -7883 324
rect -7929 -264 -7883 -252
rect -7811 324 -7765 336
rect -7811 -252 -7805 324
rect -7771 -252 -7765 324
rect -7811 -264 -7765 -252
rect -7693 324 -7647 336
rect -7693 -252 -7687 324
rect -7653 -252 -7647 324
rect -7693 -264 -7647 -252
rect -7575 324 -7529 336
rect -7575 -252 -7569 324
rect -7535 -252 -7529 324
rect -7575 -264 -7529 -252
rect -7457 324 -7411 336
rect -7457 -252 -7451 324
rect -7417 -252 -7411 324
rect -7457 -264 -7411 -252
rect -7339 324 -7293 336
rect -7339 -252 -7333 324
rect -7299 -252 -7293 324
rect -7339 -264 -7293 -252
rect -7221 324 -7175 336
rect -7221 -252 -7215 324
rect -7181 -252 -7175 324
rect -7221 -264 -7175 -252
rect -7103 324 -7057 336
rect -7103 -252 -7097 324
rect -7063 -252 -7057 324
rect -7103 -264 -7057 -252
rect -6985 324 -6939 336
rect -6985 -252 -6979 324
rect -6945 -252 -6939 324
rect -6985 -264 -6939 -252
rect -6867 324 -6821 336
rect -6867 -252 -6861 324
rect -6827 -252 -6821 324
rect -6867 -264 -6821 -252
rect -6749 324 -6703 336
rect -6749 -252 -6743 324
rect -6709 -252 -6703 324
rect -6749 -264 -6703 -252
rect -6631 324 -6585 336
rect -6631 -252 -6625 324
rect -6591 -252 -6585 324
rect -6631 -264 -6585 -252
rect -6513 324 -6467 336
rect -6513 -252 -6507 324
rect -6473 -252 -6467 324
rect -6513 -264 -6467 -252
rect -6395 324 -6349 336
rect -6395 -252 -6389 324
rect -6355 -252 -6349 324
rect -6395 -264 -6349 -252
rect -6277 324 -6231 336
rect -6277 -252 -6271 324
rect -6237 -252 -6231 324
rect -6277 -264 -6231 -252
rect -6159 324 -6113 336
rect -6159 -252 -6153 324
rect -6119 -252 -6113 324
rect -6159 -264 -6113 -252
rect -6041 324 -5995 336
rect -6041 -252 -6035 324
rect -6001 -252 -5995 324
rect -6041 -264 -5995 -252
rect -5923 324 -5877 336
rect -5923 -252 -5917 324
rect -5883 -252 -5877 324
rect -5923 -264 -5877 -252
rect -5805 324 -5759 336
rect -5805 -252 -5799 324
rect -5765 -252 -5759 324
rect -5805 -264 -5759 -252
rect -5687 324 -5641 336
rect -5687 -252 -5681 324
rect -5647 -252 -5641 324
rect -5687 -264 -5641 -252
rect -5569 324 -5523 336
rect -5569 -252 -5563 324
rect -5529 -252 -5523 324
rect -5569 -264 -5523 -252
rect -5451 324 -5405 336
rect -5451 -252 -5445 324
rect -5411 -252 -5405 324
rect -5451 -264 -5405 -252
rect -5333 324 -5287 336
rect -5333 -252 -5327 324
rect -5293 -252 -5287 324
rect -5333 -264 -5287 -252
rect -5215 324 -5169 336
rect -5215 -252 -5209 324
rect -5175 -252 -5169 324
rect -5215 -264 -5169 -252
rect -5097 324 -5051 336
rect -5097 -252 -5091 324
rect -5057 -252 -5051 324
rect -5097 -264 -5051 -252
rect -4979 324 -4933 336
rect -4979 -252 -4973 324
rect -4939 -252 -4933 324
rect -4979 -264 -4933 -252
rect -4861 324 -4815 336
rect -4861 -252 -4855 324
rect -4821 -252 -4815 324
rect -4861 -264 -4815 -252
rect -4743 324 -4697 336
rect -4743 -252 -4737 324
rect -4703 -252 -4697 324
rect -4743 -264 -4697 -252
rect -4625 324 -4579 336
rect -4625 -252 -4619 324
rect -4585 -252 -4579 324
rect -4625 -264 -4579 -252
rect -4507 324 -4461 336
rect -4507 -252 -4501 324
rect -4467 -252 -4461 324
rect -4507 -264 -4461 -252
rect -4389 324 -4343 336
rect -4389 -252 -4383 324
rect -4349 -252 -4343 324
rect -4389 -264 -4343 -252
rect -4271 324 -4225 336
rect -4271 -252 -4265 324
rect -4231 -252 -4225 324
rect -4271 -264 -4225 -252
rect -4153 324 -4107 336
rect -4153 -252 -4147 324
rect -4113 -252 -4107 324
rect -4153 -264 -4107 -252
rect -4035 324 -3989 336
rect -4035 -252 -4029 324
rect -3995 -252 -3989 324
rect -4035 -264 -3989 -252
rect -3917 324 -3871 336
rect -3917 -252 -3911 324
rect -3877 -252 -3871 324
rect -3917 -264 -3871 -252
rect -3799 324 -3753 336
rect -3799 -252 -3793 324
rect -3759 -252 -3753 324
rect -3799 -264 -3753 -252
rect -3681 324 -3635 336
rect -3681 -252 -3675 324
rect -3641 -252 -3635 324
rect -3681 -264 -3635 -252
rect -3563 324 -3517 336
rect -3563 -252 -3557 324
rect -3523 -252 -3517 324
rect -3563 -264 -3517 -252
rect -3445 324 -3399 336
rect -3445 -252 -3439 324
rect -3405 -252 -3399 324
rect -3445 -264 -3399 -252
rect -3327 324 -3281 336
rect -3327 -252 -3321 324
rect -3287 -252 -3281 324
rect -3327 -264 -3281 -252
rect -3209 324 -3163 336
rect -3209 -252 -3203 324
rect -3169 -252 -3163 324
rect -3209 -264 -3163 -252
rect -3091 324 -3045 336
rect -3091 -252 -3085 324
rect -3051 -252 -3045 324
rect -3091 -264 -3045 -252
rect -2973 324 -2927 336
rect -2973 -252 -2967 324
rect -2933 -252 -2927 324
rect -2973 -264 -2927 -252
rect -2855 324 -2809 336
rect -2855 -252 -2849 324
rect -2815 -252 -2809 324
rect -2855 -264 -2809 -252
rect -2737 324 -2691 336
rect -2737 -252 -2731 324
rect -2697 -252 -2691 324
rect -2737 -264 -2691 -252
rect -2619 324 -2573 336
rect -2619 -252 -2613 324
rect -2579 -252 -2573 324
rect -2619 -264 -2573 -252
rect -2501 324 -2455 336
rect -2501 -252 -2495 324
rect -2461 -252 -2455 324
rect -2501 -264 -2455 -252
rect -2383 324 -2337 336
rect -2383 -252 -2377 324
rect -2343 -252 -2337 324
rect -2383 -264 -2337 -252
rect -2265 324 -2219 336
rect -2265 -252 -2259 324
rect -2225 -252 -2219 324
rect -2265 -264 -2219 -252
rect -2147 324 -2101 336
rect -2147 -252 -2141 324
rect -2107 -252 -2101 324
rect -2147 -264 -2101 -252
rect -2029 324 -1983 336
rect -2029 -252 -2023 324
rect -1989 -252 -1983 324
rect -2029 -264 -1983 -252
rect -1911 324 -1865 336
rect -1911 -252 -1905 324
rect -1871 -252 -1865 324
rect -1911 -264 -1865 -252
rect -1793 324 -1747 336
rect -1793 -252 -1787 324
rect -1753 -252 -1747 324
rect -1793 -264 -1747 -252
rect -1675 324 -1629 336
rect -1675 -252 -1669 324
rect -1635 -252 -1629 324
rect -1675 -264 -1629 -252
rect -1557 324 -1511 336
rect -1557 -252 -1551 324
rect -1517 -252 -1511 324
rect -1557 -264 -1511 -252
rect -1439 324 -1393 336
rect -1439 -252 -1433 324
rect -1399 -252 -1393 324
rect -1439 -264 -1393 -252
rect -1321 324 -1275 336
rect -1321 -252 -1315 324
rect -1281 -252 -1275 324
rect -1321 -264 -1275 -252
rect -1203 324 -1157 336
rect -1203 -252 -1197 324
rect -1163 -252 -1157 324
rect -1203 -264 -1157 -252
rect -1085 324 -1039 336
rect -1085 -252 -1079 324
rect -1045 -252 -1039 324
rect -1085 -264 -1039 -252
rect -967 324 -921 336
rect -967 -252 -961 324
rect -927 -252 -921 324
rect -967 -264 -921 -252
rect -849 324 -803 336
rect -849 -252 -843 324
rect -809 -252 -803 324
rect -849 -264 -803 -252
rect -731 324 -685 336
rect -731 -252 -725 324
rect -691 -252 -685 324
rect -731 -264 -685 -252
rect -613 324 -567 336
rect -613 -252 -607 324
rect -573 -252 -567 324
rect -613 -264 -567 -252
rect -495 324 -449 336
rect -495 -252 -489 324
rect -455 -252 -449 324
rect -495 -264 -449 -252
rect -377 324 -331 336
rect -377 -252 -371 324
rect -337 -252 -331 324
rect -377 -264 -331 -252
rect -259 324 -213 336
rect -259 -252 -253 324
rect -219 -252 -213 324
rect -259 -264 -213 -252
rect -141 324 -95 336
rect -141 -252 -135 324
rect -101 -252 -95 324
rect -141 -264 -95 -252
rect -23 324 23 336
rect -23 -252 -17 324
rect 17 -252 23 324
rect -23 -264 23 -252
rect 95 324 141 336
rect 95 -252 101 324
rect 135 -252 141 324
rect 95 -264 141 -252
rect 213 324 259 336
rect 213 -252 219 324
rect 253 -252 259 324
rect 213 -264 259 -252
rect 331 324 377 336
rect 331 -252 337 324
rect 371 -252 377 324
rect 331 -264 377 -252
rect 449 324 495 336
rect 449 -252 455 324
rect 489 -252 495 324
rect 449 -264 495 -252
rect 567 324 613 336
rect 567 -252 573 324
rect 607 -252 613 324
rect 567 -264 613 -252
rect 685 324 731 336
rect 685 -252 691 324
rect 725 -252 731 324
rect 685 -264 731 -252
rect 803 324 849 336
rect 803 -252 809 324
rect 843 -252 849 324
rect 803 -264 849 -252
rect 921 324 967 336
rect 921 -252 927 324
rect 961 -252 967 324
rect 921 -264 967 -252
rect 1039 324 1085 336
rect 1039 -252 1045 324
rect 1079 -252 1085 324
rect 1039 -264 1085 -252
rect 1157 324 1203 336
rect 1157 -252 1163 324
rect 1197 -252 1203 324
rect 1157 -264 1203 -252
rect 1275 324 1321 336
rect 1275 -252 1281 324
rect 1315 -252 1321 324
rect 1275 -264 1321 -252
rect 1393 324 1439 336
rect 1393 -252 1399 324
rect 1433 -252 1439 324
rect 1393 -264 1439 -252
rect 1511 324 1557 336
rect 1511 -252 1517 324
rect 1551 -252 1557 324
rect 1511 -264 1557 -252
rect 1629 324 1675 336
rect 1629 -252 1635 324
rect 1669 -252 1675 324
rect 1629 -264 1675 -252
rect 1747 324 1793 336
rect 1747 -252 1753 324
rect 1787 -252 1793 324
rect 1747 -264 1793 -252
rect 1865 324 1911 336
rect 1865 -252 1871 324
rect 1905 -252 1911 324
rect 1865 -264 1911 -252
rect 1983 324 2029 336
rect 1983 -252 1989 324
rect 2023 -252 2029 324
rect 1983 -264 2029 -252
rect 2101 324 2147 336
rect 2101 -252 2107 324
rect 2141 -252 2147 324
rect 2101 -264 2147 -252
rect 2219 324 2265 336
rect 2219 -252 2225 324
rect 2259 -252 2265 324
rect 2219 -264 2265 -252
rect 2337 324 2383 336
rect 2337 -252 2343 324
rect 2377 -252 2383 324
rect 2337 -264 2383 -252
rect 2455 324 2501 336
rect 2455 -252 2461 324
rect 2495 -252 2501 324
rect 2455 -264 2501 -252
rect 2573 324 2619 336
rect 2573 -252 2579 324
rect 2613 -252 2619 324
rect 2573 -264 2619 -252
rect 2691 324 2737 336
rect 2691 -252 2697 324
rect 2731 -252 2737 324
rect 2691 -264 2737 -252
rect 2809 324 2855 336
rect 2809 -252 2815 324
rect 2849 -252 2855 324
rect 2809 -264 2855 -252
rect 2927 324 2973 336
rect 2927 -252 2933 324
rect 2967 -252 2973 324
rect 2927 -264 2973 -252
rect 3045 324 3091 336
rect 3045 -252 3051 324
rect 3085 -252 3091 324
rect 3045 -264 3091 -252
rect 3163 324 3209 336
rect 3163 -252 3169 324
rect 3203 -252 3209 324
rect 3163 -264 3209 -252
rect 3281 324 3327 336
rect 3281 -252 3287 324
rect 3321 -252 3327 324
rect 3281 -264 3327 -252
rect 3399 324 3445 336
rect 3399 -252 3405 324
rect 3439 -252 3445 324
rect 3399 -264 3445 -252
rect 3517 324 3563 336
rect 3517 -252 3523 324
rect 3557 -252 3563 324
rect 3517 -264 3563 -252
rect 3635 324 3681 336
rect 3635 -252 3641 324
rect 3675 -252 3681 324
rect 3635 -264 3681 -252
rect 3753 324 3799 336
rect 3753 -252 3759 324
rect 3793 -252 3799 324
rect 3753 -264 3799 -252
rect 3871 324 3917 336
rect 3871 -252 3877 324
rect 3911 -252 3917 324
rect 3871 -264 3917 -252
rect 3989 324 4035 336
rect 3989 -252 3995 324
rect 4029 -252 4035 324
rect 3989 -264 4035 -252
rect 4107 324 4153 336
rect 4107 -252 4113 324
rect 4147 -252 4153 324
rect 4107 -264 4153 -252
rect 4225 324 4271 336
rect 4225 -252 4231 324
rect 4265 -252 4271 324
rect 4225 -264 4271 -252
rect 4343 324 4389 336
rect 4343 -252 4349 324
rect 4383 -252 4389 324
rect 4343 -264 4389 -252
rect 4461 324 4507 336
rect 4461 -252 4467 324
rect 4501 -252 4507 324
rect 4461 -264 4507 -252
rect 4579 324 4625 336
rect 4579 -252 4585 324
rect 4619 -252 4625 324
rect 4579 -264 4625 -252
rect 4697 324 4743 336
rect 4697 -252 4703 324
rect 4737 -252 4743 324
rect 4697 -264 4743 -252
rect 4815 324 4861 336
rect 4815 -252 4821 324
rect 4855 -252 4861 324
rect 4815 -264 4861 -252
rect 4933 324 4979 336
rect 4933 -252 4939 324
rect 4973 -252 4979 324
rect 4933 -264 4979 -252
rect 5051 324 5097 336
rect 5051 -252 5057 324
rect 5091 -252 5097 324
rect 5051 -264 5097 -252
rect 5169 324 5215 336
rect 5169 -252 5175 324
rect 5209 -252 5215 324
rect 5169 -264 5215 -252
rect 5287 324 5333 336
rect 5287 -252 5293 324
rect 5327 -252 5333 324
rect 5287 -264 5333 -252
rect 5405 324 5451 336
rect 5405 -252 5411 324
rect 5445 -252 5451 324
rect 5405 -264 5451 -252
rect 5523 324 5569 336
rect 5523 -252 5529 324
rect 5563 -252 5569 324
rect 5523 -264 5569 -252
rect 5641 324 5687 336
rect 5641 -252 5647 324
rect 5681 -252 5687 324
rect 5641 -264 5687 -252
rect 5759 324 5805 336
rect 5759 -252 5765 324
rect 5799 -252 5805 324
rect 5759 -264 5805 -252
rect 5877 324 5923 336
rect 5877 -252 5883 324
rect 5917 -252 5923 324
rect 5877 -264 5923 -252
rect 5995 324 6041 336
rect 5995 -252 6001 324
rect 6035 -252 6041 324
rect 5995 -264 6041 -252
rect 6113 324 6159 336
rect 6113 -252 6119 324
rect 6153 -252 6159 324
rect 6113 -264 6159 -252
rect 6231 324 6277 336
rect 6231 -252 6237 324
rect 6271 -252 6277 324
rect 6231 -264 6277 -252
rect 6349 324 6395 336
rect 6349 -252 6355 324
rect 6389 -252 6395 324
rect 6349 -264 6395 -252
rect 6467 324 6513 336
rect 6467 -252 6473 324
rect 6507 -252 6513 324
rect 6467 -264 6513 -252
rect 6585 324 6631 336
rect 6585 -252 6591 324
rect 6625 -252 6631 324
rect 6585 -264 6631 -252
rect 6703 324 6749 336
rect 6703 -252 6709 324
rect 6743 -252 6749 324
rect 6703 -264 6749 -252
rect 6821 324 6867 336
rect 6821 -252 6827 324
rect 6861 -252 6867 324
rect 6821 -264 6867 -252
rect 6939 324 6985 336
rect 6939 -252 6945 324
rect 6979 -252 6985 324
rect 6939 -264 6985 -252
rect 7057 324 7103 336
rect 7057 -252 7063 324
rect 7097 -252 7103 324
rect 7057 -264 7103 -252
rect 7175 324 7221 336
rect 7175 -252 7181 324
rect 7215 -252 7221 324
rect 7175 -264 7221 -252
rect 7293 324 7339 336
rect 7293 -252 7299 324
rect 7333 -252 7339 324
rect 7293 -264 7339 -252
rect 7411 324 7457 336
rect 7411 -252 7417 324
rect 7451 -252 7457 324
rect 7411 -264 7457 -252
rect 7529 324 7575 336
rect 7529 -252 7535 324
rect 7569 -252 7575 324
rect 7529 -264 7575 -252
rect 7647 324 7693 336
rect 7647 -252 7653 324
rect 7687 -252 7693 324
rect 7647 -264 7693 -252
rect 7765 324 7811 336
rect 7765 -252 7771 324
rect 7805 -252 7811 324
rect 7765 -264 7811 -252
rect 7883 324 7929 336
rect 7883 -252 7889 324
rect 7923 -252 7929 324
rect 7883 -264 7929 -252
rect 8001 324 8047 336
rect 8001 -252 8007 324
rect 8041 -252 8047 324
rect 8001 -264 8047 -252
rect 8119 324 8165 336
rect 8119 -252 8125 324
rect 8159 -252 8165 324
rect 8119 -264 8165 -252
rect 8237 324 8283 336
rect 8237 -252 8243 324
rect 8277 -252 8283 324
rect 8237 -264 8283 -252
rect 8355 324 8401 336
rect 8355 -252 8361 324
rect 8395 -252 8401 324
rect 8355 -264 8401 -252
rect 8473 324 8519 336
rect 8473 -252 8479 324
rect 8513 -252 8519 324
rect 8473 -264 8519 -252
rect 8591 324 8637 336
rect 8591 -252 8597 324
rect 8631 -252 8637 324
rect 8591 -264 8637 -252
rect 8709 324 8755 336
rect 8709 -252 8715 324
rect 8749 -252 8755 324
rect 8709 -264 8755 -252
rect 8827 324 8873 336
rect 8827 -252 8833 324
rect 8867 -252 8873 324
rect 8827 -264 8873 -252
rect 8945 324 8991 336
rect 8945 -252 8951 324
rect 8985 -252 8991 324
rect 8945 -264 8991 -252
rect 9063 324 9109 336
rect 9063 -252 9069 324
rect 9103 -252 9109 324
rect 9063 -264 9109 -252
rect 9181 324 9227 336
rect 9181 -252 9187 324
rect 9221 -252 9227 324
rect 9181 -264 9227 -252
rect 9299 324 9345 336
rect 9299 -252 9305 324
rect 9339 -252 9345 324
rect 9299 -264 9345 -252
rect 9417 324 9463 336
rect 9417 -252 9423 324
rect 9457 -252 9463 324
rect 9417 -264 9463 -252
rect 9535 324 9581 336
rect 9535 -252 9541 324
rect 9575 -252 9581 324
rect 9535 -264 9581 -252
rect 9653 324 9699 336
rect 9653 -252 9659 324
rect 9693 -252 9699 324
rect 9653 -264 9699 -252
rect 9771 324 9817 336
rect 9771 -252 9777 324
rect 9811 -252 9817 324
rect 9771 -264 9817 -252
rect 9889 324 9935 336
rect 9889 -252 9895 324
rect 9929 -252 9935 324
rect 9889 -264 9935 -252
rect 10007 324 10053 336
rect 10007 -252 10013 324
rect 10047 -252 10053 324
rect 10007 -264 10053 -252
rect 10125 324 10171 336
rect 10125 -252 10131 324
rect 10165 -252 10171 324
rect 10125 -264 10171 -252
rect 10243 324 10289 336
rect 10243 -252 10249 324
rect 10283 -252 10289 324
rect 10243 -264 10289 -252
rect 10361 324 10407 336
rect 10361 -252 10367 324
rect 10401 -252 10407 324
rect 10361 -264 10407 -252
rect 10479 324 10525 336
rect 10479 -252 10485 324
rect 10519 -252 10525 324
rect 10479 -264 10525 -252
rect 10597 324 10643 336
rect 10597 -252 10603 324
rect 10637 -252 10643 324
rect 10597 -264 10643 -252
rect 10715 324 10761 336
rect 10715 -252 10721 324
rect 10755 -252 10761 324
rect 10715 -264 10761 -252
rect 10833 324 10879 336
rect 10833 -252 10839 324
rect 10873 -252 10879 324
rect 10833 -264 10879 -252
rect 10951 324 10997 336
rect 10951 -252 10957 324
rect 10991 -252 10997 324
rect 10951 -264 10997 -252
rect 11069 324 11115 336
rect 11069 -252 11075 324
rect 11109 -252 11115 324
rect 11069 -264 11115 -252
rect 11187 324 11233 336
rect 11187 -252 11193 324
rect 11227 -252 11233 324
rect 11187 -264 11233 -252
rect 11305 324 11351 336
rect 11305 -252 11311 324
rect 11345 -252 11351 324
rect 11305 -264 11351 -252
rect 11423 324 11469 336
rect 11423 -252 11429 324
rect 11463 -252 11469 324
rect 11423 -264 11469 -252
rect 11541 324 11587 336
rect 11541 -252 11547 324
rect 11581 -252 11587 324
rect 11541 -264 11587 -252
rect 11659 324 11705 336
rect 11659 -252 11665 324
rect 11699 -252 11705 324
rect 11659 -264 11705 -252
rect 11777 324 11823 336
rect 11777 -252 11783 324
rect 11817 -252 11823 324
rect 11777 -264 11823 -252
rect 11895 324 11941 336
rect 11895 -252 11901 324
rect 11935 -252 11941 324
rect 11895 -264 11941 -252
rect 12013 324 12059 336
rect 12013 -252 12019 324
rect 12053 -252 12059 324
rect 12013 -264 12059 -252
rect 12131 324 12177 336
rect 12131 -252 12137 324
rect 12171 -252 12177 324
rect 12131 -264 12177 -252
rect 12249 324 12295 336
rect 12249 -252 12255 324
rect 12289 -252 12295 324
rect 12249 -264 12295 -252
rect 12367 324 12413 336
rect 12367 -252 12373 324
rect 12407 -252 12413 324
rect 12367 -264 12413 -252
rect 12485 324 12531 336
rect 12485 -252 12491 324
rect 12525 -252 12531 324
rect 12485 -264 12531 -252
rect 12603 324 12649 336
rect 12603 -252 12609 324
rect 12643 -252 12649 324
rect 12603 -264 12649 -252
rect 12721 324 12767 336
rect 12721 -252 12727 324
rect 12761 -252 12767 324
rect 12721 -264 12767 -252
rect 12839 324 12885 336
rect 12839 -252 12845 324
rect 12879 -252 12885 324
rect 12839 -264 12885 -252
rect 12957 324 13003 336
rect 12957 -252 12963 324
rect 12997 -252 13003 324
rect 12957 -264 13003 -252
rect 13075 324 13121 336
rect 13075 -252 13081 324
rect 13115 -252 13121 324
rect 13075 -264 13121 -252
rect 13193 324 13239 336
rect 13193 -252 13199 324
rect 13233 -252 13239 324
rect 13193 -264 13239 -252
rect 13311 324 13357 336
rect 13311 -252 13317 324
rect 13351 -252 13357 324
rect 13311 -264 13357 -252
rect 13429 324 13475 336
rect 13429 -252 13435 324
rect 13469 -252 13475 324
rect 13429 -264 13475 -252
rect 13547 324 13593 336
rect 13547 -252 13553 324
rect 13587 -252 13593 324
rect 13547 -264 13593 -252
rect 13665 324 13711 336
rect 13665 -252 13671 324
rect 13705 -252 13711 324
rect 13665 -264 13711 -252
rect 13783 324 13829 336
rect 13783 -252 13789 324
rect 13823 -252 13829 324
rect 13783 -264 13829 -252
rect 13901 324 13947 336
rect 13901 -252 13907 324
rect 13941 -252 13947 324
rect 13901 -264 13947 -252
rect 14019 324 14065 336
rect 14019 -252 14025 324
rect 14059 -252 14065 324
rect 14019 -264 14065 -252
rect 14137 324 14183 336
rect 14137 -252 14143 324
rect 14177 -252 14183 324
rect 14137 -264 14183 -252
rect 14255 324 14301 336
rect 14255 -252 14261 324
rect 14295 -252 14301 324
rect 14255 -264 14301 -252
rect 14373 324 14419 336
rect 14373 -252 14379 324
rect 14413 -252 14419 324
rect 14373 -264 14419 -252
rect 14491 324 14537 336
rect 14491 -252 14497 324
rect 14531 -252 14537 324
rect 14491 -264 14537 -252
rect 14609 324 14655 336
rect 14609 -252 14615 324
rect 14649 -252 14655 324
rect 14609 -264 14655 -252
rect 14727 324 14773 336
rect 14727 -252 14733 324
rect 14767 -252 14773 324
rect 14727 -264 14773 -252
rect -14720 -311 -14662 -305
rect -14720 -345 -14708 -311
rect -14674 -345 -14662 -311
rect -14720 -351 -14662 -345
rect -14602 -311 -14544 -305
rect -14602 -345 -14590 -311
rect -14556 -345 -14544 -311
rect -14602 -351 -14544 -345
rect -14484 -311 -14426 -305
rect -14484 -345 -14472 -311
rect -14438 -345 -14426 -311
rect -14484 -351 -14426 -345
rect -14366 -311 -14308 -305
rect -14366 -345 -14354 -311
rect -14320 -345 -14308 -311
rect -14366 -351 -14308 -345
rect -14248 -311 -14190 -305
rect -14248 -345 -14236 -311
rect -14202 -345 -14190 -311
rect -14248 -351 -14190 -345
rect -14130 -311 -14072 -305
rect -14130 -345 -14118 -311
rect -14084 -345 -14072 -311
rect -14130 -351 -14072 -345
rect -14012 -311 -13954 -305
rect -14012 -345 -14000 -311
rect -13966 -345 -13954 -311
rect -14012 -351 -13954 -345
rect -13894 -311 -13836 -305
rect -13894 -345 -13882 -311
rect -13848 -345 -13836 -311
rect -13894 -351 -13836 -345
rect -13776 -311 -13718 -305
rect -13776 -345 -13764 -311
rect -13730 -345 -13718 -311
rect -13776 -351 -13718 -345
rect -13658 -311 -13600 -305
rect -13658 -345 -13646 -311
rect -13612 -345 -13600 -311
rect -13658 -351 -13600 -345
rect -13540 -311 -13482 -305
rect -13540 -345 -13528 -311
rect -13494 -345 -13482 -311
rect -13540 -351 -13482 -345
rect -13422 -311 -13364 -305
rect -13422 -345 -13410 -311
rect -13376 -345 -13364 -311
rect -13422 -351 -13364 -345
rect -13304 -311 -13246 -305
rect -13304 -345 -13292 -311
rect -13258 -345 -13246 -311
rect -13304 -351 -13246 -345
rect -13186 -311 -13128 -305
rect -13186 -345 -13174 -311
rect -13140 -345 -13128 -311
rect -13186 -351 -13128 -345
rect -13068 -311 -13010 -305
rect -13068 -345 -13056 -311
rect -13022 -345 -13010 -311
rect -13068 -351 -13010 -345
rect -12950 -311 -12892 -305
rect -12950 -345 -12938 -311
rect -12904 -345 -12892 -311
rect -12950 -351 -12892 -345
rect -12832 -311 -12774 -305
rect -12832 -345 -12820 -311
rect -12786 -345 -12774 -311
rect -12832 -351 -12774 -345
rect -12714 -311 -12656 -305
rect -12714 -345 -12702 -311
rect -12668 -345 -12656 -311
rect -12714 -351 -12656 -345
rect -12596 -311 -12538 -305
rect -12596 -345 -12584 -311
rect -12550 -345 -12538 -311
rect -12596 -351 -12538 -345
rect -12478 -311 -12420 -305
rect -12478 -345 -12466 -311
rect -12432 -345 -12420 -311
rect -12478 -351 -12420 -345
rect -12360 -311 -12302 -305
rect -12360 -345 -12348 -311
rect -12314 -345 -12302 -311
rect -12360 -351 -12302 -345
rect -12242 -311 -12184 -305
rect -12242 -345 -12230 -311
rect -12196 -345 -12184 -311
rect -12242 -351 -12184 -345
rect -12124 -311 -12066 -305
rect -12124 -345 -12112 -311
rect -12078 -345 -12066 -311
rect -12124 -351 -12066 -345
rect -12006 -311 -11948 -305
rect -12006 -345 -11994 -311
rect -11960 -345 -11948 -311
rect -12006 -351 -11948 -345
rect -11888 -311 -11830 -305
rect -11888 -345 -11876 -311
rect -11842 -345 -11830 -311
rect -11888 -351 -11830 -345
rect -11770 -311 -11712 -305
rect -11770 -345 -11758 -311
rect -11724 -345 -11712 -311
rect -11770 -351 -11712 -345
rect -11652 -311 -11594 -305
rect -11652 -345 -11640 -311
rect -11606 -345 -11594 -311
rect -11652 -351 -11594 -345
rect -11534 -311 -11476 -305
rect -11534 -345 -11522 -311
rect -11488 -345 -11476 -311
rect -11534 -351 -11476 -345
rect -11416 -311 -11358 -305
rect -11416 -345 -11404 -311
rect -11370 -345 -11358 -311
rect -11416 -351 -11358 -345
rect -11298 -311 -11240 -305
rect -11298 -345 -11286 -311
rect -11252 -345 -11240 -311
rect -11298 -351 -11240 -345
rect -11180 -311 -11122 -305
rect -11180 -345 -11168 -311
rect -11134 -345 -11122 -311
rect -11180 -351 -11122 -345
rect -11062 -311 -11004 -305
rect -11062 -345 -11050 -311
rect -11016 -345 -11004 -311
rect -11062 -351 -11004 -345
rect -10944 -311 -10886 -305
rect -10944 -345 -10932 -311
rect -10898 -345 -10886 -311
rect -10944 -351 -10886 -345
rect -10826 -311 -10768 -305
rect -10826 -345 -10814 -311
rect -10780 -345 -10768 -311
rect -10826 -351 -10768 -345
rect -10708 -311 -10650 -305
rect -10708 -345 -10696 -311
rect -10662 -345 -10650 -311
rect -10708 -351 -10650 -345
rect -10590 -311 -10532 -305
rect -10590 -345 -10578 -311
rect -10544 -345 -10532 -311
rect -10590 -351 -10532 -345
rect -10472 -311 -10414 -305
rect -10472 -345 -10460 -311
rect -10426 -345 -10414 -311
rect -10472 -351 -10414 -345
rect -10354 -311 -10296 -305
rect -10354 -345 -10342 -311
rect -10308 -345 -10296 -311
rect -10354 -351 -10296 -345
rect -10236 -311 -10178 -305
rect -10236 -345 -10224 -311
rect -10190 -345 -10178 -311
rect -10236 -351 -10178 -345
rect -10118 -311 -10060 -305
rect -10118 -345 -10106 -311
rect -10072 -345 -10060 -311
rect -10118 -351 -10060 -345
rect -10000 -311 -9942 -305
rect -10000 -345 -9988 -311
rect -9954 -345 -9942 -311
rect -10000 -351 -9942 -345
rect -9882 -311 -9824 -305
rect -9882 -345 -9870 -311
rect -9836 -345 -9824 -311
rect -9882 -351 -9824 -345
rect -9764 -311 -9706 -305
rect -9764 -345 -9752 -311
rect -9718 -345 -9706 -311
rect -9764 -351 -9706 -345
rect -9646 -311 -9588 -305
rect -9646 -345 -9634 -311
rect -9600 -345 -9588 -311
rect -9646 -351 -9588 -345
rect -9528 -311 -9470 -305
rect -9528 -345 -9516 -311
rect -9482 -345 -9470 -311
rect -9528 -351 -9470 -345
rect -9410 -311 -9352 -305
rect -9410 -345 -9398 -311
rect -9364 -345 -9352 -311
rect -9410 -351 -9352 -345
rect -9292 -311 -9234 -305
rect -9292 -345 -9280 -311
rect -9246 -345 -9234 -311
rect -9292 -351 -9234 -345
rect -9174 -311 -9116 -305
rect -9174 -345 -9162 -311
rect -9128 -345 -9116 -311
rect -9174 -351 -9116 -345
rect -9056 -311 -8998 -305
rect -9056 -345 -9044 -311
rect -9010 -345 -8998 -311
rect -9056 -351 -8998 -345
rect -8938 -311 -8880 -305
rect -8938 -345 -8926 -311
rect -8892 -345 -8880 -311
rect -8938 -351 -8880 -345
rect -8820 -311 -8762 -305
rect -8820 -345 -8808 -311
rect -8774 -345 -8762 -311
rect -8820 -351 -8762 -345
rect -8702 -311 -8644 -305
rect -8702 -345 -8690 -311
rect -8656 -345 -8644 -311
rect -8702 -351 -8644 -345
rect -8584 -311 -8526 -305
rect -8584 -345 -8572 -311
rect -8538 -345 -8526 -311
rect -8584 -351 -8526 -345
rect -8466 -311 -8408 -305
rect -8466 -345 -8454 -311
rect -8420 -345 -8408 -311
rect -8466 -351 -8408 -345
rect -8348 -311 -8290 -305
rect -8348 -345 -8336 -311
rect -8302 -345 -8290 -311
rect -8348 -351 -8290 -345
rect -8230 -311 -8172 -305
rect -8230 -345 -8218 -311
rect -8184 -345 -8172 -311
rect -8230 -351 -8172 -345
rect -8112 -311 -8054 -305
rect -8112 -345 -8100 -311
rect -8066 -345 -8054 -311
rect -8112 -351 -8054 -345
rect -7994 -311 -7936 -305
rect -7994 -345 -7982 -311
rect -7948 -345 -7936 -311
rect -7994 -351 -7936 -345
rect -7876 -311 -7818 -305
rect -7876 -345 -7864 -311
rect -7830 -345 -7818 -311
rect -7876 -351 -7818 -345
rect -7758 -311 -7700 -305
rect -7758 -345 -7746 -311
rect -7712 -345 -7700 -311
rect -7758 -351 -7700 -345
rect -7640 -311 -7582 -305
rect -7640 -345 -7628 -311
rect -7594 -345 -7582 -311
rect -7640 -351 -7582 -345
rect -7522 -311 -7464 -305
rect -7522 -345 -7510 -311
rect -7476 -345 -7464 -311
rect -7522 -351 -7464 -345
rect -7404 -311 -7346 -305
rect -7404 -345 -7392 -311
rect -7358 -345 -7346 -311
rect -7404 -351 -7346 -345
rect -7286 -311 -7228 -305
rect -7286 -345 -7274 -311
rect -7240 -345 -7228 -311
rect -7286 -351 -7228 -345
rect -7168 -311 -7110 -305
rect -7168 -345 -7156 -311
rect -7122 -345 -7110 -311
rect -7168 -351 -7110 -345
rect -7050 -311 -6992 -305
rect -7050 -345 -7038 -311
rect -7004 -345 -6992 -311
rect -7050 -351 -6992 -345
rect -6932 -311 -6874 -305
rect -6932 -345 -6920 -311
rect -6886 -345 -6874 -311
rect -6932 -351 -6874 -345
rect -6814 -311 -6756 -305
rect -6814 -345 -6802 -311
rect -6768 -345 -6756 -311
rect -6814 -351 -6756 -345
rect -6696 -311 -6638 -305
rect -6696 -345 -6684 -311
rect -6650 -345 -6638 -311
rect -6696 -351 -6638 -345
rect -6578 -311 -6520 -305
rect -6578 -345 -6566 -311
rect -6532 -345 -6520 -311
rect -6578 -351 -6520 -345
rect -6460 -311 -6402 -305
rect -6460 -345 -6448 -311
rect -6414 -345 -6402 -311
rect -6460 -351 -6402 -345
rect -6342 -311 -6284 -305
rect -6342 -345 -6330 -311
rect -6296 -345 -6284 -311
rect -6342 -351 -6284 -345
rect -6224 -311 -6166 -305
rect -6224 -345 -6212 -311
rect -6178 -345 -6166 -311
rect -6224 -351 -6166 -345
rect -6106 -311 -6048 -305
rect -6106 -345 -6094 -311
rect -6060 -345 -6048 -311
rect -6106 -351 -6048 -345
rect -5988 -311 -5930 -305
rect -5988 -345 -5976 -311
rect -5942 -345 -5930 -311
rect -5988 -351 -5930 -345
rect -5870 -311 -5812 -305
rect -5870 -345 -5858 -311
rect -5824 -345 -5812 -311
rect -5870 -351 -5812 -345
rect -5752 -311 -5694 -305
rect -5752 -345 -5740 -311
rect -5706 -345 -5694 -311
rect -5752 -351 -5694 -345
rect -5634 -311 -5576 -305
rect -5634 -345 -5622 -311
rect -5588 -345 -5576 -311
rect -5634 -351 -5576 -345
rect -5516 -311 -5458 -305
rect -5516 -345 -5504 -311
rect -5470 -345 -5458 -311
rect -5516 -351 -5458 -345
rect -5398 -311 -5340 -305
rect -5398 -345 -5386 -311
rect -5352 -345 -5340 -311
rect -5398 -351 -5340 -345
rect -5280 -311 -5222 -305
rect -5280 -345 -5268 -311
rect -5234 -345 -5222 -311
rect -5280 -351 -5222 -345
rect -5162 -311 -5104 -305
rect -5162 -345 -5150 -311
rect -5116 -345 -5104 -311
rect -5162 -351 -5104 -345
rect -5044 -311 -4986 -305
rect -5044 -345 -5032 -311
rect -4998 -345 -4986 -311
rect -5044 -351 -4986 -345
rect -4926 -311 -4868 -305
rect -4926 -345 -4914 -311
rect -4880 -345 -4868 -311
rect -4926 -351 -4868 -345
rect -4808 -311 -4750 -305
rect -4808 -345 -4796 -311
rect -4762 -345 -4750 -311
rect -4808 -351 -4750 -345
rect -4690 -311 -4632 -305
rect -4690 -345 -4678 -311
rect -4644 -345 -4632 -311
rect -4690 -351 -4632 -345
rect -4572 -311 -4514 -305
rect -4572 -345 -4560 -311
rect -4526 -345 -4514 -311
rect -4572 -351 -4514 -345
rect -4454 -311 -4396 -305
rect -4454 -345 -4442 -311
rect -4408 -345 -4396 -311
rect -4454 -351 -4396 -345
rect -4336 -311 -4278 -305
rect -4336 -345 -4324 -311
rect -4290 -345 -4278 -311
rect -4336 -351 -4278 -345
rect -4218 -311 -4160 -305
rect -4218 -345 -4206 -311
rect -4172 -345 -4160 -311
rect -4218 -351 -4160 -345
rect -4100 -311 -4042 -305
rect -4100 -345 -4088 -311
rect -4054 -345 -4042 -311
rect -4100 -351 -4042 -345
rect -3982 -311 -3924 -305
rect -3982 -345 -3970 -311
rect -3936 -345 -3924 -311
rect -3982 -351 -3924 -345
rect -3864 -311 -3806 -305
rect -3864 -345 -3852 -311
rect -3818 -345 -3806 -311
rect -3864 -351 -3806 -345
rect -3746 -311 -3688 -305
rect -3746 -345 -3734 -311
rect -3700 -345 -3688 -311
rect -3746 -351 -3688 -345
rect -3628 -311 -3570 -305
rect -3628 -345 -3616 -311
rect -3582 -345 -3570 -311
rect -3628 -351 -3570 -345
rect -3510 -311 -3452 -305
rect -3510 -345 -3498 -311
rect -3464 -345 -3452 -311
rect -3510 -351 -3452 -345
rect -3392 -311 -3334 -305
rect -3392 -345 -3380 -311
rect -3346 -345 -3334 -311
rect -3392 -351 -3334 -345
rect -3274 -311 -3216 -305
rect -3274 -345 -3262 -311
rect -3228 -345 -3216 -311
rect -3274 -351 -3216 -345
rect -3156 -311 -3098 -305
rect -3156 -345 -3144 -311
rect -3110 -345 -3098 -311
rect -3156 -351 -3098 -345
rect -3038 -311 -2980 -305
rect -3038 -345 -3026 -311
rect -2992 -345 -2980 -311
rect -3038 -351 -2980 -345
rect -2920 -311 -2862 -305
rect -2920 -345 -2908 -311
rect -2874 -345 -2862 -311
rect -2920 -351 -2862 -345
rect -2802 -311 -2744 -305
rect -2802 -345 -2790 -311
rect -2756 -345 -2744 -311
rect -2802 -351 -2744 -345
rect -2684 -311 -2626 -305
rect -2684 -345 -2672 -311
rect -2638 -345 -2626 -311
rect -2684 -351 -2626 -345
rect -2566 -311 -2508 -305
rect -2566 -345 -2554 -311
rect -2520 -345 -2508 -311
rect -2566 -351 -2508 -345
rect -2448 -311 -2390 -305
rect -2448 -345 -2436 -311
rect -2402 -345 -2390 -311
rect -2448 -351 -2390 -345
rect -2330 -311 -2272 -305
rect -2330 -345 -2318 -311
rect -2284 -345 -2272 -311
rect -2330 -351 -2272 -345
rect -2212 -311 -2154 -305
rect -2212 -345 -2200 -311
rect -2166 -345 -2154 -311
rect -2212 -351 -2154 -345
rect -2094 -311 -2036 -305
rect -2094 -345 -2082 -311
rect -2048 -345 -2036 -311
rect -2094 -351 -2036 -345
rect -1976 -311 -1918 -305
rect -1976 -345 -1964 -311
rect -1930 -345 -1918 -311
rect -1976 -351 -1918 -345
rect -1858 -311 -1800 -305
rect -1858 -345 -1846 -311
rect -1812 -345 -1800 -311
rect -1858 -351 -1800 -345
rect -1740 -311 -1682 -305
rect -1740 -345 -1728 -311
rect -1694 -345 -1682 -311
rect -1740 -351 -1682 -345
rect -1622 -311 -1564 -305
rect -1622 -345 -1610 -311
rect -1576 -345 -1564 -311
rect -1622 -351 -1564 -345
rect -1504 -311 -1446 -305
rect -1504 -345 -1492 -311
rect -1458 -345 -1446 -311
rect -1504 -351 -1446 -345
rect -1386 -311 -1328 -305
rect -1386 -345 -1374 -311
rect -1340 -345 -1328 -311
rect -1386 -351 -1328 -345
rect -1268 -311 -1210 -305
rect -1268 -345 -1256 -311
rect -1222 -345 -1210 -311
rect -1268 -351 -1210 -345
rect -1150 -311 -1092 -305
rect -1150 -345 -1138 -311
rect -1104 -345 -1092 -311
rect -1150 -351 -1092 -345
rect -1032 -311 -974 -305
rect -1032 -345 -1020 -311
rect -986 -345 -974 -311
rect -1032 -351 -974 -345
rect -914 -311 -856 -305
rect -914 -345 -902 -311
rect -868 -345 -856 -311
rect -914 -351 -856 -345
rect -796 -311 -738 -305
rect -796 -345 -784 -311
rect -750 -345 -738 -311
rect -796 -351 -738 -345
rect -678 -311 -620 -305
rect -678 -345 -666 -311
rect -632 -345 -620 -311
rect -678 -351 -620 -345
rect -560 -311 -502 -305
rect -560 -345 -548 -311
rect -514 -345 -502 -311
rect -560 -351 -502 -345
rect -442 -311 -384 -305
rect -442 -345 -430 -311
rect -396 -345 -384 -311
rect -442 -351 -384 -345
rect -324 -311 -266 -305
rect -324 -345 -312 -311
rect -278 -345 -266 -311
rect -324 -351 -266 -345
rect -206 -311 -148 -305
rect -206 -345 -194 -311
rect -160 -345 -148 -311
rect -206 -351 -148 -345
rect -88 -311 -30 -305
rect -88 -345 -76 -311
rect -42 -345 -30 -311
rect -88 -351 -30 -345
rect 30 -311 88 -305
rect 30 -345 42 -311
rect 76 -345 88 -311
rect 30 -351 88 -345
rect 148 -311 206 -305
rect 148 -345 160 -311
rect 194 -345 206 -311
rect 148 -351 206 -345
rect 266 -311 324 -305
rect 266 -345 278 -311
rect 312 -345 324 -311
rect 266 -351 324 -345
rect 384 -311 442 -305
rect 384 -345 396 -311
rect 430 -345 442 -311
rect 384 -351 442 -345
rect 502 -311 560 -305
rect 502 -345 514 -311
rect 548 -345 560 -311
rect 502 -351 560 -345
rect 620 -311 678 -305
rect 620 -345 632 -311
rect 666 -345 678 -311
rect 620 -351 678 -345
rect 738 -311 796 -305
rect 738 -345 750 -311
rect 784 -345 796 -311
rect 738 -351 796 -345
rect 856 -311 914 -305
rect 856 -345 868 -311
rect 902 -345 914 -311
rect 856 -351 914 -345
rect 974 -311 1032 -305
rect 974 -345 986 -311
rect 1020 -345 1032 -311
rect 974 -351 1032 -345
rect 1092 -311 1150 -305
rect 1092 -345 1104 -311
rect 1138 -345 1150 -311
rect 1092 -351 1150 -345
rect 1210 -311 1268 -305
rect 1210 -345 1222 -311
rect 1256 -345 1268 -311
rect 1210 -351 1268 -345
rect 1328 -311 1386 -305
rect 1328 -345 1340 -311
rect 1374 -345 1386 -311
rect 1328 -351 1386 -345
rect 1446 -311 1504 -305
rect 1446 -345 1458 -311
rect 1492 -345 1504 -311
rect 1446 -351 1504 -345
rect 1564 -311 1622 -305
rect 1564 -345 1576 -311
rect 1610 -345 1622 -311
rect 1564 -351 1622 -345
rect 1682 -311 1740 -305
rect 1682 -345 1694 -311
rect 1728 -345 1740 -311
rect 1682 -351 1740 -345
rect 1800 -311 1858 -305
rect 1800 -345 1812 -311
rect 1846 -345 1858 -311
rect 1800 -351 1858 -345
rect 1918 -311 1976 -305
rect 1918 -345 1930 -311
rect 1964 -345 1976 -311
rect 1918 -351 1976 -345
rect 2036 -311 2094 -305
rect 2036 -345 2048 -311
rect 2082 -345 2094 -311
rect 2036 -351 2094 -345
rect 2154 -311 2212 -305
rect 2154 -345 2166 -311
rect 2200 -345 2212 -311
rect 2154 -351 2212 -345
rect 2272 -311 2330 -305
rect 2272 -345 2284 -311
rect 2318 -345 2330 -311
rect 2272 -351 2330 -345
rect 2390 -311 2448 -305
rect 2390 -345 2402 -311
rect 2436 -345 2448 -311
rect 2390 -351 2448 -345
rect 2508 -311 2566 -305
rect 2508 -345 2520 -311
rect 2554 -345 2566 -311
rect 2508 -351 2566 -345
rect 2626 -311 2684 -305
rect 2626 -345 2638 -311
rect 2672 -345 2684 -311
rect 2626 -351 2684 -345
rect 2744 -311 2802 -305
rect 2744 -345 2756 -311
rect 2790 -345 2802 -311
rect 2744 -351 2802 -345
rect 2862 -311 2920 -305
rect 2862 -345 2874 -311
rect 2908 -345 2920 -311
rect 2862 -351 2920 -345
rect 2980 -311 3038 -305
rect 2980 -345 2992 -311
rect 3026 -345 3038 -311
rect 2980 -351 3038 -345
rect 3098 -311 3156 -305
rect 3098 -345 3110 -311
rect 3144 -345 3156 -311
rect 3098 -351 3156 -345
rect 3216 -311 3274 -305
rect 3216 -345 3228 -311
rect 3262 -345 3274 -311
rect 3216 -351 3274 -345
rect 3334 -311 3392 -305
rect 3334 -345 3346 -311
rect 3380 -345 3392 -311
rect 3334 -351 3392 -345
rect 3452 -311 3510 -305
rect 3452 -345 3464 -311
rect 3498 -345 3510 -311
rect 3452 -351 3510 -345
rect 3570 -311 3628 -305
rect 3570 -345 3582 -311
rect 3616 -345 3628 -311
rect 3570 -351 3628 -345
rect 3688 -311 3746 -305
rect 3688 -345 3700 -311
rect 3734 -345 3746 -311
rect 3688 -351 3746 -345
rect 3806 -311 3864 -305
rect 3806 -345 3818 -311
rect 3852 -345 3864 -311
rect 3806 -351 3864 -345
rect 3924 -311 3982 -305
rect 3924 -345 3936 -311
rect 3970 -345 3982 -311
rect 3924 -351 3982 -345
rect 4042 -311 4100 -305
rect 4042 -345 4054 -311
rect 4088 -345 4100 -311
rect 4042 -351 4100 -345
rect 4160 -311 4218 -305
rect 4160 -345 4172 -311
rect 4206 -345 4218 -311
rect 4160 -351 4218 -345
rect 4278 -311 4336 -305
rect 4278 -345 4290 -311
rect 4324 -345 4336 -311
rect 4278 -351 4336 -345
rect 4396 -311 4454 -305
rect 4396 -345 4408 -311
rect 4442 -345 4454 -311
rect 4396 -351 4454 -345
rect 4514 -311 4572 -305
rect 4514 -345 4526 -311
rect 4560 -345 4572 -311
rect 4514 -351 4572 -345
rect 4632 -311 4690 -305
rect 4632 -345 4644 -311
rect 4678 -345 4690 -311
rect 4632 -351 4690 -345
rect 4750 -311 4808 -305
rect 4750 -345 4762 -311
rect 4796 -345 4808 -311
rect 4750 -351 4808 -345
rect 4868 -311 4926 -305
rect 4868 -345 4880 -311
rect 4914 -345 4926 -311
rect 4868 -351 4926 -345
rect 4986 -311 5044 -305
rect 4986 -345 4998 -311
rect 5032 -345 5044 -311
rect 4986 -351 5044 -345
rect 5104 -311 5162 -305
rect 5104 -345 5116 -311
rect 5150 -345 5162 -311
rect 5104 -351 5162 -345
rect 5222 -311 5280 -305
rect 5222 -345 5234 -311
rect 5268 -345 5280 -311
rect 5222 -351 5280 -345
rect 5340 -311 5398 -305
rect 5340 -345 5352 -311
rect 5386 -345 5398 -311
rect 5340 -351 5398 -345
rect 5458 -311 5516 -305
rect 5458 -345 5470 -311
rect 5504 -345 5516 -311
rect 5458 -351 5516 -345
rect 5576 -311 5634 -305
rect 5576 -345 5588 -311
rect 5622 -345 5634 -311
rect 5576 -351 5634 -345
rect 5694 -311 5752 -305
rect 5694 -345 5706 -311
rect 5740 -345 5752 -311
rect 5694 -351 5752 -345
rect 5812 -311 5870 -305
rect 5812 -345 5824 -311
rect 5858 -345 5870 -311
rect 5812 -351 5870 -345
rect 5930 -311 5988 -305
rect 5930 -345 5942 -311
rect 5976 -345 5988 -311
rect 5930 -351 5988 -345
rect 6048 -311 6106 -305
rect 6048 -345 6060 -311
rect 6094 -345 6106 -311
rect 6048 -351 6106 -345
rect 6166 -311 6224 -305
rect 6166 -345 6178 -311
rect 6212 -345 6224 -311
rect 6166 -351 6224 -345
rect 6284 -311 6342 -305
rect 6284 -345 6296 -311
rect 6330 -345 6342 -311
rect 6284 -351 6342 -345
rect 6402 -311 6460 -305
rect 6402 -345 6414 -311
rect 6448 -345 6460 -311
rect 6402 -351 6460 -345
rect 6520 -311 6578 -305
rect 6520 -345 6532 -311
rect 6566 -345 6578 -311
rect 6520 -351 6578 -345
rect 6638 -311 6696 -305
rect 6638 -345 6650 -311
rect 6684 -345 6696 -311
rect 6638 -351 6696 -345
rect 6756 -311 6814 -305
rect 6756 -345 6768 -311
rect 6802 -345 6814 -311
rect 6756 -351 6814 -345
rect 6874 -311 6932 -305
rect 6874 -345 6886 -311
rect 6920 -345 6932 -311
rect 6874 -351 6932 -345
rect 6992 -311 7050 -305
rect 6992 -345 7004 -311
rect 7038 -345 7050 -311
rect 6992 -351 7050 -345
rect 7110 -311 7168 -305
rect 7110 -345 7122 -311
rect 7156 -345 7168 -311
rect 7110 -351 7168 -345
rect 7228 -311 7286 -305
rect 7228 -345 7240 -311
rect 7274 -345 7286 -311
rect 7228 -351 7286 -345
rect 7346 -311 7404 -305
rect 7346 -345 7358 -311
rect 7392 -345 7404 -311
rect 7346 -351 7404 -345
rect 7464 -311 7522 -305
rect 7464 -345 7476 -311
rect 7510 -345 7522 -311
rect 7464 -351 7522 -345
rect 7582 -311 7640 -305
rect 7582 -345 7594 -311
rect 7628 -345 7640 -311
rect 7582 -351 7640 -345
rect 7700 -311 7758 -305
rect 7700 -345 7712 -311
rect 7746 -345 7758 -311
rect 7700 -351 7758 -345
rect 7818 -311 7876 -305
rect 7818 -345 7830 -311
rect 7864 -345 7876 -311
rect 7818 -351 7876 -345
rect 7936 -311 7994 -305
rect 7936 -345 7948 -311
rect 7982 -345 7994 -311
rect 7936 -351 7994 -345
rect 8054 -311 8112 -305
rect 8054 -345 8066 -311
rect 8100 -345 8112 -311
rect 8054 -351 8112 -345
rect 8172 -311 8230 -305
rect 8172 -345 8184 -311
rect 8218 -345 8230 -311
rect 8172 -351 8230 -345
rect 8290 -311 8348 -305
rect 8290 -345 8302 -311
rect 8336 -345 8348 -311
rect 8290 -351 8348 -345
rect 8408 -311 8466 -305
rect 8408 -345 8420 -311
rect 8454 -345 8466 -311
rect 8408 -351 8466 -345
rect 8526 -311 8584 -305
rect 8526 -345 8538 -311
rect 8572 -345 8584 -311
rect 8526 -351 8584 -345
rect 8644 -311 8702 -305
rect 8644 -345 8656 -311
rect 8690 -345 8702 -311
rect 8644 -351 8702 -345
rect 8762 -311 8820 -305
rect 8762 -345 8774 -311
rect 8808 -345 8820 -311
rect 8762 -351 8820 -345
rect 8880 -311 8938 -305
rect 8880 -345 8892 -311
rect 8926 -345 8938 -311
rect 8880 -351 8938 -345
rect 8998 -311 9056 -305
rect 8998 -345 9010 -311
rect 9044 -345 9056 -311
rect 8998 -351 9056 -345
rect 9116 -311 9174 -305
rect 9116 -345 9128 -311
rect 9162 -345 9174 -311
rect 9116 -351 9174 -345
rect 9234 -311 9292 -305
rect 9234 -345 9246 -311
rect 9280 -345 9292 -311
rect 9234 -351 9292 -345
rect 9352 -311 9410 -305
rect 9352 -345 9364 -311
rect 9398 -345 9410 -311
rect 9352 -351 9410 -345
rect 9470 -311 9528 -305
rect 9470 -345 9482 -311
rect 9516 -345 9528 -311
rect 9470 -351 9528 -345
rect 9588 -311 9646 -305
rect 9588 -345 9600 -311
rect 9634 -345 9646 -311
rect 9588 -351 9646 -345
rect 9706 -311 9764 -305
rect 9706 -345 9718 -311
rect 9752 -345 9764 -311
rect 9706 -351 9764 -345
rect 9824 -311 9882 -305
rect 9824 -345 9836 -311
rect 9870 -345 9882 -311
rect 9824 -351 9882 -345
rect 9942 -311 10000 -305
rect 9942 -345 9954 -311
rect 9988 -345 10000 -311
rect 9942 -351 10000 -345
rect 10060 -311 10118 -305
rect 10060 -345 10072 -311
rect 10106 -345 10118 -311
rect 10060 -351 10118 -345
rect 10178 -311 10236 -305
rect 10178 -345 10190 -311
rect 10224 -345 10236 -311
rect 10178 -351 10236 -345
rect 10296 -311 10354 -305
rect 10296 -345 10308 -311
rect 10342 -345 10354 -311
rect 10296 -351 10354 -345
rect 10414 -311 10472 -305
rect 10414 -345 10426 -311
rect 10460 -345 10472 -311
rect 10414 -351 10472 -345
rect 10532 -311 10590 -305
rect 10532 -345 10544 -311
rect 10578 -345 10590 -311
rect 10532 -351 10590 -345
rect 10650 -311 10708 -305
rect 10650 -345 10662 -311
rect 10696 -345 10708 -311
rect 10650 -351 10708 -345
rect 10768 -311 10826 -305
rect 10768 -345 10780 -311
rect 10814 -345 10826 -311
rect 10768 -351 10826 -345
rect 10886 -311 10944 -305
rect 10886 -345 10898 -311
rect 10932 -345 10944 -311
rect 10886 -351 10944 -345
rect 11004 -311 11062 -305
rect 11004 -345 11016 -311
rect 11050 -345 11062 -311
rect 11004 -351 11062 -345
rect 11122 -311 11180 -305
rect 11122 -345 11134 -311
rect 11168 -345 11180 -311
rect 11122 -351 11180 -345
rect 11240 -311 11298 -305
rect 11240 -345 11252 -311
rect 11286 -345 11298 -311
rect 11240 -351 11298 -345
rect 11358 -311 11416 -305
rect 11358 -345 11370 -311
rect 11404 -345 11416 -311
rect 11358 -351 11416 -345
rect 11476 -311 11534 -305
rect 11476 -345 11488 -311
rect 11522 -345 11534 -311
rect 11476 -351 11534 -345
rect 11594 -311 11652 -305
rect 11594 -345 11606 -311
rect 11640 -345 11652 -311
rect 11594 -351 11652 -345
rect 11712 -311 11770 -305
rect 11712 -345 11724 -311
rect 11758 -345 11770 -311
rect 11712 -351 11770 -345
rect 11830 -311 11888 -305
rect 11830 -345 11842 -311
rect 11876 -345 11888 -311
rect 11830 -351 11888 -345
rect 11948 -311 12006 -305
rect 11948 -345 11960 -311
rect 11994 -345 12006 -311
rect 11948 -351 12006 -345
rect 12066 -311 12124 -305
rect 12066 -345 12078 -311
rect 12112 -345 12124 -311
rect 12066 -351 12124 -345
rect 12184 -311 12242 -305
rect 12184 -345 12196 -311
rect 12230 -345 12242 -311
rect 12184 -351 12242 -345
rect 12302 -311 12360 -305
rect 12302 -345 12314 -311
rect 12348 -345 12360 -311
rect 12302 -351 12360 -345
rect 12420 -311 12478 -305
rect 12420 -345 12432 -311
rect 12466 -345 12478 -311
rect 12420 -351 12478 -345
rect 12538 -311 12596 -305
rect 12538 -345 12550 -311
rect 12584 -345 12596 -311
rect 12538 -351 12596 -345
rect 12656 -311 12714 -305
rect 12656 -345 12668 -311
rect 12702 -345 12714 -311
rect 12656 -351 12714 -345
rect 12774 -311 12832 -305
rect 12774 -345 12786 -311
rect 12820 -345 12832 -311
rect 12774 -351 12832 -345
rect 12892 -311 12950 -305
rect 12892 -345 12904 -311
rect 12938 -345 12950 -311
rect 12892 -351 12950 -345
rect 13010 -311 13068 -305
rect 13010 -345 13022 -311
rect 13056 -345 13068 -311
rect 13010 -351 13068 -345
rect 13128 -311 13186 -305
rect 13128 -345 13140 -311
rect 13174 -345 13186 -311
rect 13128 -351 13186 -345
rect 13246 -311 13304 -305
rect 13246 -345 13258 -311
rect 13292 -345 13304 -311
rect 13246 -351 13304 -345
rect 13364 -311 13422 -305
rect 13364 -345 13376 -311
rect 13410 -345 13422 -311
rect 13364 -351 13422 -345
rect 13482 -311 13540 -305
rect 13482 -345 13494 -311
rect 13528 -345 13540 -311
rect 13482 -351 13540 -345
rect 13600 -311 13658 -305
rect 13600 -345 13612 -311
rect 13646 -345 13658 -311
rect 13600 -351 13658 -345
rect 13718 -311 13776 -305
rect 13718 -345 13730 -311
rect 13764 -345 13776 -311
rect 13718 -351 13776 -345
rect 13836 -311 13894 -305
rect 13836 -345 13848 -311
rect 13882 -345 13894 -311
rect 13836 -351 13894 -345
rect 13954 -311 14012 -305
rect 13954 -345 13966 -311
rect 14000 -345 14012 -311
rect 13954 -351 14012 -345
rect 14072 -311 14130 -305
rect 14072 -345 14084 -311
rect 14118 -345 14130 -311
rect 14072 -351 14130 -345
rect 14190 -311 14248 -305
rect 14190 -345 14202 -311
rect 14236 -345 14248 -311
rect 14190 -351 14248 -345
rect 14308 -311 14366 -305
rect 14308 -345 14320 -311
rect 14354 -345 14366 -311
rect 14308 -351 14366 -345
rect 14426 -311 14484 -305
rect 14426 -345 14438 -311
rect 14472 -345 14484 -311
rect 14426 -351 14484 -345
rect 14544 -311 14602 -305
rect 14544 -345 14556 -311
rect 14590 -345 14602 -311
rect 14544 -351 14602 -345
rect 14662 -311 14720 -305
rect 14662 -345 14674 -311
rect 14708 -345 14720 -311
rect 14662 -351 14720 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -14864 -431 14864 431
string parameters w 3 l 0.3 m 1 nf 250 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
