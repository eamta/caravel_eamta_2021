magic
tech sky130A
timestamp 1616200722
<< nwell >>
rect 2351 1361 2512 1363
rect 2265 1351 2512 1361
rect 2265 1148 2669 1351
rect 2265 1041 3811 1148
rect 2332 1039 3811 1041
rect 2350 1037 2356 1039
rect 4495 395 4765 1360
rect 4523 390 4765 395
rect 4583 336 4765 390
rect 4585 -80 4765 336
rect 2324 -409 2470 -88
rect 4585 -179 4790 -80
rect 4599 -182 4790 -179
<< pwell >>
rect 65 455 1102 567
rect -147 -3 1133 455
rect 2024 106 2146 319
rect -144 -465 33 -3
rect -144 -585 941 -465
rect -144 -1441 1088 -585
rect 2454 -1071 3486 -876
rect 1933 -1134 3486 -1071
rect 1933 -1246 3560 -1134
rect 1273 -1327 3560 -1246
rect 1273 -1385 1959 -1327
rect 2349 -1449 3560 -1327
<< poly >>
rect 2206 226 2349 285
rect 2325 -1172 2349 226
rect 2758 -1172 2953 -1084
rect 3525 -1172 3606 -1169
rect 2195 -1230 3606 -1172
rect 3523 -1240 3606 -1230
rect 3523 -1278 3543 -1240
rect 3583 -1278 3606 -1240
rect 3523 -1303 3606 -1278
rect 3525 -1304 3606 -1303
<< polycont >>
rect 3543 -1278 3583 -1240
<< locali >>
rect 3522 -1222 3603 -1221
rect 3522 -1290 3530 -1222
rect 3596 -1290 3603 -1222
<< viali >>
rect 3530 -1240 3596 -1222
rect 3530 -1278 3543 -1240
rect 3543 -1278 3583 -1240
rect 3583 -1278 3596 -1240
rect 3530 -1294 3596 -1278
<< metal1 >>
rect 4187 1360 4529 1363
rect 4187 1030 4768 1360
rect 21 472 48 1022
rect 1983 759 2025 859
rect 4120 762 4162 857
rect 4482 831 4767 1030
rect 313 472 318 474
rect 21 419 318 472
rect 313 377 318 419
rect 416 377 421 474
rect 2097 330 2235 380
rect 4239 330 4372 380
rect 2379 231 2384 306
rect 2447 231 2452 306
rect -4 63 546 65
rect -4 23 511 63
rect -4 -442 24 23
rect 506 22 511 23
rect 548 22 553 63
rect 513 -19 545 22
rect -4 -447 23 -442
rect -4 -453 74 -447
rect 76 -532 81 -416
rect 2393 -449 2423 231
rect -144 -753 329 -639
rect 1976 -688 2022 -593
rect 4378 -686 4419 -593
rect -144 -758 381 -753
rect -144 -1441 709 -758
rect 2094 -1122 2231 -1072
rect 4488 -1120 4627 -1069
rect 3523 -1222 3603 -1209
rect 3523 -1294 3530 -1222
rect 3596 -1294 3603 -1222
rect 3523 -1303 3603 -1294
<< via1 >>
rect 318 377 416 474
rect 2384 231 2447 306
rect 511 22 548 63
rect 3530 -1294 3596 -1222
<< metal2 >>
rect 329 1387 395 1490
rect 359 1023 379 1387
rect 1022 1363 2360 1364
rect 3150 1363 3195 1366
rect 1022 1330 3197 1363
rect 224 983 601 1023
rect 318 474 416 479
rect 1023 441 1045 1330
rect 2418 1021 2442 1024
rect 2418 993 2733 1021
rect 318 372 416 377
rect 348 -32 385 372
rect 2418 311 2442 993
rect 3150 511 3195 1330
rect 2384 306 2447 311
rect 2384 226 2447 231
rect 3143 173 3195 511
rect 4318 217 4769 295
rect 3143 116 3451 173
rect 511 63 548 68
rect 511 -23 548 22
rect 348 -38 384 -32
rect 349 -60 384 -38
rect 511 -59 2778 -23
rect 850 -999 1065 -930
rect 3414 -939 3451 116
rect 4692 -80 4767 217
rect 1007 -1397 1049 -999
rect 3398 -1397 3460 -939
rect 4692 -1135 4768 -80
rect 4692 -1158 4770 -1135
rect 3550 -1211 3587 -1209
rect 3530 -1217 3587 -1211
rect 3530 -1222 3596 -1217
rect 4578 -1229 4770 -1158
rect 3530 -1310 3596 -1294
rect 3530 -1359 3587 -1310
rect 1007 -1422 3460 -1397
rect 3398 -1423 3460 -1422
rect 3533 -1382 3586 -1359
rect 4692 -1382 4770 -1229
rect 3533 -1451 4770 -1382
rect 4692 -1454 4770 -1451
use part  part_0
timestamp 1616191796
transform 1 0 1592 0 1 151
box 877 -149 2935 1213
use counter1b  counter1b_0
timestamp 1616191617
transform 1 0 -545 0 1 149
box 545 -149 2935 1281
use counter1b  counter1b_1
timestamp 1616191617
transform 1 0 -548 0 1 -1300
box 545 -149 2935 1281
use counter1b  counter1b_3
timestamp 1616191617
transform 1 0 1849 0 1 -1300
box 545 -149 2935 1281
<< labels >>
rlabel pwell 2800 -1197 2912 -1101 1 CLR
rlabel metal1 4527 -1108 4571 -1078 1 Qb2
rlabel metal1 4383 -679 4411 -661 1 Q2
rlabel metal1 2123 -1107 2173 -1086 1 Qb1
rlabel metal1 2118 338 2183 369 1 Qb0
rlabel metal1 1989 769 2015 790 1 Q0
rlabel metal1 -8 -1312 267 -1063 1 VSS
rlabel metal2 850 -999 939 -935 1 CLK
rlabel metal1 1983 -680 2019 -658 1 Q1
rlabel metal2 348 1440 386 1473 1 CE
rlabel metal1 4256 1152 4472 1266 1 vdd
rlabel metal1 4126 770 4152 795 1 Q3
rlabel metal1 4255 340 4310 368 1 Qb3
<< end >>
