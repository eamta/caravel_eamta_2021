magic
tech sky130A
magscale 1 2
timestamp 1615910487
<< pwell >>
rect -1949 -2342 1949 2342
<< nmos >>
rect -1753 794 -1613 2194
rect -1555 794 -1415 2194
rect -1357 794 -1217 2194
rect -1159 794 -1019 2194
rect -961 794 -821 2194
rect -763 794 -623 2194
rect -565 794 -425 2194
rect -367 794 -227 2194
rect -169 794 -29 2194
rect 29 794 169 2194
rect 227 794 367 2194
rect 425 794 565 2194
rect 623 794 763 2194
rect 821 794 961 2194
rect 1019 794 1159 2194
rect 1217 794 1357 2194
rect 1415 794 1555 2194
rect 1613 794 1753 2194
rect -1753 -700 -1613 700
rect -1555 -700 -1415 700
rect -1357 -700 -1217 700
rect -1159 -700 -1019 700
rect -961 -700 -821 700
rect -763 -700 -623 700
rect -565 -700 -425 700
rect -367 -700 -227 700
rect -169 -700 -29 700
rect 29 -700 169 700
rect 227 -700 367 700
rect 425 -700 565 700
rect 623 -700 763 700
rect 821 -700 961 700
rect 1019 -700 1159 700
rect 1217 -700 1357 700
rect 1415 -700 1555 700
rect 1613 -700 1753 700
rect -1753 -2194 -1613 -794
rect -1555 -2194 -1415 -794
rect -1357 -2194 -1217 -794
rect -1159 -2194 -1019 -794
rect -961 -2194 -821 -794
rect -763 -2194 -623 -794
rect -565 -2194 -425 -794
rect -367 -2194 -227 -794
rect -169 -2194 -29 -794
rect 29 -2194 169 -794
rect 227 -2194 367 -794
rect 425 -2194 565 -794
rect 623 -2194 763 -794
rect 821 -2194 961 -794
rect 1019 -2194 1159 -794
rect 1217 -2194 1357 -794
rect 1415 -2194 1555 -794
rect 1613 -2194 1753 -794
<< ndiff >>
rect -1811 2182 -1753 2194
rect -1811 806 -1799 2182
rect -1765 806 -1753 2182
rect -1811 794 -1753 806
rect -1613 2182 -1555 2194
rect -1613 806 -1601 2182
rect -1567 806 -1555 2182
rect -1613 794 -1555 806
rect -1415 2182 -1357 2194
rect -1415 806 -1403 2182
rect -1369 806 -1357 2182
rect -1415 794 -1357 806
rect -1217 2182 -1159 2194
rect -1217 806 -1205 2182
rect -1171 806 -1159 2182
rect -1217 794 -1159 806
rect -1019 2182 -961 2194
rect -1019 806 -1007 2182
rect -973 806 -961 2182
rect -1019 794 -961 806
rect -821 2182 -763 2194
rect -821 806 -809 2182
rect -775 806 -763 2182
rect -821 794 -763 806
rect -623 2182 -565 2194
rect -623 806 -611 2182
rect -577 806 -565 2182
rect -623 794 -565 806
rect -425 2182 -367 2194
rect -425 806 -413 2182
rect -379 806 -367 2182
rect -425 794 -367 806
rect -227 2182 -169 2194
rect -227 806 -215 2182
rect -181 806 -169 2182
rect -227 794 -169 806
rect -29 2182 29 2194
rect -29 806 -17 2182
rect 17 806 29 2182
rect -29 794 29 806
rect 169 2182 227 2194
rect 169 806 181 2182
rect 215 806 227 2182
rect 169 794 227 806
rect 367 2182 425 2194
rect 367 806 379 2182
rect 413 806 425 2182
rect 367 794 425 806
rect 565 2182 623 2194
rect 565 806 577 2182
rect 611 806 623 2182
rect 565 794 623 806
rect 763 2182 821 2194
rect 763 806 775 2182
rect 809 806 821 2182
rect 763 794 821 806
rect 961 2182 1019 2194
rect 961 806 973 2182
rect 1007 806 1019 2182
rect 961 794 1019 806
rect 1159 2182 1217 2194
rect 1159 806 1171 2182
rect 1205 806 1217 2182
rect 1159 794 1217 806
rect 1357 2182 1415 2194
rect 1357 806 1369 2182
rect 1403 806 1415 2182
rect 1357 794 1415 806
rect 1555 2182 1613 2194
rect 1555 806 1567 2182
rect 1601 806 1613 2182
rect 1555 794 1613 806
rect 1753 2182 1811 2194
rect 1753 806 1765 2182
rect 1799 806 1811 2182
rect 1753 794 1811 806
rect -1811 688 -1753 700
rect -1811 -688 -1799 688
rect -1765 -688 -1753 688
rect -1811 -700 -1753 -688
rect -1613 688 -1555 700
rect -1613 -688 -1601 688
rect -1567 -688 -1555 688
rect -1613 -700 -1555 -688
rect -1415 688 -1357 700
rect -1415 -688 -1403 688
rect -1369 -688 -1357 688
rect -1415 -700 -1357 -688
rect -1217 688 -1159 700
rect -1217 -688 -1205 688
rect -1171 -688 -1159 688
rect -1217 -700 -1159 -688
rect -1019 688 -961 700
rect -1019 -688 -1007 688
rect -973 -688 -961 688
rect -1019 -700 -961 -688
rect -821 688 -763 700
rect -821 -688 -809 688
rect -775 -688 -763 688
rect -821 -700 -763 -688
rect -623 688 -565 700
rect -623 -688 -611 688
rect -577 -688 -565 688
rect -623 -700 -565 -688
rect -425 688 -367 700
rect -425 -688 -413 688
rect -379 -688 -367 688
rect -425 -700 -367 -688
rect -227 688 -169 700
rect -227 -688 -215 688
rect -181 -688 -169 688
rect -227 -700 -169 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 169 688 227 700
rect 169 -688 181 688
rect 215 -688 227 688
rect 169 -700 227 -688
rect 367 688 425 700
rect 367 -688 379 688
rect 413 -688 425 688
rect 367 -700 425 -688
rect 565 688 623 700
rect 565 -688 577 688
rect 611 -688 623 688
rect 565 -700 623 -688
rect 763 688 821 700
rect 763 -688 775 688
rect 809 -688 821 688
rect 763 -700 821 -688
rect 961 688 1019 700
rect 961 -688 973 688
rect 1007 -688 1019 688
rect 961 -700 1019 -688
rect 1159 688 1217 700
rect 1159 -688 1171 688
rect 1205 -688 1217 688
rect 1159 -700 1217 -688
rect 1357 688 1415 700
rect 1357 -688 1369 688
rect 1403 -688 1415 688
rect 1357 -700 1415 -688
rect 1555 688 1613 700
rect 1555 -688 1567 688
rect 1601 -688 1613 688
rect 1555 -700 1613 -688
rect 1753 688 1811 700
rect 1753 -688 1765 688
rect 1799 -688 1811 688
rect 1753 -700 1811 -688
rect -1811 -806 -1753 -794
rect -1811 -2182 -1799 -806
rect -1765 -2182 -1753 -806
rect -1811 -2194 -1753 -2182
rect -1613 -806 -1555 -794
rect -1613 -2182 -1601 -806
rect -1567 -2182 -1555 -806
rect -1613 -2194 -1555 -2182
rect -1415 -806 -1357 -794
rect -1415 -2182 -1403 -806
rect -1369 -2182 -1357 -806
rect -1415 -2194 -1357 -2182
rect -1217 -806 -1159 -794
rect -1217 -2182 -1205 -806
rect -1171 -2182 -1159 -806
rect -1217 -2194 -1159 -2182
rect -1019 -806 -961 -794
rect -1019 -2182 -1007 -806
rect -973 -2182 -961 -806
rect -1019 -2194 -961 -2182
rect -821 -806 -763 -794
rect -821 -2182 -809 -806
rect -775 -2182 -763 -806
rect -821 -2194 -763 -2182
rect -623 -806 -565 -794
rect -623 -2182 -611 -806
rect -577 -2182 -565 -806
rect -623 -2194 -565 -2182
rect -425 -806 -367 -794
rect -425 -2182 -413 -806
rect -379 -2182 -367 -806
rect -425 -2194 -367 -2182
rect -227 -806 -169 -794
rect -227 -2182 -215 -806
rect -181 -2182 -169 -806
rect -227 -2194 -169 -2182
rect -29 -806 29 -794
rect -29 -2182 -17 -806
rect 17 -2182 29 -806
rect -29 -2194 29 -2182
rect 169 -806 227 -794
rect 169 -2182 181 -806
rect 215 -2182 227 -806
rect 169 -2194 227 -2182
rect 367 -806 425 -794
rect 367 -2182 379 -806
rect 413 -2182 425 -806
rect 367 -2194 425 -2182
rect 565 -806 623 -794
rect 565 -2182 577 -806
rect 611 -2182 623 -806
rect 565 -2194 623 -2182
rect 763 -806 821 -794
rect 763 -2182 775 -806
rect 809 -2182 821 -806
rect 763 -2194 821 -2182
rect 961 -806 1019 -794
rect 961 -2182 973 -806
rect 1007 -2182 1019 -806
rect 961 -2194 1019 -2182
rect 1159 -806 1217 -794
rect 1159 -2182 1171 -806
rect 1205 -2182 1217 -806
rect 1159 -2194 1217 -2182
rect 1357 -806 1415 -794
rect 1357 -2182 1369 -806
rect 1403 -2182 1415 -806
rect 1357 -2194 1415 -2182
rect 1555 -806 1613 -794
rect 1555 -2182 1567 -806
rect 1601 -2182 1613 -806
rect 1555 -2194 1613 -2182
rect 1753 -806 1811 -794
rect 1753 -2182 1765 -806
rect 1799 -2182 1811 -806
rect 1753 -2194 1811 -2182
<< ndiffc >>
rect -1799 806 -1765 2182
rect -1601 806 -1567 2182
rect -1403 806 -1369 2182
rect -1205 806 -1171 2182
rect -1007 806 -973 2182
rect -809 806 -775 2182
rect -611 806 -577 2182
rect -413 806 -379 2182
rect -215 806 -181 2182
rect -17 806 17 2182
rect 181 806 215 2182
rect 379 806 413 2182
rect 577 806 611 2182
rect 775 806 809 2182
rect 973 806 1007 2182
rect 1171 806 1205 2182
rect 1369 806 1403 2182
rect 1567 806 1601 2182
rect 1765 806 1799 2182
rect -1799 -688 -1765 688
rect -1601 -688 -1567 688
rect -1403 -688 -1369 688
rect -1205 -688 -1171 688
rect -1007 -688 -973 688
rect -809 -688 -775 688
rect -611 -688 -577 688
rect -413 -688 -379 688
rect -215 -688 -181 688
rect -17 -688 17 688
rect 181 -688 215 688
rect 379 -688 413 688
rect 577 -688 611 688
rect 775 -688 809 688
rect 973 -688 1007 688
rect 1171 -688 1205 688
rect 1369 -688 1403 688
rect 1567 -688 1601 688
rect 1765 -688 1799 688
rect -1799 -2182 -1765 -806
rect -1601 -2182 -1567 -806
rect -1403 -2182 -1369 -806
rect -1205 -2182 -1171 -806
rect -1007 -2182 -973 -806
rect -809 -2182 -775 -806
rect -611 -2182 -577 -806
rect -413 -2182 -379 -806
rect -215 -2182 -181 -806
rect -17 -2182 17 -806
rect 181 -2182 215 -806
rect 379 -2182 413 -806
rect 577 -2182 611 -806
rect 775 -2182 809 -806
rect 973 -2182 1007 -806
rect 1171 -2182 1205 -806
rect 1369 -2182 1403 -806
rect 1567 -2182 1601 -806
rect 1765 -2182 1799 -806
<< psubdiff >>
rect -1913 2272 -1817 2306
rect 1817 2272 1913 2306
rect -1913 2210 -1879 2272
rect 1879 2210 1913 2272
rect -1913 -2272 -1879 -2210
rect 1879 -2272 1913 -2210
rect -1913 -2306 -1817 -2272
rect 1817 -2306 1913 -2272
<< psubdiffcont >>
rect -1817 2272 1817 2306
rect -1913 -2210 -1879 2210
rect 1879 -2210 1913 2210
rect -1817 -2306 1817 -2272
<< poly >>
rect -1753 2194 -1613 2220
rect -1555 2194 -1415 2220
rect -1357 2194 -1217 2220
rect -1159 2194 -1019 2220
rect -961 2194 -821 2220
rect -763 2194 -623 2220
rect -565 2194 -425 2220
rect -367 2194 -227 2220
rect -169 2194 -29 2220
rect 29 2194 169 2220
rect 227 2194 367 2220
rect 425 2194 565 2220
rect 623 2194 763 2220
rect 821 2194 961 2220
rect 1019 2194 1159 2220
rect 1217 2194 1357 2220
rect 1415 2194 1555 2220
rect 1613 2194 1753 2220
rect -1753 768 -1613 794
rect -1555 768 -1415 794
rect -1357 768 -1217 794
rect -1159 768 -1019 794
rect -961 768 -821 794
rect -763 768 -623 794
rect -565 768 -425 794
rect -367 768 -227 794
rect -169 768 -29 794
rect 29 768 169 794
rect 227 768 367 794
rect 425 768 565 794
rect 623 768 763 794
rect 821 768 961 794
rect 1019 768 1159 794
rect 1217 768 1357 794
rect 1415 768 1555 794
rect 1613 768 1753 794
rect -1753 700 -1613 726
rect -1555 700 -1415 726
rect -1357 700 -1217 726
rect -1159 700 -1019 726
rect -961 700 -821 726
rect -763 700 -623 726
rect -565 700 -425 726
rect -367 700 -227 726
rect -169 700 -29 726
rect 29 700 169 726
rect 227 700 367 726
rect 425 700 565 726
rect 623 700 763 726
rect 821 700 961 726
rect 1019 700 1159 726
rect 1217 700 1357 726
rect 1415 700 1555 726
rect 1613 700 1753 726
rect -1753 -726 -1613 -700
rect -1555 -726 -1415 -700
rect -1357 -726 -1217 -700
rect -1159 -726 -1019 -700
rect -961 -726 -821 -700
rect -763 -726 -623 -700
rect -565 -726 -425 -700
rect -367 -726 -227 -700
rect -169 -726 -29 -700
rect 29 -726 169 -700
rect 227 -726 367 -700
rect 425 -726 565 -700
rect 623 -726 763 -700
rect 821 -726 961 -700
rect 1019 -726 1159 -700
rect 1217 -726 1357 -700
rect 1415 -726 1555 -700
rect 1613 -726 1753 -700
rect -1753 -794 -1613 -768
rect -1555 -794 -1415 -768
rect -1357 -794 -1217 -768
rect -1159 -794 -1019 -768
rect -961 -794 -821 -768
rect -763 -794 -623 -768
rect -565 -794 -425 -768
rect -367 -794 -227 -768
rect -169 -794 -29 -768
rect 29 -794 169 -768
rect 227 -794 367 -768
rect 425 -794 565 -768
rect 623 -794 763 -768
rect 821 -794 961 -768
rect 1019 -794 1159 -768
rect 1217 -794 1357 -768
rect 1415 -794 1555 -768
rect 1613 -794 1753 -768
rect -1753 -2220 -1613 -2194
rect -1555 -2220 -1415 -2194
rect -1357 -2220 -1217 -2194
rect -1159 -2220 -1019 -2194
rect -961 -2220 -821 -2194
rect -763 -2220 -623 -2194
rect -565 -2220 -425 -2194
rect -367 -2220 -227 -2194
rect -169 -2220 -29 -2194
rect 29 -2220 169 -2194
rect 227 -2220 367 -2194
rect 425 -2220 565 -2194
rect 623 -2220 763 -2194
rect 821 -2220 961 -2194
rect 1019 -2220 1159 -2194
rect 1217 -2220 1357 -2194
rect 1415 -2220 1555 -2194
rect 1613 -2220 1753 -2194
<< locali >>
rect -1913 2272 -1817 2306
rect 1817 2272 1913 2306
rect -1913 2210 -1879 2272
rect 1879 2210 1913 2272
rect -1799 2182 -1765 2198
rect -1799 790 -1765 806
rect -1601 2182 -1567 2198
rect -1601 790 -1567 806
rect -1403 2182 -1369 2198
rect -1403 790 -1369 806
rect -1205 2182 -1171 2198
rect -1205 790 -1171 806
rect -1007 2182 -973 2198
rect -1007 790 -973 806
rect -809 2182 -775 2198
rect -809 790 -775 806
rect -611 2182 -577 2198
rect -611 790 -577 806
rect -413 2182 -379 2198
rect -413 790 -379 806
rect -215 2182 -181 2198
rect -215 790 -181 806
rect -17 2182 17 2198
rect -17 790 17 806
rect 181 2182 215 2198
rect 181 790 215 806
rect 379 2182 413 2198
rect 379 790 413 806
rect 577 2182 611 2198
rect 577 790 611 806
rect 775 2182 809 2198
rect 775 790 809 806
rect 973 2182 1007 2198
rect 973 790 1007 806
rect 1171 2182 1205 2198
rect 1171 790 1205 806
rect 1369 2182 1403 2198
rect 1369 790 1403 806
rect 1567 2182 1601 2198
rect 1567 790 1601 806
rect 1765 2182 1799 2198
rect 1765 790 1799 806
rect -1799 688 -1765 704
rect -1799 -704 -1765 -688
rect -1601 688 -1567 704
rect -1601 -704 -1567 -688
rect -1403 688 -1369 704
rect -1403 -704 -1369 -688
rect -1205 688 -1171 704
rect -1205 -704 -1171 -688
rect -1007 688 -973 704
rect -1007 -704 -973 -688
rect -809 688 -775 704
rect -809 -704 -775 -688
rect -611 688 -577 704
rect -611 -704 -577 -688
rect -413 688 -379 704
rect -413 -704 -379 -688
rect -215 688 -181 704
rect -215 -704 -181 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 181 688 215 704
rect 181 -704 215 -688
rect 379 688 413 704
rect 379 -704 413 -688
rect 577 688 611 704
rect 577 -704 611 -688
rect 775 688 809 704
rect 775 -704 809 -688
rect 973 688 1007 704
rect 973 -704 1007 -688
rect 1171 688 1205 704
rect 1171 -704 1205 -688
rect 1369 688 1403 704
rect 1369 -704 1403 -688
rect 1567 688 1601 704
rect 1567 -704 1601 -688
rect 1765 688 1799 704
rect 1765 -704 1799 -688
rect -1799 -806 -1765 -790
rect -1799 -2198 -1765 -2182
rect -1601 -806 -1567 -790
rect -1601 -2198 -1567 -2182
rect -1403 -806 -1369 -790
rect -1403 -2198 -1369 -2182
rect -1205 -806 -1171 -790
rect -1205 -2198 -1171 -2182
rect -1007 -806 -973 -790
rect -1007 -2198 -973 -2182
rect -809 -806 -775 -790
rect -809 -2198 -775 -2182
rect -611 -806 -577 -790
rect -611 -2198 -577 -2182
rect -413 -806 -379 -790
rect -413 -2198 -379 -2182
rect -215 -806 -181 -790
rect -215 -2198 -181 -2182
rect -17 -806 17 -790
rect -17 -2198 17 -2182
rect 181 -806 215 -790
rect 181 -2198 215 -2182
rect 379 -806 413 -790
rect 379 -2198 413 -2182
rect 577 -806 611 -790
rect 577 -2198 611 -2182
rect 775 -806 809 -790
rect 775 -2198 809 -2182
rect 973 -806 1007 -790
rect 973 -2198 1007 -2182
rect 1171 -806 1205 -790
rect 1171 -2198 1205 -2182
rect 1369 -806 1403 -790
rect 1369 -2198 1403 -2182
rect 1567 -806 1601 -790
rect 1567 -2198 1601 -2182
rect 1765 -806 1799 -790
rect 1765 -2198 1799 -2182
rect -1913 -2272 -1879 -2210
rect 1879 -2272 1913 -2210
rect -1913 -2306 -1817 -2272
rect 1817 -2306 1913 -2272
<< viali >>
rect -1799 806 -1765 2182
rect -1601 806 -1567 2182
rect -1403 806 -1369 2182
rect -1205 806 -1171 2182
rect -1007 806 -973 2182
rect -809 806 -775 2182
rect -611 806 -577 2182
rect -413 806 -379 2182
rect -215 806 -181 2182
rect -17 806 17 2182
rect 181 806 215 2182
rect 379 806 413 2182
rect 577 806 611 2182
rect 775 806 809 2182
rect 973 806 1007 2182
rect 1171 806 1205 2182
rect 1369 806 1403 2182
rect 1567 806 1601 2182
rect 1765 806 1799 2182
rect -1799 -688 -1765 688
rect -1601 -688 -1567 688
rect -1403 -688 -1369 688
rect -1205 -688 -1171 688
rect -1007 -688 -973 688
rect -809 -688 -775 688
rect -611 -688 -577 688
rect -413 -688 -379 688
rect -215 -688 -181 688
rect -17 -688 17 688
rect 181 -688 215 688
rect 379 -688 413 688
rect 577 -688 611 688
rect 775 -688 809 688
rect 973 -688 1007 688
rect 1171 -688 1205 688
rect 1369 -688 1403 688
rect 1567 -688 1601 688
rect 1765 -688 1799 688
rect -1799 -2182 -1765 -806
rect -1601 -2182 -1567 -806
rect -1403 -2182 -1369 -806
rect -1205 -2182 -1171 -806
rect -1007 -2182 -973 -806
rect -809 -2182 -775 -806
rect -611 -2182 -577 -806
rect -413 -2182 -379 -806
rect -215 -2182 -181 -806
rect -17 -2182 17 -806
rect 181 -2182 215 -806
rect 379 -2182 413 -806
rect 577 -2182 611 -806
rect 775 -2182 809 -806
rect 973 -2182 1007 -806
rect 1171 -2182 1205 -806
rect 1369 -2182 1403 -806
rect 1567 -2182 1601 -806
rect 1765 -2182 1799 -806
<< metal1 >>
rect -1805 2182 -1759 2194
rect -1805 806 -1799 2182
rect -1765 806 -1759 2182
rect -1805 794 -1759 806
rect -1607 2182 -1561 2194
rect -1607 806 -1601 2182
rect -1567 806 -1561 2182
rect -1607 794 -1561 806
rect -1409 2182 -1363 2194
rect -1409 806 -1403 2182
rect -1369 806 -1363 2182
rect -1409 794 -1363 806
rect -1211 2182 -1165 2194
rect -1211 806 -1205 2182
rect -1171 806 -1165 2182
rect -1211 794 -1165 806
rect -1013 2182 -967 2194
rect -1013 806 -1007 2182
rect -973 806 -967 2182
rect -1013 794 -967 806
rect -815 2182 -769 2194
rect -815 806 -809 2182
rect -775 806 -769 2182
rect -815 794 -769 806
rect -617 2182 -571 2194
rect -617 806 -611 2182
rect -577 806 -571 2182
rect -617 794 -571 806
rect -419 2182 -373 2194
rect -419 806 -413 2182
rect -379 806 -373 2182
rect -419 794 -373 806
rect -221 2182 -175 2194
rect -221 806 -215 2182
rect -181 806 -175 2182
rect -221 794 -175 806
rect -23 2182 23 2194
rect -23 806 -17 2182
rect 17 806 23 2182
rect -23 794 23 806
rect 175 2182 221 2194
rect 175 806 181 2182
rect 215 806 221 2182
rect 175 794 221 806
rect 373 2182 419 2194
rect 373 806 379 2182
rect 413 806 419 2182
rect 373 794 419 806
rect 571 2182 617 2194
rect 571 806 577 2182
rect 611 806 617 2182
rect 571 794 617 806
rect 769 2182 815 2194
rect 769 806 775 2182
rect 809 806 815 2182
rect 769 794 815 806
rect 967 2182 1013 2194
rect 967 806 973 2182
rect 1007 806 1013 2182
rect 967 794 1013 806
rect 1165 2182 1211 2194
rect 1165 806 1171 2182
rect 1205 806 1211 2182
rect 1165 794 1211 806
rect 1363 2182 1409 2194
rect 1363 806 1369 2182
rect 1403 806 1409 2182
rect 1363 794 1409 806
rect 1561 2182 1607 2194
rect 1561 806 1567 2182
rect 1601 806 1607 2182
rect 1561 794 1607 806
rect 1759 2182 1805 2194
rect 1759 806 1765 2182
rect 1799 806 1805 2182
rect 1759 794 1805 806
rect -1805 688 -1759 700
rect -1805 -688 -1799 688
rect -1765 -688 -1759 688
rect -1805 -700 -1759 -688
rect -1607 688 -1561 700
rect -1607 -688 -1601 688
rect -1567 -688 -1561 688
rect -1607 -700 -1561 -688
rect -1409 688 -1363 700
rect -1409 -688 -1403 688
rect -1369 -688 -1363 688
rect -1409 -700 -1363 -688
rect -1211 688 -1165 700
rect -1211 -688 -1205 688
rect -1171 -688 -1165 688
rect -1211 -700 -1165 -688
rect -1013 688 -967 700
rect -1013 -688 -1007 688
rect -973 -688 -967 688
rect -1013 -700 -967 -688
rect -815 688 -769 700
rect -815 -688 -809 688
rect -775 -688 -769 688
rect -815 -700 -769 -688
rect -617 688 -571 700
rect -617 -688 -611 688
rect -577 -688 -571 688
rect -617 -700 -571 -688
rect -419 688 -373 700
rect -419 -688 -413 688
rect -379 -688 -373 688
rect -419 -700 -373 -688
rect -221 688 -175 700
rect -221 -688 -215 688
rect -181 -688 -175 688
rect -221 -700 -175 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 175 688 221 700
rect 175 -688 181 688
rect 215 -688 221 688
rect 175 -700 221 -688
rect 373 688 419 700
rect 373 -688 379 688
rect 413 -688 419 688
rect 373 -700 419 -688
rect 571 688 617 700
rect 571 -688 577 688
rect 611 -688 617 688
rect 571 -700 617 -688
rect 769 688 815 700
rect 769 -688 775 688
rect 809 -688 815 688
rect 769 -700 815 -688
rect 967 688 1013 700
rect 967 -688 973 688
rect 1007 -688 1013 688
rect 967 -700 1013 -688
rect 1165 688 1211 700
rect 1165 -688 1171 688
rect 1205 -688 1211 688
rect 1165 -700 1211 -688
rect 1363 688 1409 700
rect 1363 -688 1369 688
rect 1403 -688 1409 688
rect 1363 -700 1409 -688
rect 1561 688 1607 700
rect 1561 -688 1567 688
rect 1601 -688 1607 688
rect 1561 -700 1607 -688
rect 1759 688 1805 700
rect 1759 -688 1765 688
rect 1799 -688 1805 688
rect 1759 -700 1805 -688
rect -1805 -806 -1759 -794
rect -1805 -2182 -1799 -806
rect -1765 -2182 -1759 -806
rect -1805 -2194 -1759 -2182
rect -1607 -806 -1561 -794
rect -1607 -2182 -1601 -806
rect -1567 -2182 -1561 -806
rect -1607 -2194 -1561 -2182
rect -1409 -806 -1363 -794
rect -1409 -2182 -1403 -806
rect -1369 -2182 -1363 -806
rect -1409 -2194 -1363 -2182
rect -1211 -806 -1165 -794
rect -1211 -2182 -1205 -806
rect -1171 -2182 -1165 -806
rect -1211 -2194 -1165 -2182
rect -1013 -806 -967 -794
rect -1013 -2182 -1007 -806
rect -973 -2182 -967 -806
rect -1013 -2194 -967 -2182
rect -815 -806 -769 -794
rect -815 -2182 -809 -806
rect -775 -2182 -769 -806
rect -815 -2194 -769 -2182
rect -617 -806 -571 -794
rect -617 -2182 -611 -806
rect -577 -2182 -571 -806
rect -617 -2194 -571 -2182
rect -419 -806 -373 -794
rect -419 -2182 -413 -806
rect -379 -2182 -373 -806
rect -419 -2194 -373 -2182
rect -221 -806 -175 -794
rect -221 -2182 -215 -806
rect -181 -2182 -175 -806
rect -221 -2194 -175 -2182
rect -23 -806 23 -794
rect -23 -2182 -17 -806
rect 17 -2182 23 -806
rect -23 -2194 23 -2182
rect 175 -806 221 -794
rect 175 -2182 181 -806
rect 215 -2182 221 -806
rect 175 -2194 221 -2182
rect 373 -806 419 -794
rect 373 -2182 379 -806
rect 413 -2182 419 -806
rect 373 -2194 419 -2182
rect 571 -806 617 -794
rect 571 -2182 577 -806
rect 611 -2182 617 -806
rect 571 -2194 617 -2182
rect 769 -806 815 -794
rect 769 -2182 775 -806
rect 809 -2182 815 -806
rect 769 -2194 815 -2182
rect 967 -806 1013 -794
rect 967 -2182 973 -806
rect 1007 -2182 1013 -806
rect 967 -2194 1013 -2182
rect 1165 -806 1211 -794
rect 1165 -2182 1171 -806
rect 1205 -2182 1211 -806
rect 1165 -2194 1211 -2182
rect 1363 -806 1409 -794
rect 1363 -2182 1369 -806
rect 1403 -2182 1409 -806
rect 1363 -2194 1409 -2182
rect 1561 -806 1607 -794
rect 1561 -2182 1567 -806
rect 1601 -2182 1607 -806
rect 1561 -2194 1607 -2182
rect 1759 -806 1805 -794
rect 1759 -2182 1765 -806
rect 1799 -2182 1805 -806
rect 1759 -2194 1805 -2182
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1896 -2289 1896 2289
string parameters w 7 l 0.7 m 3 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
