magic
tech sky130A
magscale 1 2
timestamp 1623247083
<< error_p >>
rect -845 1572 -787 1578
rect -653 1572 -595 1578
rect -461 1572 -403 1578
rect -269 1572 -211 1578
rect -77 1572 -19 1578
rect 115 1572 173 1578
rect 307 1572 365 1578
rect 499 1572 557 1578
rect 691 1572 749 1578
rect 883 1572 941 1578
rect -845 1538 -833 1572
rect -653 1538 -641 1572
rect -461 1538 -449 1572
rect -269 1538 -257 1572
rect -77 1538 -65 1572
rect 115 1538 127 1572
rect 307 1538 319 1572
rect 499 1538 511 1572
rect 691 1538 703 1572
rect 883 1538 895 1572
rect -845 1532 -787 1538
rect -653 1532 -595 1538
rect -461 1532 -403 1538
rect -269 1532 -211 1538
rect -77 1532 -19 1538
rect 115 1532 173 1538
rect 307 1532 365 1538
rect 499 1532 557 1538
rect 691 1532 749 1538
rect 883 1532 941 1538
rect -941 -1538 -883 -1532
rect -749 -1538 -691 -1532
rect -557 -1538 -499 -1532
rect -365 -1538 -307 -1532
rect -173 -1538 -115 -1532
rect 19 -1538 77 -1532
rect 211 -1538 269 -1532
rect 403 -1538 461 -1532
rect 595 -1538 653 -1532
rect 787 -1538 845 -1532
rect -941 -1572 -929 -1538
rect -749 -1572 -737 -1538
rect -557 -1572 -545 -1538
rect -365 -1572 -353 -1538
rect -173 -1572 -161 -1538
rect 19 -1572 31 -1538
rect 211 -1572 223 -1538
rect 403 -1572 415 -1538
rect 595 -1572 607 -1538
rect 787 -1572 799 -1538
rect -941 -1578 -883 -1572
rect -749 -1578 -691 -1572
rect -557 -1578 -499 -1572
rect -365 -1578 -307 -1572
rect -173 -1578 -115 -1572
rect 19 -1578 77 -1572
rect 211 -1578 269 -1572
rect 403 -1578 461 -1572
rect 595 -1578 653 -1572
rect 787 -1578 845 -1572
<< pwell >>
rect -1127 -1710 1127 1710
<< nmoslvt >>
rect -927 -1500 -897 1500
rect -831 -1500 -801 1500
rect -735 -1500 -705 1500
rect -639 -1500 -609 1500
rect -543 -1500 -513 1500
rect -447 -1500 -417 1500
rect -351 -1500 -321 1500
rect -255 -1500 -225 1500
rect -159 -1500 -129 1500
rect -63 -1500 -33 1500
rect 33 -1500 63 1500
rect 129 -1500 159 1500
rect 225 -1500 255 1500
rect 321 -1500 351 1500
rect 417 -1500 447 1500
rect 513 -1500 543 1500
rect 609 -1500 639 1500
rect 705 -1500 735 1500
rect 801 -1500 831 1500
rect 897 -1500 927 1500
<< ndiff >>
rect -989 1488 -927 1500
rect -989 -1488 -977 1488
rect -943 -1488 -927 1488
rect -989 -1500 -927 -1488
rect -897 1488 -831 1500
rect -897 -1488 -881 1488
rect -847 -1488 -831 1488
rect -897 -1500 -831 -1488
rect -801 1488 -735 1500
rect -801 -1488 -785 1488
rect -751 -1488 -735 1488
rect -801 -1500 -735 -1488
rect -705 1488 -639 1500
rect -705 -1488 -689 1488
rect -655 -1488 -639 1488
rect -705 -1500 -639 -1488
rect -609 1488 -543 1500
rect -609 -1488 -593 1488
rect -559 -1488 -543 1488
rect -609 -1500 -543 -1488
rect -513 1488 -447 1500
rect -513 -1488 -497 1488
rect -463 -1488 -447 1488
rect -513 -1500 -447 -1488
rect -417 1488 -351 1500
rect -417 -1488 -401 1488
rect -367 -1488 -351 1488
rect -417 -1500 -351 -1488
rect -321 1488 -255 1500
rect -321 -1488 -305 1488
rect -271 -1488 -255 1488
rect -321 -1500 -255 -1488
rect -225 1488 -159 1500
rect -225 -1488 -209 1488
rect -175 -1488 -159 1488
rect -225 -1500 -159 -1488
rect -129 1488 -63 1500
rect -129 -1488 -113 1488
rect -79 -1488 -63 1488
rect -129 -1500 -63 -1488
rect -33 1488 33 1500
rect -33 -1488 -17 1488
rect 17 -1488 33 1488
rect -33 -1500 33 -1488
rect 63 1488 129 1500
rect 63 -1488 79 1488
rect 113 -1488 129 1488
rect 63 -1500 129 -1488
rect 159 1488 225 1500
rect 159 -1488 175 1488
rect 209 -1488 225 1488
rect 159 -1500 225 -1488
rect 255 1488 321 1500
rect 255 -1488 271 1488
rect 305 -1488 321 1488
rect 255 -1500 321 -1488
rect 351 1488 417 1500
rect 351 -1488 367 1488
rect 401 -1488 417 1488
rect 351 -1500 417 -1488
rect 447 1488 513 1500
rect 447 -1488 463 1488
rect 497 -1488 513 1488
rect 447 -1500 513 -1488
rect 543 1488 609 1500
rect 543 -1488 559 1488
rect 593 -1488 609 1488
rect 543 -1500 609 -1488
rect 639 1488 705 1500
rect 639 -1488 655 1488
rect 689 -1488 705 1488
rect 639 -1500 705 -1488
rect 735 1488 801 1500
rect 735 -1488 751 1488
rect 785 -1488 801 1488
rect 735 -1500 801 -1488
rect 831 1488 897 1500
rect 831 -1488 847 1488
rect 881 -1488 897 1488
rect 831 -1500 897 -1488
rect 927 1488 989 1500
rect 927 -1488 943 1488
rect 977 -1488 989 1488
rect 927 -1500 989 -1488
<< ndiffc >>
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
<< psubdiff >>
rect -1091 1640 -995 1674
rect 995 1640 1091 1674
rect -1091 -1640 -1057 1640
rect 1057 1578 1091 1640
rect 1057 -1640 1091 -1578
rect -1091 -1674 1091 -1640
<< psubdiffcont >>
rect -995 1640 995 1674
rect 1057 -1578 1091 1578
<< poly >>
rect -849 1572 -783 1588
rect -849 1538 -833 1572
rect -799 1538 -783 1572
rect -927 1500 -897 1526
rect -849 1522 -783 1538
rect -657 1572 -591 1588
rect -657 1538 -641 1572
rect -607 1538 -591 1572
rect -831 1500 -801 1522
rect -735 1500 -705 1526
rect -657 1522 -591 1538
rect -465 1572 -399 1588
rect -465 1538 -449 1572
rect -415 1538 -399 1572
rect -639 1500 -609 1522
rect -543 1500 -513 1526
rect -465 1522 -399 1538
rect -273 1572 -207 1588
rect -273 1538 -257 1572
rect -223 1538 -207 1572
rect -447 1500 -417 1522
rect -351 1500 -321 1526
rect -273 1522 -207 1538
rect -81 1572 -15 1588
rect -81 1538 -65 1572
rect -31 1538 -15 1572
rect -255 1500 -225 1522
rect -159 1500 -129 1526
rect -81 1522 -15 1538
rect 111 1572 177 1588
rect 111 1538 127 1572
rect 161 1538 177 1572
rect -63 1500 -33 1522
rect 33 1500 63 1526
rect 111 1522 177 1538
rect 303 1572 369 1588
rect 303 1538 319 1572
rect 353 1538 369 1572
rect 129 1500 159 1522
rect 225 1500 255 1526
rect 303 1522 369 1538
rect 495 1572 561 1588
rect 495 1538 511 1572
rect 545 1538 561 1572
rect 321 1500 351 1522
rect 417 1500 447 1526
rect 495 1522 561 1538
rect 687 1572 753 1588
rect 687 1538 703 1572
rect 737 1538 753 1572
rect 513 1500 543 1522
rect 609 1500 639 1526
rect 687 1522 753 1538
rect 879 1572 945 1588
rect 879 1538 895 1572
rect 929 1538 945 1572
rect 705 1500 735 1522
rect 801 1500 831 1526
rect 879 1522 945 1538
rect 897 1500 927 1522
rect -927 -1522 -897 -1500
rect -945 -1538 -879 -1522
rect -831 -1526 -801 -1500
rect -735 -1522 -705 -1500
rect -945 -1572 -929 -1538
rect -895 -1572 -879 -1538
rect -945 -1588 -879 -1572
rect -753 -1538 -687 -1522
rect -639 -1526 -609 -1500
rect -543 -1522 -513 -1500
rect -753 -1572 -737 -1538
rect -703 -1572 -687 -1538
rect -753 -1588 -687 -1572
rect -561 -1538 -495 -1522
rect -447 -1526 -417 -1500
rect -351 -1522 -321 -1500
rect -561 -1572 -545 -1538
rect -511 -1572 -495 -1538
rect -561 -1588 -495 -1572
rect -369 -1538 -303 -1522
rect -255 -1526 -225 -1500
rect -159 -1522 -129 -1500
rect -369 -1572 -353 -1538
rect -319 -1572 -303 -1538
rect -369 -1588 -303 -1572
rect -177 -1538 -111 -1522
rect -63 -1526 -33 -1500
rect 33 -1522 63 -1500
rect -177 -1572 -161 -1538
rect -127 -1572 -111 -1538
rect -177 -1588 -111 -1572
rect 15 -1538 81 -1522
rect 129 -1526 159 -1500
rect 225 -1522 255 -1500
rect 15 -1572 31 -1538
rect 65 -1572 81 -1538
rect 15 -1588 81 -1572
rect 207 -1538 273 -1522
rect 321 -1526 351 -1500
rect 417 -1522 447 -1500
rect 207 -1572 223 -1538
rect 257 -1572 273 -1538
rect 207 -1588 273 -1572
rect 399 -1538 465 -1522
rect 513 -1526 543 -1500
rect 609 -1522 639 -1500
rect 399 -1572 415 -1538
rect 449 -1572 465 -1538
rect 399 -1588 465 -1572
rect 591 -1538 657 -1522
rect 705 -1526 735 -1500
rect 801 -1522 831 -1500
rect 591 -1572 607 -1538
rect 641 -1572 657 -1538
rect 591 -1588 657 -1572
rect 783 -1538 849 -1522
rect 897 -1526 927 -1500
rect 783 -1572 799 -1538
rect 833 -1572 849 -1538
rect 783 -1588 849 -1572
<< polycont >>
rect -833 1538 -799 1572
rect -641 1538 -607 1572
rect -449 1538 -415 1572
rect -257 1538 -223 1572
rect -65 1538 -31 1572
rect 127 1538 161 1572
rect 319 1538 353 1572
rect 511 1538 545 1572
rect 703 1538 737 1572
rect 895 1538 929 1572
rect -929 -1572 -895 -1538
rect -737 -1572 -703 -1538
rect -545 -1572 -511 -1538
rect -353 -1572 -319 -1538
rect -161 -1572 -127 -1538
rect 31 -1572 65 -1538
rect 223 -1572 257 -1538
rect 415 -1572 449 -1538
rect 607 -1572 641 -1538
rect 799 -1572 833 -1538
<< locali >>
rect -1091 1640 -995 1674
rect 995 1640 1091 1674
rect -1091 -1640 -1057 1640
rect 1057 1578 1091 1640
rect -849 1538 -833 1572
rect -799 1538 -783 1572
rect -657 1538 -641 1572
rect -607 1538 -591 1572
rect -465 1538 -449 1572
rect -415 1538 -399 1572
rect -273 1538 -257 1572
rect -223 1538 -207 1572
rect -81 1538 -65 1572
rect -31 1538 -15 1572
rect 111 1538 127 1572
rect 161 1538 177 1572
rect 303 1538 319 1572
rect 353 1538 369 1572
rect 495 1538 511 1572
rect 545 1538 561 1572
rect 687 1538 703 1572
rect 737 1538 753 1572
rect 879 1538 895 1572
rect 929 1538 945 1572
rect -977 1488 -943 1504
rect -977 -1504 -943 -1488
rect -881 1488 -847 1504
rect -881 -1504 -847 -1488
rect -785 1488 -751 1504
rect -785 -1504 -751 -1488
rect -689 1488 -655 1504
rect -689 -1504 -655 -1488
rect -593 1488 -559 1504
rect -593 -1504 -559 -1488
rect -497 1488 -463 1504
rect -497 -1504 -463 -1488
rect -401 1488 -367 1504
rect -401 -1504 -367 -1488
rect -305 1488 -271 1504
rect -305 -1504 -271 -1488
rect -209 1488 -175 1504
rect -209 -1504 -175 -1488
rect -113 1488 -79 1504
rect -113 -1504 -79 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 79 1488 113 1504
rect 79 -1504 113 -1488
rect 175 1488 209 1504
rect 175 -1504 209 -1488
rect 271 1488 305 1504
rect 271 -1504 305 -1488
rect 367 1488 401 1504
rect 367 -1504 401 -1488
rect 463 1488 497 1504
rect 463 -1504 497 -1488
rect 559 1488 593 1504
rect 559 -1504 593 -1488
rect 655 1488 689 1504
rect 655 -1504 689 -1488
rect 751 1488 785 1504
rect 751 -1504 785 -1488
rect 847 1488 881 1504
rect 847 -1504 881 -1488
rect 943 1488 977 1504
rect 943 -1504 977 -1488
rect -945 -1572 -929 -1538
rect -895 -1572 -879 -1538
rect -753 -1572 -737 -1538
rect -703 -1572 -687 -1538
rect -561 -1572 -545 -1538
rect -511 -1572 -495 -1538
rect -369 -1572 -353 -1538
rect -319 -1572 -303 -1538
rect -177 -1572 -161 -1538
rect -127 -1572 -111 -1538
rect 15 -1572 31 -1538
rect 65 -1572 81 -1538
rect 207 -1572 223 -1538
rect 257 -1572 273 -1538
rect 399 -1572 415 -1538
rect 449 -1572 465 -1538
rect 591 -1572 607 -1538
rect 641 -1572 657 -1538
rect 783 -1572 799 -1538
rect 833 -1572 849 -1538
rect 1057 -1640 1091 -1578
rect -1091 -1674 1091 -1640
<< viali >>
rect -833 1538 -799 1572
rect -641 1538 -607 1572
rect -449 1538 -415 1572
rect -257 1538 -223 1572
rect -65 1538 -31 1572
rect 127 1538 161 1572
rect 319 1538 353 1572
rect 511 1538 545 1572
rect 703 1538 737 1572
rect 895 1538 929 1572
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
rect -929 -1572 -895 -1538
rect -737 -1572 -703 -1538
rect -545 -1572 -511 -1538
rect -353 -1572 -319 -1538
rect -161 -1572 -127 -1538
rect 31 -1572 65 -1538
rect 223 -1572 257 -1538
rect 415 -1572 449 -1538
rect 607 -1572 641 -1538
rect 799 -1572 833 -1538
<< metal1 >>
rect -845 1572 -787 1578
rect -845 1538 -833 1572
rect -799 1538 -787 1572
rect -845 1532 -787 1538
rect -653 1572 -595 1578
rect -653 1538 -641 1572
rect -607 1538 -595 1572
rect -653 1532 -595 1538
rect -461 1572 -403 1578
rect -461 1538 -449 1572
rect -415 1538 -403 1572
rect -461 1532 -403 1538
rect -269 1572 -211 1578
rect -269 1538 -257 1572
rect -223 1538 -211 1572
rect -269 1532 -211 1538
rect -77 1572 -19 1578
rect -77 1538 -65 1572
rect -31 1538 -19 1572
rect -77 1532 -19 1538
rect 115 1572 173 1578
rect 115 1538 127 1572
rect 161 1538 173 1572
rect 115 1532 173 1538
rect 307 1572 365 1578
rect 307 1538 319 1572
rect 353 1538 365 1572
rect 307 1532 365 1538
rect 499 1572 557 1578
rect 499 1538 511 1572
rect 545 1538 557 1572
rect 499 1532 557 1538
rect 691 1572 749 1578
rect 691 1538 703 1572
rect 737 1538 749 1572
rect 691 1532 749 1538
rect 883 1572 941 1578
rect 883 1538 895 1572
rect 929 1538 941 1572
rect 883 1532 941 1538
rect -983 1488 -937 1500
rect -983 -1488 -977 1488
rect -943 -1488 -937 1488
rect -983 -1500 -937 -1488
rect -887 1488 -841 1500
rect -887 -1488 -881 1488
rect -847 -1488 -841 1488
rect -887 -1500 -841 -1488
rect -791 1488 -745 1500
rect -791 -1488 -785 1488
rect -751 -1488 -745 1488
rect -791 -1500 -745 -1488
rect -695 1488 -649 1500
rect -695 -1488 -689 1488
rect -655 -1488 -649 1488
rect -695 -1500 -649 -1488
rect -599 1488 -553 1500
rect -599 -1488 -593 1488
rect -559 -1488 -553 1488
rect -599 -1500 -553 -1488
rect -503 1488 -457 1500
rect -503 -1488 -497 1488
rect -463 -1488 -457 1488
rect -503 -1500 -457 -1488
rect -407 1488 -361 1500
rect -407 -1488 -401 1488
rect -367 -1488 -361 1488
rect -407 -1500 -361 -1488
rect -311 1488 -265 1500
rect -311 -1488 -305 1488
rect -271 -1488 -265 1488
rect -311 -1500 -265 -1488
rect -215 1488 -169 1500
rect -215 -1488 -209 1488
rect -175 -1488 -169 1488
rect -215 -1500 -169 -1488
rect -119 1488 -73 1500
rect -119 -1488 -113 1488
rect -79 -1488 -73 1488
rect -119 -1500 -73 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 73 1488 119 1500
rect 73 -1488 79 1488
rect 113 -1488 119 1488
rect 73 -1500 119 -1488
rect 169 1488 215 1500
rect 169 -1488 175 1488
rect 209 -1488 215 1488
rect 169 -1500 215 -1488
rect 265 1488 311 1500
rect 265 -1488 271 1488
rect 305 -1488 311 1488
rect 265 -1500 311 -1488
rect 361 1488 407 1500
rect 361 -1488 367 1488
rect 401 -1488 407 1488
rect 361 -1500 407 -1488
rect 457 1488 503 1500
rect 457 -1488 463 1488
rect 497 -1488 503 1488
rect 457 -1500 503 -1488
rect 553 1488 599 1500
rect 553 -1488 559 1488
rect 593 -1488 599 1488
rect 553 -1500 599 -1488
rect 649 1488 695 1500
rect 649 -1488 655 1488
rect 689 -1488 695 1488
rect 649 -1500 695 -1488
rect 745 1488 791 1500
rect 745 -1488 751 1488
rect 785 -1488 791 1488
rect 745 -1500 791 -1488
rect 841 1488 887 1500
rect 841 -1488 847 1488
rect 881 -1488 887 1488
rect 841 -1500 887 -1488
rect 937 1488 983 1500
rect 937 -1488 943 1488
rect 977 -1488 983 1488
rect 937 -1500 983 -1488
rect -941 -1538 -883 -1532
rect -941 -1572 -929 -1538
rect -895 -1572 -883 -1538
rect -941 -1578 -883 -1572
rect -749 -1538 -691 -1532
rect -749 -1572 -737 -1538
rect -703 -1572 -691 -1538
rect -749 -1578 -691 -1572
rect -557 -1538 -499 -1532
rect -557 -1572 -545 -1538
rect -511 -1572 -499 -1538
rect -557 -1578 -499 -1572
rect -365 -1538 -307 -1532
rect -365 -1572 -353 -1538
rect -319 -1572 -307 -1538
rect -365 -1578 -307 -1572
rect -173 -1538 -115 -1532
rect -173 -1572 -161 -1538
rect -127 -1572 -115 -1538
rect -173 -1578 -115 -1572
rect 19 -1538 77 -1532
rect 19 -1572 31 -1538
rect 65 -1572 77 -1538
rect 19 -1578 77 -1572
rect 211 -1538 269 -1532
rect 211 -1572 223 -1538
rect 257 -1572 269 -1538
rect 211 -1578 269 -1572
rect 403 -1538 461 -1532
rect 403 -1572 415 -1538
rect 449 -1572 461 -1538
rect 403 -1578 461 -1572
rect 595 -1538 653 -1532
rect 595 -1572 607 -1538
rect 641 -1572 653 -1538
rect 595 -1578 653 -1572
rect 787 -1538 845 -1532
rect 787 -1572 799 -1538
rect 833 -1572 845 -1538
rect 787 -1578 845 -1572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1074 -1657 1074 1657
string parameters w 15 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
