magic
tech sky130A
magscale 1 2
timestamp 1615928575
<< nmos >>
rect -2274 -1531 -1674 1469
rect -1616 -1531 -1016 1469
rect -958 -1531 -358 1469
rect -300 -1531 300 1469
rect 358 -1531 958 1469
rect 1016 -1531 1616 1469
rect 1674 -1531 2274 1469
<< ndiff >>
rect -2332 1457 -2274 1469
rect -2332 -1519 -2320 1457
rect -2286 -1519 -2274 1457
rect -2332 -1531 -2274 -1519
rect -1674 1457 -1616 1469
rect -1674 -1519 -1662 1457
rect -1628 -1519 -1616 1457
rect -1674 -1531 -1616 -1519
rect -1016 1457 -958 1469
rect -1016 -1519 -1004 1457
rect -970 -1519 -958 1457
rect -1016 -1531 -958 -1519
rect -358 1457 -300 1469
rect -358 -1519 -346 1457
rect -312 -1519 -300 1457
rect -358 -1531 -300 -1519
rect 300 1457 358 1469
rect 300 -1519 312 1457
rect 346 -1519 358 1457
rect 300 -1531 358 -1519
rect 958 1457 1016 1469
rect 958 -1519 970 1457
rect 1004 -1519 1016 1457
rect 958 -1531 1016 -1519
rect 1616 1457 1674 1469
rect 1616 -1519 1628 1457
rect 1662 -1519 1674 1457
rect 1616 -1531 1674 -1519
rect 2274 1457 2332 1469
rect 2274 -1519 2286 1457
rect 2320 -1519 2332 1457
rect 2274 -1531 2332 -1519
<< ndiffc >>
rect -2320 -1519 -2286 1457
rect -1662 -1519 -1628 1457
rect -1004 -1519 -970 1457
rect -346 -1519 -312 1457
rect 312 -1519 346 1457
rect 970 -1519 1004 1457
rect 1628 -1519 1662 1457
rect 2286 -1519 2320 1457
<< poly >>
rect -2274 1541 -1674 1557
rect -2274 1507 -2258 1541
rect -1690 1507 -1674 1541
rect -2274 1469 -1674 1507
rect -1616 1541 -1016 1557
rect -1616 1507 -1600 1541
rect -1032 1507 -1016 1541
rect -1616 1469 -1016 1507
rect -958 1541 -358 1557
rect -958 1507 -942 1541
rect -374 1507 -358 1541
rect -958 1469 -358 1507
rect -300 1541 300 1557
rect -300 1507 -284 1541
rect 284 1507 300 1541
rect -300 1469 300 1507
rect 358 1541 958 1557
rect 358 1507 374 1541
rect 942 1507 958 1541
rect 358 1469 958 1507
rect 1016 1541 1616 1557
rect 1016 1507 1032 1541
rect 1600 1507 1616 1541
rect 1016 1469 1616 1507
rect 1674 1541 2274 1557
rect 1674 1507 1690 1541
rect 2258 1507 2274 1541
rect 1674 1469 2274 1507
rect -2274 -1557 -1674 -1531
rect -1616 -1557 -1016 -1531
rect -958 -1557 -358 -1531
rect -300 -1557 300 -1531
rect 358 -1557 958 -1531
rect 1016 -1557 1616 -1531
rect 1674 -1557 2274 -1531
<< polycont >>
rect -2258 1507 -1690 1541
rect -1600 1507 -1032 1541
rect -942 1507 -374 1541
rect -284 1507 284 1541
rect 374 1507 942 1541
rect 1032 1507 1600 1541
rect 1690 1507 2258 1541
<< locali >>
rect -2274 1507 -2258 1541
rect -1690 1507 -1674 1541
rect -1616 1507 -1600 1541
rect -1032 1507 -1016 1541
rect -958 1507 -942 1541
rect -374 1507 -358 1541
rect -300 1507 -284 1541
rect 284 1507 300 1541
rect 358 1507 374 1541
rect 942 1507 958 1541
rect 1016 1507 1032 1541
rect 1600 1507 1616 1541
rect 1674 1507 1690 1541
rect 2258 1507 2274 1541
rect -2320 1457 -2286 1473
rect -2320 -1535 -2286 -1519
rect -1662 1457 -1628 1473
rect -1662 -1535 -1628 -1519
rect -1004 1457 -970 1473
rect -1004 -1535 -970 -1519
rect -346 1457 -312 1473
rect -346 -1535 -312 -1519
rect 312 1457 346 1473
rect 312 -1535 346 -1519
rect 970 1457 1004 1473
rect 970 -1535 1004 -1519
rect 1628 1457 1662 1473
rect 1628 -1535 1662 -1519
rect 2286 1457 2320 1473
rect 2286 -1535 2320 -1519
<< viali >>
rect -2258 1507 -1690 1541
rect -1600 1507 -1032 1541
rect -942 1507 -374 1541
rect -284 1507 284 1541
rect 374 1507 942 1541
rect 1032 1507 1600 1541
rect 1690 1507 2258 1541
rect -2320 -1519 -2286 1457
rect -1662 -1519 -1628 1457
rect -1004 -1519 -970 1457
rect -346 -1519 -312 1457
rect 312 -1519 346 1457
rect 970 -1519 1004 1457
rect 1628 -1519 1662 1457
rect 2286 -1519 2320 1457
<< metal1 >>
rect -2270 1541 -1678 1547
rect -2270 1507 -2258 1541
rect -1690 1507 -1678 1541
rect -2270 1501 -1678 1507
rect -1612 1541 -1020 1547
rect -1612 1507 -1600 1541
rect -1032 1507 -1020 1541
rect -1612 1501 -1020 1507
rect -954 1541 -362 1547
rect -954 1507 -942 1541
rect -374 1507 -362 1541
rect -954 1501 -362 1507
rect -296 1541 296 1547
rect -296 1507 -284 1541
rect 284 1507 296 1541
rect -296 1501 296 1507
rect 362 1541 954 1547
rect 362 1507 374 1541
rect 942 1507 954 1541
rect 362 1501 954 1507
rect 1020 1541 1612 1547
rect 1020 1507 1032 1541
rect 1600 1507 1612 1541
rect 1020 1501 1612 1507
rect 1678 1541 2270 1547
rect 1678 1507 1690 1541
rect 2258 1507 2270 1541
rect 1678 1501 2270 1507
rect -2326 1457 -2280 1469
rect -2326 -1519 -2320 1457
rect -2286 -1519 -2280 1457
rect -2326 -1531 -2280 -1519
rect -1668 1457 -1622 1469
rect -1668 -1519 -1662 1457
rect -1628 -1519 -1622 1457
rect -1668 -1531 -1622 -1519
rect -1010 1457 -964 1469
rect -1010 -1519 -1004 1457
rect -970 -1519 -964 1457
rect -1010 -1531 -964 -1519
rect -352 1457 -306 1469
rect -352 -1519 -346 1457
rect -312 -1519 -306 1457
rect -352 -1531 -306 -1519
rect 306 1457 352 1469
rect 306 -1519 312 1457
rect 346 -1519 352 1457
rect 306 -1531 352 -1519
rect 964 1457 1010 1469
rect 964 -1519 970 1457
rect 1004 -1519 1010 1457
rect 964 -1531 1010 -1519
rect 1622 1457 1668 1469
rect 1622 -1519 1628 1457
rect 1662 -1519 1668 1457
rect 1622 -1531 1668 -1519
rect 2280 1457 2326 1469
rect 2280 -1519 2286 1457
rect 2320 -1519 2326 1457
rect 2280 -1531 2326 -1519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 15 l 3 m 1 nf 7 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
