magic
tech sky130A
magscale 1 2
timestamp 1615944125
<< pwell >>
rect -1701 -448 1701 448
<< nmos >>
rect -1505 -300 -1445 300
rect -1387 -300 -1327 300
rect -1269 -300 -1209 300
rect -1151 -300 -1091 300
rect -1033 -300 -973 300
rect -915 -300 -855 300
rect -797 -300 -737 300
rect -679 -300 -619 300
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect 619 -300 679 300
rect 737 -300 797 300
rect 855 -300 915 300
rect 973 -300 1033 300
rect 1091 -300 1151 300
rect 1209 -300 1269 300
rect 1327 -300 1387 300
rect 1445 -300 1505 300
<< ndiff >>
rect -1563 288 -1505 300
rect -1563 -288 -1551 288
rect -1517 -288 -1505 288
rect -1563 -300 -1505 -288
rect -1445 288 -1387 300
rect -1445 -288 -1433 288
rect -1399 -288 -1387 288
rect -1445 -300 -1387 -288
rect -1327 288 -1269 300
rect -1327 -288 -1315 288
rect -1281 -288 -1269 288
rect -1327 -300 -1269 -288
rect -1209 288 -1151 300
rect -1209 -288 -1197 288
rect -1163 -288 -1151 288
rect -1209 -300 -1151 -288
rect -1091 288 -1033 300
rect -1091 -288 -1079 288
rect -1045 -288 -1033 288
rect -1091 -300 -1033 -288
rect -973 288 -915 300
rect -973 -288 -961 288
rect -927 -288 -915 288
rect -973 -300 -915 -288
rect -855 288 -797 300
rect -855 -288 -843 288
rect -809 -288 -797 288
rect -855 -300 -797 -288
rect -737 288 -679 300
rect -737 -288 -725 288
rect -691 -288 -679 288
rect -737 -300 -679 -288
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect 679 288 737 300
rect 679 -288 691 288
rect 725 -288 737 288
rect 679 -300 737 -288
rect 797 288 855 300
rect 797 -288 809 288
rect 843 -288 855 288
rect 797 -300 855 -288
rect 915 288 973 300
rect 915 -288 927 288
rect 961 -288 973 288
rect 915 -300 973 -288
rect 1033 288 1091 300
rect 1033 -288 1045 288
rect 1079 -288 1091 288
rect 1033 -300 1091 -288
rect 1151 288 1209 300
rect 1151 -288 1163 288
rect 1197 -288 1209 288
rect 1151 -300 1209 -288
rect 1269 288 1327 300
rect 1269 -288 1281 288
rect 1315 -288 1327 288
rect 1269 -300 1327 -288
rect 1387 288 1445 300
rect 1387 -288 1399 288
rect 1433 -288 1445 288
rect 1387 -300 1445 -288
rect 1505 288 1563 300
rect 1505 -288 1517 288
rect 1551 -288 1563 288
rect 1505 -300 1563 -288
<< ndiffc >>
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
<< psubdiff >>
rect -1665 378 -1569 412
rect 1569 378 1665 412
rect -1665 316 -1631 378
rect 1631 316 1665 378
rect -1665 -378 -1631 -316
rect 1631 -378 1665 -316
rect -1665 -412 -1569 -378
rect 1569 -412 1665 -378
<< psubdiffcont >>
rect -1569 378 1569 412
rect -1665 -316 -1631 316
rect 1631 -316 1665 316
rect -1569 -412 1569 -378
<< poly >>
rect -1505 300 -1445 326
rect -1387 300 -1327 326
rect -1269 300 -1209 326
rect -1151 300 -1091 326
rect -1033 300 -973 326
rect -915 300 -855 326
rect -797 300 -737 326
rect -679 300 -619 326
rect -561 300 -501 326
rect -443 300 -383 326
rect -325 300 -265 326
rect -207 300 -147 326
rect -89 300 -29 326
rect 29 300 89 326
rect 147 300 207 326
rect 265 300 325 326
rect 383 300 443 326
rect 501 300 561 326
rect 619 300 679 326
rect 737 300 797 326
rect 855 300 915 326
rect 973 300 1033 326
rect 1091 300 1151 326
rect 1209 300 1269 326
rect 1327 300 1387 326
rect 1445 300 1505 326
rect -1505 -326 -1445 -300
rect -1387 -326 -1327 -300
rect -1269 -326 -1209 -300
rect -1151 -326 -1091 -300
rect -1033 -326 -973 -300
rect -915 -326 -855 -300
rect -797 -326 -737 -300
rect -679 -326 -619 -300
rect -561 -326 -501 -300
rect -443 -326 -383 -300
rect -325 -326 -265 -300
rect -207 -326 -147 -300
rect -89 -326 -29 -300
rect 29 -326 89 -300
rect 147 -326 207 -300
rect 265 -326 325 -300
rect 383 -326 443 -300
rect 501 -326 561 -300
rect 619 -326 679 -300
rect 737 -326 797 -300
rect 855 -326 915 -300
rect 973 -326 1033 -300
rect 1091 -326 1151 -300
rect 1209 -326 1269 -300
rect 1327 -326 1387 -300
rect 1445 -326 1505 -300
<< locali >>
rect -1665 378 -1569 412
rect 1569 378 1665 412
rect -1665 316 -1631 378
rect 1631 316 1665 378
rect -1551 288 -1517 304
rect -1551 -304 -1517 -288
rect -1433 288 -1399 304
rect -1433 -304 -1399 -288
rect -1315 288 -1281 304
rect -1315 -304 -1281 -288
rect -1197 288 -1163 304
rect -1197 -304 -1163 -288
rect -1079 288 -1045 304
rect -1079 -304 -1045 -288
rect -961 288 -927 304
rect -961 -304 -927 -288
rect -843 288 -809 304
rect -843 -304 -809 -288
rect -725 288 -691 304
rect -725 -304 -691 -288
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect 691 288 725 304
rect 691 -304 725 -288
rect 809 288 843 304
rect 809 -304 843 -288
rect 927 288 961 304
rect 927 -304 961 -288
rect 1045 288 1079 304
rect 1045 -304 1079 -288
rect 1163 288 1197 304
rect 1163 -304 1197 -288
rect 1281 288 1315 304
rect 1281 -304 1315 -288
rect 1399 288 1433 304
rect 1399 -304 1433 -288
rect 1517 288 1551 304
rect 1517 -304 1551 -288
rect -1665 -378 -1631 -316
rect 1631 -378 1665 -316
rect -1665 -412 -1569 -378
rect 1569 -412 1665 -378
<< viali >>
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
<< metal1 >>
rect -1557 288 -1511 300
rect -1557 -288 -1551 288
rect -1517 -288 -1511 288
rect -1557 -300 -1511 -288
rect -1439 288 -1393 300
rect -1439 -288 -1433 288
rect -1399 -288 -1393 288
rect -1439 -300 -1393 -288
rect -1321 288 -1275 300
rect -1321 -288 -1315 288
rect -1281 -288 -1275 288
rect -1321 -300 -1275 -288
rect -1203 288 -1157 300
rect -1203 -288 -1197 288
rect -1163 -288 -1157 288
rect -1203 -300 -1157 -288
rect -1085 288 -1039 300
rect -1085 -288 -1079 288
rect -1045 -288 -1039 288
rect -1085 -300 -1039 -288
rect -967 288 -921 300
rect -967 -288 -961 288
rect -927 -288 -921 288
rect -967 -300 -921 -288
rect -849 288 -803 300
rect -849 -288 -843 288
rect -809 -288 -803 288
rect -849 -300 -803 -288
rect -731 288 -685 300
rect -731 -288 -725 288
rect -691 -288 -685 288
rect -731 -300 -685 -288
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect 685 288 731 300
rect 685 -288 691 288
rect 725 -288 731 288
rect 685 -300 731 -288
rect 803 288 849 300
rect 803 -288 809 288
rect 843 -288 849 288
rect 803 -300 849 -288
rect 921 288 967 300
rect 921 -288 927 288
rect 961 -288 967 288
rect 921 -300 967 -288
rect 1039 288 1085 300
rect 1039 -288 1045 288
rect 1079 -288 1085 288
rect 1039 -300 1085 -288
rect 1157 288 1203 300
rect 1157 -288 1163 288
rect 1197 -288 1203 288
rect 1157 -300 1203 -288
rect 1275 288 1321 300
rect 1275 -288 1281 288
rect 1315 -288 1321 288
rect 1275 -300 1321 -288
rect 1393 288 1439 300
rect 1393 -288 1399 288
rect 1433 -288 1439 288
rect 1393 -300 1439 -288
rect 1511 288 1557 300
rect 1511 -288 1517 288
rect 1551 -288 1557 288
rect 1511 -300 1557 -288
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1648 -395 1648 395
string parameters w 3 l 0.3 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
