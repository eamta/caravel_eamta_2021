magic
tech sky130A
magscale 1 2
timestamp 1615949206
<< metal1 >>
rect 5629 1891 5935 1915
rect 5629 1812 5694 1891
rect 5869 1812 5935 1891
rect 5629 1683 5935 1812
rect 5419 1637 6145 1683
rect 5363 -92 5409 1605
rect 5548 77 5558 1593
rect 5610 77 5620 1593
rect 5759 -92 5805 1605
rect 5944 77 5954 1593
rect 6006 77 6016 1593
rect 6155 -92 6201 1605
<< via1 >>
rect 5694 1812 5869 1891
rect 5558 77 5610 1593
rect 5954 77 6006 1593
<< metal2 >>
rect 5558 2049 6006 2059
rect 5558 1989 5669 2049
rect 5729 1989 5761 2049
rect 5821 1989 5855 2049
rect 5915 1989 6006 2049
rect 5558 1979 6006 1989
rect 5558 1593 5610 1979
rect 5694 1891 5869 1901
rect 5694 1802 5869 1812
rect 5558 67 5610 77
rect 5954 1593 6006 1979
rect 5954 67 6006 77
<< via2 >>
rect 5669 1989 5729 2049
rect 5761 1989 5821 2049
rect 5855 1989 5915 2049
rect 5694 1812 5869 1891
<< metal3 >>
rect 5657 2049 6116 2059
rect 5657 1989 5669 2049
rect 5729 1989 5761 2049
rect 5821 1989 5855 2049
rect 5915 1989 6116 2049
rect 5657 1979 6116 1989
rect 4940 1891 5883 1915
rect 4940 1812 5694 1891
rect 5869 1812 5883 1891
rect 4940 1788 5883 1812
use sky130_fd_pr__nfet_01v8_MXMZMC  sky130_fd_pr__nfet_01v8_MXMZMC_0
timestamp 1615949206
transform 1 0 5782 0 1 866
box -563 -949 563 949
<< end >>
