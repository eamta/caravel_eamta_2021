magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 298 1095 333 1129
rect 299 1076 333 1095
rect 129 1027 187 1033
rect 129 993 141 1027
rect 129 987 187 993
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 318 583 333 1076
rect 352 1042 387 1076
rect 667 1042 702 1076
rect 352 583 386 1042
rect 668 1023 702 1042
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 352 549 367 583
rect 687 530 702 1023
rect 721 989 756 1023
rect 1036 989 1071 1023
rect 721 646 755 989
rect 1037 970 1071 989
rect 1056 927 1071 970
rect 867 921 925 927
rect 867 887 879 921
rect 867 881 925 887
rect 835 770 869 804
rect 923 770 957 804
rect 1037 770 1071 927
rect 1090 936 1125 970
rect 1405 936 1440 953
rect 1090 770 1124 936
rect 1406 935 1440 936
rect 1406 899 1476 935
rect 1423 874 1494 899
rect 1236 868 1294 874
rect 1236 836 1248 868
rect 1406 865 1494 874
rect 1774 865 1809 899
rect 1236 828 1294 836
rect 1406 808 1493 865
rect 1775 846 1809 865
rect 1208 804 1322 808
rect 1204 800 1326 804
rect 1204 770 1238 800
rect 1292 770 1326 800
rect 1406 770 1756 808
rect 762 736 1756 770
rect 823 660 881 700
rect 888 660 969 700
rect 923 656 957 660
rect 721 530 756 646
rect 866 631 888 646
rect 881 629 888 631
rect 863 619 888 629
rect 942 634 960 646
rect 942 622 988 634
rect 863 613 925 619
rect 863 579 888 613
rect 920 579 929 613
rect 942 579 963 622
rect 863 573 925 579
rect 863 563 888 573
rect 873 548 888 563
rect 942 548 944 579
rect 954 545 963 579
rect 1037 568 1076 736
rect 721 496 736 530
rect 742 511 755 530
rect 1037 511 1071 568
rect 742 477 888 511
rect 942 477 1071 511
rect 1090 512 1124 736
rect 1192 665 1230 700
rect 1130 534 1158 634
rect 1165 618 1176 646
rect 1192 632 1246 665
rect 1192 607 1250 632
rect 1292 619 1326 652
rect 1327 646 1338 687
rect 1200 582 1250 607
rect 1284 594 1329 607
rect 1212 568 1246 582
rect 1284 568 1330 594
rect 1284 566 1329 568
rect 1236 560 1329 566
rect 1232 534 1329 560
rect 1236 526 1248 534
rect 1284 526 1329 534
rect 1236 520 1298 526
rect 1284 512 1298 520
rect 1406 512 1756 736
rect 1090 466 1176 512
rect 1284 466 1342 512
rect 1372 466 1756 512
rect 1090 435 1118 466
rect 1406 458 1756 466
rect 1124 441 1176 458
rect 1201 447 1257 458
rect 1284 452 1406 458
rect 1284 448 1410 452
rect 1423 448 1756 458
rect 1212 435 1246 447
rect 1284 441 1756 448
rect 1090 424 1129 435
rect 1201 424 1257 435
rect 1288 430 1756 441
rect 1288 424 1476 430
rect 1423 414 1476 424
rect 1020 380 1024 414
rect 1322 390 1476 414
rect 1555 394 1673 405
rect 1423 388 1476 390
rect 1459 382 1460 388
rect 1566 382 1662 394
rect 1459 376 1471 382
rect 1555 376 1673 382
rect 1459 371 1674 376
rect 1794 371 1809 846
rect 1828 812 1863 846
rect 2143 812 2178 846
rect 1828 371 1862 812
rect 2144 793 2178 812
rect 1974 744 2032 750
rect 1974 710 1986 744
rect 1974 704 2032 710
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1130 308 1132 342
rect 1425 337 1674 342
rect 1828 337 1843 371
rect 2163 318 2178 793
rect 2197 759 2232 793
rect 2512 759 2547 793
rect 2197 318 2231 759
rect 2513 740 2547 759
rect 2899 740 2952 741
rect 2343 691 2401 697
rect 2343 657 2355 691
rect 2343 651 2401 657
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 904 238 908 272
rect 1462 244 1464 272
rect 2532 265 2547 740
rect 2566 706 2601 740
rect 2881 706 2952 740
rect 2566 265 2600 706
rect 2882 705 2952 706
rect 2899 671 2970 705
rect 3250 671 3285 705
rect 2712 638 2770 644
rect 2712 604 2724 638
rect 2712 598 2770 604
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 1430 238 1464 244
rect 2566 231 2581 265
rect 2899 212 2969 671
rect 3251 652 3285 671
rect 3081 603 3139 609
rect 3081 569 3093 603
rect 3081 563 3139 569
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2899 176 2952 212
rect 3270 159 3285 652
rect 3304 618 3339 652
rect 3304 159 3338 618
rect 3450 550 3508 556
rect 3450 516 3462 550
rect 3620 527 3654 545
rect 3450 510 3508 516
rect 3620 491 3690 527
rect 3637 457 3708 491
rect 3988 457 4023 491
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 1174 90 1176 128
rect 3304 125 3319 159
rect 3637 106 3707 457
rect 3989 438 4023 457
rect 3819 389 3877 395
rect 3819 355 3831 389
rect 3819 349 3877 355
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 1212 54 1214 90
rect 3637 70 3690 106
rect 4008 53 4023 438
rect 4042 404 4077 438
rect 4042 53 4076 404
rect 4188 336 4246 342
rect 4188 302 4200 336
rect 4188 296 4246 302
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
<< nwell >>
rect 706 430 1756 808
<< nmos >>
rect 800 28 830 118
rect 1000 26 1030 206
rect 1088 26 1118 206
rect 1342 26 1372 206
rect 1430 26 1460 206
rect 1632 28 1662 118
<< pmos >>
rect 800 466 830 646
rect 1000 466 1030 646
rect 1088 466 1118 646
rect 1342 466 1372 646
rect 1430 466 1460 646
rect 1632 466 1662 646
<< ndiff >>
rect 742 88 800 118
rect 742 54 754 88
rect 788 54 800 88
rect 742 28 800 54
rect 830 88 888 118
rect 830 54 842 88
rect 876 54 888 88
rect 830 28 888 54
rect 942 88 1000 206
rect 942 54 954 88
rect 988 54 1000 88
rect 942 26 1000 54
rect 1030 88 1088 206
rect 1030 54 1042 88
rect 1076 54 1088 88
rect 1030 26 1088 54
rect 1118 88 1176 206
rect 1118 54 1130 88
rect 1164 54 1176 88
rect 1118 26 1176 54
rect 1284 88 1342 206
rect 1284 54 1296 88
rect 1330 54 1342 88
rect 1284 26 1342 54
rect 1372 26 1430 206
rect 1460 88 1518 206
rect 1460 54 1472 88
rect 1506 54 1518 88
rect 1460 26 1518 54
rect 1574 88 1632 118
rect 1574 54 1586 88
rect 1620 54 1632 88
rect 1574 28 1632 54
rect 1662 88 1720 118
rect 1662 54 1674 88
rect 1708 54 1720 88
rect 1662 28 1720 54
<< pdiff >>
rect 742 618 800 646
rect 742 584 754 618
rect 788 584 800 618
rect 742 466 800 584
rect 830 618 888 646
rect 830 584 842 618
rect 876 584 888 618
rect 830 466 888 584
rect 942 618 1000 646
rect 942 584 954 618
rect 988 584 1000 618
rect 942 466 1000 584
rect 1030 618 1088 646
rect 1030 584 1042 618
rect 1076 584 1088 618
rect 1030 466 1088 584
rect 1118 618 1176 646
rect 1118 584 1130 618
rect 1164 584 1176 618
rect 1118 466 1176 584
rect 1284 618 1342 646
rect 1284 584 1296 618
rect 1330 584 1342 618
rect 1284 466 1342 584
rect 1372 618 1430 646
rect 1372 584 1384 618
rect 1418 584 1430 618
rect 1372 466 1430 584
rect 1460 618 1518 646
rect 1460 584 1472 618
rect 1506 584 1518 618
rect 1460 466 1518 584
rect 1574 618 1632 646
rect 1574 584 1586 618
rect 1620 584 1632 618
rect 1574 466 1632 584
rect 1662 618 1720 646
rect 1662 584 1674 618
rect 1708 584 1720 618
rect 1662 466 1720 584
<< ndiffc >>
rect 754 54 788 88
rect 842 54 876 88
rect 954 54 988 88
rect 1042 54 1076 88
rect 1130 54 1164 88
rect 1296 54 1330 88
rect 1472 54 1506 88
rect 1586 54 1620 88
rect 1674 54 1708 88
<< pdiffc >>
rect 754 584 788 618
rect 842 584 876 618
rect 954 584 988 618
rect 1042 584 1076 618
rect 1130 584 1164 618
rect 1296 584 1330 618
rect 1384 584 1418 618
rect 1472 584 1506 618
rect 1586 584 1620 618
rect 1674 584 1708 618
<< psubdiff >>
rect 762 -64 786 -30
rect 1678 -64 1702 -30
<< nsubdiff >>
rect 762 736 786 770
rect 1676 736 1700 770
<< psubdiffcont >>
rect 786 -64 1678 -30
<< nsubdiffcont >>
rect 786 736 1676 770
<< poly >>
rect 800 646 830 672
rect 1000 646 1030 672
rect 1088 646 1118 672
rect 1342 646 1372 672
rect 1430 646 1460 672
rect 1632 646 1662 672
rect 1196 618 1262 632
rect 1196 584 1212 618
rect 1246 584 1262 618
rect 1196 566 1262 584
rect 800 288 830 466
rect 1000 430 1030 466
rect 970 414 1038 430
rect 970 380 990 414
rect 1020 380 1038 414
rect 970 364 1038 380
rect 800 272 922 288
rect 800 238 874 272
rect 904 238 922 272
rect 800 222 922 238
rect 800 118 830 222
rect 1000 206 1030 364
rect 1088 358 1118 466
rect 1080 342 1146 358
rect 1080 308 1098 342
rect 1130 308 1146 342
rect 1080 292 1146 308
rect 1088 206 1118 292
rect 800 2 830 28
rect 1212 104 1246 566
rect 1342 430 1372 466
rect 1322 414 1388 430
rect 1322 380 1338 414
rect 1372 380 1388 414
rect 1322 364 1388 380
rect 1342 206 1372 364
rect 1430 288 1460 466
rect 1632 430 1662 466
rect 1566 414 1662 430
rect 1566 380 1582 414
rect 1616 380 1662 414
rect 1566 364 1662 380
rect 1414 272 1478 288
rect 1414 238 1430 272
rect 1462 238 1478 272
rect 1414 222 1478 238
rect 1430 206 1460 222
rect 1196 90 1262 104
rect 1196 54 1212 90
rect 1246 54 1262 90
rect 1196 38 1262 54
rect 1632 118 1662 364
rect 1000 0 1030 26
rect 1088 0 1118 26
rect 1342 0 1372 26
rect 1430 0 1460 26
rect 1632 2 1662 28
<< polycont >>
rect 1212 584 1246 618
rect 990 380 1020 414
rect 874 238 904 272
rect 1098 308 1130 342
rect 1338 380 1372 414
rect 1582 380 1616 414
rect 1430 238 1462 272
rect 1212 54 1246 90
<< locali >>
rect 754 736 786 770
rect 1676 736 1692 770
rect 754 618 788 634
rect 754 414 788 584
rect 842 618 876 736
rect 842 568 876 584
rect 954 618 988 634
rect 954 534 988 584
rect 1042 618 1076 736
rect 1212 668 1506 702
rect 1042 568 1076 584
rect 1130 618 1164 634
rect 1130 534 1164 584
rect 1212 618 1246 668
rect 1212 568 1246 584
rect 1296 618 1330 668
rect 1296 568 1330 584
rect 1384 618 1418 634
rect 1384 534 1418 584
rect 1472 618 1506 668
rect 1472 568 1506 584
rect 1586 618 1620 736
rect 1586 568 1620 584
rect 1674 618 1708 634
rect 954 500 1418 534
rect 754 380 990 414
rect 1020 380 1040 414
rect 1322 380 1338 414
rect 1372 380 1582 414
rect 1616 380 1632 414
rect 754 88 788 380
rect 1674 342 1708 584
rect 1080 308 1098 342
rect 1130 308 1708 342
rect 854 238 874 272
rect 904 238 1428 272
rect 1462 238 1478 272
rect 754 38 788 54
rect 842 88 876 104
rect 842 -30 876 54
rect 954 88 988 104
rect 954 -30 988 54
rect 1042 88 1088 104
rect 1076 54 1088 88
rect 1042 38 1088 54
rect 1130 90 1330 104
rect 1130 88 1212 90
rect 1164 54 1212 88
rect 1246 88 1330 90
rect 1246 54 1296 88
rect 1130 38 1330 54
rect 1472 88 1506 104
rect 1472 -30 1506 54
rect 1586 88 1620 104
rect 1586 -30 1620 54
rect 1674 88 1708 308
rect 1674 38 1708 54
rect 754 -64 786 -30
rect 1678 -64 1694 -30
<< viali >>
rect 786 736 1676 770
rect 1338 380 1372 414
rect 1428 238 1430 272
rect 1430 238 1462 272
rect 1212 54 1246 90
rect 786 -64 1676 -30
<< metal1 >>
rect 706 770 1756 808
rect 706 736 786 770
rect 1676 736 1756 770
rect 706 698 1756 736
rect 1322 414 1388 430
rect 1322 380 1338 414
rect 1372 380 1388 414
rect 1322 364 1388 380
rect 1414 272 1478 288
rect 1414 238 1428 272
rect 1462 238 1478 272
rect 1414 222 1478 238
rect 0 0 200 200
rect 1196 90 1262 104
rect 1196 54 1212 90
rect 1246 54 1262 90
rect 1196 38 1262 54
rect 706 -30 1756 8
rect 706 -64 786 -30
rect 1676 -64 1756 -30
rect 706 -102 1756 -64
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use sky130_fd_pr__pfet_01v8_XSLFBL  XM0
timestamp 1624053917
transform 1 0 158 0 1 856
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM3
timestamp 1624053917
transform 1 0 1265 0 1 697
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_L9ESED  XM4
timestamp 1624053917
transform 1 0 1634 0 1 635
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM5
timestamp 1624053917
transform 1 0 2003 0 1 582
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM6
timestamp 1624053917
transform 1 0 2372 0 1 529
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM7
timestamp 1624053917
transform 1 0 2741 0 1 476
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_XSLFBL  XM8
timestamp 1624053917
transform 1 0 3110 0 1 432
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM10
timestamp 1624053917
transform 1 0 3479 0 1 379
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM11
timestamp 1624053917
transform 1 0 4217 0 1 219
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3848 0 1 272
box -211 -255 211 255
<< labels >>
rlabel metal1 1196 38 1262 54 5 Z
rlabel metal1 1228 808 1228 808 1 VDD
rlabel metal1 1228 -102 1228 -102 5 VSS
rlabel metal1 1446 222 1446 222 5 B
rlabel metal1 1322 364 1388 380 5 A
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 B
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Z
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 VDD
port 7 nsew
<< end >>
