magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -19085 222 -19027 228
rect -18893 222 -18835 228
rect -18701 222 -18643 228
rect -18509 222 -18451 228
rect -18317 222 -18259 228
rect -18125 222 -18067 228
rect -17933 222 -17875 228
rect -17741 222 -17683 228
rect -17549 222 -17491 228
rect -17357 222 -17299 228
rect -17165 222 -17107 228
rect -16973 222 -16915 228
rect -16781 222 -16723 228
rect -16589 222 -16531 228
rect -16397 222 -16339 228
rect -16205 222 -16147 228
rect -16013 222 -15955 228
rect -15821 222 -15763 228
rect -15629 222 -15571 228
rect -15437 222 -15379 228
rect -15245 222 -15187 228
rect -15053 222 -14995 228
rect -14861 222 -14803 228
rect -14669 222 -14611 228
rect -14477 222 -14419 228
rect -14285 222 -14227 228
rect -14093 222 -14035 228
rect -13901 222 -13843 228
rect -13709 222 -13651 228
rect -13517 222 -13459 228
rect -13325 222 -13267 228
rect -13133 222 -13075 228
rect -12941 222 -12883 228
rect -12749 222 -12691 228
rect -12557 222 -12499 228
rect -12365 222 -12307 228
rect -12173 222 -12115 228
rect -11981 222 -11923 228
rect -11789 222 -11731 228
rect -11597 222 -11539 228
rect -11405 222 -11347 228
rect -11213 222 -11155 228
rect -11021 222 -10963 228
rect -10829 222 -10771 228
rect -10637 222 -10579 228
rect -10445 222 -10387 228
rect -10253 222 -10195 228
rect -10061 222 -10003 228
rect -9869 222 -9811 228
rect -9677 222 -9619 228
rect -9485 222 -9427 228
rect -9293 222 -9235 228
rect -9101 222 -9043 228
rect -8909 222 -8851 228
rect -8717 222 -8659 228
rect -8525 222 -8467 228
rect -8333 222 -8275 228
rect -8141 222 -8083 228
rect -7949 222 -7891 228
rect -7757 222 -7699 228
rect -7565 222 -7507 228
rect -7373 222 -7315 228
rect -7181 222 -7123 228
rect -6989 222 -6931 228
rect -6797 222 -6739 228
rect -6605 222 -6547 228
rect -6413 222 -6355 228
rect -6221 222 -6163 228
rect -6029 222 -5971 228
rect -5837 222 -5779 228
rect -5645 222 -5587 228
rect -5453 222 -5395 228
rect -5261 222 -5203 228
rect -5069 222 -5011 228
rect -4877 222 -4819 228
rect -4685 222 -4627 228
rect -4493 222 -4435 228
rect -4301 222 -4243 228
rect -4109 222 -4051 228
rect -3917 222 -3859 228
rect -3725 222 -3667 228
rect -3533 222 -3475 228
rect -3341 222 -3283 228
rect -3149 222 -3091 228
rect -2957 222 -2899 228
rect -2765 222 -2707 228
rect -2573 222 -2515 228
rect -2381 222 -2323 228
rect -2189 222 -2131 228
rect -1997 222 -1939 228
rect -1805 222 -1747 228
rect -1613 222 -1555 228
rect -1421 222 -1363 228
rect -1229 222 -1171 228
rect -1037 222 -979 228
rect -845 222 -787 228
rect -653 222 -595 228
rect -461 222 -403 228
rect -269 222 -211 228
rect -77 222 -19 228
rect 115 222 173 228
rect 307 222 365 228
rect 499 222 557 228
rect 691 222 749 228
rect 883 222 941 228
rect 1075 222 1133 228
rect 1267 222 1325 228
rect 1459 222 1517 228
rect 1651 222 1709 228
rect 1843 222 1901 228
rect 2035 222 2093 228
rect 2227 222 2285 228
rect 2419 222 2477 228
rect 2611 222 2669 228
rect 2803 222 2861 228
rect 2995 222 3053 228
rect 3187 222 3245 228
rect 3379 222 3437 228
rect 3571 222 3629 228
rect 3763 222 3821 228
rect 3955 222 4013 228
rect 4147 222 4205 228
rect 4339 222 4397 228
rect 4531 222 4589 228
rect 4723 222 4781 228
rect 4915 222 4973 228
rect 5107 222 5165 228
rect 5299 222 5357 228
rect 5491 222 5549 228
rect 5683 222 5741 228
rect 5875 222 5933 228
rect 6067 222 6125 228
rect 6259 222 6317 228
rect 6451 222 6509 228
rect 6643 222 6701 228
rect 6835 222 6893 228
rect 7027 222 7085 228
rect 7219 222 7277 228
rect 7411 222 7469 228
rect 7603 222 7661 228
rect 7795 222 7853 228
rect 7987 222 8045 228
rect 8179 222 8237 228
rect 8371 222 8429 228
rect 8563 222 8621 228
rect 8755 222 8813 228
rect 8947 222 9005 228
rect 9139 222 9197 228
rect 9331 222 9389 228
rect 9523 222 9581 228
rect 9715 222 9773 228
rect 9907 222 9965 228
rect 10099 222 10157 228
rect 10291 222 10349 228
rect 10483 222 10541 228
rect 10675 222 10733 228
rect 10867 222 10925 228
rect 11059 222 11117 228
rect 11251 222 11309 228
rect 11443 222 11501 228
rect 11635 222 11693 228
rect 11827 222 11885 228
rect 12019 222 12077 228
rect 12211 222 12269 228
rect 12403 222 12461 228
rect 12595 222 12653 228
rect 12787 222 12845 228
rect 12979 222 13037 228
rect 13171 222 13229 228
rect 13363 222 13421 228
rect 13555 222 13613 228
rect 13747 222 13805 228
rect 13939 222 13997 228
rect 14131 222 14189 228
rect 14323 222 14381 228
rect 14515 222 14573 228
rect 14707 222 14765 228
rect 14899 222 14957 228
rect 15091 222 15149 228
rect 15283 222 15341 228
rect 15475 222 15533 228
rect 15667 222 15725 228
rect 15859 222 15917 228
rect 16051 222 16109 228
rect 16243 222 16301 228
rect 16435 222 16493 228
rect 16627 222 16685 228
rect 16819 222 16877 228
rect 17011 222 17069 228
rect 17203 222 17261 228
rect 17395 222 17453 228
rect 17587 222 17645 228
rect 17779 222 17837 228
rect 17971 222 18029 228
rect 18163 222 18221 228
rect 18355 222 18413 228
rect 18547 222 18605 228
rect 18739 222 18797 228
rect 18931 222 18989 228
rect 19123 222 19181 228
rect -19085 188 -19073 222
rect -18893 188 -18881 222
rect -18701 188 -18689 222
rect -18509 188 -18497 222
rect -18317 188 -18305 222
rect -18125 188 -18113 222
rect -17933 188 -17921 222
rect -17741 188 -17729 222
rect -17549 188 -17537 222
rect -17357 188 -17345 222
rect -17165 188 -17153 222
rect -16973 188 -16961 222
rect -16781 188 -16769 222
rect -16589 188 -16577 222
rect -16397 188 -16385 222
rect -16205 188 -16193 222
rect -16013 188 -16001 222
rect -15821 188 -15809 222
rect -15629 188 -15617 222
rect -15437 188 -15425 222
rect -15245 188 -15233 222
rect -15053 188 -15041 222
rect -14861 188 -14849 222
rect -14669 188 -14657 222
rect -14477 188 -14465 222
rect -14285 188 -14273 222
rect -14093 188 -14081 222
rect -13901 188 -13889 222
rect -13709 188 -13697 222
rect -13517 188 -13505 222
rect -13325 188 -13313 222
rect -13133 188 -13121 222
rect -12941 188 -12929 222
rect -12749 188 -12737 222
rect -12557 188 -12545 222
rect -12365 188 -12353 222
rect -12173 188 -12161 222
rect -11981 188 -11969 222
rect -11789 188 -11777 222
rect -11597 188 -11585 222
rect -11405 188 -11393 222
rect -11213 188 -11201 222
rect -11021 188 -11009 222
rect -10829 188 -10817 222
rect -10637 188 -10625 222
rect -10445 188 -10433 222
rect -10253 188 -10241 222
rect -10061 188 -10049 222
rect -9869 188 -9857 222
rect -9677 188 -9665 222
rect -9485 188 -9473 222
rect -9293 188 -9281 222
rect -9101 188 -9089 222
rect -8909 188 -8897 222
rect -8717 188 -8705 222
rect -8525 188 -8513 222
rect -8333 188 -8321 222
rect -8141 188 -8129 222
rect -7949 188 -7937 222
rect -7757 188 -7745 222
rect -7565 188 -7553 222
rect -7373 188 -7361 222
rect -7181 188 -7169 222
rect -6989 188 -6977 222
rect -6797 188 -6785 222
rect -6605 188 -6593 222
rect -6413 188 -6401 222
rect -6221 188 -6209 222
rect -6029 188 -6017 222
rect -5837 188 -5825 222
rect -5645 188 -5633 222
rect -5453 188 -5441 222
rect -5261 188 -5249 222
rect -5069 188 -5057 222
rect -4877 188 -4865 222
rect -4685 188 -4673 222
rect -4493 188 -4481 222
rect -4301 188 -4289 222
rect -4109 188 -4097 222
rect -3917 188 -3905 222
rect -3725 188 -3713 222
rect -3533 188 -3521 222
rect -3341 188 -3329 222
rect -3149 188 -3137 222
rect -2957 188 -2945 222
rect -2765 188 -2753 222
rect -2573 188 -2561 222
rect -2381 188 -2369 222
rect -2189 188 -2177 222
rect -1997 188 -1985 222
rect -1805 188 -1793 222
rect -1613 188 -1601 222
rect -1421 188 -1409 222
rect -1229 188 -1217 222
rect -1037 188 -1025 222
rect -845 188 -833 222
rect -653 188 -641 222
rect -461 188 -449 222
rect -269 188 -257 222
rect -77 188 -65 222
rect 115 188 127 222
rect 307 188 319 222
rect 499 188 511 222
rect 691 188 703 222
rect 883 188 895 222
rect 1075 188 1087 222
rect 1267 188 1279 222
rect 1459 188 1471 222
rect 1651 188 1663 222
rect 1843 188 1855 222
rect 2035 188 2047 222
rect 2227 188 2239 222
rect 2419 188 2431 222
rect 2611 188 2623 222
rect 2803 188 2815 222
rect 2995 188 3007 222
rect 3187 188 3199 222
rect 3379 188 3391 222
rect 3571 188 3583 222
rect 3763 188 3775 222
rect 3955 188 3967 222
rect 4147 188 4159 222
rect 4339 188 4351 222
rect 4531 188 4543 222
rect 4723 188 4735 222
rect 4915 188 4927 222
rect 5107 188 5119 222
rect 5299 188 5311 222
rect 5491 188 5503 222
rect 5683 188 5695 222
rect 5875 188 5887 222
rect 6067 188 6079 222
rect 6259 188 6271 222
rect 6451 188 6463 222
rect 6643 188 6655 222
rect 6835 188 6847 222
rect 7027 188 7039 222
rect 7219 188 7231 222
rect 7411 188 7423 222
rect 7603 188 7615 222
rect 7795 188 7807 222
rect 7987 188 7999 222
rect 8179 188 8191 222
rect 8371 188 8383 222
rect 8563 188 8575 222
rect 8755 188 8767 222
rect 8947 188 8959 222
rect 9139 188 9151 222
rect 9331 188 9343 222
rect 9523 188 9535 222
rect 9715 188 9727 222
rect 9907 188 9919 222
rect 10099 188 10111 222
rect 10291 188 10303 222
rect 10483 188 10495 222
rect 10675 188 10687 222
rect 10867 188 10879 222
rect 11059 188 11071 222
rect 11251 188 11263 222
rect 11443 188 11455 222
rect 11635 188 11647 222
rect 11827 188 11839 222
rect 12019 188 12031 222
rect 12211 188 12223 222
rect 12403 188 12415 222
rect 12595 188 12607 222
rect 12787 188 12799 222
rect 12979 188 12991 222
rect 13171 188 13183 222
rect 13363 188 13375 222
rect 13555 188 13567 222
rect 13747 188 13759 222
rect 13939 188 13951 222
rect 14131 188 14143 222
rect 14323 188 14335 222
rect 14515 188 14527 222
rect 14707 188 14719 222
rect 14899 188 14911 222
rect 15091 188 15103 222
rect 15283 188 15295 222
rect 15475 188 15487 222
rect 15667 188 15679 222
rect 15859 188 15871 222
rect 16051 188 16063 222
rect 16243 188 16255 222
rect 16435 188 16447 222
rect 16627 188 16639 222
rect 16819 188 16831 222
rect 17011 188 17023 222
rect 17203 188 17215 222
rect 17395 188 17407 222
rect 17587 188 17599 222
rect 17779 188 17791 222
rect 17971 188 17983 222
rect 18163 188 18175 222
rect 18355 188 18367 222
rect 18547 188 18559 222
rect 18739 188 18751 222
rect 18931 188 18943 222
rect 19123 188 19135 222
rect -19085 182 -19027 188
rect -18893 182 -18835 188
rect -18701 182 -18643 188
rect -18509 182 -18451 188
rect -18317 182 -18259 188
rect -18125 182 -18067 188
rect -17933 182 -17875 188
rect -17741 182 -17683 188
rect -17549 182 -17491 188
rect -17357 182 -17299 188
rect -17165 182 -17107 188
rect -16973 182 -16915 188
rect -16781 182 -16723 188
rect -16589 182 -16531 188
rect -16397 182 -16339 188
rect -16205 182 -16147 188
rect -16013 182 -15955 188
rect -15821 182 -15763 188
rect -15629 182 -15571 188
rect -15437 182 -15379 188
rect -15245 182 -15187 188
rect -15053 182 -14995 188
rect -14861 182 -14803 188
rect -14669 182 -14611 188
rect -14477 182 -14419 188
rect -14285 182 -14227 188
rect -14093 182 -14035 188
rect -13901 182 -13843 188
rect -13709 182 -13651 188
rect -13517 182 -13459 188
rect -13325 182 -13267 188
rect -13133 182 -13075 188
rect -12941 182 -12883 188
rect -12749 182 -12691 188
rect -12557 182 -12499 188
rect -12365 182 -12307 188
rect -12173 182 -12115 188
rect -11981 182 -11923 188
rect -11789 182 -11731 188
rect -11597 182 -11539 188
rect -11405 182 -11347 188
rect -11213 182 -11155 188
rect -11021 182 -10963 188
rect -10829 182 -10771 188
rect -10637 182 -10579 188
rect -10445 182 -10387 188
rect -10253 182 -10195 188
rect -10061 182 -10003 188
rect -9869 182 -9811 188
rect -9677 182 -9619 188
rect -9485 182 -9427 188
rect -9293 182 -9235 188
rect -9101 182 -9043 188
rect -8909 182 -8851 188
rect -8717 182 -8659 188
rect -8525 182 -8467 188
rect -8333 182 -8275 188
rect -8141 182 -8083 188
rect -7949 182 -7891 188
rect -7757 182 -7699 188
rect -7565 182 -7507 188
rect -7373 182 -7315 188
rect -7181 182 -7123 188
rect -6989 182 -6931 188
rect -6797 182 -6739 188
rect -6605 182 -6547 188
rect -6413 182 -6355 188
rect -6221 182 -6163 188
rect -6029 182 -5971 188
rect -5837 182 -5779 188
rect -5645 182 -5587 188
rect -5453 182 -5395 188
rect -5261 182 -5203 188
rect -5069 182 -5011 188
rect -4877 182 -4819 188
rect -4685 182 -4627 188
rect -4493 182 -4435 188
rect -4301 182 -4243 188
rect -4109 182 -4051 188
rect -3917 182 -3859 188
rect -3725 182 -3667 188
rect -3533 182 -3475 188
rect -3341 182 -3283 188
rect -3149 182 -3091 188
rect -2957 182 -2899 188
rect -2765 182 -2707 188
rect -2573 182 -2515 188
rect -2381 182 -2323 188
rect -2189 182 -2131 188
rect -1997 182 -1939 188
rect -1805 182 -1747 188
rect -1613 182 -1555 188
rect -1421 182 -1363 188
rect -1229 182 -1171 188
rect -1037 182 -979 188
rect -845 182 -787 188
rect -653 182 -595 188
rect -461 182 -403 188
rect -269 182 -211 188
rect -77 182 -19 188
rect 115 182 173 188
rect 307 182 365 188
rect 499 182 557 188
rect 691 182 749 188
rect 883 182 941 188
rect 1075 182 1133 188
rect 1267 182 1325 188
rect 1459 182 1517 188
rect 1651 182 1709 188
rect 1843 182 1901 188
rect 2035 182 2093 188
rect 2227 182 2285 188
rect 2419 182 2477 188
rect 2611 182 2669 188
rect 2803 182 2861 188
rect 2995 182 3053 188
rect 3187 182 3245 188
rect 3379 182 3437 188
rect 3571 182 3629 188
rect 3763 182 3821 188
rect 3955 182 4013 188
rect 4147 182 4205 188
rect 4339 182 4397 188
rect 4531 182 4589 188
rect 4723 182 4781 188
rect 4915 182 4973 188
rect 5107 182 5165 188
rect 5299 182 5357 188
rect 5491 182 5549 188
rect 5683 182 5741 188
rect 5875 182 5933 188
rect 6067 182 6125 188
rect 6259 182 6317 188
rect 6451 182 6509 188
rect 6643 182 6701 188
rect 6835 182 6893 188
rect 7027 182 7085 188
rect 7219 182 7277 188
rect 7411 182 7469 188
rect 7603 182 7661 188
rect 7795 182 7853 188
rect 7987 182 8045 188
rect 8179 182 8237 188
rect 8371 182 8429 188
rect 8563 182 8621 188
rect 8755 182 8813 188
rect 8947 182 9005 188
rect 9139 182 9197 188
rect 9331 182 9389 188
rect 9523 182 9581 188
rect 9715 182 9773 188
rect 9907 182 9965 188
rect 10099 182 10157 188
rect 10291 182 10349 188
rect 10483 182 10541 188
rect 10675 182 10733 188
rect 10867 182 10925 188
rect 11059 182 11117 188
rect 11251 182 11309 188
rect 11443 182 11501 188
rect 11635 182 11693 188
rect 11827 182 11885 188
rect 12019 182 12077 188
rect 12211 182 12269 188
rect 12403 182 12461 188
rect 12595 182 12653 188
rect 12787 182 12845 188
rect 12979 182 13037 188
rect 13171 182 13229 188
rect 13363 182 13421 188
rect 13555 182 13613 188
rect 13747 182 13805 188
rect 13939 182 13997 188
rect 14131 182 14189 188
rect 14323 182 14381 188
rect 14515 182 14573 188
rect 14707 182 14765 188
rect 14899 182 14957 188
rect 15091 182 15149 188
rect 15283 182 15341 188
rect 15475 182 15533 188
rect 15667 182 15725 188
rect 15859 182 15917 188
rect 16051 182 16109 188
rect 16243 182 16301 188
rect 16435 182 16493 188
rect 16627 182 16685 188
rect 16819 182 16877 188
rect 17011 182 17069 188
rect 17203 182 17261 188
rect 17395 182 17453 188
rect 17587 182 17645 188
rect 17779 182 17837 188
rect 17971 182 18029 188
rect 18163 182 18221 188
rect 18355 182 18413 188
rect 18547 182 18605 188
rect 18739 182 18797 188
rect 18931 182 18989 188
rect 19123 182 19181 188
rect -19181 -188 -19123 -182
rect -18989 -188 -18931 -182
rect -18797 -188 -18739 -182
rect -18605 -188 -18547 -182
rect -18413 -188 -18355 -182
rect -18221 -188 -18163 -182
rect -18029 -188 -17971 -182
rect -17837 -188 -17779 -182
rect -17645 -188 -17587 -182
rect -17453 -188 -17395 -182
rect -17261 -188 -17203 -182
rect -17069 -188 -17011 -182
rect -16877 -188 -16819 -182
rect -16685 -188 -16627 -182
rect -16493 -188 -16435 -182
rect -16301 -188 -16243 -182
rect -16109 -188 -16051 -182
rect -15917 -188 -15859 -182
rect -15725 -188 -15667 -182
rect -15533 -188 -15475 -182
rect -15341 -188 -15283 -182
rect -15149 -188 -15091 -182
rect -14957 -188 -14899 -182
rect -14765 -188 -14707 -182
rect -14573 -188 -14515 -182
rect -14381 -188 -14323 -182
rect -14189 -188 -14131 -182
rect -13997 -188 -13939 -182
rect -13805 -188 -13747 -182
rect -13613 -188 -13555 -182
rect -13421 -188 -13363 -182
rect -13229 -188 -13171 -182
rect -13037 -188 -12979 -182
rect -12845 -188 -12787 -182
rect -12653 -188 -12595 -182
rect -12461 -188 -12403 -182
rect -12269 -188 -12211 -182
rect -12077 -188 -12019 -182
rect -11885 -188 -11827 -182
rect -11693 -188 -11635 -182
rect -11501 -188 -11443 -182
rect -11309 -188 -11251 -182
rect -11117 -188 -11059 -182
rect -10925 -188 -10867 -182
rect -10733 -188 -10675 -182
rect -10541 -188 -10483 -182
rect -10349 -188 -10291 -182
rect -10157 -188 -10099 -182
rect -9965 -188 -9907 -182
rect -9773 -188 -9715 -182
rect -9581 -188 -9523 -182
rect -9389 -188 -9331 -182
rect -9197 -188 -9139 -182
rect -9005 -188 -8947 -182
rect -8813 -188 -8755 -182
rect -8621 -188 -8563 -182
rect -8429 -188 -8371 -182
rect -8237 -188 -8179 -182
rect -8045 -188 -7987 -182
rect -7853 -188 -7795 -182
rect -7661 -188 -7603 -182
rect -7469 -188 -7411 -182
rect -7277 -188 -7219 -182
rect -7085 -188 -7027 -182
rect -6893 -188 -6835 -182
rect -6701 -188 -6643 -182
rect -6509 -188 -6451 -182
rect -6317 -188 -6259 -182
rect -6125 -188 -6067 -182
rect -5933 -188 -5875 -182
rect -5741 -188 -5683 -182
rect -5549 -188 -5491 -182
rect -5357 -188 -5299 -182
rect -5165 -188 -5107 -182
rect -4973 -188 -4915 -182
rect -4781 -188 -4723 -182
rect -4589 -188 -4531 -182
rect -4397 -188 -4339 -182
rect -4205 -188 -4147 -182
rect -4013 -188 -3955 -182
rect -3821 -188 -3763 -182
rect -3629 -188 -3571 -182
rect -3437 -188 -3379 -182
rect -3245 -188 -3187 -182
rect -3053 -188 -2995 -182
rect -2861 -188 -2803 -182
rect -2669 -188 -2611 -182
rect -2477 -188 -2419 -182
rect -2285 -188 -2227 -182
rect -2093 -188 -2035 -182
rect -1901 -188 -1843 -182
rect -1709 -188 -1651 -182
rect -1517 -188 -1459 -182
rect -1325 -188 -1267 -182
rect -1133 -188 -1075 -182
rect -941 -188 -883 -182
rect -749 -188 -691 -182
rect -557 -188 -499 -182
rect -365 -188 -307 -182
rect -173 -188 -115 -182
rect 19 -188 77 -182
rect 211 -188 269 -182
rect 403 -188 461 -182
rect 595 -188 653 -182
rect 787 -188 845 -182
rect 979 -188 1037 -182
rect 1171 -188 1229 -182
rect 1363 -188 1421 -182
rect 1555 -188 1613 -182
rect 1747 -188 1805 -182
rect 1939 -188 1997 -182
rect 2131 -188 2189 -182
rect 2323 -188 2381 -182
rect 2515 -188 2573 -182
rect 2707 -188 2765 -182
rect 2899 -188 2957 -182
rect 3091 -188 3149 -182
rect 3283 -188 3341 -182
rect 3475 -188 3533 -182
rect 3667 -188 3725 -182
rect 3859 -188 3917 -182
rect 4051 -188 4109 -182
rect 4243 -188 4301 -182
rect 4435 -188 4493 -182
rect 4627 -188 4685 -182
rect 4819 -188 4877 -182
rect 5011 -188 5069 -182
rect 5203 -188 5261 -182
rect 5395 -188 5453 -182
rect 5587 -188 5645 -182
rect 5779 -188 5837 -182
rect 5971 -188 6029 -182
rect 6163 -188 6221 -182
rect 6355 -188 6413 -182
rect 6547 -188 6605 -182
rect 6739 -188 6797 -182
rect 6931 -188 6989 -182
rect 7123 -188 7181 -182
rect 7315 -188 7373 -182
rect 7507 -188 7565 -182
rect 7699 -188 7757 -182
rect 7891 -188 7949 -182
rect 8083 -188 8141 -182
rect 8275 -188 8333 -182
rect 8467 -188 8525 -182
rect 8659 -188 8717 -182
rect 8851 -188 8909 -182
rect 9043 -188 9101 -182
rect 9235 -188 9293 -182
rect 9427 -188 9485 -182
rect 9619 -188 9677 -182
rect 9811 -188 9869 -182
rect 10003 -188 10061 -182
rect 10195 -188 10253 -182
rect 10387 -188 10445 -182
rect 10579 -188 10637 -182
rect 10771 -188 10829 -182
rect 10963 -188 11021 -182
rect 11155 -188 11213 -182
rect 11347 -188 11405 -182
rect 11539 -188 11597 -182
rect 11731 -188 11789 -182
rect 11923 -188 11981 -182
rect 12115 -188 12173 -182
rect 12307 -188 12365 -182
rect 12499 -188 12557 -182
rect 12691 -188 12749 -182
rect 12883 -188 12941 -182
rect 13075 -188 13133 -182
rect 13267 -188 13325 -182
rect 13459 -188 13517 -182
rect 13651 -188 13709 -182
rect 13843 -188 13901 -182
rect 14035 -188 14093 -182
rect 14227 -188 14285 -182
rect 14419 -188 14477 -182
rect 14611 -188 14669 -182
rect 14803 -188 14861 -182
rect 14995 -188 15053 -182
rect 15187 -188 15245 -182
rect 15379 -188 15437 -182
rect 15571 -188 15629 -182
rect 15763 -188 15821 -182
rect 15955 -188 16013 -182
rect 16147 -188 16205 -182
rect 16339 -188 16397 -182
rect 16531 -188 16589 -182
rect 16723 -188 16781 -182
rect 16915 -188 16973 -182
rect 17107 -188 17165 -182
rect 17299 -188 17357 -182
rect 17491 -188 17549 -182
rect 17683 -188 17741 -182
rect 17875 -188 17933 -182
rect 18067 -188 18125 -182
rect 18259 -188 18317 -182
rect 18451 -188 18509 -182
rect 18643 -188 18701 -182
rect 18835 -188 18893 -182
rect 19027 -188 19085 -182
rect -19181 -222 -19169 -188
rect -18989 -222 -18977 -188
rect -18797 -222 -18785 -188
rect -18605 -222 -18593 -188
rect -18413 -222 -18401 -188
rect -18221 -222 -18209 -188
rect -18029 -222 -18017 -188
rect -17837 -222 -17825 -188
rect -17645 -222 -17633 -188
rect -17453 -222 -17441 -188
rect -17261 -222 -17249 -188
rect -17069 -222 -17057 -188
rect -16877 -222 -16865 -188
rect -16685 -222 -16673 -188
rect -16493 -222 -16481 -188
rect -16301 -222 -16289 -188
rect -16109 -222 -16097 -188
rect -15917 -222 -15905 -188
rect -15725 -222 -15713 -188
rect -15533 -222 -15521 -188
rect -15341 -222 -15329 -188
rect -15149 -222 -15137 -188
rect -14957 -222 -14945 -188
rect -14765 -222 -14753 -188
rect -14573 -222 -14561 -188
rect -14381 -222 -14369 -188
rect -14189 -222 -14177 -188
rect -13997 -222 -13985 -188
rect -13805 -222 -13793 -188
rect -13613 -222 -13601 -188
rect -13421 -222 -13409 -188
rect -13229 -222 -13217 -188
rect -13037 -222 -13025 -188
rect -12845 -222 -12833 -188
rect -12653 -222 -12641 -188
rect -12461 -222 -12449 -188
rect -12269 -222 -12257 -188
rect -12077 -222 -12065 -188
rect -11885 -222 -11873 -188
rect -11693 -222 -11681 -188
rect -11501 -222 -11489 -188
rect -11309 -222 -11297 -188
rect -11117 -222 -11105 -188
rect -10925 -222 -10913 -188
rect -10733 -222 -10721 -188
rect -10541 -222 -10529 -188
rect -10349 -222 -10337 -188
rect -10157 -222 -10145 -188
rect -9965 -222 -9953 -188
rect -9773 -222 -9761 -188
rect -9581 -222 -9569 -188
rect -9389 -222 -9377 -188
rect -9197 -222 -9185 -188
rect -9005 -222 -8993 -188
rect -8813 -222 -8801 -188
rect -8621 -222 -8609 -188
rect -8429 -222 -8417 -188
rect -8237 -222 -8225 -188
rect -8045 -222 -8033 -188
rect -7853 -222 -7841 -188
rect -7661 -222 -7649 -188
rect -7469 -222 -7457 -188
rect -7277 -222 -7265 -188
rect -7085 -222 -7073 -188
rect -6893 -222 -6881 -188
rect -6701 -222 -6689 -188
rect -6509 -222 -6497 -188
rect -6317 -222 -6305 -188
rect -6125 -222 -6113 -188
rect -5933 -222 -5921 -188
rect -5741 -222 -5729 -188
rect -5549 -222 -5537 -188
rect -5357 -222 -5345 -188
rect -5165 -222 -5153 -188
rect -4973 -222 -4961 -188
rect -4781 -222 -4769 -188
rect -4589 -222 -4577 -188
rect -4397 -222 -4385 -188
rect -4205 -222 -4193 -188
rect -4013 -222 -4001 -188
rect -3821 -222 -3809 -188
rect -3629 -222 -3617 -188
rect -3437 -222 -3425 -188
rect -3245 -222 -3233 -188
rect -3053 -222 -3041 -188
rect -2861 -222 -2849 -188
rect -2669 -222 -2657 -188
rect -2477 -222 -2465 -188
rect -2285 -222 -2273 -188
rect -2093 -222 -2081 -188
rect -1901 -222 -1889 -188
rect -1709 -222 -1697 -188
rect -1517 -222 -1505 -188
rect -1325 -222 -1313 -188
rect -1133 -222 -1121 -188
rect -941 -222 -929 -188
rect -749 -222 -737 -188
rect -557 -222 -545 -188
rect -365 -222 -353 -188
rect -173 -222 -161 -188
rect 19 -222 31 -188
rect 211 -222 223 -188
rect 403 -222 415 -188
rect 595 -222 607 -188
rect 787 -222 799 -188
rect 979 -222 991 -188
rect 1171 -222 1183 -188
rect 1363 -222 1375 -188
rect 1555 -222 1567 -188
rect 1747 -222 1759 -188
rect 1939 -222 1951 -188
rect 2131 -222 2143 -188
rect 2323 -222 2335 -188
rect 2515 -222 2527 -188
rect 2707 -222 2719 -188
rect 2899 -222 2911 -188
rect 3091 -222 3103 -188
rect 3283 -222 3295 -188
rect 3475 -222 3487 -188
rect 3667 -222 3679 -188
rect 3859 -222 3871 -188
rect 4051 -222 4063 -188
rect 4243 -222 4255 -188
rect 4435 -222 4447 -188
rect 4627 -222 4639 -188
rect 4819 -222 4831 -188
rect 5011 -222 5023 -188
rect 5203 -222 5215 -188
rect 5395 -222 5407 -188
rect 5587 -222 5599 -188
rect 5779 -222 5791 -188
rect 5971 -222 5983 -188
rect 6163 -222 6175 -188
rect 6355 -222 6367 -188
rect 6547 -222 6559 -188
rect 6739 -222 6751 -188
rect 6931 -222 6943 -188
rect 7123 -222 7135 -188
rect 7315 -222 7327 -188
rect 7507 -222 7519 -188
rect 7699 -222 7711 -188
rect 7891 -222 7903 -188
rect 8083 -222 8095 -188
rect 8275 -222 8287 -188
rect 8467 -222 8479 -188
rect 8659 -222 8671 -188
rect 8851 -222 8863 -188
rect 9043 -222 9055 -188
rect 9235 -222 9247 -188
rect 9427 -222 9439 -188
rect 9619 -222 9631 -188
rect 9811 -222 9823 -188
rect 10003 -222 10015 -188
rect 10195 -222 10207 -188
rect 10387 -222 10399 -188
rect 10579 -222 10591 -188
rect 10771 -222 10783 -188
rect 10963 -222 10975 -188
rect 11155 -222 11167 -188
rect 11347 -222 11359 -188
rect 11539 -222 11551 -188
rect 11731 -222 11743 -188
rect 11923 -222 11935 -188
rect 12115 -222 12127 -188
rect 12307 -222 12319 -188
rect 12499 -222 12511 -188
rect 12691 -222 12703 -188
rect 12883 -222 12895 -188
rect 13075 -222 13087 -188
rect 13267 -222 13279 -188
rect 13459 -222 13471 -188
rect 13651 -222 13663 -188
rect 13843 -222 13855 -188
rect 14035 -222 14047 -188
rect 14227 -222 14239 -188
rect 14419 -222 14431 -188
rect 14611 -222 14623 -188
rect 14803 -222 14815 -188
rect 14995 -222 15007 -188
rect 15187 -222 15199 -188
rect 15379 -222 15391 -188
rect 15571 -222 15583 -188
rect 15763 -222 15775 -188
rect 15955 -222 15967 -188
rect 16147 -222 16159 -188
rect 16339 -222 16351 -188
rect 16531 -222 16543 -188
rect 16723 -222 16735 -188
rect 16915 -222 16927 -188
rect 17107 -222 17119 -188
rect 17299 -222 17311 -188
rect 17491 -222 17503 -188
rect 17683 -222 17695 -188
rect 17875 -222 17887 -188
rect 18067 -222 18079 -188
rect 18259 -222 18271 -188
rect 18451 -222 18463 -188
rect 18643 -222 18655 -188
rect 18835 -222 18847 -188
rect 19027 -222 19039 -188
rect -19181 -228 -19123 -222
rect -18989 -228 -18931 -222
rect -18797 -228 -18739 -222
rect -18605 -228 -18547 -222
rect -18413 -228 -18355 -222
rect -18221 -228 -18163 -222
rect -18029 -228 -17971 -222
rect -17837 -228 -17779 -222
rect -17645 -228 -17587 -222
rect -17453 -228 -17395 -222
rect -17261 -228 -17203 -222
rect -17069 -228 -17011 -222
rect -16877 -228 -16819 -222
rect -16685 -228 -16627 -222
rect -16493 -228 -16435 -222
rect -16301 -228 -16243 -222
rect -16109 -228 -16051 -222
rect -15917 -228 -15859 -222
rect -15725 -228 -15667 -222
rect -15533 -228 -15475 -222
rect -15341 -228 -15283 -222
rect -15149 -228 -15091 -222
rect -14957 -228 -14899 -222
rect -14765 -228 -14707 -222
rect -14573 -228 -14515 -222
rect -14381 -228 -14323 -222
rect -14189 -228 -14131 -222
rect -13997 -228 -13939 -222
rect -13805 -228 -13747 -222
rect -13613 -228 -13555 -222
rect -13421 -228 -13363 -222
rect -13229 -228 -13171 -222
rect -13037 -228 -12979 -222
rect -12845 -228 -12787 -222
rect -12653 -228 -12595 -222
rect -12461 -228 -12403 -222
rect -12269 -228 -12211 -222
rect -12077 -228 -12019 -222
rect -11885 -228 -11827 -222
rect -11693 -228 -11635 -222
rect -11501 -228 -11443 -222
rect -11309 -228 -11251 -222
rect -11117 -228 -11059 -222
rect -10925 -228 -10867 -222
rect -10733 -228 -10675 -222
rect -10541 -228 -10483 -222
rect -10349 -228 -10291 -222
rect -10157 -228 -10099 -222
rect -9965 -228 -9907 -222
rect -9773 -228 -9715 -222
rect -9581 -228 -9523 -222
rect -9389 -228 -9331 -222
rect -9197 -228 -9139 -222
rect -9005 -228 -8947 -222
rect -8813 -228 -8755 -222
rect -8621 -228 -8563 -222
rect -8429 -228 -8371 -222
rect -8237 -228 -8179 -222
rect -8045 -228 -7987 -222
rect -7853 -228 -7795 -222
rect -7661 -228 -7603 -222
rect -7469 -228 -7411 -222
rect -7277 -228 -7219 -222
rect -7085 -228 -7027 -222
rect -6893 -228 -6835 -222
rect -6701 -228 -6643 -222
rect -6509 -228 -6451 -222
rect -6317 -228 -6259 -222
rect -6125 -228 -6067 -222
rect -5933 -228 -5875 -222
rect -5741 -228 -5683 -222
rect -5549 -228 -5491 -222
rect -5357 -228 -5299 -222
rect -5165 -228 -5107 -222
rect -4973 -228 -4915 -222
rect -4781 -228 -4723 -222
rect -4589 -228 -4531 -222
rect -4397 -228 -4339 -222
rect -4205 -228 -4147 -222
rect -4013 -228 -3955 -222
rect -3821 -228 -3763 -222
rect -3629 -228 -3571 -222
rect -3437 -228 -3379 -222
rect -3245 -228 -3187 -222
rect -3053 -228 -2995 -222
rect -2861 -228 -2803 -222
rect -2669 -228 -2611 -222
rect -2477 -228 -2419 -222
rect -2285 -228 -2227 -222
rect -2093 -228 -2035 -222
rect -1901 -228 -1843 -222
rect -1709 -228 -1651 -222
rect -1517 -228 -1459 -222
rect -1325 -228 -1267 -222
rect -1133 -228 -1075 -222
rect -941 -228 -883 -222
rect -749 -228 -691 -222
rect -557 -228 -499 -222
rect -365 -228 -307 -222
rect -173 -228 -115 -222
rect 19 -228 77 -222
rect 211 -228 269 -222
rect 403 -228 461 -222
rect 595 -228 653 -222
rect 787 -228 845 -222
rect 979 -228 1037 -222
rect 1171 -228 1229 -222
rect 1363 -228 1421 -222
rect 1555 -228 1613 -222
rect 1747 -228 1805 -222
rect 1939 -228 1997 -222
rect 2131 -228 2189 -222
rect 2323 -228 2381 -222
rect 2515 -228 2573 -222
rect 2707 -228 2765 -222
rect 2899 -228 2957 -222
rect 3091 -228 3149 -222
rect 3283 -228 3341 -222
rect 3475 -228 3533 -222
rect 3667 -228 3725 -222
rect 3859 -228 3917 -222
rect 4051 -228 4109 -222
rect 4243 -228 4301 -222
rect 4435 -228 4493 -222
rect 4627 -228 4685 -222
rect 4819 -228 4877 -222
rect 5011 -228 5069 -222
rect 5203 -228 5261 -222
rect 5395 -228 5453 -222
rect 5587 -228 5645 -222
rect 5779 -228 5837 -222
rect 5971 -228 6029 -222
rect 6163 -228 6221 -222
rect 6355 -228 6413 -222
rect 6547 -228 6605 -222
rect 6739 -228 6797 -222
rect 6931 -228 6989 -222
rect 7123 -228 7181 -222
rect 7315 -228 7373 -222
rect 7507 -228 7565 -222
rect 7699 -228 7757 -222
rect 7891 -228 7949 -222
rect 8083 -228 8141 -222
rect 8275 -228 8333 -222
rect 8467 -228 8525 -222
rect 8659 -228 8717 -222
rect 8851 -228 8909 -222
rect 9043 -228 9101 -222
rect 9235 -228 9293 -222
rect 9427 -228 9485 -222
rect 9619 -228 9677 -222
rect 9811 -228 9869 -222
rect 10003 -228 10061 -222
rect 10195 -228 10253 -222
rect 10387 -228 10445 -222
rect 10579 -228 10637 -222
rect 10771 -228 10829 -222
rect 10963 -228 11021 -222
rect 11155 -228 11213 -222
rect 11347 -228 11405 -222
rect 11539 -228 11597 -222
rect 11731 -228 11789 -222
rect 11923 -228 11981 -222
rect 12115 -228 12173 -222
rect 12307 -228 12365 -222
rect 12499 -228 12557 -222
rect 12691 -228 12749 -222
rect 12883 -228 12941 -222
rect 13075 -228 13133 -222
rect 13267 -228 13325 -222
rect 13459 -228 13517 -222
rect 13651 -228 13709 -222
rect 13843 -228 13901 -222
rect 14035 -228 14093 -222
rect 14227 -228 14285 -222
rect 14419 -228 14477 -222
rect 14611 -228 14669 -222
rect 14803 -228 14861 -222
rect 14995 -228 15053 -222
rect 15187 -228 15245 -222
rect 15379 -228 15437 -222
rect 15571 -228 15629 -222
rect 15763 -228 15821 -222
rect 15955 -228 16013 -222
rect 16147 -228 16205 -222
rect 16339 -228 16397 -222
rect 16531 -228 16589 -222
rect 16723 -228 16781 -222
rect 16915 -228 16973 -222
rect 17107 -228 17165 -222
rect 17299 -228 17357 -222
rect 17491 -228 17549 -222
rect 17683 -228 17741 -222
rect 17875 -228 17933 -222
rect 18067 -228 18125 -222
rect 18259 -228 18317 -222
rect 18451 -228 18509 -222
rect 18643 -228 18701 -222
rect 18835 -228 18893 -222
rect 19027 -228 19085 -222
<< pwell >>
rect -19367 -360 19367 360
<< nmos >>
rect -19167 -150 -19137 150
rect -19071 -150 -19041 150
rect -18975 -150 -18945 150
rect -18879 -150 -18849 150
rect -18783 -150 -18753 150
rect -18687 -150 -18657 150
rect -18591 -150 -18561 150
rect -18495 -150 -18465 150
rect -18399 -150 -18369 150
rect -18303 -150 -18273 150
rect -18207 -150 -18177 150
rect -18111 -150 -18081 150
rect -18015 -150 -17985 150
rect -17919 -150 -17889 150
rect -17823 -150 -17793 150
rect -17727 -150 -17697 150
rect -17631 -150 -17601 150
rect -17535 -150 -17505 150
rect -17439 -150 -17409 150
rect -17343 -150 -17313 150
rect -17247 -150 -17217 150
rect -17151 -150 -17121 150
rect -17055 -150 -17025 150
rect -16959 -150 -16929 150
rect -16863 -150 -16833 150
rect -16767 -150 -16737 150
rect -16671 -150 -16641 150
rect -16575 -150 -16545 150
rect -16479 -150 -16449 150
rect -16383 -150 -16353 150
rect -16287 -150 -16257 150
rect -16191 -150 -16161 150
rect -16095 -150 -16065 150
rect -15999 -150 -15969 150
rect -15903 -150 -15873 150
rect -15807 -150 -15777 150
rect -15711 -150 -15681 150
rect -15615 -150 -15585 150
rect -15519 -150 -15489 150
rect -15423 -150 -15393 150
rect -15327 -150 -15297 150
rect -15231 -150 -15201 150
rect -15135 -150 -15105 150
rect -15039 -150 -15009 150
rect -14943 -150 -14913 150
rect -14847 -150 -14817 150
rect -14751 -150 -14721 150
rect -14655 -150 -14625 150
rect -14559 -150 -14529 150
rect -14463 -150 -14433 150
rect -14367 -150 -14337 150
rect -14271 -150 -14241 150
rect -14175 -150 -14145 150
rect -14079 -150 -14049 150
rect -13983 -150 -13953 150
rect -13887 -150 -13857 150
rect -13791 -150 -13761 150
rect -13695 -150 -13665 150
rect -13599 -150 -13569 150
rect -13503 -150 -13473 150
rect -13407 -150 -13377 150
rect -13311 -150 -13281 150
rect -13215 -150 -13185 150
rect -13119 -150 -13089 150
rect -13023 -150 -12993 150
rect -12927 -150 -12897 150
rect -12831 -150 -12801 150
rect -12735 -150 -12705 150
rect -12639 -150 -12609 150
rect -12543 -150 -12513 150
rect -12447 -150 -12417 150
rect -12351 -150 -12321 150
rect -12255 -150 -12225 150
rect -12159 -150 -12129 150
rect -12063 -150 -12033 150
rect -11967 -150 -11937 150
rect -11871 -150 -11841 150
rect -11775 -150 -11745 150
rect -11679 -150 -11649 150
rect -11583 -150 -11553 150
rect -11487 -150 -11457 150
rect -11391 -150 -11361 150
rect -11295 -150 -11265 150
rect -11199 -150 -11169 150
rect -11103 -150 -11073 150
rect -11007 -150 -10977 150
rect -10911 -150 -10881 150
rect -10815 -150 -10785 150
rect -10719 -150 -10689 150
rect -10623 -150 -10593 150
rect -10527 -150 -10497 150
rect -10431 -150 -10401 150
rect -10335 -150 -10305 150
rect -10239 -150 -10209 150
rect -10143 -150 -10113 150
rect -10047 -150 -10017 150
rect -9951 -150 -9921 150
rect -9855 -150 -9825 150
rect -9759 -150 -9729 150
rect -9663 -150 -9633 150
rect -9567 -150 -9537 150
rect -9471 -150 -9441 150
rect -9375 -150 -9345 150
rect -9279 -150 -9249 150
rect -9183 -150 -9153 150
rect -9087 -150 -9057 150
rect -8991 -150 -8961 150
rect -8895 -150 -8865 150
rect -8799 -150 -8769 150
rect -8703 -150 -8673 150
rect -8607 -150 -8577 150
rect -8511 -150 -8481 150
rect -8415 -150 -8385 150
rect -8319 -150 -8289 150
rect -8223 -150 -8193 150
rect -8127 -150 -8097 150
rect -8031 -150 -8001 150
rect -7935 -150 -7905 150
rect -7839 -150 -7809 150
rect -7743 -150 -7713 150
rect -7647 -150 -7617 150
rect -7551 -150 -7521 150
rect -7455 -150 -7425 150
rect -7359 -150 -7329 150
rect -7263 -150 -7233 150
rect -7167 -150 -7137 150
rect -7071 -150 -7041 150
rect -6975 -150 -6945 150
rect -6879 -150 -6849 150
rect -6783 -150 -6753 150
rect -6687 -150 -6657 150
rect -6591 -150 -6561 150
rect -6495 -150 -6465 150
rect -6399 -150 -6369 150
rect -6303 -150 -6273 150
rect -6207 -150 -6177 150
rect -6111 -150 -6081 150
rect -6015 -150 -5985 150
rect -5919 -150 -5889 150
rect -5823 -150 -5793 150
rect -5727 -150 -5697 150
rect -5631 -150 -5601 150
rect -5535 -150 -5505 150
rect -5439 -150 -5409 150
rect -5343 -150 -5313 150
rect -5247 -150 -5217 150
rect -5151 -150 -5121 150
rect -5055 -150 -5025 150
rect -4959 -150 -4929 150
rect -4863 -150 -4833 150
rect -4767 -150 -4737 150
rect -4671 -150 -4641 150
rect -4575 -150 -4545 150
rect -4479 -150 -4449 150
rect -4383 -150 -4353 150
rect -4287 -150 -4257 150
rect -4191 -150 -4161 150
rect -4095 -150 -4065 150
rect -3999 -150 -3969 150
rect -3903 -150 -3873 150
rect -3807 -150 -3777 150
rect -3711 -150 -3681 150
rect -3615 -150 -3585 150
rect -3519 -150 -3489 150
rect -3423 -150 -3393 150
rect -3327 -150 -3297 150
rect -3231 -150 -3201 150
rect -3135 -150 -3105 150
rect -3039 -150 -3009 150
rect -2943 -150 -2913 150
rect -2847 -150 -2817 150
rect -2751 -150 -2721 150
rect -2655 -150 -2625 150
rect -2559 -150 -2529 150
rect -2463 -150 -2433 150
rect -2367 -150 -2337 150
rect -2271 -150 -2241 150
rect -2175 -150 -2145 150
rect -2079 -150 -2049 150
rect -1983 -150 -1953 150
rect -1887 -150 -1857 150
rect -1791 -150 -1761 150
rect -1695 -150 -1665 150
rect -1599 -150 -1569 150
rect -1503 -150 -1473 150
rect -1407 -150 -1377 150
rect -1311 -150 -1281 150
rect -1215 -150 -1185 150
rect -1119 -150 -1089 150
rect -1023 -150 -993 150
rect -927 -150 -897 150
rect -831 -150 -801 150
rect -735 -150 -705 150
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
rect 705 -150 735 150
rect 801 -150 831 150
rect 897 -150 927 150
rect 993 -150 1023 150
rect 1089 -150 1119 150
rect 1185 -150 1215 150
rect 1281 -150 1311 150
rect 1377 -150 1407 150
rect 1473 -150 1503 150
rect 1569 -150 1599 150
rect 1665 -150 1695 150
rect 1761 -150 1791 150
rect 1857 -150 1887 150
rect 1953 -150 1983 150
rect 2049 -150 2079 150
rect 2145 -150 2175 150
rect 2241 -150 2271 150
rect 2337 -150 2367 150
rect 2433 -150 2463 150
rect 2529 -150 2559 150
rect 2625 -150 2655 150
rect 2721 -150 2751 150
rect 2817 -150 2847 150
rect 2913 -150 2943 150
rect 3009 -150 3039 150
rect 3105 -150 3135 150
rect 3201 -150 3231 150
rect 3297 -150 3327 150
rect 3393 -150 3423 150
rect 3489 -150 3519 150
rect 3585 -150 3615 150
rect 3681 -150 3711 150
rect 3777 -150 3807 150
rect 3873 -150 3903 150
rect 3969 -150 3999 150
rect 4065 -150 4095 150
rect 4161 -150 4191 150
rect 4257 -150 4287 150
rect 4353 -150 4383 150
rect 4449 -150 4479 150
rect 4545 -150 4575 150
rect 4641 -150 4671 150
rect 4737 -150 4767 150
rect 4833 -150 4863 150
rect 4929 -150 4959 150
rect 5025 -150 5055 150
rect 5121 -150 5151 150
rect 5217 -150 5247 150
rect 5313 -150 5343 150
rect 5409 -150 5439 150
rect 5505 -150 5535 150
rect 5601 -150 5631 150
rect 5697 -150 5727 150
rect 5793 -150 5823 150
rect 5889 -150 5919 150
rect 5985 -150 6015 150
rect 6081 -150 6111 150
rect 6177 -150 6207 150
rect 6273 -150 6303 150
rect 6369 -150 6399 150
rect 6465 -150 6495 150
rect 6561 -150 6591 150
rect 6657 -150 6687 150
rect 6753 -150 6783 150
rect 6849 -150 6879 150
rect 6945 -150 6975 150
rect 7041 -150 7071 150
rect 7137 -150 7167 150
rect 7233 -150 7263 150
rect 7329 -150 7359 150
rect 7425 -150 7455 150
rect 7521 -150 7551 150
rect 7617 -150 7647 150
rect 7713 -150 7743 150
rect 7809 -150 7839 150
rect 7905 -150 7935 150
rect 8001 -150 8031 150
rect 8097 -150 8127 150
rect 8193 -150 8223 150
rect 8289 -150 8319 150
rect 8385 -150 8415 150
rect 8481 -150 8511 150
rect 8577 -150 8607 150
rect 8673 -150 8703 150
rect 8769 -150 8799 150
rect 8865 -150 8895 150
rect 8961 -150 8991 150
rect 9057 -150 9087 150
rect 9153 -150 9183 150
rect 9249 -150 9279 150
rect 9345 -150 9375 150
rect 9441 -150 9471 150
rect 9537 -150 9567 150
rect 9633 -150 9663 150
rect 9729 -150 9759 150
rect 9825 -150 9855 150
rect 9921 -150 9951 150
rect 10017 -150 10047 150
rect 10113 -150 10143 150
rect 10209 -150 10239 150
rect 10305 -150 10335 150
rect 10401 -150 10431 150
rect 10497 -150 10527 150
rect 10593 -150 10623 150
rect 10689 -150 10719 150
rect 10785 -150 10815 150
rect 10881 -150 10911 150
rect 10977 -150 11007 150
rect 11073 -150 11103 150
rect 11169 -150 11199 150
rect 11265 -150 11295 150
rect 11361 -150 11391 150
rect 11457 -150 11487 150
rect 11553 -150 11583 150
rect 11649 -150 11679 150
rect 11745 -150 11775 150
rect 11841 -150 11871 150
rect 11937 -150 11967 150
rect 12033 -150 12063 150
rect 12129 -150 12159 150
rect 12225 -150 12255 150
rect 12321 -150 12351 150
rect 12417 -150 12447 150
rect 12513 -150 12543 150
rect 12609 -150 12639 150
rect 12705 -150 12735 150
rect 12801 -150 12831 150
rect 12897 -150 12927 150
rect 12993 -150 13023 150
rect 13089 -150 13119 150
rect 13185 -150 13215 150
rect 13281 -150 13311 150
rect 13377 -150 13407 150
rect 13473 -150 13503 150
rect 13569 -150 13599 150
rect 13665 -150 13695 150
rect 13761 -150 13791 150
rect 13857 -150 13887 150
rect 13953 -150 13983 150
rect 14049 -150 14079 150
rect 14145 -150 14175 150
rect 14241 -150 14271 150
rect 14337 -150 14367 150
rect 14433 -150 14463 150
rect 14529 -150 14559 150
rect 14625 -150 14655 150
rect 14721 -150 14751 150
rect 14817 -150 14847 150
rect 14913 -150 14943 150
rect 15009 -150 15039 150
rect 15105 -150 15135 150
rect 15201 -150 15231 150
rect 15297 -150 15327 150
rect 15393 -150 15423 150
rect 15489 -150 15519 150
rect 15585 -150 15615 150
rect 15681 -150 15711 150
rect 15777 -150 15807 150
rect 15873 -150 15903 150
rect 15969 -150 15999 150
rect 16065 -150 16095 150
rect 16161 -150 16191 150
rect 16257 -150 16287 150
rect 16353 -150 16383 150
rect 16449 -150 16479 150
rect 16545 -150 16575 150
rect 16641 -150 16671 150
rect 16737 -150 16767 150
rect 16833 -150 16863 150
rect 16929 -150 16959 150
rect 17025 -150 17055 150
rect 17121 -150 17151 150
rect 17217 -150 17247 150
rect 17313 -150 17343 150
rect 17409 -150 17439 150
rect 17505 -150 17535 150
rect 17601 -150 17631 150
rect 17697 -150 17727 150
rect 17793 -150 17823 150
rect 17889 -150 17919 150
rect 17985 -150 18015 150
rect 18081 -150 18111 150
rect 18177 -150 18207 150
rect 18273 -150 18303 150
rect 18369 -150 18399 150
rect 18465 -150 18495 150
rect 18561 -150 18591 150
rect 18657 -150 18687 150
rect 18753 -150 18783 150
rect 18849 -150 18879 150
rect 18945 -150 18975 150
rect 19041 -150 19071 150
rect 19137 -150 19167 150
<< ndiff >>
rect -19229 138 -19167 150
rect -19229 -138 -19217 138
rect -19183 -138 -19167 138
rect -19229 -150 -19167 -138
rect -19137 138 -19071 150
rect -19137 -138 -19121 138
rect -19087 -138 -19071 138
rect -19137 -150 -19071 -138
rect -19041 138 -18975 150
rect -19041 -138 -19025 138
rect -18991 -138 -18975 138
rect -19041 -150 -18975 -138
rect -18945 138 -18879 150
rect -18945 -138 -18929 138
rect -18895 -138 -18879 138
rect -18945 -150 -18879 -138
rect -18849 138 -18783 150
rect -18849 -138 -18833 138
rect -18799 -138 -18783 138
rect -18849 -150 -18783 -138
rect -18753 138 -18687 150
rect -18753 -138 -18737 138
rect -18703 -138 -18687 138
rect -18753 -150 -18687 -138
rect -18657 138 -18591 150
rect -18657 -138 -18641 138
rect -18607 -138 -18591 138
rect -18657 -150 -18591 -138
rect -18561 138 -18495 150
rect -18561 -138 -18545 138
rect -18511 -138 -18495 138
rect -18561 -150 -18495 -138
rect -18465 138 -18399 150
rect -18465 -138 -18449 138
rect -18415 -138 -18399 138
rect -18465 -150 -18399 -138
rect -18369 138 -18303 150
rect -18369 -138 -18353 138
rect -18319 -138 -18303 138
rect -18369 -150 -18303 -138
rect -18273 138 -18207 150
rect -18273 -138 -18257 138
rect -18223 -138 -18207 138
rect -18273 -150 -18207 -138
rect -18177 138 -18111 150
rect -18177 -138 -18161 138
rect -18127 -138 -18111 138
rect -18177 -150 -18111 -138
rect -18081 138 -18015 150
rect -18081 -138 -18065 138
rect -18031 -138 -18015 138
rect -18081 -150 -18015 -138
rect -17985 138 -17919 150
rect -17985 -138 -17969 138
rect -17935 -138 -17919 138
rect -17985 -150 -17919 -138
rect -17889 138 -17823 150
rect -17889 -138 -17873 138
rect -17839 -138 -17823 138
rect -17889 -150 -17823 -138
rect -17793 138 -17727 150
rect -17793 -138 -17777 138
rect -17743 -138 -17727 138
rect -17793 -150 -17727 -138
rect -17697 138 -17631 150
rect -17697 -138 -17681 138
rect -17647 -138 -17631 138
rect -17697 -150 -17631 -138
rect -17601 138 -17535 150
rect -17601 -138 -17585 138
rect -17551 -138 -17535 138
rect -17601 -150 -17535 -138
rect -17505 138 -17439 150
rect -17505 -138 -17489 138
rect -17455 -138 -17439 138
rect -17505 -150 -17439 -138
rect -17409 138 -17343 150
rect -17409 -138 -17393 138
rect -17359 -138 -17343 138
rect -17409 -150 -17343 -138
rect -17313 138 -17247 150
rect -17313 -138 -17297 138
rect -17263 -138 -17247 138
rect -17313 -150 -17247 -138
rect -17217 138 -17151 150
rect -17217 -138 -17201 138
rect -17167 -138 -17151 138
rect -17217 -150 -17151 -138
rect -17121 138 -17055 150
rect -17121 -138 -17105 138
rect -17071 -138 -17055 138
rect -17121 -150 -17055 -138
rect -17025 138 -16959 150
rect -17025 -138 -17009 138
rect -16975 -138 -16959 138
rect -17025 -150 -16959 -138
rect -16929 138 -16863 150
rect -16929 -138 -16913 138
rect -16879 -138 -16863 138
rect -16929 -150 -16863 -138
rect -16833 138 -16767 150
rect -16833 -138 -16817 138
rect -16783 -138 -16767 138
rect -16833 -150 -16767 -138
rect -16737 138 -16671 150
rect -16737 -138 -16721 138
rect -16687 -138 -16671 138
rect -16737 -150 -16671 -138
rect -16641 138 -16575 150
rect -16641 -138 -16625 138
rect -16591 -138 -16575 138
rect -16641 -150 -16575 -138
rect -16545 138 -16479 150
rect -16545 -138 -16529 138
rect -16495 -138 -16479 138
rect -16545 -150 -16479 -138
rect -16449 138 -16383 150
rect -16449 -138 -16433 138
rect -16399 -138 -16383 138
rect -16449 -150 -16383 -138
rect -16353 138 -16287 150
rect -16353 -138 -16337 138
rect -16303 -138 -16287 138
rect -16353 -150 -16287 -138
rect -16257 138 -16191 150
rect -16257 -138 -16241 138
rect -16207 -138 -16191 138
rect -16257 -150 -16191 -138
rect -16161 138 -16095 150
rect -16161 -138 -16145 138
rect -16111 -138 -16095 138
rect -16161 -150 -16095 -138
rect -16065 138 -15999 150
rect -16065 -138 -16049 138
rect -16015 -138 -15999 138
rect -16065 -150 -15999 -138
rect -15969 138 -15903 150
rect -15969 -138 -15953 138
rect -15919 -138 -15903 138
rect -15969 -150 -15903 -138
rect -15873 138 -15807 150
rect -15873 -138 -15857 138
rect -15823 -138 -15807 138
rect -15873 -150 -15807 -138
rect -15777 138 -15711 150
rect -15777 -138 -15761 138
rect -15727 -138 -15711 138
rect -15777 -150 -15711 -138
rect -15681 138 -15615 150
rect -15681 -138 -15665 138
rect -15631 -138 -15615 138
rect -15681 -150 -15615 -138
rect -15585 138 -15519 150
rect -15585 -138 -15569 138
rect -15535 -138 -15519 138
rect -15585 -150 -15519 -138
rect -15489 138 -15423 150
rect -15489 -138 -15473 138
rect -15439 -138 -15423 138
rect -15489 -150 -15423 -138
rect -15393 138 -15327 150
rect -15393 -138 -15377 138
rect -15343 -138 -15327 138
rect -15393 -150 -15327 -138
rect -15297 138 -15231 150
rect -15297 -138 -15281 138
rect -15247 -138 -15231 138
rect -15297 -150 -15231 -138
rect -15201 138 -15135 150
rect -15201 -138 -15185 138
rect -15151 -138 -15135 138
rect -15201 -150 -15135 -138
rect -15105 138 -15039 150
rect -15105 -138 -15089 138
rect -15055 -138 -15039 138
rect -15105 -150 -15039 -138
rect -15009 138 -14943 150
rect -15009 -138 -14993 138
rect -14959 -138 -14943 138
rect -15009 -150 -14943 -138
rect -14913 138 -14847 150
rect -14913 -138 -14897 138
rect -14863 -138 -14847 138
rect -14913 -150 -14847 -138
rect -14817 138 -14751 150
rect -14817 -138 -14801 138
rect -14767 -138 -14751 138
rect -14817 -150 -14751 -138
rect -14721 138 -14655 150
rect -14721 -138 -14705 138
rect -14671 -138 -14655 138
rect -14721 -150 -14655 -138
rect -14625 138 -14559 150
rect -14625 -138 -14609 138
rect -14575 -138 -14559 138
rect -14625 -150 -14559 -138
rect -14529 138 -14463 150
rect -14529 -138 -14513 138
rect -14479 -138 -14463 138
rect -14529 -150 -14463 -138
rect -14433 138 -14367 150
rect -14433 -138 -14417 138
rect -14383 -138 -14367 138
rect -14433 -150 -14367 -138
rect -14337 138 -14271 150
rect -14337 -138 -14321 138
rect -14287 -138 -14271 138
rect -14337 -150 -14271 -138
rect -14241 138 -14175 150
rect -14241 -138 -14225 138
rect -14191 -138 -14175 138
rect -14241 -150 -14175 -138
rect -14145 138 -14079 150
rect -14145 -138 -14129 138
rect -14095 -138 -14079 138
rect -14145 -150 -14079 -138
rect -14049 138 -13983 150
rect -14049 -138 -14033 138
rect -13999 -138 -13983 138
rect -14049 -150 -13983 -138
rect -13953 138 -13887 150
rect -13953 -138 -13937 138
rect -13903 -138 -13887 138
rect -13953 -150 -13887 -138
rect -13857 138 -13791 150
rect -13857 -138 -13841 138
rect -13807 -138 -13791 138
rect -13857 -150 -13791 -138
rect -13761 138 -13695 150
rect -13761 -138 -13745 138
rect -13711 -138 -13695 138
rect -13761 -150 -13695 -138
rect -13665 138 -13599 150
rect -13665 -138 -13649 138
rect -13615 -138 -13599 138
rect -13665 -150 -13599 -138
rect -13569 138 -13503 150
rect -13569 -138 -13553 138
rect -13519 -138 -13503 138
rect -13569 -150 -13503 -138
rect -13473 138 -13407 150
rect -13473 -138 -13457 138
rect -13423 -138 -13407 138
rect -13473 -150 -13407 -138
rect -13377 138 -13311 150
rect -13377 -138 -13361 138
rect -13327 -138 -13311 138
rect -13377 -150 -13311 -138
rect -13281 138 -13215 150
rect -13281 -138 -13265 138
rect -13231 -138 -13215 138
rect -13281 -150 -13215 -138
rect -13185 138 -13119 150
rect -13185 -138 -13169 138
rect -13135 -138 -13119 138
rect -13185 -150 -13119 -138
rect -13089 138 -13023 150
rect -13089 -138 -13073 138
rect -13039 -138 -13023 138
rect -13089 -150 -13023 -138
rect -12993 138 -12927 150
rect -12993 -138 -12977 138
rect -12943 -138 -12927 138
rect -12993 -150 -12927 -138
rect -12897 138 -12831 150
rect -12897 -138 -12881 138
rect -12847 -138 -12831 138
rect -12897 -150 -12831 -138
rect -12801 138 -12735 150
rect -12801 -138 -12785 138
rect -12751 -138 -12735 138
rect -12801 -150 -12735 -138
rect -12705 138 -12639 150
rect -12705 -138 -12689 138
rect -12655 -138 -12639 138
rect -12705 -150 -12639 -138
rect -12609 138 -12543 150
rect -12609 -138 -12593 138
rect -12559 -138 -12543 138
rect -12609 -150 -12543 -138
rect -12513 138 -12447 150
rect -12513 -138 -12497 138
rect -12463 -138 -12447 138
rect -12513 -150 -12447 -138
rect -12417 138 -12351 150
rect -12417 -138 -12401 138
rect -12367 -138 -12351 138
rect -12417 -150 -12351 -138
rect -12321 138 -12255 150
rect -12321 -138 -12305 138
rect -12271 -138 -12255 138
rect -12321 -150 -12255 -138
rect -12225 138 -12159 150
rect -12225 -138 -12209 138
rect -12175 -138 -12159 138
rect -12225 -150 -12159 -138
rect -12129 138 -12063 150
rect -12129 -138 -12113 138
rect -12079 -138 -12063 138
rect -12129 -150 -12063 -138
rect -12033 138 -11967 150
rect -12033 -138 -12017 138
rect -11983 -138 -11967 138
rect -12033 -150 -11967 -138
rect -11937 138 -11871 150
rect -11937 -138 -11921 138
rect -11887 -138 -11871 138
rect -11937 -150 -11871 -138
rect -11841 138 -11775 150
rect -11841 -138 -11825 138
rect -11791 -138 -11775 138
rect -11841 -150 -11775 -138
rect -11745 138 -11679 150
rect -11745 -138 -11729 138
rect -11695 -138 -11679 138
rect -11745 -150 -11679 -138
rect -11649 138 -11583 150
rect -11649 -138 -11633 138
rect -11599 -138 -11583 138
rect -11649 -150 -11583 -138
rect -11553 138 -11487 150
rect -11553 -138 -11537 138
rect -11503 -138 -11487 138
rect -11553 -150 -11487 -138
rect -11457 138 -11391 150
rect -11457 -138 -11441 138
rect -11407 -138 -11391 138
rect -11457 -150 -11391 -138
rect -11361 138 -11295 150
rect -11361 -138 -11345 138
rect -11311 -138 -11295 138
rect -11361 -150 -11295 -138
rect -11265 138 -11199 150
rect -11265 -138 -11249 138
rect -11215 -138 -11199 138
rect -11265 -150 -11199 -138
rect -11169 138 -11103 150
rect -11169 -138 -11153 138
rect -11119 -138 -11103 138
rect -11169 -150 -11103 -138
rect -11073 138 -11007 150
rect -11073 -138 -11057 138
rect -11023 -138 -11007 138
rect -11073 -150 -11007 -138
rect -10977 138 -10911 150
rect -10977 -138 -10961 138
rect -10927 -138 -10911 138
rect -10977 -150 -10911 -138
rect -10881 138 -10815 150
rect -10881 -138 -10865 138
rect -10831 -138 -10815 138
rect -10881 -150 -10815 -138
rect -10785 138 -10719 150
rect -10785 -138 -10769 138
rect -10735 -138 -10719 138
rect -10785 -150 -10719 -138
rect -10689 138 -10623 150
rect -10689 -138 -10673 138
rect -10639 -138 -10623 138
rect -10689 -150 -10623 -138
rect -10593 138 -10527 150
rect -10593 -138 -10577 138
rect -10543 -138 -10527 138
rect -10593 -150 -10527 -138
rect -10497 138 -10431 150
rect -10497 -138 -10481 138
rect -10447 -138 -10431 138
rect -10497 -150 -10431 -138
rect -10401 138 -10335 150
rect -10401 -138 -10385 138
rect -10351 -138 -10335 138
rect -10401 -150 -10335 -138
rect -10305 138 -10239 150
rect -10305 -138 -10289 138
rect -10255 -138 -10239 138
rect -10305 -150 -10239 -138
rect -10209 138 -10143 150
rect -10209 -138 -10193 138
rect -10159 -138 -10143 138
rect -10209 -150 -10143 -138
rect -10113 138 -10047 150
rect -10113 -138 -10097 138
rect -10063 -138 -10047 138
rect -10113 -150 -10047 -138
rect -10017 138 -9951 150
rect -10017 -138 -10001 138
rect -9967 -138 -9951 138
rect -10017 -150 -9951 -138
rect -9921 138 -9855 150
rect -9921 -138 -9905 138
rect -9871 -138 -9855 138
rect -9921 -150 -9855 -138
rect -9825 138 -9759 150
rect -9825 -138 -9809 138
rect -9775 -138 -9759 138
rect -9825 -150 -9759 -138
rect -9729 138 -9663 150
rect -9729 -138 -9713 138
rect -9679 -138 -9663 138
rect -9729 -150 -9663 -138
rect -9633 138 -9567 150
rect -9633 -138 -9617 138
rect -9583 -138 -9567 138
rect -9633 -150 -9567 -138
rect -9537 138 -9471 150
rect -9537 -138 -9521 138
rect -9487 -138 -9471 138
rect -9537 -150 -9471 -138
rect -9441 138 -9375 150
rect -9441 -138 -9425 138
rect -9391 -138 -9375 138
rect -9441 -150 -9375 -138
rect -9345 138 -9279 150
rect -9345 -138 -9329 138
rect -9295 -138 -9279 138
rect -9345 -150 -9279 -138
rect -9249 138 -9183 150
rect -9249 -138 -9233 138
rect -9199 -138 -9183 138
rect -9249 -150 -9183 -138
rect -9153 138 -9087 150
rect -9153 -138 -9137 138
rect -9103 -138 -9087 138
rect -9153 -150 -9087 -138
rect -9057 138 -8991 150
rect -9057 -138 -9041 138
rect -9007 -138 -8991 138
rect -9057 -150 -8991 -138
rect -8961 138 -8895 150
rect -8961 -138 -8945 138
rect -8911 -138 -8895 138
rect -8961 -150 -8895 -138
rect -8865 138 -8799 150
rect -8865 -138 -8849 138
rect -8815 -138 -8799 138
rect -8865 -150 -8799 -138
rect -8769 138 -8703 150
rect -8769 -138 -8753 138
rect -8719 -138 -8703 138
rect -8769 -150 -8703 -138
rect -8673 138 -8607 150
rect -8673 -138 -8657 138
rect -8623 -138 -8607 138
rect -8673 -150 -8607 -138
rect -8577 138 -8511 150
rect -8577 -138 -8561 138
rect -8527 -138 -8511 138
rect -8577 -150 -8511 -138
rect -8481 138 -8415 150
rect -8481 -138 -8465 138
rect -8431 -138 -8415 138
rect -8481 -150 -8415 -138
rect -8385 138 -8319 150
rect -8385 -138 -8369 138
rect -8335 -138 -8319 138
rect -8385 -150 -8319 -138
rect -8289 138 -8223 150
rect -8289 -138 -8273 138
rect -8239 -138 -8223 138
rect -8289 -150 -8223 -138
rect -8193 138 -8127 150
rect -8193 -138 -8177 138
rect -8143 -138 -8127 138
rect -8193 -150 -8127 -138
rect -8097 138 -8031 150
rect -8097 -138 -8081 138
rect -8047 -138 -8031 138
rect -8097 -150 -8031 -138
rect -8001 138 -7935 150
rect -8001 -138 -7985 138
rect -7951 -138 -7935 138
rect -8001 -150 -7935 -138
rect -7905 138 -7839 150
rect -7905 -138 -7889 138
rect -7855 -138 -7839 138
rect -7905 -150 -7839 -138
rect -7809 138 -7743 150
rect -7809 -138 -7793 138
rect -7759 -138 -7743 138
rect -7809 -150 -7743 -138
rect -7713 138 -7647 150
rect -7713 -138 -7697 138
rect -7663 -138 -7647 138
rect -7713 -150 -7647 -138
rect -7617 138 -7551 150
rect -7617 -138 -7601 138
rect -7567 -138 -7551 138
rect -7617 -150 -7551 -138
rect -7521 138 -7455 150
rect -7521 -138 -7505 138
rect -7471 -138 -7455 138
rect -7521 -150 -7455 -138
rect -7425 138 -7359 150
rect -7425 -138 -7409 138
rect -7375 -138 -7359 138
rect -7425 -150 -7359 -138
rect -7329 138 -7263 150
rect -7329 -138 -7313 138
rect -7279 -138 -7263 138
rect -7329 -150 -7263 -138
rect -7233 138 -7167 150
rect -7233 -138 -7217 138
rect -7183 -138 -7167 138
rect -7233 -150 -7167 -138
rect -7137 138 -7071 150
rect -7137 -138 -7121 138
rect -7087 -138 -7071 138
rect -7137 -150 -7071 -138
rect -7041 138 -6975 150
rect -7041 -138 -7025 138
rect -6991 -138 -6975 138
rect -7041 -150 -6975 -138
rect -6945 138 -6879 150
rect -6945 -138 -6929 138
rect -6895 -138 -6879 138
rect -6945 -150 -6879 -138
rect -6849 138 -6783 150
rect -6849 -138 -6833 138
rect -6799 -138 -6783 138
rect -6849 -150 -6783 -138
rect -6753 138 -6687 150
rect -6753 -138 -6737 138
rect -6703 -138 -6687 138
rect -6753 -150 -6687 -138
rect -6657 138 -6591 150
rect -6657 -138 -6641 138
rect -6607 -138 -6591 138
rect -6657 -150 -6591 -138
rect -6561 138 -6495 150
rect -6561 -138 -6545 138
rect -6511 -138 -6495 138
rect -6561 -150 -6495 -138
rect -6465 138 -6399 150
rect -6465 -138 -6449 138
rect -6415 -138 -6399 138
rect -6465 -150 -6399 -138
rect -6369 138 -6303 150
rect -6369 -138 -6353 138
rect -6319 -138 -6303 138
rect -6369 -150 -6303 -138
rect -6273 138 -6207 150
rect -6273 -138 -6257 138
rect -6223 -138 -6207 138
rect -6273 -150 -6207 -138
rect -6177 138 -6111 150
rect -6177 -138 -6161 138
rect -6127 -138 -6111 138
rect -6177 -150 -6111 -138
rect -6081 138 -6015 150
rect -6081 -138 -6065 138
rect -6031 -138 -6015 138
rect -6081 -150 -6015 -138
rect -5985 138 -5919 150
rect -5985 -138 -5969 138
rect -5935 -138 -5919 138
rect -5985 -150 -5919 -138
rect -5889 138 -5823 150
rect -5889 -138 -5873 138
rect -5839 -138 -5823 138
rect -5889 -150 -5823 -138
rect -5793 138 -5727 150
rect -5793 -138 -5777 138
rect -5743 -138 -5727 138
rect -5793 -150 -5727 -138
rect -5697 138 -5631 150
rect -5697 -138 -5681 138
rect -5647 -138 -5631 138
rect -5697 -150 -5631 -138
rect -5601 138 -5535 150
rect -5601 -138 -5585 138
rect -5551 -138 -5535 138
rect -5601 -150 -5535 -138
rect -5505 138 -5439 150
rect -5505 -138 -5489 138
rect -5455 -138 -5439 138
rect -5505 -150 -5439 -138
rect -5409 138 -5343 150
rect -5409 -138 -5393 138
rect -5359 -138 -5343 138
rect -5409 -150 -5343 -138
rect -5313 138 -5247 150
rect -5313 -138 -5297 138
rect -5263 -138 -5247 138
rect -5313 -150 -5247 -138
rect -5217 138 -5151 150
rect -5217 -138 -5201 138
rect -5167 -138 -5151 138
rect -5217 -150 -5151 -138
rect -5121 138 -5055 150
rect -5121 -138 -5105 138
rect -5071 -138 -5055 138
rect -5121 -150 -5055 -138
rect -5025 138 -4959 150
rect -5025 -138 -5009 138
rect -4975 -138 -4959 138
rect -5025 -150 -4959 -138
rect -4929 138 -4863 150
rect -4929 -138 -4913 138
rect -4879 -138 -4863 138
rect -4929 -150 -4863 -138
rect -4833 138 -4767 150
rect -4833 -138 -4817 138
rect -4783 -138 -4767 138
rect -4833 -150 -4767 -138
rect -4737 138 -4671 150
rect -4737 -138 -4721 138
rect -4687 -138 -4671 138
rect -4737 -150 -4671 -138
rect -4641 138 -4575 150
rect -4641 -138 -4625 138
rect -4591 -138 -4575 138
rect -4641 -150 -4575 -138
rect -4545 138 -4479 150
rect -4545 -138 -4529 138
rect -4495 -138 -4479 138
rect -4545 -150 -4479 -138
rect -4449 138 -4383 150
rect -4449 -138 -4433 138
rect -4399 -138 -4383 138
rect -4449 -150 -4383 -138
rect -4353 138 -4287 150
rect -4353 -138 -4337 138
rect -4303 -138 -4287 138
rect -4353 -150 -4287 -138
rect -4257 138 -4191 150
rect -4257 -138 -4241 138
rect -4207 -138 -4191 138
rect -4257 -150 -4191 -138
rect -4161 138 -4095 150
rect -4161 -138 -4145 138
rect -4111 -138 -4095 138
rect -4161 -150 -4095 -138
rect -4065 138 -3999 150
rect -4065 -138 -4049 138
rect -4015 -138 -3999 138
rect -4065 -150 -3999 -138
rect -3969 138 -3903 150
rect -3969 -138 -3953 138
rect -3919 -138 -3903 138
rect -3969 -150 -3903 -138
rect -3873 138 -3807 150
rect -3873 -138 -3857 138
rect -3823 -138 -3807 138
rect -3873 -150 -3807 -138
rect -3777 138 -3711 150
rect -3777 -138 -3761 138
rect -3727 -138 -3711 138
rect -3777 -150 -3711 -138
rect -3681 138 -3615 150
rect -3681 -138 -3665 138
rect -3631 -138 -3615 138
rect -3681 -150 -3615 -138
rect -3585 138 -3519 150
rect -3585 -138 -3569 138
rect -3535 -138 -3519 138
rect -3585 -150 -3519 -138
rect -3489 138 -3423 150
rect -3489 -138 -3473 138
rect -3439 -138 -3423 138
rect -3489 -150 -3423 -138
rect -3393 138 -3327 150
rect -3393 -138 -3377 138
rect -3343 -138 -3327 138
rect -3393 -150 -3327 -138
rect -3297 138 -3231 150
rect -3297 -138 -3281 138
rect -3247 -138 -3231 138
rect -3297 -150 -3231 -138
rect -3201 138 -3135 150
rect -3201 -138 -3185 138
rect -3151 -138 -3135 138
rect -3201 -150 -3135 -138
rect -3105 138 -3039 150
rect -3105 -138 -3089 138
rect -3055 -138 -3039 138
rect -3105 -150 -3039 -138
rect -3009 138 -2943 150
rect -3009 -138 -2993 138
rect -2959 -138 -2943 138
rect -3009 -150 -2943 -138
rect -2913 138 -2847 150
rect -2913 -138 -2897 138
rect -2863 -138 -2847 138
rect -2913 -150 -2847 -138
rect -2817 138 -2751 150
rect -2817 -138 -2801 138
rect -2767 -138 -2751 138
rect -2817 -150 -2751 -138
rect -2721 138 -2655 150
rect -2721 -138 -2705 138
rect -2671 -138 -2655 138
rect -2721 -150 -2655 -138
rect -2625 138 -2559 150
rect -2625 -138 -2609 138
rect -2575 -138 -2559 138
rect -2625 -150 -2559 -138
rect -2529 138 -2463 150
rect -2529 -138 -2513 138
rect -2479 -138 -2463 138
rect -2529 -150 -2463 -138
rect -2433 138 -2367 150
rect -2433 -138 -2417 138
rect -2383 -138 -2367 138
rect -2433 -150 -2367 -138
rect -2337 138 -2271 150
rect -2337 -138 -2321 138
rect -2287 -138 -2271 138
rect -2337 -150 -2271 -138
rect -2241 138 -2175 150
rect -2241 -138 -2225 138
rect -2191 -138 -2175 138
rect -2241 -150 -2175 -138
rect -2145 138 -2079 150
rect -2145 -138 -2129 138
rect -2095 -138 -2079 138
rect -2145 -150 -2079 -138
rect -2049 138 -1983 150
rect -2049 -138 -2033 138
rect -1999 -138 -1983 138
rect -2049 -150 -1983 -138
rect -1953 138 -1887 150
rect -1953 -138 -1937 138
rect -1903 -138 -1887 138
rect -1953 -150 -1887 -138
rect -1857 138 -1791 150
rect -1857 -138 -1841 138
rect -1807 -138 -1791 138
rect -1857 -150 -1791 -138
rect -1761 138 -1695 150
rect -1761 -138 -1745 138
rect -1711 -138 -1695 138
rect -1761 -150 -1695 -138
rect -1665 138 -1599 150
rect -1665 -138 -1649 138
rect -1615 -138 -1599 138
rect -1665 -150 -1599 -138
rect -1569 138 -1503 150
rect -1569 -138 -1553 138
rect -1519 -138 -1503 138
rect -1569 -150 -1503 -138
rect -1473 138 -1407 150
rect -1473 -138 -1457 138
rect -1423 -138 -1407 138
rect -1473 -150 -1407 -138
rect -1377 138 -1311 150
rect -1377 -138 -1361 138
rect -1327 -138 -1311 138
rect -1377 -150 -1311 -138
rect -1281 138 -1215 150
rect -1281 -138 -1265 138
rect -1231 -138 -1215 138
rect -1281 -150 -1215 -138
rect -1185 138 -1119 150
rect -1185 -138 -1169 138
rect -1135 -138 -1119 138
rect -1185 -150 -1119 -138
rect -1089 138 -1023 150
rect -1089 -138 -1073 138
rect -1039 -138 -1023 138
rect -1089 -150 -1023 -138
rect -993 138 -927 150
rect -993 -138 -977 138
rect -943 -138 -927 138
rect -993 -150 -927 -138
rect -897 138 -831 150
rect -897 -138 -881 138
rect -847 -138 -831 138
rect -897 -150 -831 -138
rect -801 138 -735 150
rect -801 -138 -785 138
rect -751 -138 -735 138
rect -801 -150 -735 -138
rect -705 138 -639 150
rect -705 -138 -689 138
rect -655 -138 -639 138
rect -705 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 705 150
rect 639 -138 655 138
rect 689 -138 705 138
rect 639 -150 705 -138
rect 735 138 801 150
rect 735 -138 751 138
rect 785 -138 801 138
rect 735 -150 801 -138
rect 831 138 897 150
rect 831 -138 847 138
rect 881 -138 897 138
rect 831 -150 897 -138
rect 927 138 993 150
rect 927 -138 943 138
rect 977 -138 993 138
rect 927 -150 993 -138
rect 1023 138 1089 150
rect 1023 -138 1039 138
rect 1073 -138 1089 138
rect 1023 -150 1089 -138
rect 1119 138 1185 150
rect 1119 -138 1135 138
rect 1169 -138 1185 138
rect 1119 -150 1185 -138
rect 1215 138 1281 150
rect 1215 -138 1231 138
rect 1265 -138 1281 138
rect 1215 -150 1281 -138
rect 1311 138 1377 150
rect 1311 -138 1327 138
rect 1361 -138 1377 138
rect 1311 -150 1377 -138
rect 1407 138 1473 150
rect 1407 -138 1423 138
rect 1457 -138 1473 138
rect 1407 -150 1473 -138
rect 1503 138 1569 150
rect 1503 -138 1519 138
rect 1553 -138 1569 138
rect 1503 -150 1569 -138
rect 1599 138 1665 150
rect 1599 -138 1615 138
rect 1649 -138 1665 138
rect 1599 -150 1665 -138
rect 1695 138 1761 150
rect 1695 -138 1711 138
rect 1745 -138 1761 138
rect 1695 -150 1761 -138
rect 1791 138 1857 150
rect 1791 -138 1807 138
rect 1841 -138 1857 138
rect 1791 -150 1857 -138
rect 1887 138 1953 150
rect 1887 -138 1903 138
rect 1937 -138 1953 138
rect 1887 -150 1953 -138
rect 1983 138 2049 150
rect 1983 -138 1999 138
rect 2033 -138 2049 138
rect 1983 -150 2049 -138
rect 2079 138 2145 150
rect 2079 -138 2095 138
rect 2129 -138 2145 138
rect 2079 -150 2145 -138
rect 2175 138 2241 150
rect 2175 -138 2191 138
rect 2225 -138 2241 138
rect 2175 -150 2241 -138
rect 2271 138 2337 150
rect 2271 -138 2287 138
rect 2321 -138 2337 138
rect 2271 -150 2337 -138
rect 2367 138 2433 150
rect 2367 -138 2383 138
rect 2417 -138 2433 138
rect 2367 -150 2433 -138
rect 2463 138 2529 150
rect 2463 -138 2479 138
rect 2513 -138 2529 138
rect 2463 -150 2529 -138
rect 2559 138 2625 150
rect 2559 -138 2575 138
rect 2609 -138 2625 138
rect 2559 -150 2625 -138
rect 2655 138 2721 150
rect 2655 -138 2671 138
rect 2705 -138 2721 138
rect 2655 -150 2721 -138
rect 2751 138 2817 150
rect 2751 -138 2767 138
rect 2801 -138 2817 138
rect 2751 -150 2817 -138
rect 2847 138 2913 150
rect 2847 -138 2863 138
rect 2897 -138 2913 138
rect 2847 -150 2913 -138
rect 2943 138 3009 150
rect 2943 -138 2959 138
rect 2993 -138 3009 138
rect 2943 -150 3009 -138
rect 3039 138 3105 150
rect 3039 -138 3055 138
rect 3089 -138 3105 138
rect 3039 -150 3105 -138
rect 3135 138 3201 150
rect 3135 -138 3151 138
rect 3185 -138 3201 138
rect 3135 -150 3201 -138
rect 3231 138 3297 150
rect 3231 -138 3247 138
rect 3281 -138 3297 138
rect 3231 -150 3297 -138
rect 3327 138 3393 150
rect 3327 -138 3343 138
rect 3377 -138 3393 138
rect 3327 -150 3393 -138
rect 3423 138 3489 150
rect 3423 -138 3439 138
rect 3473 -138 3489 138
rect 3423 -150 3489 -138
rect 3519 138 3585 150
rect 3519 -138 3535 138
rect 3569 -138 3585 138
rect 3519 -150 3585 -138
rect 3615 138 3681 150
rect 3615 -138 3631 138
rect 3665 -138 3681 138
rect 3615 -150 3681 -138
rect 3711 138 3777 150
rect 3711 -138 3727 138
rect 3761 -138 3777 138
rect 3711 -150 3777 -138
rect 3807 138 3873 150
rect 3807 -138 3823 138
rect 3857 -138 3873 138
rect 3807 -150 3873 -138
rect 3903 138 3969 150
rect 3903 -138 3919 138
rect 3953 -138 3969 138
rect 3903 -150 3969 -138
rect 3999 138 4065 150
rect 3999 -138 4015 138
rect 4049 -138 4065 138
rect 3999 -150 4065 -138
rect 4095 138 4161 150
rect 4095 -138 4111 138
rect 4145 -138 4161 138
rect 4095 -150 4161 -138
rect 4191 138 4257 150
rect 4191 -138 4207 138
rect 4241 -138 4257 138
rect 4191 -150 4257 -138
rect 4287 138 4353 150
rect 4287 -138 4303 138
rect 4337 -138 4353 138
rect 4287 -150 4353 -138
rect 4383 138 4449 150
rect 4383 -138 4399 138
rect 4433 -138 4449 138
rect 4383 -150 4449 -138
rect 4479 138 4545 150
rect 4479 -138 4495 138
rect 4529 -138 4545 138
rect 4479 -150 4545 -138
rect 4575 138 4641 150
rect 4575 -138 4591 138
rect 4625 -138 4641 138
rect 4575 -150 4641 -138
rect 4671 138 4737 150
rect 4671 -138 4687 138
rect 4721 -138 4737 138
rect 4671 -150 4737 -138
rect 4767 138 4833 150
rect 4767 -138 4783 138
rect 4817 -138 4833 138
rect 4767 -150 4833 -138
rect 4863 138 4929 150
rect 4863 -138 4879 138
rect 4913 -138 4929 138
rect 4863 -150 4929 -138
rect 4959 138 5025 150
rect 4959 -138 4975 138
rect 5009 -138 5025 138
rect 4959 -150 5025 -138
rect 5055 138 5121 150
rect 5055 -138 5071 138
rect 5105 -138 5121 138
rect 5055 -150 5121 -138
rect 5151 138 5217 150
rect 5151 -138 5167 138
rect 5201 -138 5217 138
rect 5151 -150 5217 -138
rect 5247 138 5313 150
rect 5247 -138 5263 138
rect 5297 -138 5313 138
rect 5247 -150 5313 -138
rect 5343 138 5409 150
rect 5343 -138 5359 138
rect 5393 -138 5409 138
rect 5343 -150 5409 -138
rect 5439 138 5505 150
rect 5439 -138 5455 138
rect 5489 -138 5505 138
rect 5439 -150 5505 -138
rect 5535 138 5601 150
rect 5535 -138 5551 138
rect 5585 -138 5601 138
rect 5535 -150 5601 -138
rect 5631 138 5697 150
rect 5631 -138 5647 138
rect 5681 -138 5697 138
rect 5631 -150 5697 -138
rect 5727 138 5793 150
rect 5727 -138 5743 138
rect 5777 -138 5793 138
rect 5727 -150 5793 -138
rect 5823 138 5889 150
rect 5823 -138 5839 138
rect 5873 -138 5889 138
rect 5823 -150 5889 -138
rect 5919 138 5985 150
rect 5919 -138 5935 138
rect 5969 -138 5985 138
rect 5919 -150 5985 -138
rect 6015 138 6081 150
rect 6015 -138 6031 138
rect 6065 -138 6081 138
rect 6015 -150 6081 -138
rect 6111 138 6177 150
rect 6111 -138 6127 138
rect 6161 -138 6177 138
rect 6111 -150 6177 -138
rect 6207 138 6273 150
rect 6207 -138 6223 138
rect 6257 -138 6273 138
rect 6207 -150 6273 -138
rect 6303 138 6369 150
rect 6303 -138 6319 138
rect 6353 -138 6369 138
rect 6303 -150 6369 -138
rect 6399 138 6465 150
rect 6399 -138 6415 138
rect 6449 -138 6465 138
rect 6399 -150 6465 -138
rect 6495 138 6561 150
rect 6495 -138 6511 138
rect 6545 -138 6561 138
rect 6495 -150 6561 -138
rect 6591 138 6657 150
rect 6591 -138 6607 138
rect 6641 -138 6657 138
rect 6591 -150 6657 -138
rect 6687 138 6753 150
rect 6687 -138 6703 138
rect 6737 -138 6753 138
rect 6687 -150 6753 -138
rect 6783 138 6849 150
rect 6783 -138 6799 138
rect 6833 -138 6849 138
rect 6783 -150 6849 -138
rect 6879 138 6945 150
rect 6879 -138 6895 138
rect 6929 -138 6945 138
rect 6879 -150 6945 -138
rect 6975 138 7041 150
rect 6975 -138 6991 138
rect 7025 -138 7041 138
rect 6975 -150 7041 -138
rect 7071 138 7137 150
rect 7071 -138 7087 138
rect 7121 -138 7137 138
rect 7071 -150 7137 -138
rect 7167 138 7233 150
rect 7167 -138 7183 138
rect 7217 -138 7233 138
rect 7167 -150 7233 -138
rect 7263 138 7329 150
rect 7263 -138 7279 138
rect 7313 -138 7329 138
rect 7263 -150 7329 -138
rect 7359 138 7425 150
rect 7359 -138 7375 138
rect 7409 -138 7425 138
rect 7359 -150 7425 -138
rect 7455 138 7521 150
rect 7455 -138 7471 138
rect 7505 -138 7521 138
rect 7455 -150 7521 -138
rect 7551 138 7617 150
rect 7551 -138 7567 138
rect 7601 -138 7617 138
rect 7551 -150 7617 -138
rect 7647 138 7713 150
rect 7647 -138 7663 138
rect 7697 -138 7713 138
rect 7647 -150 7713 -138
rect 7743 138 7809 150
rect 7743 -138 7759 138
rect 7793 -138 7809 138
rect 7743 -150 7809 -138
rect 7839 138 7905 150
rect 7839 -138 7855 138
rect 7889 -138 7905 138
rect 7839 -150 7905 -138
rect 7935 138 8001 150
rect 7935 -138 7951 138
rect 7985 -138 8001 138
rect 7935 -150 8001 -138
rect 8031 138 8097 150
rect 8031 -138 8047 138
rect 8081 -138 8097 138
rect 8031 -150 8097 -138
rect 8127 138 8193 150
rect 8127 -138 8143 138
rect 8177 -138 8193 138
rect 8127 -150 8193 -138
rect 8223 138 8289 150
rect 8223 -138 8239 138
rect 8273 -138 8289 138
rect 8223 -150 8289 -138
rect 8319 138 8385 150
rect 8319 -138 8335 138
rect 8369 -138 8385 138
rect 8319 -150 8385 -138
rect 8415 138 8481 150
rect 8415 -138 8431 138
rect 8465 -138 8481 138
rect 8415 -150 8481 -138
rect 8511 138 8577 150
rect 8511 -138 8527 138
rect 8561 -138 8577 138
rect 8511 -150 8577 -138
rect 8607 138 8673 150
rect 8607 -138 8623 138
rect 8657 -138 8673 138
rect 8607 -150 8673 -138
rect 8703 138 8769 150
rect 8703 -138 8719 138
rect 8753 -138 8769 138
rect 8703 -150 8769 -138
rect 8799 138 8865 150
rect 8799 -138 8815 138
rect 8849 -138 8865 138
rect 8799 -150 8865 -138
rect 8895 138 8961 150
rect 8895 -138 8911 138
rect 8945 -138 8961 138
rect 8895 -150 8961 -138
rect 8991 138 9057 150
rect 8991 -138 9007 138
rect 9041 -138 9057 138
rect 8991 -150 9057 -138
rect 9087 138 9153 150
rect 9087 -138 9103 138
rect 9137 -138 9153 138
rect 9087 -150 9153 -138
rect 9183 138 9249 150
rect 9183 -138 9199 138
rect 9233 -138 9249 138
rect 9183 -150 9249 -138
rect 9279 138 9345 150
rect 9279 -138 9295 138
rect 9329 -138 9345 138
rect 9279 -150 9345 -138
rect 9375 138 9441 150
rect 9375 -138 9391 138
rect 9425 -138 9441 138
rect 9375 -150 9441 -138
rect 9471 138 9537 150
rect 9471 -138 9487 138
rect 9521 -138 9537 138
rect 9471 -150 9537 -138
rect 9567 138 9633 150
rect 9567 -138 9583 138
rect 9617 -138 9633 138
rect 9567 -150 9633 -138
rect 9663 138 9729 150
rect 9663 -138 9679 138
rect 9713 -138 9729 138
rect 9663 -150 9729 -138
rect 9759 138 9825 150
rect 9759 -138 9775 138
rect 9809 -138 9825 138
rect 9759 -150 9825 -138
rect 9855 138 9921 150
rect 9855 -138 9871 138
rect 9905 -138 9921 138
rect 9855 -150 9921 -138
rect 9951 138 10017 150
rect 9951 -138 9967 138
rect 10001 -138 10017 138
rect 9951 -150 10017 -138
rect 10047 138 10113 150
rect 10047 -138 10063 138
rect 10097 -138 10113 138
rect 10047 -150 10113 -138
rect 10143 138 10209 150
rect 10143 -138 10159 138
rect 10193 -138 10209 138
rect 10143 -150 10209 -138
rect 10239 138 10305 150
rect 10239 -138 10255 138
rect 10289 -138 10305 138
rect 10239 -150 10305 -138
rect 10335 138 10401 150
rect 10335 -138 10351 138
rect 10385 -138 10401 138
rect 10335 -150 10401 -138
rect 10431 138 10497 150
rect 10431 -138 10447 138
rect 10481 -138 10497 138
rect 10431 -150 10497 -138
rect 10527 138 10593 150
rect 10527 -138 10543 138
rect 10577 -138 10593 138
rect 10527 -150 10593 -138
rect 10623 138 10689 150
rect 10623 -138 10639 138
rect 10673 -138 10689 138
rect 10623 -150 10689 -138
rect 10719 138 10785 150
rect 10719 -138 10735 138
rect 10769 -138 10785 138
rect 10719 -150 10785 -138
rect 10815 138 10881 150
rect 10815 -138 10831 138
rect 10865 -138 10881 138
rect 10815 -150 10881 -138
rect 10911 138 10977 150
rect 10911 -138 10927 138
rect 10961 -138 10977 138
rect 10911 -150 10977 -138
rect 11007 138 11073 150
rect 11007 -138 11023 138
rect 11057 -138 11073 138
rect 11007 -150 11073 -138
rect 11103 138 11169 150
rect 11103 -138 11119 138
rect 11153 -138 11169 138
rect 11103 -150 11169 -138
rect 11199 138 11265 150
rect 11199 -138 11215 138
rect 11249 -138 11265 138
rect 11199 -150 11265 -138
rect 11295 138 11361 150
rect 11295 -138 11311 138
rect 11345 -138 11361 138
rect 11295 -150 11361 -138
rect 11391 138 11457 150
rect 11391 -138 11407 138
rect 11441 -138 11457 138
rect 11391 -150 11457 -138
rect 11487 138 11553 150
rect 11487 -138 11503 138
rect 11537 -138 11553 138
rect 11487 -150 11553 -138
rect 11583 138 11649 150
rect 11583 -138 11599 138
rect 11633 -138 11649 138
rect 11583 -150 11649 -138
rect 11679 138 11745 150
rect 11679 -138 11695 138
rect 11729 -138 11745 138
rect 11679 -150 11745 -138
rect 11775 138 11841 150
rect 11775 -138 11791 138
rect 11825 -138 11841 138
rect 11775 -150 11841 -138
rect 11871 138 11937 150
rect 11871 -138 11887 138
rect 11921 -138 11937 138
rect 11871 -150 11937 -138
rect 11967 138 12033 150
rect 11967 -138 11983 138
rect 12017 -138 12033 138
rect 11967 -150 12033 -138
rect 12063 138 12129 150
rect 12063 -138 12079 138
rect 12113 -138 12129 138
rect 12063 -150 12129 -138
rect 12159 138 12225 150
rect 12159 -138 12175 138
rect 12209 -138 12225 138
rect 12159 -150 12225 -138
rect 12255 138 12321 150
rect 12255 -138 12271 138
rect 12305 -138 12321 138
rect 12255 -150 12321 -138
rect 12351 138 12417 150
rect 12351 -138 12367 138
rect 12401 -138 12417 138
rect 12351 -150 12417 -138
rect 12447 138 12513 150
rect 12447 -138 12463 138
rect 12497 -138 12513 138
rect 12447 -150 12513 -138
rect 12543 138 12609 150
rect 12543 -138 12559 138
rect 12593 -138 12609 138
rect 12543 -150 12609 -138
rect 12639 138 12705 150
rect 12639 -138 12655 138
rect 12689 -138 12705 138
rect 12639 -150 12705 -138
rect 12735 138 12801 150
rect 12735 -138 12751 138
rect 12785 -138 12801 138
rect 12735 -150 12801 -138
rect 12831 138 12897 150
rect 12831 -138 12847 138
rect 12881 -138 12897 138
rect 12831 -150 12897 -138
rect 12927 138 12993 150
rect 12927 -138 12943 138
rect 12977 -138 12993 138
rect 12927 -150 12993 -138
rect 13023 138 13089 150
rect 13023 -138 13039 138
rect 13073 -138 13089 138
rect 13023 -150 13089 -138
rect 13119 138 13185 150
rect 13119 -138 13135 138
rect 13169 -138 13185 138
rect 13119 -150 13185 -138
rect 13215 138 13281 150
rect 13215 -138 13231 138
rect 13265 -138 13281 138
rect 13215 -150 13281 -138
rect 13311 138 13377 150
rect 13311 -138 13327 138
rect 13361 -138 13377 138
rect 13311 -150 13377 -138
rect 13407 138 13473 150
rect 13407 -138 13423 138
rect 13457 -138 13473 138
rect 13407 -150 13473 -138
rect 13503 138 13569 150
rect 13503 -138 13519 138
rect 13553 -138 13569 138
rect 13503 -150 13569 -138
rect 13599 138 13665 150
rect 13599 -138 13615 138
rect 13649 -138 13665 138
rect 13599 -150 13665 -138
rect 13695 138 13761 150
rect 13695 -138 13711 138
rect 13745 -138 13761 138
rect 13695 -150 13761 -138
rect 13791 138 13857 150
rect 13791 -138 13807 138
rect 13841 -138 13857 138
rect 13791 -150 13857 -138
rect 13887 138 13953 150
rect 13887 -138 13903 138
rect 13937 -138 13953 138
rect 13887 -150 13953 -138
rect 13983 138 14049 150
rect 13983 -138 13999 138
rect 14033 -138 14049 138
rect 13983 -150 14049 -138
rect 14079 138 14145 150
rect 14079 -138 14095 138
rect 14129 -138 14145 138
rect 14079 -150 14145 -138
rect 14175 138 14241 150
rect 14175 -138 14191 138
rect 14225 -138 14241 138
rect 14175 -150 14241 -138
rect 14271 138 14337 150
rect 14271 -138 14287 138
rect 14321 -138 14337 138
rect 14271 -150 14337 -138
rect 14367 138 14433 150
rect 14367 -138 14383 138
rect 14417 -138 14433 138
rect 14367 -150 14433 -138
rect 14463 138 14529 150
rect 14463 -138 14479 138
rect 14513 -138 14529 138
rect 14463 -150 14529 -138
rect 14559 138 14625 150
rect 14559 -138 14575 138
rect 14609 -138 14625 138
rect 14559 -150 14625 -138
rect 14655 138 14721 150
rect 14655 -138 14671 138
rect 14705 -138 14721 138
rect 14655 -150 14721 -138
rect 14751 138 14817 150
rect 14751 -138 14767 138
rect 14801 -138 14817 138
rect 14751 -150 14817 -138
rect 14847 138 14913 150
rect 14847 -138 14863 138
rect 14897 -138 14913 138
rect 14847 -150 14913 -138
rect 14943 138 15009 150
rect 14943 -138 14959 138
rect 14993 -138 15009 138
rect 14943 -150 15009 -138
rect 15039 138 15105 150
rect 15039 -138 15055 138
rect 15089 -138 15105 138
rect 15039 -150 15105 -138
rect 15135 138 15201 150
rect 15135 -138 15151 138
rect 15185 -138 15201 138
rect 15135 -150 15201 -138
rect 15231 138 15297 150
rect 15231 -138 15247 138
rect 15281 -138 15297 138
rect 15231 -150 15297 -138
rect 15327 138 15393 150
rect 15327 -138 15343 138
rect 15377 -138 15393 138
rect 15327 -150 15393 -138
rect 15423 138 15489 150
rect 15423 -138 15439 138
rect 15473 -138 15489 138
rect 15423 -150 15489 -138
rect 15519 138 15585 150
rect 15519 -138 15535 138
rect 15569 -138 15585 138
rect 15519 -150 15585 -138
rect 15615 138 15681 150
rect 15615 -138 15631 138
rect 15665 -138 15681 138
rect 15615 -150 15681 -138
rect 15711 138 15777 150
rect 15711 -138 15727 138
rect 15761 -138 15777 138
rect 15711 -150 15777 -138
rect 15807 138 15873 150
rect 15807 -138 15823 138
rect 15857 -138 15873 138
rect 15807 -150 15873 -138
rect 15903 138 15969 150
rect 15903 -138 15919 138
rect 15953 -138 15969 138
rect 15903 -150 15969 -138
rect 15999 138 16065 150
rect 15999 -138 16015 138
rect 16049 -138 16065 138
rect 15999 -150 16065 -138
rect 16095 138 16161 150
rect 16095 -138 16111 138
rect 16145 -138 16161 138
rect 16095 -150 16161 -138
rect 16191 138 16257 150
rect 16191 -138 16207 138
rect 16241 -138 16257 138
rect 16191 -150 16257 -138
rect 16287 138 16353 150
rect 16287 -138 16303 138
rect 16337 -138 16353 138
rect 16287 -150 16353 -138
rect 16383 138 16449 150
rect 16383 -138 16399 138
rect 16433 -138 16449 138
rect 16383 -150 16449 -138
rect 16479 138 16545 150
rect 16479 -138 16495 138
rect 16529 -138 16545 138
rect 16479 -150 16545 -138
rect 16575 138 16641 150
rect 16575 -138 16591 138
rect 16625 -138 16641 138
rect 16575 -150 16641 -138
rect 16671 138 16737 150
rect 16671 -138 16687 138
rect 16721 -138 16737 138
rect 16671 -150 16737 -138
rect 16767 138 16833 150
rect 16767 -138 16783 138
rect 16817 -138 16833 138
rect 16767 -150 16833 -138
rect 16863 138 16929 150
rect 16863 -138 16879 138
rect 16913 -138 16929 138
rect 16863 -150 16929 -138
rect 16959 138 17025 150
rect 16959 -138 16975 138
rect 17009 -138 17025 138
rect 16959 -150 17025 -138
rect 17055 138 17121 150
rect 17055 -138 17071 138
rect 17105 -138 17121 138
rect 17055 -150 17121 -138
rect 17151 138 17217 150
rect 17151 -138 17167 138
rect 17201 -138 17217 138
rect 17151 -150 17217 -138
rect 17247 138 17313 150
rect 17247 -138 17263 138
rect 17297 -138 17313 138
rect 17247 -150 17313 -138
rect 17343 138 17409 150
rect 17343 -138 17359 138
rect 17393 -138 17409 138
rect 17343 -150 17409 -138
rect 17439 138 17505 150
rect 17439 -138 17455 138
rect 17489 -138 17505 138
rect 17439 -150 17505 -138
rect 17535 138 17601 150
rect 17535 -138 17551 138
rect 17585 -138 17601 138
rect 17535 -150 17601 -138
rect 17631 138 17697 150
rect 17631 -138 17647 138
rect 17681 -138 17697 138
rect 17631 -150 17697 -138
rect 17727 138 17793 150
rect 17727 -138 17743 138
rect 17777 -138 17793 138
rect 17727 -150 17793 -138
rect 17823 138 17889 150
rect 17823 -138 17839 138
rect 17873 -138 17889 138
rect 17823 -150 17889 -138
rect 17919 138 17985 150
rect 17919 -138 17935 138
rect 17969 -138 17985 138
rect 17919 -150 17985 -138
rect 18015 138 18081 150
rect 18015 -138 18031 138
rect 18065 -138 18081 138
rect 18015 -150 18081 -138
rect 18111 138 18177 150
rect 18111 -138 18127 138
rect 18161 -138 18177 138
rect 18111 -150 18177 -138
rect 18207 138 18273 150
rect 18207 -138 18223 138
rect 18257 -138 18273 138
rect 18207 -150 18273 -138
rect 18303 138 18369 150
rect 18303 -138 18319 138
rect 18353 -138 18369 138
rect 18303 -150 18369 -138
rect 18399 138 18465 150
rect 18399 -138 18415 138
rect 18449 -138 18465 138
rect 18399 -150 18465 -138
rect 18495 138 18561 150
rect 18495 -138 18511 138
rect 18545 -138 18561 138
rect 18495 -150 18561 -138
rect 18591 138 18657 150
rect 18591 -138 18607 138
rect 18641 -138 18657 138
rect 18591 -150 18657 -138
rect 18687 138 18753 150
rect 18687 -138 18703 138
rect 18737 -138 18753 138
rect 18687 -150 18753 -138
rect 18783 138 18849 150
rect 18783 -138 18799 138
rect 18833 -138 18849 138
rect 18783 -150 18849 -138
rect 18879 138 18945 150
rect 18879 -138 18895 138
rect 18929 -138 18945 138
rect 18879 -150 18945 -138
rect 18975 138 19041 150
rect 18975 -138 18991 138
rect 19025 -138 19041 138
rect 18975 -150 19041 -138
rect 19071 138 19137 150
rect 19071 -138 19087 138
rect 19121 -138 19137 138
rect 19071 -150 19137 -138
rect 19167 138 19229 150
rect 19167 -138 19183 138
rect 19217 -138 19229 138
rect 19167 -150 19229 -138
<< ndiffc >>
rect -19217 -138 -19183 138
rect -19121 -138 -19087 138
rect -19025 -138 -18991 138
rect -18929 -138 -18895 138
rect -18833 -138 -18799 138
rect -18737 -138 -18703 138
rect -18641 -138 -18607 138
rect -18545 -138 -18511 138
rect -18449 -138 -18415 138
rect -18353 -138 -18319 138
rect -18257 -138 -18223 138
rect -18161 -138 -18127 138
rect -18065 -138 -18031 138
rect -17969 -138 -17935 138
rect -17873 -138 -17839 138
rect -17777 -138 -17743 138
rect -17681 -138 -17647 138
rect -17585 -138 -17551 138
rect -17489 -138 -17455 138
rect -17393 -138 -17359 138
rect -17297 -138 -17263 138
rect -17201 -138 -17167 138
rect -17105 -138 -17071 138
rect -17009 -138 -16975 138
rect -16913 -138 -16879 138
rect -16817 -138 -16783 138
rect -16721 -138 -16687 138
rect -16625 -138 -16591 138
rect -16529 -138 -16495 138
rect -16433 -138 -16399 138
rect -16337 -138 -16303 138
rect -16241 -138 -16207 138
rect -16145 -138 -16111 138
rect -16049 -138 -16015 138
rect -15953 -138 -15919 138
rect -15857 -138 -15823 138
rect -15761 -138 -15727 138
rect -15665 -138 -15631 138
rect -15569 -138 -15535 138
rect -15473 -138 -15439 138
rect -15377 -138 -15343 138
rect -15281 -138 -15247 138
rect -15185 -138 -15151 138
rect -15089 -138 -15055 138
rect -14993 -138 -14959 138
rect -14897 -138 -14863 138
rect -14801 -138 -14767 138
rect -14705 -138 -14671 138
rect -14609 -138 -14575 138
rect -14513 -138 -14479 138
rect -14417 -138 -14383 138
rect -14321 -138 -14287 138
rect -14225 -138 -14191 138
rect -14129 -138 -14095 138
rect -14033 -138 -13999 138
rect -13937 -138 -13903 138
rect -13841 -138 -13807 138
rect -13745 -138 -13711 138
rect -13649 -138 -13615 138
rect -13553 -138 -13519 138
rect -13457 -138 -13423 138
rect -13361 -138 -13327 138
rect -13265 -138 -13231 138
rect -13169 -138 -13135 138
rect -13073 -138 -13039 138
rect -12977 -138 -12943 138
rect -12881 -138 -12847 138
rect -12785 -138 -12751 138
rect -12689 -138 -12655 138
rect -12593 -138 -12559 138
rect -12497 -138 -12463 138
rect -12401 -138 -12367 138
rect -12305 -138 -12271 138
rect -12209 -138 -12175 138
rect -12113 -138 -12079 138
rect -12017 -138 -11983 138
rect -11921 -138 -11887 138
rect -11825 -138 -11791 138
rect -11729 -138 -11695 138
rect -11633 -138 -11599 138
rect -11537 -138 -11503 138
rect -11441 -138 -11407 138
rect -11345 -138 -11311 138
rect -11249 -138 -11215 138
rect -11153 -138 -11119 138
rect -11057 -138 -11023 138
rect -10961 -138 -10927 138
rect -10865 -138 -10831 138
rect -10769 -138 -10735 138
rect -10673 -138 -10639 138
rect -10577 -138 -10543 138
rect -10481 -138 -10447 138
rect -10385 -138 -10351 138
rect -10289 -138 -10255 138
rect -10193 -138 -10159 138
rect -10097 -138 -10063 138
rect -10001 -138 -9967 138
rect -9905 -138 -9871 138
rect -9809 -138 -9775 138
rect -9713 -138 -9679 138
rect -9617 -138 -9583 138
rect -9521 -138 -9487 138
rect -9425 -138 -9391 138
rect -9329 -138 -9295 138
rect -9233 -138 -9199 138
rect -9137 -138 -9103 138
rect -9041 -138 -9007 138
rect -8945 -138 -8911 138
rect -8849 -138 -8815 138
rect -8753 -138 -8719 138
rect -8657 -138 -8623 138
rect -8561 -138 -8527 138
rect -8465 -138 -8431 138
rect -8369 -138 -8335 138
rect -8273 -138 -8239 138
rect -8177 -138 -8143 138
rect -8081 -138 -8047 138
rect -7985 -138 -7951 138
rect -7889 -138 -7855 138
rect -7793 -138 -7759 138
rect -7697 -138 -7663 138
rect -7601 -138 -7567 138
rect -7505 -138 -7471 138
rect -7409 -138 -7375 138
rect -7313 -138 -7279 138
rect -7217 -138 -7183 138
rect -7121 -138 -7087 138
rect -7025 -138 -6991 138
rect -6929 -138 -6895 138
rect -6833 -138 -6799 138
rect -6737 -138 -6703 138
rect -6641 -138 -6607 138
rect -6545 -138 -6511 138
rect -6449 -138 -6415 138
rect -6353 -138 -6319 138
rect -6257 -138 -6223 138
rect -6161 -138 -6127 138
rect -6065 -138 -6031 138
rect -5969 -138 -5935 138
rect -5873 -138 -5839 138
rect -5777 -138 -5743 138
rect -5681 -138 -5647 138
rect -5585 -138 -5551 138
rect -5489 -138 -5455 138
rect -5393 -138 -5359 138
rect -5297 -138 -5263 138
rect -5201 -138 -5167 138
rect -5105 -138 -5071 138
rect -5009 -138 -4975 138
rect -4913 -138 -4879 138
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
rect 4879 -138 4913 138
rect 4975 -138 5009 138
rect 5071 -138 5105 138
rect 5167 -138 5201 138
rect 5263 -138 5297 138
rect 5359 -138 5393 138
rect 5455 -138 5489 138
rect 5551 -138 5585 138
rect 5647 -138 5681 138
rect 5743 -138 5777 138
rect 5839 -138 5873 138
rect 5935 -138 5969 138
rect 6031 -138 6065 138
rect 6127 -138 6161 138
rect 6223 -138 6257 138
rect 6319 -138 6353 138
rect 6415 -138 6449 138
rect 6511 -138 6545 138
rect 6607 -138 6641 138
rect 6703 -138 6737 138
rect 6799 -138 6833 138
rect 6895 -138 6929 138
rect 6991 -138 7025 138
rect 7087 -138 7121 138
rect 7183 -138 7217 138
rect 7279 -138 7313 138
rect 7375 -138 7409 138
rect 7471 -138 7505 138
rect 7567 -138 7601 138
rect 7663 -138 7697 138
rect 7759 -138 7793 138
rect 7855 -138 7889 138
rect 7951 -138 7985 138
rect 8047 -138 8081 138
rect 8143 -138 8177 138
rect 8239 -138 8273 138
rect 8335 -138 8369 138
rect 8431 -138 8465 138
rect 8527 -138 8561 138
rect 8623 -138 8657 138
rect 8719 -138 8753 138
rect 8815 -138 8849 138
rect 8911 -138 8945 138
rect 9007 -138 9041 138
rect 9103 -138 9137 138
rect 9199 -138 9233 138
rect 9295 -138 9329 138
rect 9391 -138 9425 138
rect 9487 -138 9521 138
rect 9583 -138 9617 138
rect 9679 -138 9713 138
rect 9775 -138 9809 138
rect 9871 -138 9905 138
rect 9967 -138 10001 138
rect 10063 -138 10097 138
rect 10159 -138 10193 138
rect 10255 -138 10289 138
rect 10351 -138 10385 138
rect 10447 -138 10481 138
rect 10543 -138 10577 138
rect 10639 -138 10673 138
rect 10735 -138 10769 138
rect 10831 -138 10865 138
rect 10927 -138 10961 138
rect 11023 -138 11057 138
rect 11119 -138 11153 138
rect 11215 -138 11249 138
rect 11311 -138 11345 138
rect 11407 -138 11441 138
rect 11503 -138 11537 138
rect 11599 -138 11633 138
rect 11695 -138 11729 138
rect 11791 -138 11825 138
rect 11887 -138 11921 138
rect 11983 -138 12017 138
rect 12079 -138 12113 138
rect 12175 -138 12209 138
rect 12271 -138 12305 138
rect 12367 -138 12401 138
rect 12463 -138 12497 138
rect 12559 -138 12593 138
rect 12655 -138 12689 138
rect 12751 -138 12785 138
rect 12847 -138 12881 138
rect 12943 -138 12977 138
rect 13039 -138 13073 138
rect 13135 -138 13169 138
rect 13231 -138 13265 138
rect 13327 -138 13361 138
rect 13423 -138 13457 138
rect 13519 -138 13553 138
rect 13615 -138 13649 138
rect 13711 -138 13745 138
rect 13807 -138 13841 138
rect 13903 -138 13937 138
rect 13999 -138 14033 138
rect 14095 -138 14129 138
rect 14191 -138 14225 138
rect 14287 -138 14321 138
rect 14383 -138 14417 138
rect 14479 -138 14513 138
rect 14575 -138 14609 138
rect 14671 -138 14705 138
rect 14767 -138 14801 138
rect 14863 -138 14897 138
rect 14959 -138 14993 138
rect 15055 -138 15089 138
rect 15151 -138 15185 138
rect 15247 -138 15281 138
rect 15343 -138 15377 138
rect 15439 -138 15473 138
rect 15535 -138 15569 138
rect 15631 -138 15665 138
rect 15727 -138 15761 138
rect 15823 -138 15857 138
rect 15919 -138 15953 138
rect 16015 -138 16049 138
rect 16111 -138 16145 138
rect 16207 -138 16241 138
rect 16303 -138 16337 138
rect 16399 -138 16433 138
rect 16495 -138 16529 138
rect 16591 -138 16625 138
rect 16687 -138 16721 138
rect 16783 -138 16817 138
rect 16879 -138 16913 138
rect 16975 -138 17009 138
rect 17071 -138 17105 138
rect 17167 -138 17201 138
rect 17263 -138 17297 138
rect 17359 -138 17393 138
rect 17455 -138 17489 138
rect 17551 -138 17585 138
rect 17647 -138 17681 138
rect 17743 -138 17777 138
rect 17839 -138 17873 138
rect 17935 -138 17969 138
rect 18031 -138 18065 138
rect 18127 -138 18161 138
rect 18223 -138 18257 138
rect 18319 -138 18353 138
rect 18415 -138 18449 138
rect 18511 -138 18545 138
rect 18607 -138 18641 138
rect 18703 -138 18737 138
rect 18799 -138 18833 138
rect 18895 -138 18929 138
rect 18991 -138 19025 138
rect 19087 -138 19121 138
rect 19183 -138 19217 138
<< psubdiff >>
rect -19331 290 -19235 324
rect 19235 290 19331 324
rect -19331 228 -19297 290
rect 19297 228 19331 290
rect -19331 -290 -19297 -228
rect 19297 -290 19331 -228
rect -19331 -324 -19235 -290
rect 19235 -324 19331 -290
<< psubdiffcont >>
rect -19235 290 19235 324
rect -19331 -228 -19297 228
rect 19297 -228 19331 228
rect -19235 -324 19235 -290
<< poly >>
rect -19089 222 -19023 238
rect -19089 188 -19073 222
rect -19039 188 -19023 222
rect -19167 150 -19137 176
rect -19089 172 -19023 188
rect -18897 222 -18831 238
rect -18897 188 -18881 222
rect -18847 188 -18831 222
rect -19071 150 -19041 172
rect -18975 150 -18945 176
rect -18897 172 -18831 188
rect -18705 222 -18639 238
rect -18705 188 -18689 222
rect -18655 188 -18639 222
rect -18879 150 -18849 172
rect -18783 150 -18753 176
rect -18705 172 -18639 188
rect -18513 222 -18447 238
rect -18513 188 -18497 222
rect -18463 188 -18447 222
rect -18687 150 -18657 172
rect -18591 150 -18561 176
rect -18513 172 -18447 188
rect -18321 222 -18255 238
rect -18321 188 -18305 222
rect -18271 188 -18255 222
rect -18495 150 -18465 172
rect -18399 150 -18369 176
rect -18321 172 -18255 188
rect -18129 222 -18063 238
rect -18129 188 -18113 222
rect -18079 188 -18063 222
rect -18303 150 -18273 172
rect -18207 150 -18177 176
rect -18129 172 -18063 188
rect -17937 222 -17871 238
rect -17937 188 -17921 222
rect -17887 188 -17871 222
rect -18111 150 -18081 172
rect -18015 150 -17985 176
rect -17937 172 -17871 188
rect -17745 222 -17679 238
rect -17745 188 -17729 222
rect -17695 188 -17679 222
rect -17919 150 -17889 172
rect -17823 150 -17793 176
rect -17745 172 -17679 188
rect -17553 222 -17487 238
rect -17553 188 -17537 222
rect -17503 188 -17487 222
rect -17727 150 -17697 172
rect -17631 150 -17601 176
rect -17553 172 -17487 188
rect -17361 222 -17295 238
rect -17361 188 -17345 222
rect -17311 188 -17295 222
rect -17535 150 -17505 172
rect -17439 150 -17409 176
rect -17361 172 -17295 188
rect -17169 222 -17103 238
rect -17169 188 -17153 222
rect -17119 188 -17103 222
rect -17343 150 -17313 172
rect -17247 150 -17217 176
rect -17169 172 -17103 188
rect -16977 222 -16911 238
rect -16977 188 -16961 222
rect -16927 188 -16911 222
rect -17151 150 -17121 172
rect -17055 150 -17025 176
rect -16977 172 -16911 188
rect -16785 222 -16719 238
rect -16785 188 -16769 222
rect -16735 188 -16719 222
rect -16959 150 -16929 172
rect -16863 150 -16833 176
rect -16785 172 -16719 188
rect -16593 222 -16527 238
rect -16593 188 -16577 222
rect -16543 188 -16527 222
rect -16767 150 -16737 172
rect -16671 150 -16641 176
rect -16593 172 -16527 188
rect -16401 222 -16335 238
rect -16401 188 -16385 222
rect -16351 188 -16335 222
rect -16575 150 -16545 172
rect -16479 150 -16449 176
rect -16401 172 -16335 188
rect -16209 222 -16143 238
rect -16209 188 -16193 222
rect -16159 188 -16143 222
rect -16383 150 -16353 172
rect -16287 150 -16257 176
rect -16209 172 -16143 188
rect -16017 222 -15951 238
rect -16017 188 -16001 222
rect -15967 188 -15951 222
rect -16191 150 -16161 172
rect -16095 150 -16065 176
rect -16017 172 -15951 188
rect -15825 222 -15759 238
rect -15825 188 -15809 222
rect -15775 188 -15759 222
rect -15999 150 -15969 172
rect -15903 150 -15873 176
rect -15825 172 -15759 188
rect -15633 222 -15567 238
rect -15633 188 -15617 222
rect -15583 188 -15567 222
rect -15807 150 -15777 172
rect -15711 150 -15681 176
rect -15633 172 -15567 188
rect -15441 222 -15375 238
rect -15441 188 -15425 222
rect -15391 188 -15375 222
rect -15615 150 -15585 172
rect -15519 150 -15489 176
rect -15441 172 -15375 188
rect -15249 222 -15183 238
rect -15249 188 -15233 222
rect -15199 188 -15183 222
rect -15423 150 -15393 172
rect -15327 150 -15297 176
rect -15249 172 -15183 188
rect -15057 222 -14991 238
rect -15057 188 -15041 222
rect -15007 188 -14991 222
rect -15231 150 -15201 172
rect -15135 150 -15105 176
rect -15057 172 -14991 188
rect -14865 222 -14799 238
rect -14865 188 -14849 222
rect -14815 188 -14799 222
rect -15039 150 -15009 172
rect -14943 150 -14913 176
rect -14865 172 -14799 188
rect -14673 222 -14607 238
rect -14673 188 -14657 222
rect -14623 188 -14607 222
rect -14847 150 -14817 172
rect -14751 150 -14721 176
rect -14673 172 -14607 188
rect -14481 222 -14415 238
rect -14481 188 -14465 222
rect -14431 188 -14415 222
rect -14655 150 -14625 172
rect -14559 150 -14529 176
rect -14481 172 -14415 188
rect -14289 222 -14223 238
rect -14289 188 -14273 222
rect -14239 188 -14223 222
rect -14463 150 -14433 172
rect -14367 150 -14337 176
rect -14289 172 -14223 188
rect -14097 222 -14031 238
rect -14097 188 -14081 222
rect -14047 188 -14031 222
rect -14271 150 -14241 172
rect -14175 150 -14145 176
rect -14097 172 -14031 188
rect -13905 222 -13839 238
rect -13905 188 -13889 222
rect -13855 188 -13839 222
rect -14079 150 -14049 172
rect -13983 150 -13953 176
rect -13905 172 -13839 188
rect -13713 222 -13647 238
rect -13713 188 -13697 222
rect -13663 188 -13647 222
rect -13887 150 -13857 172
rect -13791 150 -13761 176
rect -13713 172 -13647 188
rect -13521 222 -13455 238
rect -13521 188 -13505 222
rect -13471 188 -13455 222
rect -13695 150 -13665 172
rect -13599 150 -13569 176
rect -13521 172 -13455 188
rect -13329 222 -13263 238
rect -13329 188 -13313 222
rect -13279 188 -13263 222
rect -13503 150 -13473 172
rect -13407 150 -13377 176
rect -13329 172 -13263 188
rect -13137 222 -13071 238
rect -13137 188 -13121 222
rect -13087 188 -13071 222
rect -13311 150 -13281 172
rect -13215 150 -13185 176
rect -13137 172 -13071 188
rect -12945 222 -12879 238
rect -12945 188 -12929 222
rect -12895 188 -12879 222
rect -13119 150 -13089 172
rect -13023 150 -12993 176
rect -12945 172 -12879 188
rect -12753 222 -12687 238
rect -12753 188 -12737 222
rect -12703 188 -12687 222
rect -12927 150 -12897 172
rect -12831 150 -12801 176
rect -12753 172 -12687 188
rect -12561 222 -12495 238
rect -12561 188 -12545 222
rect -12511 188 -12495 222
rect -12735 150 -12705 172
rect -12639 150 -12609 176
rect -12561 172 -12495 188
rect -12369 222 -12303 238
rect -12369 188 -12353 222
rect -12319 188 -12303 222
rect -12543 150 -12513 172
rect -12447 150 -12417 176
rect -12369 172 -12303 188
rect -12177 222 -12111 238
rect -12177 188 -12161 222
rect -12127 188 -12111 222
rect -12351 150 -12321 172
rect -12255 150 -12225 176
rect -12177 172 -12111 188
rect -11985 222 -11919 238
rect -11985 188 -11969 222
rect -11935 188 -11919 222
rect -12159 150 -12129 172
rect -12063 150 -12033 176
rect -11985 172 -11919 188
rect -11793 222 -11727 238
rect -11793 188 -11777 222
rect -11743 188 -11727 222
rect -11967 150 -11937 172
rect -11871 150 -11841 176
rect -11793 172 -11727 188
rect -11601 222 -11535 238
rect -11601 188 -11585 222
rect -11551 188 -11535 222
rect -11775 150 -11745 172
rect -11679 150 -11649 176
rect -11601 172 -11535 188
rect -11409 222 -11343 238
rect -11409 188 -11393 222
rect -11359 188 -11343 222
rect -11583 150 -11553 172
rect -11487 150 -11457 176
rect -11409 172 -11343 188
rect -11217 222 -11151 238
rect -11217 188 -11201 222
rect -11167 188 -11151 222
rect -11391 150 -11361 172
rect -11295 150 -11265 176
rect -11217 172 -11151 188
rect -11025 222 -10959 238
rect -11025 188 -11009 222
rect -10975 188 -10959 222
rect -11199 150 -11169 172
rect -11103 150 -11073 176
rect -11025 172 -10959 188
rect -10833 222 -10767 238
rect -10833 188 -10817 222
rect -10783 188 -10767 222
rect -11007 150 -10977 172
rect -10911 150 -10881 176
rect -10833 172 -10767 188
rect -10641 222 -10575 238
rect -10641 188 -10625 222
rect -10591 188 -10575 222
rect -10815 150 -10785 172
rect -10719 150 -10689 176
rect -10641 172 -10575 188
rect -10449 222 -10383 238
rect -10449 188 -10433 222
rect -10399 188 -10383 222
rect -10623 150 -10593 172
rect -10527 150 -10497 176
rect -10449 172 -10383 188
rect -10257 222 -10191 238
rect -10257 188 -10241 222
rect -10207 188 -10191 222
rect -10431 150 -10401 172
rect -10335 150 -10305 176
rect -10257 172 -10191 188
rect -10065 222 -9999 238
rect -10065 188 -10049 222
rect -10015 188 -9999 222
rect -10239 150 -10209 172
rect -10143 150 -10113 176
rect -10065 172 -9999 188
rect -9873 222 -9807 238
rect -9873 188 -9857 222
rect -9823 188 -9807 222
rect -10047 150 -10017 172
rect -9951 150 -9921 176
rect -9873 172 -9807 188
rect -9681 222 -9615 238
rect -9681 188 -9665 222
rect -9631 188 -9615 222
rect -9855 150 -9825 172
rect -9759 150 -9729 176
rect -9681 172 -9615 188
rect -9489 222 -9423 238
rect -9489 188 -9473 222
rect -9439 188 -9423 222
rect -9663 150 -9633 172
rect -9567 150 -9537 176
rect -9489 172 -9423 188
rect -9297 222 -9231 238
rect -9297 188 -9281 222
rect -9247 188 -9231 222
rect -9471 150 -9441 172
rect -9375 150 -9345 176
rect -9297 172 -9231 188
rect -9105 222 -9039 238
rect -9105 188 -9089 222
rect -9055 188 -9039 222
rect -9279 150 -9249 172
rect -9183 150 -9153 176
rect -9105 172 -9039 188
rect -8913 222 -8847 238
rect -8913 188 -8897 222
rect -8863 188 -8847 222
rect -9087 150 -9057 172
rect -8991 150 -8961 176
rect -8913 172 -8847 188
rect -8721 222 -8655 238
rect -8721 188 -8705 222
rect -8671 188 -8655 222
rect -8895 150 -8865 172
rect -8799 150 -8769 176
rect -8721 172 -8655 188
rect -8529 222 -8463 238
rect -8529 188 -8513 222
rect -8479 188 -8463 222
rect -8703 150 -8673 172
rect -8607 150 -8577 176
rect -8529 172 -8463 188
rect -8337 222 -8271 238
rect -8337 188 -8321 222
rect -8287 188 -8271 222
rect -8511 150 -8481 172
rect -8415 150 -8385 176
rect -8337 172 -8271 188
rect -8145 222 -8079 238
rect -8145 188 -8129 222
rect -8095 188 -8079 222
rect -8319 150 -8289 172
rect -8223 150 -8193 176
rect -8145 172 -8079 188
rect -7953 222 -7887 238
rect -7953 188 -7937 222
rect -7903 188 -7887 222
rect -8127 150 -8097 172
rect -8031 150 -8001 176
rect -7953 172 -7887 188
rect -7761 222 -7695 238
rect -7761 188 -7745 222
rect -7711 188 -7695 222
rect -7935 150 -7905 172
rect -7839 150 -7809 176
rect -7761 172 -7695 188
rect -7569 222 -7503 238
rect -7569 188 -7553 222
rect -7519 188 -7503 222
rect -7743 150 -7713 172
rect -7647 150 -7617 176
rect -7569 172 -7503 188
rect -7377 222 -7311 238
rect -7377 188 -7361 222
rect -7327 188 -7311 222
rect -7551 150 -7521 172
rect -7455 150 -7425 176
rect -7377 172 -7311 188
rect -7185 222 -7119 238
rect -7185 188 -7169 222
rect -7135 188 -7119 222
rect -7359 150 -7329 172
rect -7263 150 -7233 176
rect -7185 172 -7119 188
rect -6993 222 -6927 238
rect -6993 188 -6977 222
rect -6943 188 -6927 222
rect -7167 150 -7137 172
rect -7071 150 -7041 176
rect -6993 172 -6927 188
rect -6801 222 -6735 238
rect -6801 188 -6785 222
rect -6751 188 -6735 222
rect -6975 150 -6945 172
rect -6879 150 -6849 176
rect -6801 172 -6735 188
rect -6609 222 -6543 238
rect -6609 188 -6593 222
rect -6559 188 -6543 222
rect -6783 150 -6753 172
rect -6687 150 -6657 176
rect -6609 172 -6543 188
rect -6417 222 -6351 238
rect -6417 188 -6401 222
rect -6367 188 -6351 222
rect -6591 150 -6561 172
rect -6495 150 -6465 176
rect -6417 172 -6351 188
rect -6225 222 -6159 238
rect -6225 188 -6209 222
rect -6175 188 -6159 222
rect -6399 150 -6369 172
rect -6303 150 -6273 176
rect -6225 172 -6159 188
rect -6033 222 -5967 238
rect -6033 188 -6017 222
rect -5983 188 -5967 222
rect -6207 150 -6177 172
rect -6111 150 -6081 176
rect -6033 172 -5967 188
rect -5841 222 -5775 238
rect -5841 188 -5825 222
rect -5791 188 -5775 222
rect -6015 150 -5985 172
rect -5919 150 -5889 176
rect -5841 172 -5775 188
rect -5649 222 -5583 238
rect -5649 188 -5633 222
rect -5599 188 -5583 222
rect -5823 150 -5793 172
rect -5727 150 -5697 176
rect -5649 172 -5583 188
rect -5457 222 -5391 238
rect -5457 188 -5441 222
rect -5407 188 -5391 222
rect -5631 150 -5601 172
rect -5535 150 -5505 176
rect -5457 172 -5391 188
rect -5265 222 -5199 238
rect -5265 188 -5249 222
rect -5215 188 -5199 222
rect -5439 150 -5409 172
rect -5343 150 -5313 176
rect -5265 172 -5199 188
rect -5073 222 -5007 238
rect -5073 188 -5057 222
rect -5023 188 -5007 222
rect -5247 150 -5217 172
rect -5151 150 -5121 176
rect -5073 172 -5007 188
rect -4881 222 -4815 238
rect -4881 188 -4865 222
rect -4831 188 -4815 222
rect -5055 150 -5025 172
rect -4959 150 -4929 176
rect -4881 172 -4815 188
rect -4689 222 -4623 238
rect -4689 188 -4673 222
rect -4639 188 -4623 222
rect -4863 150 -4833 172
rect -4767 150 -4737 176
rect -4689 172 -4623 188
rect -4497 222 -4431 238
rect -4497 188 -4481 222
rect -4447 188 -4431 222
rect -4671 150 -4641 172
rect -4575 150 -4545 176
rect -4497 172 -4431 188
rect -4305 222 -4239 238
rect -4305 188 -4289 222
rect -4255 188 -4239 222
rect -4479 150 -4449 172
rect -4383 150 -4353 176
rect -4305 172 -4239 188
rect -4113 222 -4047 238
rect -4113 188 -4097 222
rect -4063 188 -4047 222
rect -4287 150 -4257 172
rect -4191 150 -4161 176
rect -4113 172 -4047 188
rect -3921 222 -3855 238
rect -3921 188 -3905 222
rect -3871 188 -3855 222
rect -4095 150 -4065 172
rect -3999 150 -3969 176
rect -3921 172 -3855 188
rect -3729 222 -3663 238
rect -3729 188 -3713 222
rect -3679 188 -3663 222
rect -3903 150 -3873 172
rect -3807 150 -3777 176
rect -3729 172 -3663 188
rect -3537 222 -3471 238
rect -3537 188 -3521 222
rect -3487 188 -3471 222
rect -3711 150 -3681 172
rect -3615 150 -3585 176
rect -3537 172 -3471 188
rect -3345 222 -3279 238
rect -3345 188 -3329 222
rect -3295 188 -3279 222
rect -3519 150 -3489 172
rect -3423 150 -3393 176
rect -3345 172 -3279 188
rect -3153 222 -3087 238
rect -3153 188 -3137 222
rect -3103 188 -3087 222
rect -3327 150 -3297 172
rect -3231 150 -3201 176
rect -3153 172 -3087 188
rect -2961 222 -2895 238
rect -2961 188 -2945 222
rect -2911 188 -2895 222
rect -3135 150 -3105 172
rect -3039 150 -3009 176
rect -2961 172 -2895 188
rect -2769 222 -2703 238
rect -2769 188 -2753 222
rect -2719 188 -2703 222
rect -2943 150 -2913 172
rect -2847 150 -2817 176
rect -2769 172 -2703 188
rect -2577 222 -2511 238
rect -2577 188 -2561 222
rect -2527 188 -2511 222
rect -2751 150 -2721 172
rect -2655 150 -2625 176
rect -2577 172 -2511 188
rect -2385 222 -2319 238
rect -2385 188 -2369 222
rect -2335 188 -2319 222
rect -2559 150 -2529 172
rect -2463 150 -2433 176
rect -2385 172 -2319 188
rect -2193 222 -2127 238
rect -2193 188 -2177 222
rect -2143 188 -2127 222
rect -2367 150 -2337 172
rect -2271 150 -2241 176
rect -2193 172 -2127 188
rect -2001 222 -1935 238
rect -2001 188 -1985 222
rect -1951 188 -1935 222
rect -2175 150 -2145 172
rect -2079 150 -2049 176
rect -2001 172 -1935 188
rect -1809 222 -1743 238
rect -1809 188 -1793 222
rect -1759 188 -1743 222
rect -1983 150 -1953 172
rect -1887 150 -1857 176
rect -1809 172 -1743 188
rect -1617 222 -1551 238
rect -1617 188 -1601 222
rect -1567 188 -1551 222
rect -1791 150 -1761 172
rect -1695 150 -1665 176
rect -1617 172 -1551 188
rect -1425 222 -1359 238
rect -1425 188 -1409 222
rect -1375 188 -1359 222
rect -1599 150 -1569 172
rect -1503 150 -1473 176
rect -1425 172 -1359 188
rect -1233 222 -1167 238
rect -1233 188 -1217 222
rect -1183 188 -1167 222
rect -1407 150 -1377 172
rect -1311 150 -1281 176
rect -1233 172 -1167 188
rect -1041 222 -975 238
rect -1041 188 -1025 222
rect -991 188 -975 222
rect -1215 150 -1185 172
rect -1119 150 -1089 176
rect -1041 172 -975 188
rect -849 222 -783 238
rect -849 188 -833 222
rect -799 188 -783 222
rect -1023 150 -993 172
rect -927 150 -897 176
rect -849 172 -783 188
rect -657 222 -591 238
rect -657 188 -641 222
rect -607 188 -591 222
rect -831 150 -801 172
rect -735 150 -705 176
rect -657 172 -591 188
rect -465 222 -399 238
rect -465 188 -449 222
rect -415 188 -399 222
rect -639 150 -609 172
rect -543 150 -513 176
rect -465 172 -399 188
rect -273 222 -207 238
rect -273 188 -257 222
rect -223 188 -207 222
rect -447 150 -417 172
rect -351 150 -321 176
rect -273 172 -207 188
rect -81 222 -15 238
rect -81 188 -65 222
rect -31 188 -15 222
rect -255 150 -225 172
rect -159 150 -129 176
rect -81 172 -15 188
rect 111 222 177 238
rect 111 188 127 222
rect 161 188 177 222
rect -63 150 -33 172
rect 33 150 63 176
rect 111 172 177 188
rect 303 222 369 238
rect 303 188 319 222
rect 353 188 369 222
rect 129 150 159 172
rect 225 150 255 176
rect 303 172 369 188
rect 495 222 561 238
rect 495 188 511 222
rect 545 188 561 222
rect 321 150 351 172
rect 417 150 447 176
rect 495 172 561 188
rect 687 222 753 238
rect 687 188 703 222
rect 737 188 753 222
rect 513 150 543 172
rect 609 150 639 176
rect 687 172 753 188
rect 879 222 945 238
rect 879 188 895 222
rect 929 188 945 222
rect 705 150 735 172
rect 801 150 831 176
rect 879 172 945 188
rect 1071 222 1137 238
rect 1071 188 1087 222
rect 1121 188 1137 222
rect 897 150 927 172
rect 993 150 1023 176
rect 1071 172 1137 188
rect 1263 222 1329 238
rect 1263 188 1279 222
rect 1313 188 1329 222
rect 1089 150 1119 172
rect 1185 150 1215 176
rect 1263 172 1329 188
rect 1455 222 1521 238
rect 1455 188 1471 222
rect 1505 188 1521 222
rect 1281 150 1311 172
rect 1377 150 1407 176
rect 1455 172 1521 188
rect 1647 222 1713 238
rect 1647 188 1663 222
rect 1697 188 1713 222
rect 1473 150 1503 172
rect 1569 150 1599 176
rect 1647 172 1713 188
rect 1839 222 1905 238
rect 1839 188 1855 222
rect 1889 188 1905 222
rect 1665 150 1695 172
rect 1761 150 1791 176
rect 1839 172 1905 188
rect 2031 222 2097 238
rect 2031 188 2047 222
rect 2081 188 2097 222
rect 1857 150 1887 172
rect 1953 150 1983 176
rect 2031 172 2097 188
rect 2223 222 2289 238
rect 2223 188 2239 222
rect 2273 188 2289 222
rect 2049 150 2079 172
rect 2145 150 2175 176
rect 2223 172 2289 188
rect 2415 222 2481 238
rect 2415 188 2431 222
rect 2465 188 2481 222
rect 2241 150 2271 172
rect 2337 150 2367 176
rect 2415 172 2481 188
rect 2607 222 2673 238
rect 2607 188 2623 222
rect 2657 188 2673 222
rect 2433 150 2463 172
rect 2529 150 2559 176
rect 2607 172 2673 188
rect 2799 222 2865 238
rect 2799 188 2815 222
rect 2849 188 2865 222
rect 2625 150 2655 172
rect 2721 150 2751 176
rect 2799 172 2865 188
rect 2991 222 3057 238
rect 2991 188 3007 222
rect 3041 188 3057 222
rect 2817 150 2847 172
rect 2913 150 2943 176
rect 2991 172 3057 188
rect 3183 222 3249 238
rect 3183 188 3199 222
rect 3233 188 3249 222
rect 3009 150 3039 172
rect 3105 150 3135 176
rect 3183 172 3249 188
rect 3375 222 3441 238
rect 3375 188 3391 222
rect 3425 188 3441 222
rect 3201 150 3231 172
rect 3297 150 3327 176
rect 3375 172 3441 188
rect 3567 222 3633 238
rect 3567 188 3583 222
rect 3617 188 3633 222
rect 3393 150 3423 172
rect 3489 150 3519 176
rect 3567 172 3633 188
rect 3759 222 3825 238
rect 3759 188 3775 222
rect 3809 188 3825 222
rect 3585 150 3615 172
rect 3681 150 3711 176
rect 3759 172 3825 188
rect 3951 222 4017 238
rect 3951 188 3967 222
rect 4001 188 4017 222
rect 3777 150 3807 172
rect 3873 150 3903 176
rect 3951 172 4017 188
rect 4143 222 4209 238
rect 4143 188 4159 222
rect 4193 188 4209 222
rect 3969 150 3999 172
rect 4065 150 4095 176
rect 4143 172 4209 188
rect 4335 222 4401 238
rect 4335 188 4351 222
rect 4385 188 4401 222
rect 4161 150 4191 172
rect 4257 150 4287 176
rect 4335 172 4401 188
rect 4527 222 4593 238
rect 4527 188 4543 222
rect 4577 188 4593 222
rect 4353 150 4383 172
rect 4449 150 4479 176
rect 4527 172 4593 188
rect 4719 222 4785 238
rect 4719 188 4735 222
rect 4769 188 4785 222
rect 4545 150 4575 172
rect 4641 150 4671 176
rect 4719 172 4785 188
rect 4911 222 4977 238
rect 4911 188 4927 222
rect 4961 188 4977 222
rect 4737 150 4767 172
rect 4833 150 4863 176
rect 4911 172 4977 188
rect 5103 222 5169 238
rect 5103 188 5119 222
rect 5153 188 5169 222
rect 4929 150 4959 172
rect 5025 150 5055 176
rect 5103 172 5169 188
rect 5295 222 5361 238
rect 5295 188 5311 222
rect 5345 188 5361 222
rect 5121 150 5151 172
rect 5217 150 5247 176
rect 5295 172 5361 188
rect 5487 222 5553 238
rect 5487 188 5503 222
rect 5537 188 5553 222
rect 5313 150 5343 172
rect 5409 150 5439 176
rect 5487 172 5553 188
rect 5679 222 5745 238
rect 5679 188 5695 222
rect 5729 188 5745 222
rect 5505 150 5535 172
rect 5601 150 5631 176
rect 5679 172 5745 188
rect 5871 222 5937 238
rect 5871 188 5887 222
rect 5921 188 5937 222
rect 5697 150 5727 172
rect 5793 150 5823 176
rect 5871 172 5937 188
rect 6063 222 6129 238
rect 6063 188 6079 222
rect 6113 188 6129 222
rect 5889 150 5919 172
rect 5985 150 6015 176
rect 6063 172 6129 188
rect 6255 222 6321 238
rect 6255 188 6271 222
rect 6305 188 6321 222
rect 6081 150 6111 172
rect 6177 150 6207 176
rect 6255 172 6321 188
rect 6447 222 6513 238
rect 6447 188 6463 222
rect 6497 188 6513 222
rect 6273 150 6303 172
rect 6369 150 6399 176
rect 6447 172 6513 188
rect 6639 222 6705 238
rect 6639 188 6655 222
rect 6689 188 6705 222
rect 6465 150 6495 172
rect 6561 150 6591 176
rect 6639 172 6705 188
rect 6831 222 6897 238
rect 6831 188 6847 222
rect 6881 188 6897 222
rect 6657 150 6687 172
rect 6753 150 6783 176
rect 6831 172 6897 188
rect 7023 222 7089 238
rect 7023 188 7039 222
rect 7073 188 7089 222
rect 6849 150 6879 172
rect 6945 150 6975 176
rect 7023 172 7089 188
rect 7215 222 7281 238
rect 7215 188 7231 222
rect 7265 188 7281 222
rect 7041 150 7071 172
rect 7137 150 7167 176
rect 7215 172 7281 188
rect 7407 222 7473 238
rect 7407 188 7423 222
rect 7457 188 7473 222
rect 7233 150 7263 172
rect 7329 150 7359 176
rect 7407 172 7473 188
rect 7599 222 7665 238
rect 7599 188 7615 222
rect 7649 188 7665 222
rect 7425 150 7455 172
rect 7521 150 7551 176
rect 7599 172 7665 188
rect 7791 222 7857 238
rect 7791 188 7807 222
rect 7841 188 7857 222
rect 7617 150 7647 172
rect 7713 150 7743 176
rect 7791 172 7857 188
rect 7983 222 8049 238
rect 7983 188 7999 222
rect 8033 188 8049 222
rect 7809 150 7839 172
rect 7905 150 7935 176
rect 7983 172 8049 188
rect 8175 222 8241 238
rect 8175 188 8191 222
rect 8225 188 8241 222
rect 8001 150 8031 172
rect 8097 150 8127 176
rect 8175 172 8241 188
rect 8367 222 8433 238
rect 8367 188 8383 222
rect 8417 188 8433 222
rect 8193 150 8223 172
rect 8289 150 8319 176
rect 8367 172 8433 188
rect 8559 222 8625 238
rect 8559 188 8575 222
rect 8609 188 8625 222
rect 8385 150 8415 172
rect 8481 150 8511 176
rect 8559 172 8625 188
rect 8751 222 8817 238
rect 8751 188 8767 222
rect 8801 188 8817 222
rect 8577 150 8607 172
rect 8673 150 8703 176
rect 8751 172 8817 188
rect 8943 222 9009 238
rect 8943 188 8959 222
rect 8993 188 9009 222
rect 8769 150 8799 172
rect 8865 150 8895 176
rect 8943 172 9009 188
rect 9135 222 9201 238
rect 9135 188 9151 222
rect 9185 188 9201 222
rect 8961 150 8991 172
rect 9057 150 9087 176
rect 9135 172 9201 188
rect 9327 222 9393 238
rect 9327 188 9343 222
rect 9377 188 9393 222
rect 9153 150 9183 172
rect 9249 150 9279 176
rect 9327 172 9393 188
rect 9519 222 9585 238
rect 9519 188 9535 222
rect 9569 188 9585 222
rect 9345 150 9375 172
rect 9441 150 9471 176
rect 9519 172 9585 188
rect 9711 222 9777 238
rect 9711 188 9727 222
rect 9761 188 9777 222
rect 9537 150 9567 172
rect 9633 150 9663 176
rect 9711 172 9777 188
rect 9903 222 9969 238
rect 9903 188 9919 222
rect 9953 188 9969 222
rect 9729 150 9759 172
rect 9825 150 9855 176
rect 9903 172 9969 188
rect 10095 222 10161 238
rect 10095 188 10111 222
rect 10145 188 10161 222
rect 9921 150 9951 172
rect 10017 150 10047 176
rect 10095 172 10161 188
rect 10287 222 10353 238
rect 10287 188 10303 222
rect 10337 188 10353 222
rect 10113 150 10143 172
rect 10209 150 10239 176
rect 10287 172 10353 188
rect 10479 222 10545 238
rect 10479 188 10495 222
rect 10529 188 10545 222
rect 10305 150 10335 172
rect 10401 150 10431 176
rect 10479 172 10545 188
rect 10671 222 10737 238
rect 10671 188 10687 222
rect 10721 188 10737 222
rect 10497 150 10527 172
rect 10593 150 10623 176
rect 10671 172 10737 188
rect 10863 222 10929 238
rect 10863 188 10879 222
rect 10913 188 10929 222
rect 10689 150 10719 172
rect 10785 150 10815 176
rect 10863 172 10929 188
rect 11055 222 11121 238
rect 11055 188 11071 222
rect 11105 188 11121 222
rect 10881 150 10911 172
rect 10977 150 11007 176
rect 11055 172 11121 188
rect 11247 222 11313 238
rect 11247 188 11263 222
rect 11297 188 11313 222
rect 11073 150 11103 172
rect 11169 150 11199 176
rect 11247 172 11313 188
rect 11439 222 11505 238
rect 11439 188 11455 222
rect 11489 188 11505 222
rect 11265 150 11295 172
rect 11361 150 11391 176
rect 11439 172 11505 188
rect 11631 222 11697 238
rect 11631 188 11647 222
rect 11681 188 11697 222
rect 11457 150 11487 172
rect 11553 150 11583 176
rect 11631 172 11697 188
rect 11823 222 11889 238
rect 11823 188 11839 222
rect 11873 188 11889 222
rect 11649 150 11679 172
rect 11745 150 11775 176
rect 11823 172 11889 188
rect 12015 222 12081 238
rect 12015 188 12031 222
rect 12065 188 12081 222
rect 11841 150 11871 172
rect 11937 150 11967 176
rect 12015 172 12081 188
rect 12207 222 12273 238
rect 12207 188 12223 222
rect 12257 188 12273 222
rect 12033 150 12063 172
rect 12129 150 12159 176
rect 12207 172 12273 188
rect 12399 222 12465 238
rect 12399 188 12415 222
rect 12449 188 12465 222
rect 12225 150 12255 172
rect 12321 150 12351 176
rect 12399 172 12465 188
rect 12591 222 12657 238
rect 12591 188 12607 222
rect 12641 188 12657 222
rect 12417 150 12447 172
rect 12513 150 12543 176
rect 12591 172 12657 188
rect 12783 222 12849 238
rect 12783 188 12799 222
rect 12833 188 12849 222
rect 12609 150 12639 172
rect 12705 150 12735 176
rect 12783 172 12849 188
rect 12975 222 13041 238
rect 12975 188 12991 222
rect 13025 188 13041 222
rect 12801 150 12831 172
rect 12897 150 12927 176
rect 12975 172 13041 188
rect 13167 222 13233 238
rect 13167 188 13183 222
rect 13217 188 13233 222
rect 12993 150 13023 172
rect 13089 150 13119 176
rect 13167 172 13233 188
rect 13359 222 13425 238
rect 13359 188 13375 222
rect 13409 188 13425 222
rect 13185 150 13215 172
rect 13281 150 13311 176
rect 13359 172 13425 188
rect 13551 222 13617 238
rect 13551 188 13567 222
rect 13601 188 13617 222
rect 13377 150 13407 172
rect 13473 150 13503 176
rect 13551 172 13617 188
rect 13743 222 13809 238
rect 13743 188 13759 222
rect 13793 188 13809 222
rect 13569 150 13599 172
rect 13665 150 13695 176
rect 13743 172 13809 188
rect 13935 222 14001 238
rect 13935 188 13951 222
rect 13985 188 14001 222
rect 13761 150 13791 172
rect 13857 150 13887 176
rect 13935 172 14001 188
rect 14127 222 14193 238
rect 14127 188 14143 222
rect 14177 188 14193 222
rect 13953 150 13983 172
rect 14049 150 14079 176
rect 14127 172 14193 188
rect 14319 222 14385 238
rect 14319 188 14335 222
rect 14369 188 14385 222
rect 14145 150 14175 172
rect 14241 150 14271 176
rect 14319 172 14385 188
rect 14511 222 14577 238
rect 14511 188 14527 222
rect 14561 188 14577 222
rect 14337 150 14367 172
rect 14433 150 14463 176
rect 14511 172 14577 188
rect 14703 222 14769 238
rect 14703 188 14719 222
rect 14753 188 14769 222
rect 14529 150 14559 172
rect 14625 150 14655 176
rect 14703 172 14769 188
rect 14895 222 14961 238
rect 14895 188 14911 222
rect 14945 188 14961 222
rect 14721 150 14751 172
rect 14817 150 14847 176
rect 14895 172 14961 188
rect 15087 222 15153 238
rect 15087 188 15103 222
rect 15137 188 15153 222
rect 14913 150 14943 172
rect 15009 150 15039 176
rect 15087 172 15153 188
rect 15279 222 15345 238
rect 15279 188 15295 222
rect 15329 188 15345 222
rect 15105 150 15135 172
rect 15201 150 15231 176
rect 15279 172 15345 188
rect 15471 222 15537 238
rect 15471 188 15487 222
rect 15521 188 15537 222
rect 15297 150 15327 172
rect 15393 150 15423 176
rect 15471 172 15537 188
rect 15663 222 15729 238
rect 15663 188 15679 222
rect 15713 188 15729 222
rect 15489 150 15519 172
rect 15585 150 15615 176
rect 15663 172 15729 188
rect 15855 222 15921 238
rect 15855 188 15871 222
rect 15905 188 15921 222
rect 15681 150 15711 172
rect 15777 150 15807 176
rect 15855 172 15921 188
rect 16047 222 16113 238
rect 16047 188 16063 222
rect 16097 188 16113 222
rect 15873 150 15903 172
rect 15969 150 15999 176
rect 16047 172 16113 188
rect 16239 222 16305 238
rect 16239 188 16255 222
rect 16289 188 16305 222
rect 16065 150 16095 172
rect 16161 150 16191 176
rect 16239 172 16305 188
rect 16431 222 16497 238
rect 16431 188 16447 222
rect 16481 188 16497 222
rect 16257 150 16287 172
rect 16353 150 16383 176
rect 16431 172 16497 188
rect 16623 222 16689 238
rect 16623 188 16639 222
rect 16673 188 16689 222
rect 16449 150 16479 172
rect 16545 150 16575 176
rect 16623 172 16689 188
rect 16815 222 16881 238
rect 16815 188 16831 222
rect 16865 188 16881 222
rect 16641 150 16671 172
rect 16737 150 16767 176
rect 16815 172 16881 188
rect 17007 222 17073 238
rect 17007 188 17023 222
rect 17057 188 17073 222
rect 16833 150 16863 172
rect 16929 150 16959 176
rect 17007 172 17073 188
rect 17199 222 17265 238
rect 17199 188 17215 222
rect 17249 188 17265 222
rect 17025 150 17055 172
rect 17121 150 17151 176
rect 17199 172 17265 188
rect 17391 222 17457 238
rect 17391 188 17407 222
rect 17441 188 17457 222
rect 17217 150 17247 172
rect 17313 150 17343 176
rect 17391 172 17457 188
rect 17583 222 17649 238
rect 17583 188 17599 222
rect 17633 188 17649 222
rect 17409 150 17439 172
rect 17505 150 17535 176
rect 17583 172 17649 188
rect 17775 222 17841 238
rect 17775 188 17791 222
rect 17825 188 17841 222
rect 17601 150 17631 172
rect 17697 150 17727 176
rect 17775 172 17841 188
rect 17967 222 18033 238
rect 17967 188 17983 222
rect 18017 188 18033 222
rect 17793 150 17823 172
rect 17889 150 17919 176
rect 17967 172 18033 188
rect 18159 222 18225 238
rect 18159 188 18175 222
rect 18209 188 18225 222
rect 17985 150 18015 172
rect 18081 150 18111 176
rect 18159 172 18225 188
rect 18351 222 18417 238
rect 18351 188 18367 222
rect 18401 188 18417 222
rect 18177 150 18207 172
rect 18273 150 18303 176
rect 18351 172 18417 188
rect 18543 222 18609 238
rect 18543 188 18559 222
rect 18593 188 18609 222
rect 18369 150 18399 172
rect 18465 150 18495 176
rect 18543 172 18609 188
rect 18735 222 18801 238
rect 18735 188 18751 222
rect 18785 188 18801 222
rect 18561 150 18591 172
rect 18657 150 18687 176
rect 18735 172 18801 188
rect 18927 222 18993 238
rect 18927 188 18943 222
rect 18977 188 18993 222
rect 18753 150 18783 172
rect 18849 150 18879 176
rect 18927 172 18993 188
rect 19119 222 19185 238
rect 19119 188 19135 222
rect 19169 188 19185 222
rect 18945 150 18975 172
rect 19041 150 19071 176
rect 19119 172 19185 188
rect 19137 150 19167 172
rect -19167 -172 -19137 -150
rect -19185 -188 -19119 -172
rect -19071 -176 -19041 -150
rect -18975 -172 -18945 -150
rect -19185 -222 -19169 -188
rect -19135 -222 -19119 -188
rect -19185 -238 -19119 -222
rect -18993 -188 -18927 -172
rect -18879 -176 -18849 -150
rect -18783 -172 -18753 -150
rect -18993 -222 -18977 -188
rect -18943 -222 -18927 -188
rect -18993 -238 -18927 -222
rect -18801 -188 -18735 -172
rect -18687 -176 -18657 -150
rect -18591 -172 -18561 -150
rect -18801 -222 -18785 -188
rect -18751 -222 -18735 -188
rect -18801 -238 -18735 -222
rect -18609 -188 -18543 -172
rect -18495 -176 -18465 -150
rect -18399 -172 -18369 -150
rect -18609 -222 -18593 -188
rect -18559 -222 -18543 -188
rect -18609 -238 -18543 -222
rect -18417 -188 -18351 -172
rect -18303 -176 -18273 -150
rect -18207 -172 -18177 -150
rect -18417 -222 -18401 -188
rect -18367 -222 -18351 -188
rect -18417 -238 -18351 -222
rect -18225 -188 -18159 -172
rect -18111 -176 -18081 -150
rect -18015 -172 -17985 -150
rect -18225 -222 -18209 -188
rect -18175 -222 -18159 -188
rect -18225 -238 -18159 -222
rect -18033 -188 -17967 -172
rect -17919 -176 -17889 -150
rect -17823 -172 -17793 -150
rect -18033 -222 -18017 -188
rect -17983 -222 -17967 -188
rect -18033 -238 -17967 -222
rect -17841 -188 -17775 -172
rect -17727 -176 -17697 -150
rect -17631 -172 -17601 -150
rect -17841 -222 -17825 -188
rect -17791 -222 -17775 -188
rect -17841 -238 -17775 -222
rect -17649 -188 -17583 -172
rect -17535 -176 -17505 -150
rect -17439 -172 -17409 -150
rect -17649 -222 -17633 -188
rect -17599 -222 -17583 -188
rect -17649 -238 -17583 -222
rect -17457 -188 -17391 -172
rect -17343 -176 -17313 -150
rect -17247 -172 -17217 -150
rect -17457 -222 -17441 -188
rect -17407 -222 -17391 -188
rect -17457 -238 -17391 -222
rect -17265 -188 -17199 -172
rect -17151 -176 -17121 -150
rect -17055 -172 -17025 -150
rect -17265 -222 -17249 -188
rect -17215 -222 -17199 -188
rect -17265 -238 -17199 -222
rect -17073 -188 -17007 -172
rect -16959 -176 -16929 -150
rect -16863 -172 -16833 -150
rect -17073 -222 -17057 -188
rect -17023 -222 -17007 -188
rect -17073 -238 -17007 -222
rect -16881 -188 -16815 -172
rect -16767 -176 -16737 -150
rect -16671 -172 -16641 -150
rect -16881 -222 -16865 -188
rect -16831 -222 -16815 -188
rect -16881 -238 -16815 -222
rect -16689 -188 -16623 -172
rect -16575 -176 -16545 -150
rect -16479 -172 -16449 -150
rect -16689 -222 -16673 -188
rect -16639 -222 -16623 -188
rect -16689 -238 -16623 -222
rect -16497 -188 -16431 -172
rect -16383 -176 -16353 -150
rect -16287 -172 -16257 -150
rect -16497 -222 -16481 -188
rect -16447 -222 -16431 -188
rect -16497 -238 -16431 -222
rect -16305 -188 -16239 -172
rect -16191 -176 -16161 -150
rect -16095 -172 -16065 -150
rect -16305 -222 -16289 -188
rect -16255 -222 -16239 -188
rect -16305 -238 -16239 -222
rect -16113 -188 -16047 -172
rect -15999 -176 -15969 -150
rect -15903 -172 -15873 -150
rect -16113 -222 -16097 -188
rect -16063 -222 -16047 -188
rect -16113 -238 -16047 -222
rect -15921 -188 -15855 -172
rect -15807 -176 -15777 -150
rect -15711 -172 -15681 -150
rect -15921 -222 -15905 -188
rect -15871 -222 -15855 -188
rect -15921 -238 -15855 -222
rect -15729 -188 -15663 -172
rect -15615 -176 -15585 -150
rect -15519 -172 -15489 -150
rect -15729 -222 -15713 -188
rect -15679 -222 -15663 -188
rect -15729 -238 -15663 -222
rect -15537 -188 -15471 -172
rect -15423 -176 -15393 -150
rect -15327 -172 -15297 -150
rect -15537 -222 -15521 -188
rect -15487 -222 -15471 -188
rect -15537 -238 -15471 -222
rect -15345 -188 -15279 -172
rect -15231 -176 -15201 -150
rect -15135 -172 -15105 -150
rect -15345 -222 -15329 -188
rect -15295 -222 -15279 -188
rect -15345 -238 -15279 -222
rect -15153 -188 -15087 -172
rect -15039 -176 -15009 -150
rect -14943 -172 -14913 -150
rect -15153 -222 -15137 -188
rect -15103 -222 -15087 -188
rect -15153 -238 -15087 -222
rect -14961 -188 -14895 -172
rect -14847 -176 -14817 -150
rect -14751 -172 -14721 -150
rect -14961 -222 -14945 -188
rect -14911 -222 -14895 -188
rect -14961 -238 -14895 -222
rect -14769 -188 -14703 -172
rect -14655 -176 -14625 -150
rect -14559 -172 -14529 -150
rect -14769 -222 -14753 -188
rect -14719 -222 -14703 -188
rect -14769 -238 -14703 -222
rect -14577 -188 -14511 -172
rect -14463 -176 -14433 -150
rect -14367 -172 -14337 -150
rect -14577 -222 -14561 -188
rect -14527 -222 -14511 -188
rect -14577 -238 -14511 -222
rect -14385 -188 -14319 -172
rect -14271 -176 -14241 -150
rect -14175 -172 -14145 -150
rect -14385 -222 -14369 -188
rect -14335 -222 -14319 -188
rect -14385 -238 -14319 -222
rect -14193 -188 -14127 -172
rect -14079 -176 -14049 -150
rect -13983 -172 -13953 -150
rect -14193 -222 -14177 -188
rect -14143 -222 -14127 -188
rect -14193 -238 -14127 -222
rect -14001 -188 -13935 -172
rect -13887 -176 -13857 -150
rect -13791 -172 -13761 -150
rect -14001 -222 -13985 -188
rect -13951 -222 -13935 -188
rect -14001 -238 -13935 -222
rect -13809 -188 -13743 -172
rect -13695 -176 -13665 -150
rect -13599 -172 -13569 -150
rect -13809 -222 -13793 -188
rect -13759 -222 -13743 -188
rect -13809 -238 -13743 -222
rect -13617 -188 -13551 -172
rect -13503 -176 -13473 -150
rect -13407 -172 -13377 -150
rect -13617 -222 -13601 -188
rect -13567 -222 -13551 -188
rect -13617 -238 -13551 -222
rect -13425 -188 -13359 -172
rect -13311 -176 -13281 -150
rect -13215 -172 -13185 -150
rect -13425 -222 -13409 -188
rect -13375 -222 -13359 -188
rect -13425 -238 -13359 -222
rect -13233 -188 -13167 -172
rect -13119 -176 -13089 -150
rect -13023 -172 -12993 -150
rect -13233 -222 -13217 -188
rect -13183 -222 -13167 -188
rect -13233 -238 -13167 -222
rect -13041 -188 -12975 -172
rect -12927 -176 -12897 -150
rect -12831 -172 -12801 -150
rect -13041 -222 -13025 -188
rect -12991 -222 -12975 -188
rect -13041 -238 -12975 -222
rect -12849 -188 -12783 -172
rect -12735 -176 -12705 -150
rect -12639 -172 -12609 -150
rect -12849 -222 -12833 -188
rect -12799 -222 -12783 -188
rect -12849 -238 -12783 -222
rect -12657 -188 -12591 -172
rect -12543 -176 -12513 -150
rect -12447 -172 -12417 -150
rect -12657 -222 -12641 -188
rect -12607 -222 -12591 -188
rect -12657 -238 -12591 -222
rect -12465 -188 -12399 -172
rect -12351 -176 -12321 -150
rect -12255 -172 -12225 -150
rect -12465 -222 -12449 -188
rect -12415 -222 -12399 -188
rect -12465 -238 -12399 -222
rect -12273 -188 -12207 -172
rect -12159 -176 -12129 -150
rect -12063 -172 -12033 -150
rect -12273 -222 -12257 -188
rect -12223 -222 -12207 -188
rect -12273 -238 -12207 -222
rect -12081 -188 -12015 -172
rect -11967 -176 -11937 -150
rect -11871 -172 -11841 -150
rect -12081 -222 -12065 -188
rect -12031 -222 -12015 -188
rect -12081 -238 -12015 -222
rect -11889 -188 -11823 -172
rect -11775 -176 -11745 -150
rect -11679 -172 -11649 -150
rect -11889 -222 -11873 -188
rect -11839 -222 -11823 -188
rect -11889 -238 -11823 -222
rect -11697 -188 -11631 -172
rect -11583 -176 -11553 -150
rect -11487 -172 -11457 -150
rect -11697 -222 -11681 -188
rect -11647 -222 -11631 -188
rect -11697 -238 -11631 -222
rect -11505 -188 -11439 -172
rect -11391 -176 -11361 -150
rect -11295 -172 -11265 -150
rect -11505 -222 -11489 -188
rect -11455 -222 -11439 -188
rect -11505 -238 -11439 -222
rect -11313 -188 -11247 -172
rect -11199 -176 -11169 -150
rect -11103 -172 -11073 -150
rect -11313 -222 -11297 -188
rect -11263 -222 -11247 -188
rect -11313 -238 -11247 -222
rect -11121 -188 -11055 -172
rect -11007 -176 -10977 -150
rect -10911 -172 -10881 -150
rect -11121 -222 -11105 -188
rect -11071 -222 -11055 -188
rect -11121 -238 -11055 -222
rect -10929 -188 -10863 -172
rect -10815 -176 -10785 -150
rect -10719 -172 -10689 -150
rect -10929 -222 -10913 -188
rect -10879 -222 -10863 -188
rect -10929 -238 -10863 -222
rect -10737 -188 -10671 -172
rect -10623 -176 -10593 -150
rect -10527 -172 -10497 -150
rect -10737 -222 -10721 -188
rect -10687 -222 -10671 -188
rect -10737 -238 -10671 -222
rect -10545 -188 -10479 -172
rect -10431 -176 -10401 -150
rect -10335 -172 -10305 -150
rect -10545 -222 -10529 -188
rect -10495 -222 -10479 -188
rect -10545 -238 -10479 -222
rect -10353 -188 -10287 -172
rect -10239 -176 -10209 -150
rect -10143 -172 -10113 -150
rect -10353 -222 -10337 -188
rect -10303 -222 -10287 -188
rect -10353 -238 -10287 -222
rect -10161 -188 -10095 -172
rect -10047 -176 -10017 -150
rect -9951 -172 -9921 -150
rect -10161 -222 -10145 -188
rect -10111 -222 -10095 -188
rect -10161 -238 -10095 -222
rect -9969 -188 -9903 -172
rect -9855 -176 -9825 -150
rect -9759 -172 -9729 -150
rect -9969 -222 -9953 -188
rect -9919 -222 -9903 -188
rect -9969 -238 -9903 -222
rect -9777 -188 -9711 -172
rect -9663 -176 -9633 -150
rect -9567 -172 -9537 -150
rect -9777 -222 -9761 -188
rect -9727 -222 -9711 -188
rect -9777 -238 -9711 -222
rect -9585 -188 -9519 -172
rect -9471 -176 -9441 -150
rect -9375 -172 -9345 -150
rect -9585 -222 -9569 -188
rect -9535 -222 -9519 -188
rect -9585 -238 -9519 -222
rect -9393 -188 -9327 -172
rect -9279 -176 -9249 -150
rect -9183 -172 -9153 -150
rect -9393 -222 -9377 -188
rect -9343 -222 -9327 -188
rect -9393 -238 -9327 -222
rect -9201 -188 -9135 -172
rect -9087 -176 -9057 -150
rect -8991 -172 -8961 -150
rect -9201 -222 -9185 -188
rect -9151 -222 -9135 -188
rect -9201 -238 -9135 -222
rect -9009 -188 -8943 -172
rect -8895 -176 -8865 -150
rect -8799 -172 -8769 -150
rect -9009 -222 -8993 -188
rect -8959 -222 -8943 -188
rect -9009 -238 -8943 -222
rect -8817 -188 -8751 -172
rect -8703 -176 -8673 -150
rect -8607 -172 -8577 -150
rect -8817 -222 -8801 -188
rect -8767 -222 -8751 -188
rect -8817 -238 -8751 -222
rect -8625 -188 -8559 -172
rect -8511 -176 -8481 -150
rect -8415 -172 -8385 -150
rect -8625 -222 -8609 -188
rect -8575 -222 -8559 -188
rect -8625 -238 -8559 -222
rect -8433 -188 -8367 -172
rect -8319 -176 -8289 -150
rect -8223 -172 -8193 -150
rect -8433 -222 -8417 -188
rect -8383 -222 -8367 -188
rect -8433 -238 -8367 -222
rect -8241 -188 -8175 -172
rect -8127 -176 -8097 -150
rect -8031 -172 -8001 -150
rect -8241 -222 -8225 -188
rect -8191 -222 -8175 -188
rect -8241 -238 -8175 -222
rect -8049 -188 -7983 -172
rect -7935 -176 -7905 -150
rect -7839 -172 -7809 -150
rect -8049 -222 -8033 -188
rect -7999 -222 -7983 -188
rect -8049 -238 -7983 -222
rect -7857 -188 -7791 -172
rect -7743 -176 -7713 -150
rect -7647 -172 -7617 -150
rect -7857 -222 -7841 -188
rect -7807 -222 -7791 -188
rect -7857 -238 -7791 -222
rect -7665 -188 -7599 -172
rect -7551 -176 -7521 -150
rect -7455 -172 -7425 -150
rect -7665 -222 -7649 -188
rect -7615 -222 -7599 -188
rect -7665 -238 -7599 -222
rect -7473 -188 -7407 -172
rect -7359 -176 -7329 -150
rect -7263 -172 -7233 -150
rect -7473 -222 -7457 -188
rect -7423 -222 -7407 -188
rect -7473 -238 -7407 -222
rect -7281 -188 -7215 -172
rect -7167 -176 -7137 -150
rect -7071 -172 -7041 -150
rect -7281 -222 -7265 -188
rect -7231 -222 -7215 -188
rect -7281 -238 -7215 -222
rect -7089 -188 -7023 -172
rect -6975 -176 -6945 -150
rect -6879 -172 -6849 -150
rect -7089 -222 -7073 -188
rect -7039 -222 -7023 -188
rect -7089 -238 -7023 -222
rect -6897 -188 -6831 -172
rect -6783 -176 -6753 -150
rect -6687 -172 -6657 -150
rect -6897 -222 -6881 -188
rect -6847 -222 -6831 -188
rect -6897 -238 -6831 -222
rect -6705 -188 -6639 -172
rect -6591 -176 -6561 -150
rect -6495 -172 -6465 -150
rect -6705 -222 -6689 -188
rect -6655 -222 -6639 -188
rect -6705 -238 -6639 -222
rect -6513 -188 -6447 -172
rect -6399 -176 -6369 -150
rect -6303 -172 -6273 -150
rect -6513 -222 -6497 -188
rect -6463 -222 -6447 -188
rect -6513 -238 -6447 -222
rect -6321 -188 -6255 -172
rect -6207 -176 -6177 -150
rect -6111 -172 -6081 -150
rect -6321 -222 -6305 -188
rect -6271 -222 -6255 -188
rect -6321 -238 -6255 -222
rect -6129 -188 -6063 -172
rect -6015 -176 -5985 -150
rect -5919 -172 -5889 -150
rect -6129 -222 -6113 -188
rect -6079 -222 -6063 -188
rect -6129 -238 -6063 -222
rect -5937 -188 -5871 -172
rect -5823 -176 -5793 -150
rect -5727 -172 -5697 -150
rect -5937 -222 -5921 -188
rect -5887 -222 -5871 -188
rect -5937 -238 -5871 -222
rect -5745 -188 -5679 -172
rect -5631 -176 -5601 -150
rect -5535 -172 -5505 -150
rect -5745 -222 -5729 -188
rect -5695 -222 -5679 -188
rect -5745 -238 -5679 -222
rect -5553 -188 -5487 -172
rect -5439 -176 -5409 -150
rect -5343 -172 -5313 -150
rect -5553 -222 -5537 -188
rect -5503 -222 -5487 -188
rect -5553 -238 -5487 -222
rect -5361 -188 -5295 -172
rect -5247 -176 -5217 -150
rect -5151 -172 -5121 -150
rect -5361 -222 -5345 -188
rect -5311 -222 -5295 -188
rect -5361 -238 -5295 -222
rect -5169 -188 -5103 -172
rect -5055 -176 -5025 -150
rect -4959 -172 -4929 -150
rect -5169 -222 -5153 -188
rect -5119 -222 -5103 -188
rect -5169 -238 -5103 -222
rect -4977 -188 -4911 -172
rect -4863 -176 -4833 -150
rect -4767 -172 -4737 -150
rect -4977 -222 -4961 -188
rect -4927 -222 -4911 -188
rect -4977 -238 -4911 -222
rect -4785 -188 -4719 -172
rect -4671 -176 -4641 -150
rect -4575 -172 -4545 -150
rect -4785 -222 -4769 -188
rect -4735 -222 -4719 -188
rect -4785 -238 -4719 -222
rect -4593 -188 -4527 -172
rect -4479 -176 -4449 -150
rect -4383 -172 -4353 -150
rect -4593 -222 -4577 -188
rect -4543 -222 -4527 -188
rect -4593 -238 -4527 -222
rect -4401 -188 -4335 -172
rect -4287 -176 -4257 -150
rect -4191 -172 -4161 -150
rect -4401 -222 -4385 -188
rect -4351 -222 -4335 -188
rect -4401 -238 -4335 -222
rect -4209 -188 -4143 -172
rect -4095 -176 -4065 -150
rect -3999 -172 -3969 -150
rect -4209 -222 -4193 -188
rect -4159 -222 -4143 -188
rect -4209 -238 -4143 -222
rect -4017 -188 -3951 -172
rect -3903 -176 -3873 -150
rect -3807 -172 -3777 -150
rect -4017 -222 -4001 -188
rect -3967 -222 -3951 -188
rect -4017 -238 -3951 -222
rect -3825 -188 -3759 -172
rect -3711 -176 -3681 -150
rect -3615 -172 -3585 -150
rect -3825 -222 -3809 -188
rect -3775 -222 -3759 -188
rect -3825 -238 -3759 -222
rect -3633 -188 -3567 -172
rect -3519 -176 -3489 -150
rect -3423 -172 -3393 -150
rect -3633 -222 -3617 -188
rect -3583 -222 -3567 -188
rect -3633 -238 -3567 -222
rect -3441 -188 -3375 -172
rect -3327 -176 -3297 -150
rect -3231 -172 -3201 -150
rect -3441 -222 -3425 -188
rect -3391 -222 -3375 -188
rect -3441 -238 -3375 -222
rect -3249 -188 -3183 -172
rect -3135 -176 -3105 -150
rect -3039 -172 -3009 -150
rect -3249 -222 -3233 -188
rect -3199 -222 -3183 -188
rect -3249 -238 -3183 -222
rect -3057 -188 -2991 -172
rect -2943 -176 -2913 -150
rect -2847 -172 -2817 -150
rect -3057 -222 -3041 -188
rect -3007 -222 -2991 -188
rect -3057 -238 -2991 -222
rect -2865 -188 -2799 -172
rect -2751 -176 -2721 -150
rect -2655 -172 -2625 -150
rect -2865 -222 -2849 -188
rect -2815 -222 -2799 -188
rect -2865 -238 -2799 -222
rect -2673 -188 -2607 -172
rect -2559 -176 -2529 -150
rect -2463 -172 -2433 -150
rect -2673 -222 -2657 -188
rect -2623 -222 -2607 -188
rect -2673 -238 -2607 -222
rect -2481 -188 -2415 -172
rect -2367 -176 -2337 -150
rect -2271 -172 -2241 -150
rect -2481 -222 -2465 -188
rect -2431 -222 -2415 -188
rect -2481 -238 -2415 -222
rect -2289 -188 -2223 -172
rect -2175 -176 -2145 -150
rect -2079 -172 -2049 -150
rect -2289 -222 -2273 -188
rect -2239 -222 -2223 -188
rect -2289 -238 -2223 -222
rect -2097 -188 -2031 -172
rect -1983 -176 -1953 -150
rect -1887 -172 -1857 -150
rect -2097 -222 -2081 -188
rect -2047 -222 -2031 -188
rect -2097 -238 -2031 -222
rect -1905 -188 -1839 -172
rect -1791 -176 -1761 -150
rect -1695 -172 -1665 -150
rect -1905 -222 -1889 -188
rect -1855 -222 -1839 -188
rect -1905 -238 -1839 -222
rect -1713 -188 -1647 -172
rect -1599 -176 -1569 -150
rect -1503 -172 -1473 -150
rect -1713 -222 -1697 -188
rect -1663 -222 -1647 -188
rect -1713 -238 -1647 -222
rect -1521 -188 -1455 -172
rect -1407 -176 -1377 -150
rect -1311 -172 -1281 -150
rect -1521 -222 -1505 -188
rect -1471 -222 -1455 -188
rect -1521 -238 -1455 -222
rect -1329 -188 -1263 -172
rect -1215 -176 -1185 -150
rect -1119 -172 -1089 -150
rect -1329 -222 -1313 -188
rect -1279 -222 -1263 -188
rect -1329 -238 -1263 -222
rect -1137 -188 -1071 -172
rect -1023 -176 -993 -150
rect -927 -172 -897 -150
rect -1137 -222 -1121 -188
rect -1087 -222 -1071 -188
rect -1137 -238 -1071 -222
rect -945 -188 -879 -172
rect -831 -176 -801 -150
rect -735 -172 -705 -150
rect -945 -222 -929 -188
rect -895 -222 -879 -188
rect -945 -238 -879 -222
rect -753 -188 -687 -172
rect -639 -176 -609 -150
rect -543 -172 -513 -150
rect -753 -222 -737 -188
rect -703 -222 -687 -188
rect -753 -238 -687 -222
rect -561 -188 -495 -172
rect -447 -176 -417 -150
rect -351 -172 -321 -150
rect -561 -222 -545 -188
rect -511 -222 -495 -188
rect -561 -238 -495 -222
rect -369 -188 -303 -172
rect -255 -176 -225 -150
rect -159 -172 -129 -150
rect -369 -222 -353 -188
rect -319 -222 -303 -188
rect -369 -238 -303 -222
rect -177 -188 -111 -172
rect -63 -176 -33 -150
rect 33 -172 63 -150
rect -177 -222 -161 -188
rect -127 -222 -111 -188
rect -177 -238 -111 -222
rect 15 -188 81 -172
rect 129 -176 159 -150
rect 225 -172 255 -150
rect 15 -222 31 -188
rect 65 -222 81 -188
rect 15 -238 81 -222
rect 207 -188 273 -172
rect 321 -176 351 -150
rect 417 -172 447 -150
rect 207 -222 223 -188
rect 257 -222 273 -188
rect 207 -238 273 -222
rect 399 -188 465 -172
rect 513 -176 543 -150
rect 609 -172 639 -150
rect 399 -222 415 -188
rect 449 -222 465 -188
rect 399 -238 465 -222
rect 591 -188 657 -172
rect 705 -176 735 -150
rect 801 -172 831 -150
rect 591 -222 607 -188
rect 641 -222 657 -188
rect 591 -238 657 -222
rect 783 -188 849 -172
rect 897 -176 927 -150
rect 993 -172 1023 -150
rect 783 -222 799 -188
rect 833 -222 849 -188
rect 783 -238 849 -222
rect 975 -188 1041 -172
rect 1089 -176 1119 -150
rect 1185 -172 1215 -150
rect 975 -222 991 -188
rect 1025 -222 1041 -188
rect 975 -238 1041 -222
rect 1167 -188 1233 -172
rect 1281 -176 1311 -150
rect 1377 -172 1407 -150
rect 1167 -222 1183 -188
rect 1217 -222 1233 -188
rect 1167 -238 1233 -222
rect 1359 -188 1425 -172
rect 1473 -176 1503 -150
rect 1569 -172 1599 -150
rect 1359 -222 1375 -188
rect 1409 -222 1425 -188
rect 1359 -238 1425 -222
rect 1551 -188 1617 -172
rect 1665 -176 1695 -150
rect 1761 -172 1791 -150
rect 1551 -222 1567 -188
rect 1601 -222 1617 -188
rect 1551 -238 1617 -222
rect 1743 -188 1809 -172
rect 1857 -176 1887 -150
rect 1953 -172 1983 -150
rect 1743 -222 1759 -188
rect 1793 -222 1809 -188
rect 1743 -238 1809 -222
rect 1935 -188 2001 -172
rect 2049 -176 2079 -150
rect 2145 -172 2175 -150
rect 1935 -222 1951 -188
rect 1985 -222 2001 -188
rect 1935 -238 2001 -222
rect 2127 -188 2193 -172
rect 2241 -176 2271 -150
rect 2337 -172 2367 -150
rect 2127 -222 2143 -188
rect 2177 -222 2193 -188
rect 2127 -238 2193 -222
rect 2319 -188 2385 -172
rect 2433 -176 2463 -150
rect 2529 -172 2559 -150
rect 2319 -222 2335 -188
rect 2369 -222 2385 -188
rect 2319 -238 2385 -222
rect 2511 -188 2577 -172
rect 2625 -176 2655 -150
rect 2721 -172 2751 -150
rect 2511 -222 2527 -188
rect 2561 -222 2577 -188
rect 2511 -238 2577 -222
rect 2703 -188 2769 -172
rect 2817 -176 2847 -150
rect 2913 -172 2943 -150
rect 2703 -222 2719 -188
rect 2753 -222 2769 -188
rect 2703 -238 2769 -222
rect 2895 -188 2961 -172
rect 3009 -176 3039 -150
rect 3105 -172 3135 -150
rect 2895 -222 2911 -188
rect 2945 -222 2961 -188
rect 2895 -238 2961 -222
rect 3087 -188 3153 -172
rect 3201 -176 3231 -150
rect 3297 -172 3327 -150
rect 3087 -222 3103 -188
rect 3137 -222 3153 -188
rect 3087 -238 3153 -222
rect 3279 -188 3345 -172
rect 3393 -176 3423 -150
rect 3489 -172 3519 -150
rect 3279 -222 3295 -188
rect 3329 -222 3345 -188
rect 3279 -238 3345 -222
rect 3471 -188 3537 -172
rect 3585 -176 3615 -150
rect 3681 -172 3711 -150
rect 3471 -222 3487 -188
rect 3521 -222 3537 -188
rect 3471 -238 3537 -222
rect 3663 -188 3729 -172
rect 3777 -176 3807 -150
rect 3873 -172 3903 -150
rect 3663 -222 3679 -188
rect 3713 -222 3729 -188
rect 3663 -238 3729 -222
rect 3855 -188 3921 -172
rect 3969 -176 3999 -150
rect 4065 -172 4095 -150
rect 3855 -222 3871 -188
rect 3905 -222 3921 -188
rect 3855 -238 3921 -222
rect 4047 -188 4113 -172
rect 4161 -176 4191 -150
rect 4257 -172 4287 -150
rect 4047 -222 4063 -188
rect 4097 -222 4113 -188
rect 4047 -238 4113 -222
rect 4239 -188 4305 -172
rect 4353 -176 4383 -150
rect 4449 -172 4479 -150
rect 4239 -222 4255 -188
rect 4289 -222 4305 -188
rect 4239 -238 4305 -222
rect 4431 -188 4497 -172
rect 4545 -176 4575 -150
rect 4641 -172 4671 -150
rect 4431 -222 4447 -188
rect 4481 -222 4497 -188
rect 4431 -238 4497 -222
rect 4623 -188 4689 -172
rect 4737 -176 4767 -150
rect 4833 -172 4863 -150
rect 4623 -222 4639 -188
rect 4673 -222 4689 -188
rect 4623 -238 4689 -222
rect 4815 -188 4881 -172
rect 4929 -176 4959 -150
rect 5025 -172 5055 -150
rect 4815 -222 4831 -188
rect 4865 -222 4881 -188
rect 4815 -238 4881 -222
rect 5007 -188 5073 -172
rect 5121 -176 5151 -150
rect 5217 -172 5247 -150
rect 5007 -222 5023 -188
rect 5057 -222 5073 -188
rect 5007 -238 5073 -222
rect 5199 -188 5265 -172
rect 5313 -176 5343 -150
rect 5409 -172 5439 -150
rect 5199 -222 5215 -188
rect 5249 -222 5265 -188
rect 5199 -238 5265 -222
rect 5391 -188 5457 -172
rect 5505 -176 5535 -150
rect 5601 -172 5631 -150
rect 5391 -222 5407 -188
rect 5441 -222 5457 -188
rect 5391 -238 5457 -222
rect 5583 -188 5649 -172
rect 5697 -176 5727 -150
rect 5793 -172 5823 -150
rect 5583 -222 5599 -188
rect 5633 -222 5649 -188
rect 5583 -238 5649 -222
rect 5775 -188 5841 -172
rect 5889 -176 5919 -150
rect 5985 -172 6015 -150
rect 5775 -222 5791 -188
rect 5825 -222 5841 -188
rect 5775 -238 5841 -222
rect 5967 -188 6033 -172
rect 6081 -176 6111 -150
rect 6177 -172 6207 -150
rect 5967 -222 5983 -188
rect 6017 -222 6033 -188
rect 5967 -238 6033 -222
rect 6159 -188 6225 -172
rect 6273 -176 6303 -150
rect 6369 -172 6399 -150
rect 6159 -222 6175 -188
rect 6209 -222 6225 -188
rect 6159 -238 6225 -222
rect 6351 -188 6417 -172
rect 6465 -176 6495 -150
rect 6561 -172 6591 -150
rect 6351 -222 6367 -188
rect 6401 -222 6417 -188
rect 6351 -238 6417 -222
rect 6543 -188 6609 -172
rect 6657 -176 6687 -150
rect 6753 -172 6783 -150
rect 6543 -222 6559 -188
rect 6593 -222 6609 -188
rect 6543 -238 6609 -222
rect 6735 -188 6801 -172
rect 6849 -176 6879 -150
rect 6945 -172 6975 -150
rect 6735 -222 6751 -188
rect 6785 -222 6801 -188
rect 6735 -238 6801 -222
rect 6927 -188 6993 -172
rect 7041 -176 7071 -150
rect 7137 -172 7167 -150
rect 6927 -222 6943 -188
rect 6977 -222 6993 -188
rect 6927 -238 6993 -222
rect 7119 -188 7185 -172
rect 7233 -176 7263 -150
rect 7329 -172 7359 -150
rect 7119 -222 7135 -188
rect 7169 -222 7185 -188
rect 7119 -238 7185 -222
rect 7311 -188 7377 -172
rect 7425 -176 7455 -150
rect 7521 -172 7551 -150
rect 7311 -222 7327 -188
rect 7361 -222 7377 -188
rect 7311 -238 7377 -222
rect 7503 -188 7569 -172
rect 7617 -176 7647 -150
rect 7713 -172 7743 -150
rect 7503 -222 7519 -188
rect 7553 -222 7569 -188
rect 7503 -238 7569 -222
rect 7695 -188 7761 -172
rect 7809 -176 7839 -150
rect 7905 -172 7935 -150
rect 7695 -222 7711 -188
rect 7745 -222 7761 -188
rect 7695 -238 7761 -222
rect 7887 -188 7953 -172
rect 8001 -176 8031 -150
rect 8097 -172 8127 -150
rect 7887 -222 7903 -188
rect 7937 -222 7953 -188
rect 7887 -238 7953 -222
rect 8079 -188 8145 -172
rect 8193 -176 8223 -150
rect 8289 -172 8319 -150
rect 8079 -222 8095 -188
rect 8129 -222 8145 -188
rect 8079 -238 8145 -222
rect 8271 -188 8337 -172
rect 8385 -176 8415 -150
rect 8481 -172 8511 -150
rect 8271 -222 8287 -188
rect 8321 -222 8337 -188
rect 8271 -238 8337 -222
rect 8463 -188 8529 -172
rect 8577 -176 8607 -150
rect 8673 -172 8703 -150
rect 8463 -222 8479 -188
rect 8513 -222 8529 -188
rect 8463 -238 8529 -222
rect 8655 -188 8721 -172
rect 8769 -176 8799 -150
rect 8865 -172 8895 -150
rect 8655 -222 8671 -188
rect 8705 -222 8721 -188
rect 8655 -238 8721 -222
rect 8847 -188 8913 -172
rect 8961 -176 8991 -150
rect 9057 -172 9087 -150
rect 8847 -222 8863 -188
rect 8897 -222 8913 -188
rect 8847 -238 8913 -222
rect 9039 -188 9105 -172
rect 9153 -176 9183 -150
rect 9249 -172 9279 -150
rect 9039 -222 9055 -188
rect 9089 -222 9105 -188
rect 9039 -238 9105 -222
rect 9231 -188 9297 -172
rect 9345 -176 9375 -150
rect 9441 -172 9471 -150
rect 9231 -222 9247 -188
rect 9281 -222 9297 -188
rect 9231 -238 9297 -222
rect 9423 -188 9489 -172
rect 9537 -176 9567 -150
rect 9633 -172 9663 -150
rect 9423 -222 9439 -188
rect 9473 -222 9489 -188
rect 9423 -238 9489 -222
rect 9615 -188 9681 -172
rect 9729 -176 9759 -150
rect 9825 -172 9855 -150
rect 9615 -222 9631 -188
rect 9665 -222 9681 -188
rect 9615 -238 9681 -222
rect 9807 -188 9873 -172
rect 9921 -176 9951 -150
rect 10017 -172 10047 -150
rect 9807 -222 9823 -188
rect 9857 -222 9873 -188
rect 9807 -238 9873 -222
rect 9999 -188 10065 -172
rect 10113 -176 10143 -150
rect 10209 -172 10239 -150
rect 9999 -222 10015 -188
rect 10049 -222 10065 -188
rect 9999 -238 10065 -222
rect 10191 -188 10257 -172
rect 10305 -176 10335 -150
rect 10401 -172 10431 -150
rect 10191 -222 10207 -188
rect 10241 -222 10257 -188
rect 10191 -238 10257 -222
rect 10383 -188 10449 -172
rect 10497 -176 10527 -150
rect 10593 -172 10623 -150
rect 10383 -222 10399 -188
rect 10433 -222 10449 -188
rect 10383 -238 10449 -222
rect 10575 -188 10641 -172
rect 10689 -176 10719 -150
rect 10785 -172 10815 -150
rect 10575 -222 10591 -188
rect 10625 -222 10641 -188
rect 10575 -238 10641 -222
rect 10767 -188 10833 -172
rect 10881 -176 10911 -150
rect 10977 -172 11007 -150
rect 10767 -222 10783 -188
rect 10817 -222 10833 -188
rect 10767 -238 10833 -222
rect 10959 -188 11025 -172
rect 11073 -176 11103 -150
rect 11169 -172 11199 -150
rect 10959 -222 10975 -188
rect 11009 -222 11025 -188
rect 10959 -238 11025 -222
rect 11151 -188 11217 -172
rect 11265 -176 11295 -150
rect 11361 -172 11391 -150
rect 11151 -222 11167 -188
rect 11201 -222 11217 -188
rect 11151 -238 11217 -222
rect 11343 -188 11409 -172
rect 11457 -176 11487 -150
rect 11553 -172 11583 -150
rect 11343 -222 11359 -188
rect 11393 -222 11409 -188
rect 11343 -238 11409 -222
rect 11535 -188 11601 -172
rect 11649 -176 11679 -150
rect 11745 -172 11775 -150
rect 11535 -222 11551 -188
rect 11585 -222 11601 -188
rect 11535 -238 11601 -222
rect 11727 -188 11793 -172
rect 11841 -176 11871 -150
rect 11937 -172 11967 -150
rect 11727 -222 11743 -188
rect 11777 -222 11793 -188
rect 11727 -238 11793 -222
rect 11919 -188 11985 -172
rect 12033 -176 12063 -150
rect 12129 -172 12159 -150
rect 11919 -222 11935 -188
rect 11969 -222 11985 -188
rect 11919 -238 11985 -222
rect 12111 -188 12177 -172
rect 12225 -176 12255 -150
rect 12321 -172 12351 -150
rect 12111 -222 12127 -188
rect 12161 -222 12177 -188
rect 12111 -238 12177 -222
rect 12303 -188 12369 -172
rect 12417 -176 12447 -150
rect 12513 -172 12543 -150
rect 12303 -222 12319 -188
rect 12353 -222 12369 -188
rect 12303 -238 12369 -222
rect 12495 -188 12561 -172
rect 12609 -176 12639 -150
rect 12705 -172 12735 -150
rect 12495 -222 12511 -188
rect 12545 -222 12561 -188
rect 12495 -238 12561 -222
rect 12687 -188 12753 -172
rect 12801 -176 12831 -150
rect 12897 -172 12927 -150
rect 12687 -222 12703 -188
rect 12737 -222 12753 -188
rect 12687 -238 12753 -222
rect 12879 -188 12945 -172
rect 12993 -176 13023 -150
rect 13089 -172 13119 -150
rect 12879 -222 12895 -188
rect 12929 -222 12945 -188
rect 12879 -238 12945 -222
rect 13071 -188 13137 -172
rect 13185 -176 13215 -150
rect 13281 -172 13311 -150
rect 13071 -222 13087 -188
rect 13121 -222 13137 -188
rect 13071 -238 13137 -222
rect 13263 -188 13329 -172
rect 13377 -176 13407 -150
rect 13473 -172 13503 -150
rect 13263 -222 13279 -188
rect 13313 -222 13329 -188
rect 13263 -238 13329 -222
rect 13455 -188 13521 -172
rect 13569 -176 13599 -150
rect 13665 -172 13695 -150
rect 13455 -222 13471 -188
rect 13505 -222 13521 -188
rect 13455 -238 13521 -222
rect 13647 -188 13713 -172
rect 13761 -176 13791 -150
rect 13857 -172 13887 -150
rect 13647 -222 13663 -188
rect 13697 -222 13713 -188
rect 13647 -238 13713 -222
rect 13839 -188 13905 -172
rect 13953 -176 13983 -150
rect 14049 -172 14079 -150
rect 13839 -222 13855 -188
rect 13889 -222 13905 -188
rect 13839 -238 13905 -222
rect 14031 -188 14097 -172
rect 14145 -176 14175 -150
rect 14241 -172 14271 -150
rect 14031 -222 14047 -188
rect 14081 -222 14097 -188
rect 14031 -238 14097 -222
rect 14223 -188 14289 -172
rect 14337 -176 14367 -150
rect 14433 -172 14463 -150
rect 14223 -222 14239 -188
rect 14273 -222 14289 -188
rect 14223 -238 14289 -222
rect 14415 -188 14481 -172
rect 14529 -176 14559 -150
rect 14625 -172 14655 -150
rect 14415 -222 14431 -188
rect 14465 -222 14481 -188
rect 14415 -238 14481 -222
rect 14607 -188 14673 -172
rect 14721 -176 14751 -150
rect 14817 -172 14847 -150
rect 14607 -222 14623 -188
rect 14657 -222 14673 -188
rect 14607 -238 14673 -222
rect 14799 -188 14865 -172
rect 14913 -176 14943 -150
rect 15009 -172 15039 -150
rect 14799 -222 14815 -188
rect 14849 -222 14865 -188
rect 14799 -238 14865 -222
rect 14991 -188 15057 -172
rect 15105 -176 15135 -150
rect 15201 -172 15231 -150
rect 14991 -222 15007 -188
rect 15041 -222 15057 -188
rect 14991 -238 15057 -222
rect 15183 -188 15249 -172
rect 15297 -176 15327 -150
rect 15393 -172 15423 -150
rect 15183 -222 15199 -188
rect 15233 -222 15249 -188
rect 15183 -238 15249 -222
rect 15375 -188 15441 -172
rect 15489 -176 15519 -150
rect 15585 -172 15615 -150
rect 15375 -222 15391 -188
rect 15425 -222 15441 -188
rect 15375 -238 15441 -222
rect 15567 -188 15633 -172
rect 15681 -176 15711 -150
rect 15777 -172 15807 -150
rect 15567 -222 15583 -188
rect 15617 -222 15633 -188
rect 15567 -238 15633 -222
rect 15759 -188 15825 -172
rect 15873 -176 15903 -150
rect 15969 -172 15999 -150
rect 15759 -222 15775 -188
rect 15809 -222 15825 -188
rect 15759 -238 15825 -222
rect 15951 -188 16017 -172
rect 16065 -176 16095 -150
rect 16161 -172 16191 -150
rect 15951 -222 15967 -188
rect 16001 -222 16017 -188
rect 15951 -238 16017 -222
rect 16143 -188 16209 -172
rect 16257 -176 16287 -150
rect 16353 -172 16383 -150
rect 16143 -222 16159 -188
rect 16193 -222 16209 -188
rect 16143 -238 16209 -222
rect 16335 -188 16401 -172
rect 16449 -176 16479 -150
rect 16545 -172 16575 -150
rect 16335 -222 16351 -188
rect 16385 -222 16401 -188
rect 16335 -238 16401 -222
rect 16527 -188 16593 -172
rect 16641 -176 16671 -150
rect 16737 -172 16767 -150
rect 16527 -222 16543 -188
rect 16577 -222 16593 -188
rect 16527 -238 16593 -222
rect 16719 -188 16785 -172
rect 16833 -176 16863 -150
rect 16929 -172 16959 -150
rect 16719 -222 16735 -188
rect 16769 -222 16785 -188
rect 16719 -238 16785 -222
rect 16911 -188 16977 -172
rect 17025 -176 17055 -150
rect 17121 -172 17151 -150
rect 16911 -222 16927 -188
rect 16961 -222 16977 -188
rect 16911 -238 16977 -222
rect 17103 -188 17169 -172
rect 17217 -176 17247 -150
rect 17313 -172 17343 -150
rect 17103 -222 17119 -188
rect 17153 -222 17169 -188
rect 17103 -238 17169 -222
rect 17295 -188 17361 -172
rect 17409 -176 17439 -150
rect 17505 -172 17535 -150
rect 17295 -222 17311 -188
rect 17345 -222 17361 -188
rect 17295 -238 17361 -222
rect 17487 -188 17553 -172
rect 17601 -176 17631 -150
rect 17697 -172 17727 -150
rect 17487 -222 17503 -188
rect 17537 -222 17553 -188
rect 17487 -238 17553 -222
rect 17679 -188 17745 -172
rect 17793 -176 17823 -150
rect 17889 -172 17919 -150
rect 17679 -222 17695 -188
rect 17729 -222 17745 -188
rect 17679 -238 17745 -222
rect 17871 -188 17937 -172
rect 17985 -176 18015 -150
rect 18081 -172 18111 -150
rect 17871 -222 17887 -188
rect 17921 -222 17937 -188
rect 17871 -238 17937 -222
rect 18063 -188 18129 -172
rect 18177 -176 18207 -150
rect 18273 -172 18303 -150
rect 18063 -222 18079 -188
rect 18113 -222 18129 -188
rect 18063 -238 18129 -222
rect 18255 -188 18321 -172
rect 18369 -176 18399 -150
rect 18465 -172 18495 -150
rect 18255 -222 18271 -188
rect 18305 -222 18321 -188
rect 18255 -238 18321 -222
rect 18447 -188 18513 -172
rect 18561 -176 18591 -150
rect 18657 -172 18687 -150
rect 18447 -222 18463 -188
rect 18497 -222 18513 -188
rect 18447 -238 18513 -222
rect 18639 -188 18705 -172
rect 18753 -176 18783 -150
rect 18849 -172 18879 -150
rect 18639 -222 18655 -188
rect 18689 -222 18705 -188
rect 18639 -238 18705 -222
rect 18831 -188 18897 -172
rect 18945 -176 18975 -150
rect 19041 -172 19071 -150
rect 18831 -222 18847 -188
rect 18881 -222 18897 -188
rect 18831 -238 18897 -222
rect 19023 -188 19089 -172
rect 19137 -176 19167 -150
rect 19023 -222 19039 -188
rect 19073 -222 19089 -188
rect 19023 -238 19089 -222
<< polycont >>
rect -19073 188 -19039 222
rect -18881 188 -18847 222
rect -18689 188 -18655 222
rect -18497 188 -18463 222
rect -18305 188 -18271 222
rect -18113 188 -18079 222
rect -17921 188 -17887 222
rect -17729 188 -17695 222
rect -17537 188 -17503 222
rect -17345 188 -17311 222
rect -17153 188 -17119 222
rect -16961 188 -16927 222
rect -16769 188 -16735 222
rect -16577 188 -16543 222
rect -16385 188 -16351 222
rect -16193 188 -16159 222
rect -16001 188 -15967 222
rect -15809 188 -15775 222
rect -15617 188 -15583 222
rect -15425 188 -15391 222
rect -15233 188 -15199 222
rect -15041 188 -15007 222
rect -14849 188 -14815 222
rect -14657 188 -14623 222
rect -14465 188 -14431 222
rect -14273 188 -14239 222
rect -14081 188 -14047 222
rect -13889 188 -13855 222
rect -13697 188 -13663 222
rect -13505 188 -13471 222
rect -13313 188 -13279 222
rect -13121 188 -13087 222
rect -12929 188 -12895 222
rect -12737 188 -12703 222
rect -12545 188 -12511 222
rect -12353 188 -12319 222
rect -12161 188 -12127 222
rect -11969 188 -11935 222
rect -11777 188 -11743 222
rect -11585 188 -11551 222
rect -11393 188 -11359 222
rect -11201 188 -11167 222
rect -11009 188 -10975 222
rect -10817 188 -10783 222
rect -10625 188 -10591 222
rect -10433 188 -10399 222
rect -10241 188 -10207 222
rect -10049 188 -10015 222
rect -9857 188 -9823 222
rect -9665 188 -9631 222
rect -9473 188 -9439 222
rect -9281 188 -9247 222
rect -9089 188 -9055 222
rect -8897 188 -8863 222
rect -8705 188 -8671 222
rect -8513 188 -8479 222
rect -8321 188 -8287 222
rect -8129 188 -8095 222
rect -7937 188 -7903 222
rect -7745 188 -7711 222
rect -7553 188 -7519 222
rect -7361 188 -7327 222
rect -7169 188 -7135 222
rect -6977 188 -6943 222
rect -6785 188 -6751 222
rect -6593 188 -6559 222
rect -6401 188 -6367 222
rect -6209 188 -6175 222
rect -6017 188 -5983 222
rect -5825 188 -5791 222
rect -5633 188 -5599 222
rect -5441 188 -5407 222
rect -5249 188 -5215 222
rect -5057 188 -5023 222
rect -4865 188 -4831 222
rect -4673 188 -4639 222
rect -4481 188 -4447 222
rect -4289 188 -4255 222
rect -4097 188 -4063 222
rect -3905 188 -3871 222
rect -3713 188 -3679 222
rect -3521 188 -3487 222
rect -3329 188 -3295 222
rect -3137 188 -3103 222
rect -2945 188 -2911 222
rect -2753 188 -2719 222
rect -2561 188 -2527 222
rect -2369 188 -2335 222
rect -2177 188 -2143 222
rect -1985 188 -1951 222
rect -1793 188 -1759 222
rect -1601 188 -1567 222
rect -1409 188 -1375 222
rect -1217 188 -1183 222
rect -1025 188 -991 222
rect -833 188 -799 222
rect -641 188 -607 222
rect -449 188 -415 222
rect -257 188 -223 222
rect -65 188 -31 222
rect 127 188 161 222
rect 319 188 353 222
rect 511 188 545 222
rect 703 188 737 222
rect 895 188 929 222
rect 1087 188 1121 222
rect 1279 188 1313 222
rect 1471 188 1505 222
rect 1663 188 1697 222
rect 1855 188 1889 222
rect 2047 188 2081 222
rect 2239 188 2273 222
rect 2431 188 2465 222
rect 2623 188 2657 222
rect 2815 188 2849 222
rect 3007 188 3041 222
rect 3199 188 3233 222
rect 3391 188 3425 222
rect 3583 188 3617 222
rect 3775 188 3809 222
rect 3967 188 4001 222
rect 4159 188 4193 222
rect 4351 188 4385 222
rect 4543 188 4577 222
rect 4735 188 4769 222
rect 4927 188 4961 222
rect 5119 188 5153 222
rect 5311 188 5345 222
rect 5503 188 5537 222
rect 5695 188 5729 222
rect 5887 188 5921 222
rect 6079 188 6113 222
rect 6271 188 6305 222
rect 6463 188 6497 222
rect 6655 188 6689 222
rect 6847 188 6881 222
rect 7039 188 7073 222
rect 7231 188 7265 222
rect 7423 188 7457 222
rect 7615 188 7649 222
rect 7807 188 7841 222
rect 7999 188 8033 222
rect 8191 188 8225 222
rect 8383 188 8417 222
rect 8575 188 8609 222
rect 8767 188 8801 222
rect 8959 188 8993 222
rect 9151 188 9185 222
rect 9343 188 9377 222
rect 9535 188 9569 222
rect 9727 188 9761 222
rect 9919 188 9953 222
rect 10111 188 10145 222
rect 10303 188 10337 222
rect 10495 188 10529 222
rect 10687 188 10721 222
rect 10879 188 10913 222
rect 11071 188 11105 222
rect 11263 188 11297 222
rect 11455 188 11489 222
rect 11647 188 11681 222
rect 11839 188 11873 222
rect 12031 188 12065 222
rect 12223 188 12257 222
rect 12415 188 12449 222
rect 12607 188 12641 222
rect 12799 188 12833 222
rect 12991 188 13025 222
rect 13183 188 13217 222
rect 13375 188 13409 222
rect 13567 188 13601 222
rect 13759 188 13793 222
rect 13951 188 13985 222
rect 14143 188 14177 222
rect 14335 188 14369 222
rect 14527 188 14561 222
rect 14719 188 14753 222
rect 14911 188 14945 222
rect 15103 188 15137 222
rect 15295 188 15329 222
rect 15487 188 15521 222
rect 15679 188 15713 222
rect 15871 188 15905 222
rect 16063 188 16097 222
rect 16255 188 16289 222
rect 16447 188 16481 222
rect 16639 188 16673 222
rect 16831 188 16865 222
rect 17023 188 17057 222
rect 17215 188 17249 222
rect 17407 188 17441 222
rect 17599 188 17633 222
rect 17791 188 17825 222
rect 17983 188 18017 222
rect 18175 188 18209 222
rect 18367 188 18401 222
rect 18559 188 18593 222
rect 18751 188 18785 222
rect 18943 188 18977 222
rect 19135 188 19169 222
rect -19169 -222 -19135 -188
rect -18977 -222 -18943 -188
rect -18785 -222 -18751 -188
rect -18593 -222 -18559 -188
rect -18401 -222 -18367 -188
rect -18209 -222 -18175 -188
rect -18017 -222 -17983 -188
rect -17825 -222 -17791 -188
rect -17633 -222 -17599 -188
rect -17441 -222 -17407 -188
rect -17249 -222 -17215 -188
rect -17057 -222 -17023 -188
rect -16865 -222 -16831 -188
rect -16673 -222 -16639 -188
rect -16481 -222 -16447 -188
rect -16289 -222 -16255 -188
rect -16097 -222 -16063 -188
rect -15905 -222 -15871 -188
rect -15713 -222 -15679 -188
rect -15521 -222 -15487 -188
rect -15329 -222 -15295 -188
rect -15137 -222 -15103 -188
rect -14945 -222 -14911 -188
rect -14753 -222 -14719 -188
rect -14561 -222 -14527 -188
rect -14369 -222 -14335 -188
rect -14177 -222 -14143 -188
rect -13985 -222 -13951 -188
rect -13793 -222 -13759 -188
rect -13601 -222 -13567 -188
rect -13409 -222 -13375 -188
rect -13217 -222 -13183 -188
rect -13025 -222 -12991 -188
rect -12833 -222 -12799 -188
rect -12641 -222 -12607 -188
rect -12449 -222 -12415 -188
rect -12257 -222 -12223 -188
rect -12065 -222 -12031 -188
rect -11873 -222 -11839 -188
rect -11681 -222 -11647 -188
rect -11489 -222 -11455 -188
rect -11297 -222 -11263 -188
rect -11105 -222 -11071 -188
rect -10913 -222 -10879 -188
rect -10721 -222 -10687 -188
rect -10529 -222 -10495 -188
rect -10337 -222 -10303 -188
rect -10145 -222 -10111 -188
rect -9953 -222 -9919 -188
rect -9761 -222 -9727 -188
rect -9569 -222 -9535 -188
rect -9377 -222 -9343 -188
rect -9185 -222 -9151 -188
rect -8993 -222 -8959 -188
rect -8801 -222 -8767 -188
rect -8609 -222 -8575 -188
rect -8417 -222 -8383 -188
rect -8225 -222 -8191 -188
rect -8033 -222 -7999 -188
rect -7841 -222 -7807 -188
rect -7649 -222 -7615 -188
rect -7457 -222 -7423 -188
rect -7265 -222 -7231 -188
rect -7073 -222 -7039 -188
rect -6881 -222 -6847 -188
rect -6689 -222 -6655 -188
rect -6497 -222 -6463 -188
rect -6305 -222 -6271 -188
rect -6113 -222 -6079 -188
rect -5921 -222 -5887 -188
rect -5729 -222 -5695 -188
rect -5537 -222 -5503 -188
rect -5345 -222 -5311 -188
rect -5153 -222 -5119 -188
rect -4961 -222 -4927 -188
rect -4769 -222 -4735 -188
rect -4577 -222 -4543 -188
rect -4385 -222 -4351 -188
rect -4193 -222 -4159 -188
rect -4001 -222 -3967 -188
rect -3809 -222 -3775 -188
rect -3617 -222 -3583 -188
rect -3425 -222 -3391 -188
rect -3233 -222 -3199 -188
rect -3041 -222 -3007 -188
rect -2849 -222 -2815 -188
rect -2657 -222 -2623 -188
rect -2465 -222 -2431 -188
rect -2273 -222 -2239 -188
rect -2081 -222 -2047 -188
rect -1889 -222 -1855 -188
rect -1697 -222 -1663 -188
rect -1505 -222 -1471 -188
rect -1313 -222 -1279 -188
rect -1121 -222 -1087 -188
rect -929 -222 -895 -188
rect -737 -222 -703 -188
rect -545 -222 -511 -188
rect -353 -222 -319 -188
rect -161 -222 -127 -188
rect 31 -222 65 -188
rect 223 -222 257 -188
rect 415 -222 449 -188
rect 607 -222 641 -188
rect 799 -222 833 -188
rect 991 -222 1025 -188
rect 1183 -222 1217 -188
rect 1375 -222 1409 -188
rect 1567 -222 1601 -188
rect 1759 -222 1793 -188
rect 1951 -222 1985 -188
rect 2143 -222 2177 -188
rect 2335 -222 2369 -188
rect 2527 -222 2561 -188
rect 2719 -222 2753 -188
rect 2911 -222 2945 -188
rect 3103 -222 3137 -188
rect 3295 -222 3329 -188
rect 3487 -222 3521 -188
rect 3679 -222 3713 -188
rect 3871 -222 3905 -188
rect 4063 -222 4097 -188
rect 4255 -222 4289 -188
rect 4447 -222 4481 -188
rect 4639 -222 4673 -188
rect 4831 -222 4865 -188
rect 5023 -222 5057 -188
rect 5215 -222 5249 -188
rect 5407 -222 5441 -188
rect 5599 -222 5633 -188
rect 5791 -222 5825 -188
rect 5983 -222 6017 -188
rect 6175 -222 6209 -188
rect 6367 -222 6401 -188
rect 6559 -222 6593 -188
rect 6751 -222 6785 -188
rect 6943 -222 6977 -188
rect 7135 -222 7169 -188
rect 7327 -222 7361 -188
rect 7519 -222 7553 -188
rect 7711 -222 7745 -188
rect 7903 -222 7937 -188
rect 8095 -222 8129 -188
rect 8287 -222 8321 -188
rect 8479 -222 8513 -188
rect 8671 -222 8705 -188
rect 8863 -222 8897 -188
rect 9055 -222 9089 -188
rect 9247 -222 9281 -188
rect 9439 -222 9473 -188
rect 9631 -222 9665 -188
rect 9823 -222 9857 -188
rect 10015 -222 10049 -188
rect 10207 -222 10241 -188
rect 10399 -222 10433 -188
rect 10591 -222 10625 -188
rect 10783 -222 10817 -188
rect 10975 -222 11009 -188
rect 11167 -222 11201 -188
rect 11359 -222 11393 -188
rect 11551 -222 11585 -188
rect 11743 -222 11777 -188
rect 11935 -222 11969 -188
rect 12127 -222 12161 -188
rect 12319 -222 12353 -188
rect 12511 -222 12545 -188
rect 12703 -222 12737 -188
rect 12895 -222 12929 -188
rect 13087 -222 13121 -188
rect 13279 -222 13313 -188
rect 13471 -222 13505 -188
rect 13663 -222 13697 -188
rect 13855 -222 13889 -188
rect 14047 -222 14081 -188
rect 14239 -222 14273 -188
rect 14431 -222 14465 -188
rect 14623 -222 14657 -188
rect 14815 -222 14849 -188
rect 15007 -222 15041 -188
rect 15199 -222 15233 -188
rect 15391 -222 15425 -188
rect 15583 -222 15617 -188
rect 15775 -222 15809 -188
rect 15967 -222 16001 -188
rect 16159 -222 16193 -188
rect 16351 -222 16385 -188
rect 16543 -222 16577 -188
rect 16735 -222 16769 -188
rect 16927 -222 16961 -188
rect 17119 -222 17153 -188
rect 17311 -222 17345 -188
rect 17503 -222 17537 -188
rect 17695 -222 17729 -188
rect 17887 -222 17921 -188
rect 18079 -222 18113 -188
rect 18271 -222 18305 -188
rect 18463 -222 18497 -188
rect 18655 -222 18689 -188
rect 18847 -222 18881 -188
rect 19039 -222 19073 -188
<< locali >>
rect -19331 290 -19235 324
rect 19235 290 19331 324
rect -19331 228 -19297 290
rect 19297 228 19331 290
rect -19089 188 -19073 222
rect -19039 188 -19023 222
rect -18897 188 -18881 222
rect -18847 188 -18831 222
rect -18705 188 -18689 222
rect -18655 188 -18639 222
rect -18513 188 -18497 222
rect -18463 188 -18447 222
rect -18321 188 -18305 222
rect -18271 188 -18255 222
rect -18129 188 -18113 222
rect -18079 188 -18063 222
rect -17937 188 -17921 222
rect -17887 188 -17871 222
rect -17745 188 -17729 222
rect -17695 188 -17679 222
rect -17553 188 -17537 222
rect -17503 188 -17487 222
rect -17361 188 -17345 222
rect -17311 188 -17295 222
rect -17169 188 -17153 222
rect -17119 188 -17103 222
rect -16977 188 -16961 222
rect -16927 188 -16911 222
rect -16785 188 -16769 222
rect -16735 188 -16719 222
rect -16593 188 -16577 222
rect -16543 188 -16527 222
rect -16401 188 -16385 222
rect -16351 188 -16335 222
rect -16209 188 -16193 222
rect -16159 188 -16143 222
rect -16017 188 -16001 222
rect -15967 188 -15951 222
rect -15825 188 -15809 222
rect -15775 188 -15759 222
rect -15633 188 -15617 222
rect -15583 188 -15567 222
rect -15441 188 -15425 222
rect -15391 188 -15375 222
rect -15249 188 -15233 222
rect -15199 188 -15183 222
rect -15057 188 -15041 222
rect -15007 188 -14991 222
rect -14865 188 -14849 222
rect -14815 188 -14799 222
rect -14673 188 -14657 222
rect -14623 188 -14607 222
rect -14481 188 -14465 222
rect -14431 188 -14415 222
rect -14289 188 -14273 222
rect -14239 188 -14223 222
rect -14097 188 -14081 222
rect -14047 188 -14031 222
rect -13905 188 -13889 222
rect -13855 188 -13839 222
rect -13713 188 -13697 222
rect -13663 188 -13647 222
rect -13521 188 -13505 222
rect -13471 188 -13455 222
rect -13329 188 -13313 222
rect -13279 188 -13263 222
rect -13137 188 -13121 222
rect -13087 188 -13071 222
rect -12945 188 -12929 222
rect -12895 188 -12879 222
rect -12753 188 -12737 222
rect -12703 188 -12687 222
rect -12561 188 -12545 222
rect -12511 188 -12495 222
rect -12369 188 -12353 222
rect -12319 188 -12303 222
rect -12177 188 -12161 222
rect -12127 188 -12111 222
rect -11985 188 -11969 222
rect -11935 188 -11919 222
rect -11793 188 -11777 222
rect -11743 188 -11727 222
rect -11601 188 -11585 222
rect -11551 188 -11535 222
rect -11409 188 -11393 222
rect -11359 188 -11343 222
rect -11217 188 -11201 222
rect -11167 188 -11151 222
rect -11025 188 -11009 222
rect -10975 188 -10959 222
rect -10833 188 -10817 222
rect -10783 188 -10767 222
rect -10641 188 -10625 222
rect -10591 188 -10575 222
rect -10449 188 -10433 222
rect -10399 188 -10383 222
rect -10257 188 -10241 222
rect -10207 188 -10191 222
rect -10065 188 -10049 222
rect -10015 188 -9999 222
rect -9873 188 -9857 222
rect -9823 188 -9807 222
rect -9681 188 -9665 222
rect -9631 188 -9615 222
rect -9489 188 -9473 222
rect -9439 188 -9423 222
rect -9297 188 -9281 222
rect -9247 188 -9231 222
rect -9105 188 -9089 222
rect -9055 188 -9039 222
rect -8913 188 -8897 222
rect -8863 188 -8847 222
rect -8721 188 -8705 222
rect -8671 188 -8655 222
rect -8529 188 -8513 222
rect -8479 188 -8463 222
rect -8337 188 -8321 222
rect -8287 188 -8271 222
rect -8145 188 -8129 222
rect -8095 188 -8079 222
rect -7953 188 -7937 222
rect -7903 188 -7887 222
rect -7761 188 -7745 222
rect -7711 188 -7695 222
rect -7569 188 -7553 222
rect -7519 188 -7503 222
rect -7377 188 -7361 222
rect -7327 188 -7311 222
rect -7185 188 -7169 222
rect -7135 188 -7119 222
rect -6993 188 -6977 222
rect -6943 188 -6927 222
rect -6801 188 -6785 222
rect -6751 188 -6735 222
rect -6609 188 -6593 222
rect -6559 188 -6543 222
rect -6417 188 -6401 222
rect -6367 188 -6351 222
rect -6225 188 -6209 222
rect -6175 188 -6159 222
rect -6033 188 -6017 222
rect -5983 188 -5967 222
rect -5841 188 -5825 222
rect -5791 188 -5775 222
rect -5649 188 -5633 222
rect -5599 188 -5583 222
rect -5457 188 -5441 222
rect -5407 188 -5391 222
rect -5265 188 -5249 222
rect -5215 188 -5199 222
rect -5073 188 -5057 222
rect -5023 188 -5007 222
rect -4881 188 -4865 222
rect -4831 188 -4815 222
rect -4689 188 -4673 222
rect -4639 188 -4623 222
rect -4497 188 -4481 222
rect -4447 188 -4431 222
rect -4305 188 -4289 222
rect -4255 188 -4239 222
rect -4113 188 -4097 222
rect -4063 188 -4047 222
rect -3921 188 -3905 222
rect -3871 188 -3855 222
rect -3729 188 -3713 222
rect -3679 188 -3663 222
rect -3537 188 -3521 222
rect -3487 188 -3471 222
rect -3345 188 -3329 222
rect -3295 188 -3279 222
rect -3153 188 -3137 222
rect -3103 188 -3087 222
rect -2961 188 -2945 222
rect -2911 188 -2895 222
rect -2769 188 -2753 222
rect -2719 188 -2703 222
rect -2577 188 -2561 222
rect -2527 188 -2511 222
rect -2385 188 -2369 222
rect -2335 188 -2319 222
rect -2193 188 -2177 222
rect -2143 188 -2127 222
rect -2001 188 -1985 222
rect -1951 188 -1935 222
rect -1809 188 -1793 222
rect -1759 188 -1743 222
rect -1617 188 -1601 222
rect -1567 188 -1551 222
rect -1425 188 -1409 222
rect -1375 188 -1359 222
rect -1233 188 -1217 222
rect -1183 188 -1167 222
rect -1041 188 -1025 222
rect -991 188 -975 222
rect -849 188 -833 222
rect -799 188 -783 222
rect -657 188 -641 222
rect -607 188 -591 222
rect -465 188 -449 222
rect -415 188 -399 222
rect -273 188 -257 222
rect -223 188 -207 222
rect -81 188 -65 222
rect -31 188 -15 222
rect 111 188 127 222
rect 161 188 177 222
rect 303 188 319 222
rect 353 188 369 222
rect 495 188 511 222
rect 545 188 561 222
rect 687 188 703 222
rect 737 188 753 222
rect 879 188 895 222
rect 929 188 945 222
rect 1071 188 1087 222
rect 1121 188 1137 222
rect 1263 188 1279 222
rect 1313 188 1329 222
rect 1455 188 1471 222
rect 1505 188 1521 222
rect 1647 188 1663 222
rect 1697 188 1713 222
rect 1839 188 1855 222
rect 1889 188 1905 222
rect 2031 188 2047 222
rect 2081 188 2097 222
rect 2223 188 2239 222
rect 2273 188 2289 222
rect 2415 188 2431 222
rect 2465 188 2481 222
rect 2607 188 2623 222
rect 2657 188 2673 222
rect 2799 188 2815 222
rect 2849 188 2865 222
rect 2991 188 3007 222
rect 3041 188 3057 222
rect 3183 188 3199 222
rect 3233 188 3249 222
rect 3375 188 3391 222
rect 3425 188 3441 222
rect 3567 188 3583 222
rect 3617 188 3633 222
rect 3759 188 3775 222
rect 3809 188 3825 222
rect 3951 188 3967 222
rect 4001 188 4017 222
rect 4143 188 4159 222
rect 4193 188 4209 222
rect 4335 188 4351 222
rect 4385 188 4401 222
rect 4527 188 4543 222
rect 4577 188 4593 222
rect 4719 188 4735 222
rect 4769 188 4785 222
rect 4911 188 4927 222
rect 4961 188 4977 222
rect 5103 188 5119 222
rect 5153 188 5169 222
rect 5295 188 5311 222
rect 5345 188 5361 222
rect 5487 188 5503 222
rect 5537 188 5553 222
rect 5679 188 5695 222
rect 5729 188 5745 222
rect 5871 188 5887 222
rect 5921 188 5937 222
rect 6063 188 6079 222
rect 6113 188 6129 222
rect 6255 188 6271 222
rect 6305 188 6321 222
rect 6447 188 6463 222
rect 6497 188 6513 222
rect 6639 188 6655 222
rect 6689 188 6705 222
rect 6831 188 6847 222
rect 6881 188 6897 222
rect 7023 188 7039 222
rect 7073 188 7089 222
rect 7215 188 7231 222
rect 7265 188 7281 222
rect 7407 188 7423 222
rect 7457 188 7473 222
rect 7599 188 7615 222
rect 7649 188 7665 222
rect 7791 188 7807 222
rect 7841 188 7857 222
rect 7983 188 7999 222
rect 8033 188 8049 222
rect 8175 188 8191 222
rect 8225 188 8241 222
rect 8367 188 8383 222
rect 8417 188 8433 222
rect 8559 188 8575 222
rect 8609 188 8625 222
rect 8751 188 8767 222
rect 8801 188 8817 222
rect 8943 188 8959 222
rect 8993 188 9009 222
rect 9135 188 9151 222
rect 9185 188 9201 222
rect 9327 188 9343 222
rect 9377 188 9393 222
rect 9519 188 9535 222
rect 9569 188 9585 222
rect 9711 188 9727 222
rect 9761 188 9777 222
rect 9903 188 9919 222
rect 9953 188 9969 222
rect 10095 188 10111 222
rect 10145 188 10161 222
rect 10287 188 10303 222
rect 10337 188 10353 222
rect 10479 188 10495 222
rect 10529 188 10545 222
rect 10671 188 10687 222
rect 10721 188 10737 222
rect 10863 188 10879 222
rect 10913 188 10929 222
rect 11055 188 11071 222
rect 11105 188 11121 222
rect 11247 188 11263 222
rect 11297 188 11313 222
rect 11439 188 11455 222
rect 11489 188 11505 222
rect 11631 188 11647 222
rect 11681 188 11697 222
rect 11823 188 11839 222
rect 11873 188 11889 222
rect 12015 188 12031 222
rect 12065 188 12081 222
rect 12207 188 12223 222
rect 12257 188 12273 222
rect 12399 188 12415 222
rect 12449 188 12465 222
rect 12591 188 12607 222
rect 12641 188 12657 222
rect 12783 188 12799 222
rect 12833 188 12849 222
rect 12975 188 12991 222
rect 13025 188 13041 222
rect 13167 188 13183 222
rect 13217 188 13233 222
rect 13359 188 13375 222
rect 13409 188 13425 222
rect 13551 188 13567 222
rect 13601 188 13617 222
rect 13743 188 13759 222
rect 13793 188 13809 222
rect 13935 188 13951 222
rect 13985 188 14001 222
rect 14127 188 14143 222
rect 14177 188 14193 222
rect 14319 188 14335 222
rect 14369 188 14385 222
rect 14511 188 14527 222
rect 14561 188 14577 222
rect 14703 188 14719 222
rect 14753 188 14769 222
rect 14895 188 14911 222
rect 14945 188 14961 222
rect 15087 188 15103 222
rect 15137 188 15153 222
rect 15279 188 15295 222
rect 15329 188 15345 222
rect 15471 188 15487 222
rect 15521 188 15537 222
rect 15663 188 15679 222
rect 15713 188 15729 222
rect 15855 188 15871 222
rect 15905 188 15921 222
rect 16047 188 16063 222
rect 16097 188 16113 222
rect 16239 188 16255 222
rect 16289 188 16305 222
rect 16431 188 16447 222
rect 16481 188 16497 222
rect 16623 188 16639 222
rect 16673 188 16689 222
rect 16815 188 16831 222
rect 16865 188 16881 222
rect 17007 188 17023 222
rect 17057 188 17073 222
rect 17199 188 17215 222
rect 17249 188 17265 222
rect 17391 188 17407 222
rect 17441 188 17457 222
rect 17583 188 17599 222
rect 17633 188 17649 222
rect 17775 188 17791 222
rect 17825 188 17841 222
rect 17967 188 17983 222
rect 18017 188 18033 222
rect 18159 188 18175 222
rect 18209 188 18225 222
rect 18351 188 18367 222
rect 18401 188 18417 222
rect 18543 188 18559 222
rect 18593 188 18609 222
rect 18735 188 18751 222
rect 18785 188 18801 222
rect 18927 188 18943 222
rect 18977 188 18993 222
rect 19119 188 19135 222
rect 19169 188 19185 222
rect -19217 138 -19183 154
rect -19217 -154 -19183 -138
rect -19121 138 -19087 154
rect -19121 -154 -19087 -138
rect -19025 138 -18991 154
rect -19025 -154 -18991 -138
rect -18929 138 -18895 154
rect -18929 -154 -18895 -138
rect -18833 138 -18799 154
rect -18833 -154 -18799 -138
rect -18737 138 -18703 154
rect -18737 -154 -18703 -138
rect -18641 138 -18607 154
rect -18641 -154 -18607 -138
rect -18545 138 -18511 154
rect -18545 -154 -18511 -138
rect -18449 138 -18415 154
rect -18449 -154 -18415 -138
rect -18353 138 -18319 154
rect -18353 -154 -18319 -138
rect -18257 138 -18223 154
rect -18257 -154 -18223 -138
rect -18161 138 -18127 154
rect -18161 -154 -18127 -138
rect -18065 138 -18031 154
rect -18065 -154 -18031 -138
rect -17969 138 -17935 154
rect -17969 -154 -17935 -138
rect -17873 138 -17839 154
rect -17873 -154 -17839 -138
rect -17777 138 -17743 154
rect -17777 -154 -17743 -138
rect -17681 138 -17647 154
rect -17681 -154 -17647 -138
rect -17585 138 -17551 154
rect -17585 -154 -17551 -138
rect -17489 138 -17455 154
rect -17489 -154 -17455 -138
rect -17393 138 -17359 154
rect -17393 -154 -17359 -138
rect -17297 138 -17263 154
rect -17297 -154 -17263 -138
rect -17201 138 -17167 154
rect -17201 -154 -17167 -138
rect -17105 138 -17071 154
rect -17105 -154 -17071 -138
rect -17009 138 -16975 154
rect -17009 -154 -16975 -138
rect -16913 138 -16879 154
rect -16913 -154 -16879 -138
rect -16817 138 -16783 154
rect -16817 -154 -16783 -138
rect -16721 138 -16687 154
rect -16721 -154 -16687 -138
rect -16625 138 -16591 154
rect -16625 -154 -16591 -138
rect -16529 138 -16495 154
rect -16529 -154 -16495 -138
rect -16433 138 -16399 154
rect -16433 -154 -16399 -138
rect -16337 138 -16303 154
rect -16337 -154 -16303 -138
rect -16241 138 -16207 154
rect -16241 -154 -16207 -138
rect -16145 138 -16111 154
rect -16145 -154 -16111 -138
rect -16049 138 -16015 154
rect -16049 -154 -16015 -138
rect -15953 138 -15919 154
rect -15953 -154 -15919 -138
rect -15857 138 -15823 154
rect -15857 -154 -15823 -138
rect -15761 138 -15727 154
rect -15761 -154 -15727 -138
rect -15665 138 -15631 154
rect -15665 -154 -15631 -138
rect -15569 138 -15535 154
rect -15569 -154 -15535 -138
rect -15473 138 -15439 154
rect -15473 -154 -15439 -138
rect -15377 138 -15343 154
rect -15377 -154 -15343 -138
rect -15281 138 -15247 154
rect -15281 -154 -15247 -138
rect -15185 138 -15151 154
rect -15185 -154 -15151 -138
rect -15089 138 -15055 154
rect -15089 -154 -15055 -138
rect -14993 138 -14959 154
rect -14993 -154 -14959 -138
rect -14897 138 -14863 154
rect -14897 -154 -14863 -138
rect -14801 138 -14767 154
rect -14801 -154 -14767 -138
rect -14705 138 -14671 154
rect -14705 -154 -14671 -138
rect -14609 138 -14575 154
rect -14609 -154 -14575 -138
rect -14513 138 -14479 154
rect -14513 -154 -14479 -138
rect -14417 138 -14383 154
rect -14417 -154 -14383 -138
rect -14321 138 -14287 154
rect -14321 -154 -14287 -138
rect -14225 138 -14191 154
rect -14225 -154 -14191 -138
rect -14129 138 -14095 154
rect -14129 -154 -14095 -138
rect -14033 138 -13999 154
rect -14033 -154 -13999 -138
rect -13937 138 -13903 154
rect -13937 -154 -13903 -138
rect -13841 138 -13807 154
rect -13841 -154 -13807 -138
rect -13745 138 -13711 154
rect -13745 -154 -13711 -138
rect -13649 138 -13615 154
rect -13649 -154 -13615 -138
rect -13553 138 -13519 154
rect -13553 -154 -13519 -138
rect -13457 138 -13423 154
rect -13457 -154 -13423 -138
rect -13361 138 -13327 154
rect -13361 -154 -13327 -138
rect -13265 138 -13231 154
rect -13265 -154 -13231 -138
rect -13169 138 -13135 154
rect -13169 -154 -13135 -138
rect -13073 138 -13039 154
rect -13073 -154 -13039 -138
rect -12977 138 -12943 154
rect -12977 -154 -12943 -138
rect -12881 138 -12847 154
rect -12881 -154 -12847 -138
rect -12785 138 -12751 154
rect -12785 -154 -12751 -138
rect -12689 138 -12655 154
rect -12689 -154 -12655 -138
rect -12593 138 -12559 154
rect -12593 -154 -12559 -138
rect -12497 138 -12463 154
rect -12497 -154 -12463 -138
rect -12401 138 -12367 154
rect -12401 -154 -12367 -138
rect -12305 138 -12271 154
rect -12305 -154 -12271 -138
rect -12209 138 -12175 154
rect -12209 -154 -12175 -138
rect -12113 138 -12079 154
rect -12113 -154 -12079 -138
rect -12017 138 -11983 154
rect -12017 -154 -11983 -138
rect -11921 138 -11887 154
rect -11921 -154 -11887 -138
rect -11825 138 -11791 154
rect -11825 -154 -11791 -138
rect -11729 138 -11695 154
rect -11729 -154 -11695 -138
rect -11633 138 -11599 154
rect -11633 -154 -11599 -138
rect -11537 138 -11503 154
rect -11537 -154 -11503 -138
rect -11441 138 -11407 154
rect -11441 -154 -11407 -138
rect -11345 138 -11311 154
rect -11345 -154 -11311 -138
rect -11249 138 -11215 154
rect -11249 -154 -11215 -138
rect -11153 138 -11119 154
rect -11153 -154 -11119 -138
rect -11057 138 -11023 154
rect -11057 -154 -11023 -138
rect -10961 138 -10927 154
rect -10961 -154 -10927 -138
rect -10865 138 -10831 154
rect -10865 -154 -10831 -138
rect -10769 138 -10735 154
rect -10769 -154 -10735 -138
rect -10673 138 -10639 154
rect -10673 -154 -10639 -138
rect -10577 138 -10543 154
rect -10577 -154 -10543 -138
rect -10481 138 -10447 154
rect -10481 -154 -10447 -138
rect -10385 138 -10351 154
rect -10385 -154 -10351 -138
rect -10289 138 -10255 154
rect -10289 -154 -10255 -138
rect -10193 138 -10159 154
rect -10193 -154 -10159 -138
rect -10097 138 -10063 154
rect -10097 -154 -10063 -138
rect -10001 138 -9967 154
rect -10001 -154 -9967 -138
rect -9905 138 -9871 154
rect -9905 -154 -9871 -138
rect -9809 138 -9775 154
rect -9809 -154 -9775 -138
rect -9713 138 -9679 154
rect -9713 -154 -9679 -138
rect -9617 138 -9583 154
rect -9617 -154 -9583 -138
rect -9521 138 -9487 154
rect -9521 -154 -9487 -138
rect -9425 138 -9391 154
rect -9425 -154 -9391 -138
rect -9329 138 -9295 154
rect -9329 -154 -9295 -138
rect -9233 138 -9199 154
rect -9233 -154 -9199 -138
rect -9137 138 -9103 154
rect -9137 -154 -9103 -138
rect -9041 138 -9007 154
rect -9041 -154 -9007 -138
rect -8945 138 -8911 154
rect -8945 -154 -8911 -138
rect -8849 138 -8815 154
rect -8849 -154 -8815 -138
rect -8753 138 -8719 154
rect -8753 -154 -8719 -138
rect -8657 138 -8623 154
rect -8657 -154 -8623 -138
rect -8561 138 -8527 154
rect -8561 -154 -8527 -138
rect -8465 138 -8431 154
rect -8465 -154 -8431 -138
rect -8369 138 -8335 154
rect -8369 -154 -8335 -138
rect -8273 138 -8239 154
rect -8273 -154 -8239 -138
rect -8177 138 -8143 154
rect -8177 -154 -8143 -138
rect -8081 138 -8047 154
rect -8081 -154 -8047 -138
rect -7985 138 -7951 154
rect -7985 -154 -7951 -138
rect -7889 138 -7855 154
rect -7889 -154 -7855 -138
rect -7793 138 -7759 154
rect -7793 -154 -7759 -138
rect -7697 138 -7663 154
rect -7697 -154 -7663 -138
rect -7601 138 -7567 154
rect -7601 -154 -7567 -138
rect -7505 138 -7471 154
rect -7505 -154 -7471 -138
rect -7409 138 -7375 154
rect -7409 -154 -7375 -138
rect -7313 138 -7279 154
rect -7313 -154 -7279 -138
rect -7217 138 -7183 154
rect -7217 -154 -7183 -138
rect -7121 138 -7087 154
rect -7121 -154 -7087 -138
rect -7025 138 -6991 154
rect -7025 -154 -6991 -138
rect -6929 138 -6895 154
rect -6929 -154 -6895 -138
rect -6833 138 -6799 154
rect -6833 -154 -6799 -138
rect -6737 138 -6703 154
rect -6737 -154 -6703 -138
rect -6641 138 -6607 154
rect -6641 -154 -6607 -138
rect -6545 138 -6511 154
rect -6545 -154 -6511 -138
rect -6449 138 -6415 154
rect -6449 -154 -6415 -138
rect -6353 138 -6319 154
rect -6353 -154 -6319 -138
rect -6257 138 -6223 154
rect -6257 -154 -6223 -138
rect -6161 138 -6127 154
rect -6161 -154 -6127 -138
rect -6065 138 -6031 154
rect -6065 -154 -6031 -138
rect -5969 138 -5935 154
rect -5969 -154 -5935 -138
rect -5873 138 -5839 154
rect -5873 -154 -5839 -138
rect -5777 138 -5743 154
rect -5777 -154 -5743 -138
rect -5681 138 -5647 154
rect -5681 -154 -5647 -138
rect -5585 138 -5551 154
rect -5585 -154 -5551 -138
rect -5489 138 -5455 154
rect -5489 -154 -5455 -138
rect -5393 138 -5359 154
rect -5393 -154 -5359 -138
rect -5297 138 -5263 154
rect -5297 -154 -5263 -138
rect -5201 138 -5167 154
rect -5201 -154 -5167 -138
rect -5105 138 -5071 154
rect -5105 -154 -5071 -138
rect -5009 138 -4975 154
rect -5009 -154 -4975 -138
rect -4913 138 -4879 154
rect -4913 -154 -4879 -138
rect -4817 138 -4783 154
rect -4817 -154 -4783 -138
rect -4721 138 -4687 154
rect -4721 -154 -4687 -138
rect -4625 138 -4591 154
rect -4625 -154 -4591 -138
rect -4529 138 -4495 154
rect -4529 -154 -4495 -138
rect -4433 138 -4399 154
rect -4433 -154 -4399 -138
rect -4337 138 -4303 154
rect -4337 -154 -4303 -138
rect -4241 138 -4207 154
rect -4241 -154 -4207 -138
rect -4145 138 -4111 154
rect -4145 -154 -4111 -138
rect -4049 138 -4015 154
rect -4049 -154 -4015 -138
rect -3953 138 -3919 154
rect -3953 -154 -3919 -138
rect -3857 138 -3823 154
rect -3857 -154 -3823 -138
rect -3761 138 -3727 154
rect -3761 -154 -3727 -138
rect -3665 138 -3631 154
rect -3665 -154 -3631 -138
rect -3569 138 -3535 154
rect -3569 -154 -3535 -138
rect -3473 138 -3439 154
rect -3473 -154 -3439 -138
rect -3377 138 -3343 154
rect -3377 -154 -3343 -138
rect -3281 138 -3247 154
rect -3281 -154 -3247 -138
rect -3185 138 -3151 154
rect -3185 -154 -3151 -138
rect -3089 138 -3055 154
rect -3089 -154 -3055 -138
rect -2993 138 -2959 154
rect -2993 -154 -2959 -138
rect -2897 138 -2863 154
rect -2897 -154 -2863 -138
rect -2801 138 -2767 154
rect -2801 -154 -2767 -138
rect -2705 138 -2671 154
rect -2705 -154 -2671 -138
rect -2609 138 -2575 154
rect -2609 -154 -2575 -138
rect -2513 138 -2479 154
rect -2513 -154 -2479 -138
rect -2417 138 -2383 154
rect -2417 -154 -2383 -138
rect -2321 138 -2287 154
rect -2321 -154 -2287 -138
rect -2225 138 -2191 154
rect -2225 -154 -2191 -138
rect -2129 138 -2095 154
rect -2129 -154 -2095 -138
rect -2033 138 -1999 154
rect -2033 -154 -1999 -138
rect -1937 138 -1903 154
rect -1937 -154 -1903 -138
rect -1841 138 -1807 154
rect -1841 -154 -1807 -138
rect -1745 138 -1711 154
rect -1745 -154 -1711 -138
rect -1649 138 -1615 154
rect -1649 -154 -1615 -138
rect -1553 138 -1519 154
rect -1553 -154 -1519 -138
rect -1457 138 -1423 154
rect -1457 -154 -1423 -138
rect -1361 138 -1327 154
rect -1361 -154 -1327 -138
rect -1265 138 -1231 154
rect -1265 -154 -1231 -138
rect -1169 138 -1135 154
rect -1169 -154 -1135 -138
rect -1073 138 -1039 154
rect -1073 -154 -1039 -138
rect -977 138 -943 154
rect -977 -154 -943 -138
rect -881 138 -847 154
rect -881 -154 -847 -138
rect -785 138 -751 154
rect -785 -154 -751 -138
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect 751 138 785 154
rect 751 -154 785 -138
rect 847 138 881 154
rect 847 -154 881 -138
rect 943 138 977 154
rect 943 -154 977 -138
rect 1039 138 1073 154
rect 1039 -154 1073 -138
rect 1135 138 1169 154
rect 1135 -154 1169 -138
rect 1231 138 1265 154
rect 1231 -154 1265 -138
rect 1327 138 1361 154
rect 1327 -154 1361 -138
rect 1423 138 1457 154
rect 1423 -154 1457 -138
rect 1519 138 1553 154
rect 1519 -154 1553 -138
rect 1615 138 1649 154
rect 1615 -154 1649 -138
rect 1711 138 1745 154
rect 1711 -154 1745 -138
rect 1807 138 1841 154
rect 1807 -154 1841 -138
rect 1903 138 1937 154
rect 1903 -154 1937 -138
rect 1999 138 2033 154
rect 1999 -154 2033 -138
rect 2095 138 2129 154
rect 2095 -154 2129 -138
rect 2191 138 2225 154
rect 2191 -154 2225 -138
rect 2287 138 2321 154
rect 2287 -154 2321 -138
rect 2383 138 2417 154
rect 2383 -154 2417 -138
rect 2479 138 2513 154
rect 2479 -154 2513 -138
rect 2575 138 2609 154
rect 2575 -154 2609 -138
rect 2671 138 2705 154
rect 2671 -154 2705 -138
rect 2767 138 2801 154
rect 2767 -154 2801 -138
rect 2863 138 2897 154
rect 2863 -154 2897 -138
rect 2959 138 2993 154
rect 2959 -154 2993 -138
rect 3055 138 3089 154
rect 3055 -154 3089 -138
rect 3151 138 3185 154
rect 3151 -154 3185 -138
rect 3247 138 3281 154
rect 3247 -154 3281 -138
rect 3343 138 3377 154
rect 3343 -154 3377 -138
rect 3439 138 3473 154
rect 3439 -154 3473 -138
rect 3535 138 3569 154
rect 3535 -154 3569 -138
rect 3631 138 3665 154
rect 3631 -154 3665 -138
rect 3727 138 3761 154
rect 3727 -154 3761 -138
rect 3823 138 3857 154
rect 3823 -154 3857 -138
rect 3919 138 3953 154
rect 3919 -154 3953 -138
rect 4015 138 4049 154
rect 4015 -154 4049 -138
rect 4111 138 4145 154
rect 4111 -154 4145 -138
rect 4207 138 4241 154
rect 4207 -154 4241 -138
rect 4303 138 4337 154
rect 4303 -154 4337 -138
rect 4399 138 4433 154
rect 4399 -154 4433 -138
rect 4495 138 4529 154
rect 4495 -154 4529 -138
rect 4591 138 4625 154
rect 4591 -154 4625 -138
rect 4687 138 4721 154
rect 4687 -154 4721 -138
rect 4783 138 4817 154
rect 4783 -154 4817 -138
rect 4879 138 4913 154
rect 4879 -154 4913 -138
rect 4975 138 5009 154
rect 4975 -154 5009 -138
rect 5071 138 5105 154
rect 5071 -154 5105 -138
rect 5167 138 5201 154
rect 5167 -154 5201 -138
rect 5263 138 5297 154
rect 5263 -154 5297 -138
rect 5359 138 5393 154
rect 5359 -154 5393 -138
rect 5455 138 5489 154
rect 5455 -154 5489 -138
rect 5551 138 5585 154
rect 5551 -154 5585 -138
rect 5647 138 5681 154
rect 5647 -154 5681 -138
rect 5743 138 5777 154
rect 5743 -154 5777 -138
rect 5839 138 5873 154
rect 5839 -154 5873 -138
rect 5935 138 5969 154
rect 5935 -154 5969 -138
rect 6031 138 6065 154
rect 6031 -154 6065 -138
rect 6127 138 6161 154
rect 6127 -154 6161 -138
rect 6223 138 6257 154
rect 6223 -154 6257 -138
rect 6319 138 6353 154
rect 6319 -154 6353 -138
rect 6415 138 6449 154
rect 6415 -154 6449 -138
rect 6511 138 6545 154
rect 6511 -154 6545 -138
rect 6607 138 6641 154
rect 6607 -154 6641 -138
rect 6703 138 6737 154
rect 6703 -154 6737 -138
rect 6799 138 6833 154
rect 6799 -154 6833 -138
rect 6895 138 6929 154
rect 6895 -154 6929 -138
rect 6991 138 7025 154
rect 6991 -154 7025 -138
rect 7087 138 7121 154
rect 7087 -154 7121 -138
rect 7183 138 7217 154
rect 7183 -154 7217 -138
rect 7279 138 7313 154
rect 7279 -154 7313 -138
rect 7375 138 7409 154
rect 7375 -154 7409 -138
rect 7471 138 7505 154
rect 7471 -154 7505 -138
rect 7567 138 7601 154
rect 7567 -154 7601 -138
rect 7663 138 7697 154
rect 7663 -154 7697 -138
rect 7759 138 7793 154
rect 7759 -154 7793 -138
rect 7855 138 7889 154
rect 7855 -154 7889 -138
rect 7951 138 7985 154
rect 7951 -154 7985 -138
rect 8047 138 8081 154
rect 8047 -154 8081 -138
rect 8143 138 8177 154
rect 8143 -154 8177 -138
rect 8239 138 8273 154
rect 8239 -154 8273 -138
rect 8335 138 8369 154
rect 8335 -154 8369 -138
rect 8431 138 8465 154
rect 8431 -154 8465 -138
rect 8527 138 8561 154
rect 8527 -154 8561 -138
rect 8623 138 8657 154
rect 8623 -154 8657 -138
rect 8719 138 8753 154
rect 8719 -154 8753 -138
rect 8815 138 8849 154
rect 8815 -154 8849 -138
rect 8911 138 8945 154
rect 8911 -154 8945 -138
rect 9007 138 9041 154
rect 9007 -154 9041 -138
rect 9103 138 9137 154
rect 9103 -154 9137 -138
rect 9199 138 9233 154
rect 9199 -154 9233 -138
rect 9295 138 9329 154
rect 9295 -154 9329 -138
rect 9391 138 9425 154
rect 9391 -154 9425 -138
rect 9487 138 9521 154
rect 9487 -154 9521 -138
rect 9583 138 9617 154
rect 9583 -154 9617 -138
rect 9679 138 9713 154
rect 9679 -154 9713 -138
rect 9775 138 9809 154
rect 9775 -154 9809 -138
rect 9871 138 9905 154
rect 9871 -154 9905 -138
rect 9967 138 10001 154
rect 9967 -154 10001 -138
rect 10063 138 10097 154
rect 10063 -154 10097 -138
rect 10159 138 10193 154
rect 10159 -154 10193 -138
rect 10255 138 10289 154
rect 10255 -154 10289 -138
rect 10351 138 10385 154
rect 10351 -154 10385 -138
rect 10447 138 10481 154
rect 10447 -154 10481 -138
rect 10543 138 10577 154
rect 10543 -154 10577 -138
rect 10639 138 10673 154
rect 10639 -154 10673 -138
rect 10735 138 10769 154
rect 10735 -154 10769 -138
rect 10831 138 10865 154
rect 10831 -154 10865 -138
rect 10927 138 10961 154
rect 10927 -154 10961 -138
rect 11023 138 11057 154
rect 11023 -154 11057 -138
rect 11119 138 11153 154
rect 11119 -154 11153 -138
rect 11215 138 11249 154
rect 11215 -154 11249 -138
rect 11311 138 11345 154
rect 11311 -154 11345 -138
rect 11407 138 11441 154
rect 11407 -154 11441 -138
rect 11503 138 11537 154
rect 11503 -154 11537 -138
rect 11599 138 11633 154
rect 11599 -154 11633 -138
rect 11695 138 11729 154
rect 11695 -154 11729 -138
rect 11791 138 11825 154
rect 11791 -154 11825 -138
rect 11887 138 11921 154
rect 11887 -154 11921 -138
rect 11983 138 12017 154
rect 11983 -154 12017 -138
rect 12079 138 12113 154
rect 12079 -154 12113 -138
rect 12175 138 12209 154
rect 12175 -154 12209 -138
rect 12271 138 12305 154
rect 12271 -154 12305 -138
rect 12367 138 12401 154
rect 12367 -154 12401 -138
rect 12463 138 12497 154
rect 12463 -154 12497 -138
rect 12559 138 12593 154
rect 12559 -154 12593 -138
rect 12655 138 12689 154
rect 12655 -154 12689 -138
rect 12751 138 12785 154
rect 12751 -154 12785 -138
rect 12847 138 12881 154
rect 12847 -154 12881 -138
rect 12943 138 12977 154
rect 12943 -154 12977 -138
rect 13039 138 13073 154
rect 13039 -154 13073 -138
rect 13135 138 13169 154
rect 13135 -154 13169 -138
rect 13231 138 13265 154
rect 13231 -154 13265 -138
rect 13327 138 13361 154
rect 13327 -154 13361 -138
rect 13423 138 13457 154
rect 13423 -154 13457 -138
rect 13519 138 13553 154
rect 13519 -154 13553 -138
rect 13615 138 13649 154
rect 13615 -154 13649 -138
rect 13711 138 13745 154
rect 13711 -154 13745 -138
rect 13807 138 13841 154
rect 13807 -154 13841 -138
rect 13903 138 13937 154
rect 13903 -154 13937 -138
rect 13999 138 14033 154
rect 13999 -154 14033 -138
rect 14095 138 14129 154
rect 14095 -154 14129 -138
rect 14191 138 14225 154
rect 14191 -154 14225 -138
rect 14287 138 14321 154
rect 14287 -154 14321 -138
rect 14383 138 14417 154
rect 14383 -154 14417 -138
rect 14479 138 14513 154
rect 14479 -154 14513 -138
rect 14575 138 14609 154
rect 14575 -154 14609 -138
rect 14671 138 14705 154
rect 14671 -154 14705 -138
rect 14767 138 14801 154
rect 14767 -154 14801 -138
rect 14863 138 14897 154
rect 14863 -154 14897 -138
rect 14959 138 14993 154
rect 14959 -154 14993 -138
rect 15055 138 15089 154
rect 15055 -154 15089 -138
rect 15151 138 15185 154
rect 15151 -154 15185 -138
rect 15247 138 15281 154
rect 15247 -154 15281 -138
rect 15343 138 15377 154
rect 15343 -154 15377 -138
rect 15439 138 15473 154
rect 15439 -154 15473 -138
rect 15535 138 15569 154
rect 15535 -154 15569 -138
rect 15631 138 15665 154
rect 15631 -154 15665 -138
rect 15727 138 15761 154
rect 15727 -154 15761 -138
rect 15823 138 15857 154
rect 15823 -154 15857 -138
rect 15919 138 15953 154
rect 15919 -154 15953 -138
rect 16015 138 16049 154
rect 16015 -154 16049 -138
rect 16111 138 16145 154
rect 16111 -154 16145 -138
rect 16207 138 16241 154
rect 16207 -154 16241 -138
rect 16303 138 16337 154
rect 16303 -154 16337 -138
rect 16399 138 16433 154
rect 16399 -154 16433 -138
rect 16495 138 16529 154
rect 16495 -154 16529 -138
rect 16591 138 16625 154
rect 16591 -154 16625 -138
rect 16687 138 16721 154
rect 16687 -154 16721 -138
rect 16783 138 16817 154
rect 16783 -154 16817 -138
rect 16879 138 16913 154
rect 16879 -154 16913 -138
rect 16975 138 17009 154
rect 16975 -154 17009 -138
rect 17071 138 17105 154
rect 17071 -154 17105 -138
rect 17167 138 17201 154
rect 17167 -154 17201 -138
rect 17263 138 17297 154
rect 17263 -154 17297 -138
rect 17359 138 17393 154
rect 17359 -154 17393 -138
rect 17455 138 17489 154
rect 17455 -154 17489 -138
rect 17551 138 17585 154
rect 17551 -154 17585 -138
rect 17647 138 17681 154
rect 17647 -154 17681 -138
rect 17743 138 17777 154
rect 17743 -154 17777 -138
rect 17839 138 17873 154
rect 17839 -154 17873 -138
rect 17935 138 17969 154
rect 17935 -154 17969 -138
rect 18031 138 18065 154
rect 18031 -154 18065 -138
rect 18127 138 18161 154
rect 18127 -154 18161 -138
rect 18223 138 18257 154
rect 18223 -154 18257 -138
rect 18319 138 18353 154
rect 18319 -154 18353 -138
rect 18415 138 18449 154
rect 18415 -154 18449 -138
rect 18511 138 18545 154
rect 18511 -154 18545 -138
rect 18607 138 18641 154
rect 18607 -154 18641 -138
rect 18703 138 18737 154
rect 18703 -154 18737 -138
rect 18799 138 18833 154
rect 18799 -154 18833 -138
rect 18895 138 18929 154
rect 18895 -154 18929 -138
rect 18991 138 19025 154
rect 18991 -154 19025 -138
rect 19087 138 19121 154
rect 19087 -154 19121 -138
rect 19183 138 19217 154
rect 19183 -154 19217 -138
rect -19185 -222 -19169 -188
rect -19135 -222 -19119 -188
rect -18993 -222 -18977 -188
rect -18943 -222 -18927 -188
rect -18801 -222 -18785 -188
rect -18751 -222 -18735 -188
rect -18609 -222 -18593 -188
rect -18559 -222 -18543 -188
rect -18417 -222 -18401 -188
rect -18367 -222 -18351 -188
rect -18225 -222 -18209 -188
rect -18175 -222 -18159 -188
rect -18033 -222 -18017 -188
rect -17983 -222 -17967 -188
rect -17841 -222 -17825 -188
rect -17791 -222 -17775 -188
rect -17649 -222 -17633 -188
rect -17599 -222 -17583 -188
rect -17457 -222 -17441 -188
rect -17407 -222 -17391 -188
rect -17265 -222 -17249 -188
rect -17215 -222 -17199 -188
rect -17073 -222 -17057 -188
rect -17023 -222 -17007 -188
rect -16881 -222 -16865 -188
rect -16831 -222 -16815 -188
rect -16689 -222 -16673 -188
rect -16639 -222 -16623 -188
rect -16497 -222 -16481 -188
rect -16447 -222 -16431 -188
rect -16305 -222 -16289 -188
rect -16255 -222 -16239 -188
rect -16113 -222 -16097 -188
rect -16063 -222 -16047 -188
rect -15921 -222 -15905 -188
rect -15871 -222 -15855 -188
rect -15729 -222 -15713 -188
rect -15679 -222 -15663 -188
rect -15537 -222 -15521 -188
rect -15487 -222 -15471 -188
rect -15345 -222 -15329 -188
rect -15295 -222 -15279 -188
rect -15153 -222 -15137 -188
rect -15103 -222 -15087 -188
rect -14961 -222 -14945 -188
rect -14911 -222 -14895 -188
rect -14769 -222 -14753 -188
rect -14719 -222 -14703 -188
rect -14577 -222 -14561 -188
rect -14527 -222 -14511 -188
rect -14385 -222 -14369 -188
rect -14335 -222 -14319 -188
rect -14193 -222 -14177 -188
rect -14143 -222 -14127 -188
rect -14001 -222 -13985 -188
rect -13951 -222 -13935 -188
rect -13809 -222 -13793 -188
rect -13759 -222 -13743 -188
rect -13617 -222 -13601 -188
rect -13567 -222 -13551 -188
rect -13425 -222 -13409 -188
rect -13375 -222 -13359 -188
rect -13233 -222 -13217 -188
rect -13183 -222 -13167 -188
rect -13041 -222 -13025 -188
rect -12991 -222 -12975 -188
rect -12849 -222 -12833 -188
rect -12799 -222 -12783 -188
rect -12657 -222 -12641 -188
rect -12607 -222 -12591 -188
rect -12465 -222 -12449 -188
rect -12415 -222 -12399 -188
rect -12273 -222 -12257 -188
rect -12223 -222 -12207 -188
rect -12081 -222 -12065 -188
rect -12031 -222 -12015 -188
rect -11889 -222 -11873 -188
rect -11839 -222 -11823 -188
rect -11697 -222 -11681 -188
rect -11647 -222 -11631 -188
rect -11505 -222 -11489 -188
rect -11455 -222 -11439 -188
rect -11313 -222 -11297 -188
rect -11263 -222 -11247 -188
rect -11121 -222 -11105 -188
rect -11071 -222 -11055 -188
rect -10929 -222 -10913 -188
rect -10879 -222 -10863 -188
rect -10737 -222 -10721 -188
rect -10687 -222 -10671 -188
rect -10545 -222 -10529 -188
rect -10495 -222 -10479 -188
rect -10353 -222 -10337 -188
rect -10303 -222 -10287 -188
rect -10161 -222 -10145 -188
rect -10111 -222 -10095 -188
rect -9969 -222 -9953 -188
rect -9919 -222 -9903 -188
rect -9777 -222 -9761 -188
rect -9727 -222 -9711 -188
rect -9585 -222 -9569 -188
rect -9535 -222 -9519 -188
rect -9393 -222 -9377 -188
rect -9343 -222 -9327 -188
rect -9201 -222 -9185 -188
rect -9151 -222 -9135 -188
rect -9009 -222 -8993 -188
rect -8959 -222 -8943 -188
rect -8817 -222 -8801 -188
rect -8767 -222 -8751 -188
rect -8625 -222 -8609 -188
rect -8575 -222 -8559 -188
rect -8433 -222 -8417 -188
rect -8383 -222 -8367 -188
rect -8241 -222 -8225 -188
rect -8191 -222 -8175 -188
rect -8049 -222 -8033 -188
rect -7999 -222 -7983 -188
rect -7857 -222 -7841 -188
rect -7807 -222 -7791 -188
rect -7665 -222 -7649 -188
rect -7615 -222 -7599 -188
rect -7473 -222 -7457 -188
rect -7423 -222 -7407 -188
rect -7281 -222 -7265 -188
rect -7231 -222 -7215 -188
rect -7089 -222 -7073 -188
rect -7039 -222 -7023 -188
rect -6897 -222 -6881 -188
rect -6847 -222 -6831 -188
rect -6705 -222 -6689 -188
rect -6655 -222 -6639 -188
rect -6513 -222 -6497 -188
rect -6463 -222 -6447 -188
rect -6321 -222 -6305 -188
rect -6271 -222 -6255 -188
rect -6129 -222 -6113 -188
rect -6079 -222 -6063 -188
rect -5937 -222 -5921 -188
rect -5887 -222 -5871 -188
rect -5745 -222 -5729 -188
rect -5695 -222 -5679 -188
rect -5553 -222 -5537 -188
rect -5503 -222 -5487 -188
rect -5361 -222 -5345 -188
rect -5311 -222 -5295 -188
rect -5169 -222 -5153 -188
rect -5119 -222 -5103 -188
rect -4977 -222 -4961 -188
rect -4927 -222 -4911 -188
rect -4785 -222 -4769 -188
rect -4735 -222 -4719 -188
rect -4593 -222 -4577 -188
rect -4543 -222 -4527 -188
rect -4401 -222 -4385 -188
rect -4351 -222 -4335 -188
rect -4209 -222 -4193 -188
rect -4159 -222 -4143 -188
rect -4017 -222 -4001 -188
rect -3967 -222 -3951 -188
rect -3825 -222 -3809 -188
rect -3775 -222 -3759 -188
rect -3633 -222 -3617 -188
rect -3583 -222 -3567 -188
rect -3441 -222 -3425 -188
rect -3391 -222 -3375 -188
rect -3249 -222 -3233 -188
rect -3199 -222 -3183 -188
rect -3057 -222 -3041 -188
rect -3007 -222 -2991 -188
rect -2865 -222 -2849 -188
rect -2815 -222 -2799 -188
rect -2673 -222 -2657 -188
rect -2623 -222 -2607 -188
rect -2481 -222 -2465 -188
rect -2431 -222 -2415 -188
rect -2289 -222 -2273 -188
rect -2239 -222 -2223 -188
rect -2097 -222 -2081 -188
rect -2047 -222 -2031 -188
rect -1905 -222 -1889 -188
rect -1855 -222 -1839 -188
rect -1713 -222 -1697 -188
rect -1663 -222 -1647 -188
rect -1521 -222 -1505 -188
rect -1471 -222 -1455 -188
rect -1329 -222 -1313 -188
rect -1279 -222 -1263 -188
rect -1137 -222 -1121 -188
rect -1087 -222 -1071 -188
rect -945 -222 -929 -188
rect -895 -222 -879 -188
rect -753 -222 -737 -188
rect -703 -222 -687 -188
rect -561 -222 -545 -188
rect -511 -222 -495 -188
rect -369 -222 -353 -188
rect -319 -222 -303 -188
rect -177 -222 -161 -188
rect -127 -222 -111 -188
rect 15 -222 31 -188
rect 65 -222 81 -188
rect 207 -222 223 -188
rect 257 -222 273 -188
rect 399 -222 415 -188
rect 449 -222 465 -188
rect 591 -222 607 -188
rect 641 -222 657 -188
rect 783 -222 799 -188
rect 833 -222 849 -188
rect 975 -222 991 -188
rect 1025 -222 1041 -188
rect 1167 -222 1183 -188
rect 1217 -222 1233 -188
rect 1359 -222 1375 -188
rect 1409 -222 1425 -188
rect 1551 -222 1567 -188
rect 1601 -222 1617 -188
rect 1743 -222 1759 -188
rect 1793 -222 1809 -188
rect 1935 -222 1951 -188
rect 1985 -222 2001 -188
rect 2127 -222 2143 -188
rect 2177 -222 2193 -188
rect 2319 -222 2335 -188
rect 2369 -222 2385 -188
rect 2511 -222 2527 -188
rect 2561 -222 2577 -188
rect 2703 -222 2719 -188
rect 2753 -222 2769 -188
rect 2895 -222 2911 -188
rect 2945 -222 2961 -188
rect 3087 -222 3103 -188
rect 3137 -222 3153 -188
rect 3279 -222 3295 -188
rect 3329 -222 3345 -188
rect 3471 -222 3487 -188
rect 3521 -222 3537 -188
rect 3663 -222 3679 -188
rect 3713 -222 3729 -188
rect 3855 -222 3871 -188
rect 3905 -222 3921 -188
rect 4047 -222 4063 -188
rect 4097 -222 4113 -188
rect 4239 -222 4255 -188
rect 4289 -222 4305 -188
rect 4431 -222 4447 -188
rect 4481 -222 4497 -188
rect 4623 -222 4639 -188
rect 4673 -222 4689 -188
rect 4815 -222 4831 -188
rect 4865 -222 4881 -188
rect 5007 -222 5023 -188
rect 5057 -222 5073 -188
rect 5199 -222 5215 -188
rect 5249 -222 5265 -188
rect 5391 -222 5407 -188
rect 5441 -222 5457 -188
rect 5583 -222 5599 -188
rect 5633 -222 5649 -188
rect 5775 -222 5791 -188
rect 5825 -222 5841 -188
rect 5967 -222 5983 -188
rect 6017 -222 6033 -188
rect 6159 -222 6175 -188
rect 6209 -222 6225 -188
rect 6351 -222 6367 -188
rect 6401 -222 6417 -188
rect 6543 -222 6559 -188
rect 6593 -222 6609 -188
rect 6735 -222 6751 -188
rect 6785 -222 6801 -188
rect 6927 -222 6943 -188
rect 6977 -222 6993 -188
rect 7119 -222 7135 -188
rect 7169 -222 7185 -188
rect 7311 -222 7327 -188
rect 7361 -222 7377 -188
rect 7503 -222 7519 -188
rect 7553 -222 7569 -188
rect 7695 -222 7711 -188
rect 7745 -222 7761 -188
rect 7887 -222 7903 -188
rect 7937 -222 7953 -188
rect 8079 -222 8095 -188
rect 8129 -222 8145 -188
rect 8271 -222 8287 -188
rect 8321 -222 8337 -188
rect 8463 -222 8479 -188
rect 8513 -222 8529 -188
rect 8655 -222 8671 -188
rect 8705 -222 8721 -188
rect 8847 -222 8863 -188
rect 8897 -222 8913 -188
rect 9039 -222 9055 -188
rect 9089 -222 9105 -188
rect 9231 -222 9247 -188
rect 9281 -222 9297 -188
rect 9423 -222 9439 -188
rect 9473 -222 9489 -188
rect 9615 -222 9631 -188
rect 9665 -222 9681 -188
rect 9807 -222 9823 -188
rect 9857 -222 9873 -188
rect 9999 -222 10015 -188
rect 10049 -222 10065 -188
rect 10191 -222 10207 -188
rect 10241 -222 10257 -188
rect 10383 -222 10399 -188
rect 10433 -222 10449 -188
rect 10575 -222 10591 -188
rect 10625 -222 10641 -188
rect 10767 -222 10783 -188
rect 10817 -222 10833 -188
rect 10959 -222 10975 -188
rect 11009 -222 11025 -188
rect 11151 -222 11167 -188
rect 11201 -222 11217 -188
rect 11343 -222 11359 -188
rect 11393 -222 11409 -188
rect 11535 -222 11551 -188
rect 11585 -222 11601 -188
rect 11727 -222 11743 -188
rect 11777 -222 11793 -188
rect 11919 -222 11935 -188
rect 11969 -222 11985 -188
rect 12111 -222 12127 -188
rect 12161 -222 12177 -188
rect 12303 -222 12319 -188
rect 12353 -222 12369 -188
rect 12495 -222 12511 -188
rect 12545 -222 12561 -188
rect 12687 -222 12703 -188
rect 12737 -222 12753 -188
rect 12879 -222 12895 -188
rect 12929 -222 12945 -188
rect 13071 -222 13087 -188
rect 13121 -222 13137 -188
rect 13263 -222 13279 -188
rect 13313 -222 13329 -188
rect 13455 -222 13471 -188
rect 13505 -222 13521 -188
rect 13647 -222 13663 -188
rect 13697 -222 13713 -188
rect 13839 -222 13855 -188
rect 13889 -222 13905 -188
rect 14031 -222 14047 -188
rect 14081 -222 14097 -188
rect 14223 -222 14239 -188
rect 14273 -222 14289 -188
rect 14415 -222 14431 -188
rect 14465 -222 14481 -188
rect 14607 -222 14623 -188
rect 14657 -222 14673 -188
rect 14799 -222 14815 -188
rect 14849 -222 14865 -188
rect 14991 -222 15007 -188
rect 15041 -222 15057 -188
rect 15183 -222 15199 -188
rect 15233 -222 15249 -188
rect 15375 -222 15391 -188
rect 15425 -222 15441 -188
rect 15567 -222 15583 -188
rect 15617 -222 15633 -188
rect 15759 -222 15775 -188
rect 15809 -222 15825 -188
rect 15951 -222 15967 -188
rect 16001 -222 16017 -188
rect 16143 -222 16159 -188
rect 16193 -222 16209 -188
rect 16335 -222 16351 -188
rect 16385 -222 16401 -188
rect 16527 -222 16543 -188
rect 16577 -222 16593 -188
rect 16719 -222 16735 -188
rect 16769 -222 16785 -188
rect 16911 -222 16927 -188
rect 16961 -222 16977 -188
rect 17103 -222 17119 -188
rect 17153 -222 17169 -188
rect 17295 -222 17311 -188
rect 17345 -222 17361 -188
rect 17487 -222 17503 -188
rect 17537 -222 17553 -188
rect 17679 -222 17695 -188
rect 17729 -222 17745 -188
rect 17871 -222 17887 -188
rect 17921 -222 17937 -188
rect 18063 -222 18079 -188
rect 18113 -222 18129 -188
rect 18255 -222 18271 -188
rect 18305 -222 18321 -188
rect 18447 -222 18463 -188
rect 18497 -222 18513 -188
rect 18639 -222 18655 -188
rect 18689 -222 18705 -188
rect 18831 -222 18847 -188
rect 18881 -222 18897 -188
rect 19023 -222 19039 -188
rect 19073 -222 19089 -188
rect -19331 -290 -19297 -228
rect 19297 -290 19331 -228
rect -19331 -324 -19235 -290
rect 19235 -324 19331 -290
<< viali >>
rect -19073 188 -19039 222
rect -18881 188 -18847 222
rect -18689 188 -18655 222
rect -18497 188 -18463 222
rect -18305 188 -18271 222
rect -18113 188 -18079 222
rect -17921 188 -17887 222
rect -17729 188 -17695 222
rect -17537 188 -17503 222
rect -17345 188 -17311 222
rect -17153 188 -17119 222
rect -16961 188 -16927 222
rect -16769 188 -16735 222
rect -16577 188 -16543 222
rect -16385 188 -16351 222
rect -16193 188 -16159 222
rect -16001 188 -15967 222
rect -15809 188 -15775 222
rect -15617 188 -15583 222
rect -15425 188 -15391 222
rect -15233 188 -15199 222
rect -15041 188 -15007 222
rect -14849 188 -14815 222
rect -14657 188 -14623 222
rect -14465 188 -14431 222
rect -14273 188 -14239 222
rect -14081 188 -14047 222
rect -13889 188 -13855 222
rect -13697 188 -13663 222
rect -13505 188 -13471 222
rect -13313 188 -13279 222
rect -13121 188 -13087 222
rect -12929 188 -12895 222
rect -12737 188 -12703 222
rect -12545 188 -12511 222
rect -12353 188 -12319 222
rect -12161 188 -12127 222
rect -11969 188 -11935 222
rect -11777 188 -11743 222
rect -11585 188 -11551 222
rect -11393 188 -11359 222
rect -11201 188 -11167 222
rect -11009 188 -10975 222
rect -10817 188 -10783 222
rect -10625 188 -10591 222
rect -10433 188 -10399 222
rect -10241 188 -10207 222
rect -10049 188 -10015 222
rect -9857 188 -9823 222
rect -9665 188 -9631 222
rect -9473 188 -9439 222
rect -9281 188 -9247 222
rect -9089 188 -9055 222
rect -8897 188 -8863 222
rect -8705 188 -8671 222
rect -8513 188 -8479 222
rect -8321 188 -8287 222
rect -8129 188 -8095 222
rect -7937 188 -7903 222
rect -7745 188 -7711 222
rect -7553 188 -7519 222
rect -7361 188 -7327 222
rect -7169 188 -7135 222
rect -6977 188 -6943 222
rect -6785 188 -6751 222
rect -6593 188 -6559 222
rect -6401 188 -6367 222
rect -6209 188 -6175 222
rect -6017 188 -5983 222
rect -5825 188 -5791 222
rect -5633 188 -5599 222
rect -5441 188 -5407 222
rect -5249 188 -5215 222
rect -5057 188 -5023 222
rect -4865 188 -4831 222
rect -4673 188 -4639 222
rect -4481 188 -4447 222
rect -4289 188 -4255 222
rect -4097 188 -4063 222
rect -3905 188 -3871 222
rect -3713 188 -3679 222
rect -3521 188 -3487 222
rect -3329 188 -3295 222
rect -3137 188 -3103 222
rect -2945 188 -2911 222
rect -2753 188 -2719 222
rect -2561 188 -2527 222
rect -2369 188 -2335 222
rect -2177 188 -2143 222
rect -1985 188 -1951 222
rect -1793 188 -1759 222
rect -1601 188 -1567 222
rect -1409 188 -1375 222
rect -1217 188 -1183 222
rect -1025 188 -991 222
rect -833 188 -799 222
rect -641 188 -607 222
rect -449 188 -415 222
rect -257 188 -223 222
rect -65 188 -31 222
rect 127 188 161 222
rect 319 188 353 222
rect 511 188 545 222
rect 703 188 737 222
rect 895 188 929 222
rect 1087 188 1121 222
rect 1279 188 1313 222
rect 1471 188 1505 222
rect 1663 188 1697 222
rect 1855 188 1889 222
rect 2047 188 2081 222
rect 2239 188 2273 222
rect 2431 188 2465 222
rect 2623 188 2657 222
rect 2815 188 2849 222
rect 3007 188 3041 222
rect 3199 188 3233 222
rect 3391 188 3425 222
rect 3583 188 3617 222
rect 3775 188 3809 222
rect 3967 188 4001 222
rect 4159 188 4193 222
rect 4351 188 4385 222
rect 4543 188 4577 222
rect 4735 188 4769 222
rect 4927 188 4961 222
rect 5119 188 5153 222
rect 5311 188 5345 222
rect 5503 188 5537 222
rect 5695 188 5729 222
rect 5887 188 5921 222
rect 6079 188 6113 222
rect 6271 188 6305 222
rect 6463 188 6497 222
rect 6655 188 6689 222
rect 6847 188 6881 222
rect 7039 188 7073 222
rect 7231 188 7265 222
rect 7423 188 7457 222
rect 7615 188 7649 222
rect 7807 188 7841 222
rect 7999 188 8033 222
rect 8191 188 8225 222
rect 8383 188 8417 222
rect 8575 188 8609 222
rect 8767 188 8801 222
rect 8959 188 8993 222
rect 9151 188 9185 222
rect 9343 188 9377 222
rect 9535 188 9569 222
rect 9727 188 9761 222
rect 9919 188 9953 222
rect 10111 188 10145 222
rect 10303 188 10337 222
rect 10495 188 10529 222
rect 10687 188 10721 222
rect 10879 188 10913 222
rect 11071 188 11105 222
rect 11263 188 11297 222
rect 11455 188 11489 222
rect 11647 188 11681 222
rect 11839 188 11873 222
rect 12031 188 12065 222
rect 12223 188 12257 222
rect 12415 188 12449 222
rect 12607 188 12641 222
rect 12799 188 12833 222
rect 12991 188 13025 222
rect 13183 188 13217 222
rect 13375 188 13409 222
rect 13567 188 13601 222
rect 13759 188 13793 222
rect 13951 188 13985 222
rect 14143 188 14177 222
rect 14335 188 14369 222
rect 14527 188 14561 222
rect 14719 188 14753 222
rect 14911 188 14945 222
rect 15103 188 15137 222
rect 15295 188 15329 222
rect 15487 188 15521 222
rect 15679 188 15713 222
rect 15871 188 15905 222
rect 16063 188 16097 222
rect 16255 188 16289 222
rect 16447 188 16481 222
rect 16639 188 16673 222
rect 16831 188 16865 222
rect 17023 188 17057 222
rect 17215 188 17249 222
rect 17407 188 17441 222
rect 17599 188 17633 222
rect 17791 188 17825 222
rect 17983 188 18017 222
rect 18175 188 18209 222
rect 18367 188 18401 222
rect 18559 188 18593 222
rect 18751 188 18785 222
rect 18943 188 18977 222
rect 19135 188 19169 222
rect -19217 -138 -19183 138
rect -19121 -138 -19087 138
rect -19025 -138 -18991 138
rect -18929 -138 -18895 138
rect -18833 -138 -18799 138
rect -18737 -138 -18703 138
rect -18641 -138 -18607 138
rect -18545 -138 -18511 138
rect -18449 -138 -18415 138
rect -18353 -138 -18319 138
rect -18257 -138 -18223 138
rect -18161 -138 -18127 138
rect -18065 -138 -18031 138
rect -17969 -138 -17935 138
rect -17873 -138 -17839 138
rect -17777 -138 -17743 138
rect -17681 -138 -17647 138
rect -17585 -138 -17551 138
rect -17489 -138 -17455 138
rect -17393 -138 -17359 138
rect -17297 -138 -17263 138
rect -17201 -138 -17167 138
rect -17105 -138 -17071 138
rect -17009 -138 -16975 138
rect -16913 -138 -16879 138
rect -16817 -138 -16783 138
rect -16721 -138 -16687 138
rect -16625 -138 -16591 138
rect -16529 -138 -16495 138
rect -16433 -138 -16399 138
rect -16337 -138 -16303 138
rect -16241 -138 -16207 138
rect -16145 -138 -16111 138
rect -16049 -138 -16015 138
rect -15953 -138 -15919 138
rect -15857 -138 -15823 138
rect -15761 -138 -15727 138
rect -15665 -138 -15631 138
rect -15569 -138 -15535 138
rect -15473 -138 -15439 138
rect -15377 -138 -15343 138
rect -15281 -138 -15247 138
rect -15185 -138 -15151 138
rect -15089 -138 -15055 138
rect -14993 -138 -14959 138
rect -14897 -138 -14863 138
rect -14801 -138 -14767 138
rect -14705 -138 -14671 138
rect -14609 -138 -14575 138
rect -14513 -138 -14479 138
rect -14417 -138 -14383 138
rect -14321 -138 -14287 138
rect -14225 -138 -14191 138
rect -14129 -138 -14095 138
rect -14033 -138 -13999 138
rect -13937 -138 -13903 138
rect -13841 -138 -13807 138
rect -13745 -138 -13711 138
rect -13649 -138 -13615 138
rect -13553 -138 -13519 138
rect -13457 -138 -13423 138
rect -13361 -138 -13327 138
rect -13265 -138 -13231 138
rect -13169 -138 -13135 138
rect -13073 -138 -13039 138
rect -12977 -138 -12943 138
rect -12881 -138 -12847 138
rect -12785 -138 -12751 138
rect -12689 -138 -12655 138
rect -12593 -138 -12559 138
rect -12497 -138 -12463 138
rect -12401 -138 -12367 138
rect -12305 -138 -12271 138
rect -12209 -138 -12175 138
rect -12113 -138 -12079 138
rect -12017 -138 -11983 138
rect -11921 -138 -11887 138
rect -11825 -138 -11791 138
rect -11729 -138 -11695 138
rect -11633 -138 -11599 138
rect -11537 -138 -11503 138
rect -11441 -138 -11407 138
rect -11345 -138 -11311 138
rect -11249 -138 -11215 138
rect -11153 -138 -11119 138
rect -11057 -138 -11023 138
rect -10961 -138 -10927 138
rect -10865 -138 -10831 138
rect -10769 -138 -10735 138
rect -10673 -138 -10639 138
rect -10577 -138 -10543 138
rect -10481 -138 -10447 138
rect -10385 -138 -10351 138
rect -10289 -138 -10255 138
rect -10193 -138 -10159 138
rect -10097 -138 -10063 138
rect -10001 -138 -9967 138
rect -9905 -138 -9871 138
rect -9809 -138 -9775 138
rect -9713 -138 -9679 138
rect -9617 -138 -9583 138
rect -9521 -138 -9487 138
rect -9425 -138 -9391 138
rect -9329 -138 -9295 138
rect -9233 -138 -9199 138
rect -9137 -138 -9103 138
rect -9041 -138 -9007 138
rect -8945 -138 -8911 138
rect -8849 -138 -8815 138
rect -8753 -138 -8719 138
rect -8657 -138 -8623 138
rect -8561 -138 -8527 138
rect -8465 -138 -8431 138
rect -8369 -138 -8335 138
rect -8273 -138 -8239 138
rect -8177 -138 -8143 138
rect -8081 -138 -8047 138
rect -7985 -138 -7951 138
rect -7889 -138 -7855 138
rect -7793 -138 -7759 138
rect -7697 -138 -7663 138
rect -7601 -138 -7567 138
rect -7505 -138 -7471 138
rect -7409 -138 -7375 138
rect -7313 -138 -7279 138
rect -7217 -138 -7183 138
rect -7121 -138 -7087 138
rect -7025 -138 -6991 138
rect -6929 -138 -6895 138
rect -6833 -138 -6799 138
rect -6737 -138 -6703 138
rect -6641 -138 -6607 138
rect -6545 -138 -6511 138
rect -6449 -138 -6415 138
rect -6353 -138 -6319 138
rect -6257 -138 -6223 138
rect -6161 -138 -6127 138
rect -6065 -138 -6031 138
rect -5969 -138 -5935 138
rect -5873 -138 -5839 138
rect -5777 -138 -5743 138
rect -5681 -138 -5647 138
rect -5585 -138 -5551 138
rect -5489 -138 -5455 138
rect -5393 -138 -5359 138
rect -5297 -138 -5263 138
rect -5201 -138 -5167 138
rect -5105 -138 -5071 138
rect -5009 -138 -4975 138
rect -4913 -138 -4879 138
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
rect 4879 -138 4913 138
rect 4975 -138 5009 138
rect 5071 -138 5105 138
rect 5167 -138 5201 138
rect 5263 -138 5297 138
rect 5359 -138 5393 138
rect 5455 -138 5489 138
rect 5551 -138 5585 138
rect 5647 -138 5681 138
rect 5743 -138 5777 138
rect 5839 -138 5873 138
rect 5935 -138 5969 138
rect 6031 -138 6065 138
rect 6127 -138 6161 138
rect 6223 -138 6257 138
rect 6319 -138 6353 138
rect 6415 -138 6449 138
rect 6511 -138 6545 138
rect 6607 -138 6641 138
rect 6703 -138 6737 138
rect 6799 -138 6833 138
rect 6895 -138 6929 138
rect 6991 -138 7025 138
rect 7087 -138 7121 138
rect 7183 -138 7217 138
rect 7279 -138 7313 138
rect 7375 -138 7409 138
rect 7471 -138 7505 138
rect 7567 -138 7601 138
rect 7663 -138 7697 138
rect 7759 -138 7793 138
rect 7855 -138 7889 138
rect 7951 -138 7985 138
rect 8047 -138 8081 138
rect 8143 -138 8177 138
rect 8239 -138 8273 138
rect 8335 -138 8369 138
rect 8431 -138 8465 138
rect 8527 -138 8561 138
rect 8623 -138 8657 138
rect 8719 -138 8753 138
rect 8815 -138 8849 138
rect 8911 -138 8945 138
rect 9007 -138 9041 138
rect 9103 -138 9137 138
rect 9199 -138 9233 138
rect 9295 -138 9329 138
rect 9391 -138 9425 138
rect 9487 -138 9521 138
rect 9583 -138 9617 138
rect 9679 -138 9713 138
rect 9775 -138 9809 138
rect 9871 -138 9905 138
rect 9967 -138 10001 138
rect 10063 -138 10097 138
rect 10159 -138 10193 138
rect 10255 -138 10289 138
rect 10351 -138 10385 138
rect 10447 -138 10481 138
rect 10543 -138 10577 138
rect 10639 -138 10673 138
rect 10735 -138 10769 138
rect 10831 -138 10865 138
rect 10927 -138 10961 138
rect 11023 -138 11057 138
rect 11119 -138 11153 138
rect 11215 -138 11249 138
rect 11311 -138 11345 138
rect 11407 -138 11441 138
rect 11503 -138 11537 138
rect 11599 -138 11633 138
rect 11695 -138 11729 138
rect 11791 -138 11825 138
rect 11887 -138 11921 138
rect 11983 -138 12017 138
rect 12079 -138 12113 138
rect 12175 -138 12209 138
rect 12271 -138 12305 138
rect 12367 -138 12401 138
rect 12463 -138 12497 138
rect 12559 -138 12593 138
rect 12655 -138 12689 138
rect 12751 -138 12785 138
rect 12847 -138 12881 138
rect 12943 -138 12977 138
rect 13039 -138 13073 138
rect 13135 -138 13169 138
rect 13231 -138 13265 138
rect 13327 -138 13361 138
rect 13423 -138 13457 138
rect 13519 -138 13553 138
rect 13615 -138 13649 138
rect 13711 -138 13745 138
rect 13807 -138 13841 138
rect 13903 -138 13937 138
rect 13999 -138 14033 138
rect 14095 -138 14129 138
rect 14191 -138 14225 138
rect 14287 -138 14321 138
rect 14383 -138 14417 138
rect 14479 -138 14513 138
rect 14575 -138 14609 138
rect 14671 -138 14705 138
rect 14767 -138 14801 138
rect 14863 -138 14897 138
rect 14959 -138 14993 138
rect 15055 -138 15089 138
rect 15151 -138 15185 138
rect 15247 -138 15281 138
rect 15343 -138 15377 138
rect 15439 -138 15473 138
rect 15535 -138 15569 138
rect 15631 -138 15665 138
rect 15727 -138 15761 138
rect 15823 -138 15857 138
rect 15919 -138 15953 138
rect 16015 -138 16049 138
rect 16111 -138 16145 138
rect 16207 -138 16241 138
rect 16303 -138 16337 138
rect 16399 -138 16433 138
rect 16495 -138 16529 138
rect 16591 -138 16625 138
rect 16687 -138 16721 138
rect 16783 -138 16817 138
rect 16879 -138 16913 138
rect 16975 -138 17009 138
rect 17071 -138 17105 138
rect 17167 -138 17201 138
rect 17263 -138 17297 138
rect 17359 -138 17393 138
rect 17455 -138 17489 138
rect 17551 -138 17585 138
rect 17647 -138 17681 138
rect 17743 -138 17777 138
rect 17839 -138 17873 138
rect 17935 -138 17969 138
rect 18031 -138 18065 138
rect 18127 -138 18161 138
rect 18223 -138 18257 138
rect 18319 -138 18353 138
rect 18415 -138 18449 138
rect 18511 -138 18545 138
rect 18607 -138 18641 138
rect 18703 -138 18737 138
rect 18799 -138 18833 138
rect 18895 -138 18929 138
rect 18991 -138 19025 138
rect 19087 -138 19121 138
rect 19183 -138 19217 138
rect -19169 -222 -19135 -188
rect -18977 -222 -18943 -188
rect -18785 -222 -18751 -188
rect -18593 -222 -18559 -188
rect -18401 -222 -18367 -188
rect -18209 -222 -18175 -188
rect -18017 -222 -17983 -188
rect -17825 -222 -17791 -188
rect -17633 -222 -17599 -188
rect -17441 -222 -17407 -188
rect -17249 -222 -17215 -188
rect -17057 -222 -17023 -188
rect -16865 -222 -16831 -188
rect -16673 -222 -16639 -188
rect -16481 -222 -16447 -188
rect -16289 -222 -16255 -188
rect -16097 -222 -16063 -188
rect -15905 -222 -15871 -188
rect -15713 -222 -15679 -188
rect -15521 -222 -15487 -188
rect -15329 -222 -15295 -188
rect -15137 -222 -15103 -188
rect -14945 -222 -14911 -188
rect -14753 -222 -14719 -188
rect -14561 -222 -14527 -188
rect -14369 -222 -14335 -188
rect -14177 -222 -14143 -188
rect -13985 -222 -13951 -188
rect -13793 -222 -13759 -188
rect -13601 -222 -13567 -188
rect -13409 -222 -13375 -188
rect -13217 -222 -13183 -188
rect -13025 -222 -12991 -188
rect -12833 -222 -12799 -188
rect -12641 -222 -12607 -188
rect -12449 -222 -12415 -188
rect -12257 -222 -12223 -188
rect -12065 -222 -12031 -188
rect -11873 -222 -11839 -188
rect -11681 -222 -11647 -188
rect -11489 -222 -11455 -188
rect -11297 -222 -11263 -188
rect -11105 -222 -11071 -188
rect -10913 -222 -10879 -188
rect -10721 -222 -10687 -188
rect -10529 -222 -10495 -188
rect -10337 -222 -10303 -188
rect -10145 -222 -10111 -188
rect -9953 -222 -9919 -188
rect -9761 -222 -9727 -188
rect -9569 -222 -9535 -188
rect -9377 -222 -9343 -188
rect -9185 -222 -9151 -188
rect -8993 -222 -8959 -188
rect -8801 -222 -8767 -188
rect -8609 -222 -8575 -188
rect -8417 -222 -8383 -188
rect -8225 -222 -8191 -188
rect -8033 -222 -7999 -188
rect -7841 -222 -7807 -188
rect -7649 -222 -7615 -188
rect -7457 -222 -7423 -188
rect -7265 -222 -7231 -188
rect -7073 -222 -7039 -188
rect -6881 -222 -6847 -188
rect -6689 -222 -6655 -188
rect -6497 -222 -6463 -188
rect -6305 -222 -6271 -188
rect -6113 -222 -6079 -188
rect -5921 -222 -5887 -188
rect -5729 -222 -5695 -188
rect -5537 -222 -5503 -188
rect -5345 -222 -5311 -188
rect -5153 -222 -5119 -188
rect -4961 -222 -4927 -188
rect -4769 -222 -4735 -188
rect -4577 -222 -4543 -188
rect -4385 -222 -4351 -188
rect -4193 -222 -4159 -188
rect -4001 -222 -3967 -188
rect -3809 -222 -3775 -188
rect -3617 -222 -3583 -188
rect -3425 -222 -3391 -188
rect -3233 -222 -3199 -188
rect -3041 -222 -3007 -188
rect -2849 -222 -2815 -188
rect -2657 -222 -2623 -188
rect -2465 -222 -2431 -188
rect -2273 -222 -2239 -188
rect -2081 -222 -2047 -188
rect -1889 -222 -1855 -188
rect -1697 -222 -1663 -188
rect -1505 -222 -1471 -188
rect -1313 -222 -1279 -188
rect -1121 -222 -1087 -188
rect -929 -222 -895 -188
rect -737 -222 -703 -188
rect -545 -222 -511 -188
rect -353 -222 -319 -188
rect -161 -222 -127 -188
rect 31 -222 65 -188
rect 223 -222 257 -188
rect 415 -222 449 -188
rect 607 -222 641 -188
rect 799 -222 833 -188
rect 991 -222 1025 -188
rect 1183 -222 1217 -188
rect 1375 -222 1409 -188
rect 1567 -222 1601 -188
rect 1759 -222 1793 -188
rect 1951 -222 1985 -188
rect 2143 -222 2177 -188
rect 2335 -222 2369 -188
rect 2527 -222 2561 -188
rect 2719 -222 2753 -188
rect 2911 -222 2945 -188
rect 3103 -222 3137 -188
rect 3295 -222 3329 -188
rect 3487 -222 3521 -188
rect 3679 -222 3713 -188
rect 3871 -222 3905 -188
rect 4063 -222 4097 -188
rect 4255 -222 4289 -188
rect 4447 -222 4481 -188
rect 4639 -222 4673 -188
rect 4831 -222 4865 -188
rect 5023 -222 5057 -188
rect 5215 -222 5249 -188
rect 5407 -222 5441 -188
rect 5599 -222 5633 -188
rect 5791 -222 5825 -188
rect 5983 -222 6017 -188
rect 6175 -222 6209 -188
rect 6367 -222 6401 -188
rect 6559 -222 6593 -188
rect 6751 -222 6785 -188
rect 6943 -222 6977 -188
rect 7135 -222 7169 -188
rect 7327 -222 7361 -188
rect 7519 -222 7553 -188
rect 7711 -222 7745 -188
rect 7903 -222 7937 -188
rect 8095 -222 8129 -188
rect 8287 -222 8321 -188
rect 8479 -222 8513 -188
rect 8671 -222 8705 -188
rect 8863 -222 8897 -188
rect 9055 -222 9089 -188
rect 9247 -222 9281 -188
rect 9439 -222 9473 -188
rect 9631 -222 9665 -188
rect 9823 -222 9857 -188
rect 10015 -222 10049 -188
rect 10207 -222 10241 -188
rect 10399 -222 10433 -188
rect 10591 -222 10625 -188
rect 10783 -222 10817 -188
rect 10975 -222 11009 -188
rect 11167 -222 11201 -188
rect 11359 -222 11393 -188
rect 11551 -222 11585 -188
rect 11743 -222 11777 -188
rect 11935 -222 11969 -188
rect 12127 -222 12161 -188
rect 12319 -222 12353 -188
rect 12511 -222 12545 -188
rect 12703 -222 12737 -188
rect 12895 -222 12929 -188
rect 13087 -222 13121 -188
rect 13279 -222 13313 -188
rect 13471 -222 13505 -188
rect 13663 -222 13697 -188
rect 13855 -222 13889 -188
rect 14047 -222 14081 -188
rect 14239 -222 14273 -188
rect 14431 -222 14465 -188
rect 14623 -222 14657 -188
rect 14815 -222 14849 -188
rect 15007 -222 15041 -188
rect 15199 -222 15233 -188
rect 15391 -222 15425 -188
rect 15583 -222 15617 -188
rect 15775 -222 15809 -188
rect 15967 -222 16001 -188
rect 16159 -222 16193 -188
rect 16351 -222 16385 -188
rect 16543 -222 16577 -188
rect 16735 -222 16769 -188
rect 16927 -222 16961 -188
rect 17119 -222 17153 -188
rect 17311 -222 17345 -188
rect 17503 -222 17537 -188
rect 17695 -222 17729 -188
rect 17887 -222 17921 -188
rect 18079 -222 18113 -188
rect 18271 -222 18305 -188
rect 18463 -222 18497 -188
rect 18655 -222 18689 -188
rect 18847 -222 18881 -188
rect 19039 -222 19073 -188
<< metal1 >>
rect -19085 222 -19027 228
rect -19085 188 -19073 222
rect -19039 188 -19027 222
rect -19085 182 -19027 188
rect -18893 222 -18835 228
rect -18893 188 -18881 222
rect -18847 188 -18835 222
rect -18893 182 -18835 188
rect -18701 222 -18643 228
rect -18701 188 -18689 222
rect -18655 188 -18643 222
rect -18701 182 -18643 188
rect -18509 222 -18451 228
rect -18509 188 -18497 222
rect -18463 188 -18451 222
rect -18509 182 -18451 188
rect -18317 222 -18259 228
rect -18317 188 -18305 222
rect -18271 188 -18259 222
rect -18317 182 -18259 188
rect -18125 222 -18067 228
rect -18125 188 -18113 222
rect -18079 188 -18067 222
rect -18125 182 -18067 188
rect -17933 222 -17875 228
rect -17933 188 -17921 222
rect -17887 188 -17875 222
rect -17933 182 -17875 188
rect -17741 222 -17683 228
rect -17741 188 -17729 222
rect -17695 188 -17683 222
rect -17741 182 -17683 188
rect -17549 222 -17491 228
rect -17549 188 -17537 222
rect -17503 188 -17491 222
rect -17549 182 -17491 188
rect -17357 222 -17299 228
rect -17357 188 -17345 222
rect -17311 188 -17299 222
rect -17357 182 -17299 188
rect -17165 222 -17107 228
rect -17165 188 -17153 222
rect -17119 188 -17107 222
rect -17165 182 -17107 188
rect -16973 222 -16915 228
rect -16973 188 -16961 222
rect -16927 188 -16915 222
rect -16973 182 -16915 188
rect -16781 222 -16723 228
rect -16781 188 -16769 222
rect -16735 188 -16723 222
rect -16781 182 -16723 188
rect -16589 222 -16531 228
rect -16589 188 -16577 222
rect -16543 188 -16531 222
rect -16589 182 -16531 188
rect -16397 222 -16339 228
rect -16397 188 -16385 222
rect -16351 188 -16339 222
rect -16397 182 -16339 188
rect -16205 222 -16147 228
rect -16205 188 -16193 222
rect -16159 188 -16147 222
rect -16205 182 -16147 188
rect -16013 222 -15955 228
rect -16013 188 -16001 222
rect -15967 188 -15955 222
rect -16013 182 -15955 188
rect -15821 222 -15763 228
rect -15821 188 -15809 222
rect -15775 188 -15763 222
rect -15821 182 -15763 188
rect -15629 222 -15571 228
rect -15629 188 -15617 222
rect -15583 188 -15571 222
rect -15629 182 -15571 188
rect -15437 222 -15379 228
rect -15437 188 -15425 222
rect -15391 188 -15379 222
rect -15437 182 -15379 188
rect -15245 222 -15187 228
rect -15245 188 -15233 222
rect -15199 188 -15187 222
rect -15245 182 -15187 188
rect -15053 222 -14995 228
rect -15053 188 -15041 222
rect -15007 188 -14995 222
rect -15053 182 -14995 188
rect -14861 222 -14803 228
rect -14861 188 -14849 222
rect -14815 188 -14803 222
rect -14861 182 -14803 188
rect -14669 222 -14611 228
rect -14669 188 -14657 222
rect -14623 188 -14611 222
rect -14669 182 -14611 188
rect -14477 222 -14419 228
rect -14477 188 -14465 222
rect -14431 188 -14419 222
rect -14477 182 -14419 188
rect -14285 222 -14227 228
rect -14285 188 -14273 222
rect -14239 188 -14227 222
rect -14285 182 -14227 188
rect -14093 222 -14035 228
rect -14093 188 -14081 222
rect -14047 188 -14035 222
rect -14093 182 -14035 188
rect -13901 222 -13843 228
rect -13901 188 -13889 222
rect -13855 188 -13843 222
rect -13901 182 -13843 188
rect -13709 222 -13651 228
rect -13709 188 -13697 222
rect -13663 188 -13651 222
rect -13709 182 -13651 188
rect -13517 222 -13459 228
rect -13517 188 -13505 222
rect -13471 188 -13459 222
rect -13517 182 -13459 188
rect -13325 222 -13267 228
rect -13325 188 -13313 222
rect -13279 188 -13267 222
rect -13325 182 -13267 188
rect -13133 222 -13075 228
rect -13133 188 -13121 222
rect -13087 188 -13075 222
rect -13133 182 -13075 188
rect -12941 222 -12883 228
rect -12941 188 -12929 222
rect -12895 188 -12883 222
rect -12941 182 -12883 188
rect -12749 222 -12691 228
rect -12749 188 -12737 222
rect -12703 188 -12691 222
rect -12749 182 -12691 188
rect -12557 222 -12499 228
rect -12557 188 -12545 222
rect -12511 188 -12499 222
rect -12557 182 -12499 188
rect -12365 222 -12307 228
rect -12365 188 -12353 222
rect -12319 188 -12307 222
rect -12365 182 -12307 188
rect -12173 222 -12115 228
rect -12173 188 -12161 222
rect -12127 188 -12115 222
rect -12173 182 -12115 188
rect -11981 222 -11923 228
rect -11981 188 -11969 222
rect -11935 188 -11923 222
rect -11981 182 -11923 188
rect -11789 222 -11731 228
rect -11789 188 -11777 222
rect -11743 188 -11731 222
rect -11789 182 -11731 188
rect -11597 222 -11539 228
rect -11597 188 -11585 222
rect -11551 188 -11539 222
rect -11597 182 -11539 188
rect -11405 222 -11347 228
rect -11405 188 -11393 222
rect -11359 188 -11347 222
rect -11405 182 -11347 188
rect -11213 222 -11155 228
rect -11213 188 -11201 222
rect -11167 188 -11155 222
rect -11213 182 -11155 188
rect -11021 222 -10963 228
rect -11021 188 -11009 222
rect -10975 188 -10963 222
rect -11021 182 -10963 188
rect -10829 222 -10771 228
rect -10829 188 -10817 222
rect -10783 188 -10771 222
rect -10829 182 -10771 188
rect -10637 222 -10579 228
rect -10637 188 -10625 222
rect -10591 188 -10579 222
rect -10637 182 -10579 188
rect -10445 222 -10387 228
rect -10445 188 -10433 222
rect -10399 188 -10387 222
rect -10445 182 -10387 188
rect -10253 222 -10195 228
rect -10253 188 -10241 222
rect -10207 188 -10195 222
rect -10253 182 -10195 188
rect -10061 222 -10003 228
rect -10061 188 -10049 222
rect -10015 188 -10003 222
rect -10061 182 -10003 188
rect -9869 222 -9811 228
rect -9869 188 -9857 222
rect -9823 188 -9811 222
rect -9869 182 -9811 188
rect -9677 222 -9619 228
rect -9677 188 -9665 222
rect -9631 188 -9619 222
rect -9677 182 -9619 188
rect -9485 222 -9427 228
rect -9485 188 -9473 222
rect -9439 188 -9427 222
rect -9485 182 -9427 188
rect -9293 222 -9235 228
rect -9293 188 -9281 222
rect -9247 188 -9235 222
rect -9293 182 -9235 188
rect -9101 222 -9043 228
rect -9101 188 -9089 222
rect -9055 188 -9043 222
rect -9101 182 -9043 188
rect -8909 222 -8851 228
rect -8909 188 -8897 222
rect -8863 188 -8851 222
rect -8909 182 -8851 188
rect -8717 222 -8659 228
rect -8717 188 -8705 222
rect -8671 188 -8659 222
rect -8717 182 -8659 188
rect -8525 222 -8467 228
rect -8525 188 -8513 222
rect -8479 188 -8467 222
rect -8525 182 -8467 188
rect -8333 222 -8275 228
rect -8333 188 -8321 222
rect -8287 188 -8275 222
rect -8333 182 -8275 188
rect -8141 222 -8083 228
rect -8141 188 -8129 222
rect -8095 188 -8083 222
rect -8141 182 -8083 188
rect -7949 222 -7891 228
rect -7949 188 -7937 222
rect -7903 188 -7891 222
rect -7949 182 -7891 188
rect -7757 222 -7699 228
rect -7757 188 -7745 222
rect -7711 188 -7699 222
rect -7757 182 -7699 188
rect -7565 222 -7507 228
rect -7565 188 -7553 222
rect -7519 188 -7507 222
rect -7565 182 -7507 188
rect -7373 222 -7315 228
rect -7373 188 -7361 222
rect -7327 188 -7315 222
rect -7373 182 -7315 188
rect -7181 222 -7123 228
rect -7181 188 -7169 222
rect -7135 188 -7123 222
rect -7181 182 -7123 188
rect -6989 222 -6931 228
rect -6989 188 -6977 222
rect -6943 188 -6931 222
rect -6989 182 -6931 188
rect -6797 222 -6739 228
rect -6797 188 -6785 222
rect -6751 188 -6739 222
rect -6797 182 -6739 188
rect -6605 222 -6547 228
rect -6605 188 -6593 222
rect -6559 188 -6547 222
rect -6605 182 -6547 188
rect -6413 222 -6355 228
rect -6413 188 -6401 222
rect -6367 188 -6355 222
rect -6413 182 -6355 188
rect -6221 222 -6163 228
rect -6221 188 -6209 222
rect -6175 188 -6163 222
rect -6221 182 -6163 188
rect -6029 222 -5971 228
rect -6029 188 -6017 222
rect -5983 188 -5971 222
rect -6029 182 -5971 188
rect -5837 222 -5779 228
rect -5837 188 -5825 222
rect -5791 188 -5779 222
rect -5837 182 -5779 188
rect -5645 222 -5587 228
rect -5645 188 -5633 222
rect -5599 188 -5587 222
rect -5645 182 -5587 188
rect -5453 222 -5395 228
rect -5453 188 -5441 222
rect -5407 188 -5395 222
rect -5453 182 -5395 188
rect -5261 222 -5203 228
rect -5261 188 -5249 222
rect -5215 188 -5203 222
rect -5261 182 -5203 188
rect -5069 222 -5011 228
rect -5069 188 -5057 222
rect -5023 188 -5011 222
rect -5069 182 -5011 188
rect -4877 222 -4819 228
rect -4877 188 -4865 222
rect -4831 188 -4819 222
rect -4877 182 -4819 188
rect -4685 222 -4627 228
rect -4685 188 -4673 222
rect -4639 188 -4627 222
rect -4685 182 -4627 188
rect -4493 222 -4435 228
rect -4493 188 -4481 222
rect -4447 188 -4435 222
rect -4493 182 -4435 188
rect -4301 222 -4243 228
rect -4301 188 -4289 222
rect -4255 188 -4243 222
rect -4301 182 -4243 188
rect -4109 222 -4051 228
rect -4109 188 -4097 222
rect -4063 188 -4051 222
rect -4109 182 -4051 188
rect -3917 222 -3859 228
rect -3917 188 -3905 222
rect -3871 188 -3859 222
rect -3917 182 -3859 188
rect -3725 222 -3667 228
rect -3725 188 -3713 222
rect -3679 188 -3667 222
rect -3725 182 -3667 188
rect -3533 222 -3475 228
rect -3533 188 -3521 222
rect -3487 188 -3475 222
rect -3533 182 -3475 188
rect -3341 222 -3283 228
rect -3341 188 -3329 222
rect -3295 188 -3283 222
rect -3341 182 -3283 188
rect -3149 222 -3091 228
rect -3149 188 -3137 222
rect -3103 188 -3091 222
rect -3149 182 -3091 188
rect -2957 222 -2899 228
rect -2957 188 -2945 222
rect -2911 188 -2899 222
rect -2957 182 -2899 188
rect -2765 222 -2707 228
rect -2765 188 -2753 222
rect -2719 188 -2707 222
rect -2765 182 -2707 188
rect -2573 222 -2515 228
rect -2573 188 -2561 222
rect -2527 188 -2515 222
rect -2573 182 -2515 188
rect -2381 222 -2323 228
rect -2381 188 -2369 222
rect -2335 188 -2323 222
rect -2381 182 -2323 188
rect -2189 222 -2131 228
rect -2189 188 -2177 222
rect -2143 188 -2131 222
rect -2189 182 -2131 188
rect -1997 222 -1939 228
rect -1997 188 -1985 222
rect -1951 188 -1939 222
rect -1997 182 -1939 188
rect -1805 222 -1747 228
rect -1805 188 -1793 222
rect -1759 188 -1747 222
rect -1805 182 -1747 188
rect -1613 222 -1555 228
rect -1613 188 -1601 222
rect -1567 188 -1555 222
rect -1613 182 -1555 188
rect -1421 222 -1363 228
rect -1421 188 -1409 222
rect -1375 188 -1363 222
rect -1421 182 -1363 188
rect -1229 222 -1171 228
rect -1229 188 -1217 222
rect -1183 188 -1171 222
rect -1229 182 -1171 188
rect -1037 222 -979 228
rect -1037 188 -1025 222
rect -991 188 -979 222
rect -1037 182 -979 188
rect -845 222 -787 228
rect -845 188 -833 222
rect -799 188 -787 222
rect -845 182 -787 188
rect -653 222 -595 228
rect -653 188 -641 222
rect -607 188 -595 222
rect -653 182 -595 188
rect -461 222 -403 228
rect -461 188 -449 222
rect -415 188 -403 222
rect -461 182 -403 188
rect -269 222 -211 228
rect -269 188 -257 222
rect -223 188 -211 222
rect -269 182 -211 188
rect -77 222 -19 228
rect -77 188 -65 222
rect -31 188 -19 222
rect -77 182 -19 188
rect 115 222 173 228
rect 115 188 127 222
rect 161 188 173 222
rect 115 182 173 188
rect 307 222 365 228
rect 307 188 319 222
rect 353 188 365 222
rect 307 182 365 188
rect 499 222 557 228
rect 499 188 511 222
rect 545 188 557 222
rect 499 182 557 188
rect 691 222 749 228
rect 691 188 703 222
rect 737 188 749 222
rect 691 182 749 188
rect 883 222 941 228
rect 883 188 895 222
rect 929 188 941 222
rect 883 182 941 188
rect 1075 222 1133 228
rect 1075 188 1087 222
rect 1121 188 1133 222
rect 1075 182 1133 188
rect 1267 222 1325 228
rect 1267 188 1279 222
rect 1313 188 1325 222
rect 1267 182 1325 188
rect 1459 222 1517 228
rect 1459 188 1471 222
rect 1505 188 1517 222
rect 1459 182 1517 188
rect 1651 222 1709 228
rect 1651 188 1663 222
rect 1697 188 1709 222
rect 1651 182 1709 188
rect 1843 222 1901 228
rect 1843 188 1855 222
rect 1889 188 1901 222
rect 1843 182 1901 188
rect 2035 222 2093 228
rect 2035 188 2047 222
rect 2081 188 2093 222
rect 2035 182 2093 188
rect 2227 222 2285 228
rect 2227 188 2239 222
rect 2273 188 2285 222
rect 2227 182 2285 188
rect 2419 222 2477 228
rect 2419 188 2431 222
rect 2465 188 2477 222
rect 2419 182 2477 188
rect 2611 222 2669 228
rect 2611 188 2623 222
rect 2657 188 2669 222
rect 2611 182 2669 188
rect 2803 222 2861 228
rect 2803 188 2815 222
rect 2849 188 2861 222
rect 2803 182 2861 188
rect 2995 222 3053 228
rect 2995 188 3007 222
rect 3041 188 3053 222
rect 2995 182 3053 188
rect 3187 222 3245 228
rect 3187 188 3199 222
rect 3233 188 3245 222
rect 3187 182 3245 188
rect 3379 222 3437 228
rect 3379 188 3391 222
rect 3425 188 3437 222
rect 3379 182 3437 188
rect 3571 222 3629 228
rect 3571 188 3583 222
rect 3617 188 3629 222
rect 3571 182 3629 188
rect 3763 222 3821 228
rect 3763 188 3775 222
rect 3809 188 3821 222
rect 3763 182 3821 188
rect 3955 222 4013 228
rect 3955 188 3967 222
rect 4001 188 4013 222
rect 3955 182 4013 188
rect 4147 222 4205 228
rect 4147 188 4159 222
rect 4193 188 4205 222
rect 4147 182 4205 188
rect 4339 222 4397 228
rect 4339 188 4351 222
rect 4385 188 4397 222
rect 4339 182 4397 188
rect 4531 222 4589 228
rect 4531 188 4543 222
rect 4577 188 4589 222
rect 4531 182 4589 188
rect 4723 222 4781 228
rect 4723 188 4735 222
rect 4769 188 4781 222
rect 4723 182 4781 188
rect 4915 222 4973 228
rect 4915 188 4927 222
rect 4961 188 4973 222
rect 4915 182 4973 188
rect 5107 222 5165 228
rect 5107 188 5119 222
rect 5153 188 5165 222
rect 5107 182 5165 188
rect 5299 222 5357 228
rect 5299 188 5311 222
rect 5345 188 5357 222
rect 5299 182 5357 188
rect 5491 222 5549 228
rect 5491 188 5503 222
rect 5537 188 5549 222
rect 5491 182 5549 188
rect 5683 222 5741 228
rect 5683 188 5695 222
rect 5729 188 5741 222
rect 5683 182 5741 188
rect 5875 222 5933 228
rect 5875 188 5887 222
rect 5921 188 5933 222
rect 5875 182 5933 188
rect 6067 222 6125 228
rect 6067 188 6079 222
rect 6113 188 6125 222
rect 6067 182 6125 188
rect 6259 222 6317 228
rect 6259 188 6271 222
rect 6305 188 6317 222
rect 6259 182 6317 188
rect 6451 222 6509 228
rect 6451 188 6463 222
rect 6497 188 6509 222
rect 6451 182 6509 188
rect 6643 222 6701 228
rect 6643 188 6655 222
rect 6689 188 6701 222
rect 6643 182 6701 188
rect 6835 222 6893 228
rect 6835 188 6847 222
rect 6881 188 6893 222
rect 6835 182 6893 188
rect 7027 222 7085 228
rect 7027 188 7039 222
rect 7073 188 7085 222
rect 7027 182 7085 188
rect 7219 222 7277 228
rect 7219 188 7231 222
rect 7265 188 7277 222
rect 7219 182 7277 188
rect 7411 222 7469 228
rect 7411 188 7423 222
rect 7457 188 7469 222
rect 7411 182 7469 188
rect 7603 222 7661 228
rect 7603 188 7615 222
rect 7649 188 7661 222
rect 7603 182 7661 188
rect 7795 222 7853 228
rect 7795 188 7807 222
rect 7841 188 7853 222
rect 7795 182 7853 188
rect 7987 222 8045 228
rect 7987 188 7999 222
rect 8033 188 8045 222
rect 7987 182 8045 188
rect 8179 222 8237 228
rect 8179 188 8191 222
rect 8225 188 8237 222
rect 8179 182 8237 188
rect 8371 222 8429 228
rect 8371 188 8383 222
rect 8417 188 8429 222
rect 8371 182 8429 188
rect 8563 222 8621 228
rect 8563 188 8575 222
rect 8609 188 8621 222
rect 8563 182 8621 188
rect 8755 222 8813 228
rect 8755 188 8767 222
rect 8801 188 8813 222
rect 8755 182 8813 188
rect 8947 222 9005 228
rect 8947 188 8959 222
rect 8993 188 9005 222
rect 8947 182 9005 188
rect 9139 222 9197 228
rect 9139 188 9151 222
rect 9185 188 9197 222
rect 9139 182 9197 188
rect 9331 222 9389 228
rect 9331 188 9343 222
rect 9377 188 9389 222
rect 9331 182 9389 188
rect 9523 222 9581 228
rect 9523 188 9535 222
rect 9569 188 9581 222
rect 9523 182 9581 188
rect 9715 222 9773 228
rect 9715 188 9727 222
rect 9761 188 9773 222
rect 9715 182 9773 188
rect 9907 222 9965 228
rect 9907 188 9919 222
rect 9953 188 9965 222
rect 9907 182 9965 188
rect 10099 222 10157 228
rect 10099 188 10111 222
rect 10145 188 10157 222
rect 10099 182 10157 188
rect 10291 222 10349 228
rect 10291 188 10303 222
rect 10337 188 10349 222
rect 10291 182 10349 188
rect 10483 222 10541 228
rect 10483 188 10495 222
rect 10529 188 10541 222
rect 10483 182 10541 188
rect 10675 222 10733 228
rect 10675 188 10687 222
rect 10721 188 10733 222
rect 10675 182 10733 188
rect 10867 222 10925 228
rect 10867 188 10879 222
rect 10913 188 10925 222
rect 10867 182 10925 188
rect 11059 222 11117 228
rect 11059 188 11071 222
rect 11105 188 11117 222
rect 11059 182 11117 188
rect 11251 222 11309 228
rect 11251 188 11263 222
rect 11297 188 11309 222
rect 11251 182 11309 188
rect 11443 222 11501 228
rect 11443 188 11455 222
rect 11489 188 11501 222
rect 11443 182 11501 188
rect 11635 222 11693 228
rect 11635 188 11647 222
rect 11681 188 11693 222
rect 11635 182 11693 188
rect 11827 222 11885 228
rect 11827 188 11839 222
rect 11873 188 11885 222
rect 11827 182 11885 188
rect 12019 222 12077 228
rect 12019 188 12031 222
rect 12065 188 12077 222
rect 12019 182 12077 188
rect 12211 222 12269 228
rect 12211 188 12223 222
rect 12257 188 12269 222
rect 12211 182 12269 188
rect 12403 222 12461 228
rect 12403 188 12415 222
rect 12449 188 12461 222
rect 12403 182 12461 188
rect 12595 222 12653 228
rect 12595 188 12607 222
rect 12641 188 12653 222
rect 12595 182 12653 188
rect 12787 222 12845 228
rect 12787 188 12799 222
rect 12833 188 12845 222
rect 12787 182 12845 188
rect 12979 222 13037 228
rect 12979 188 12991 222
rect 13025 188 13037 222
rect 12979 182 13037 188
rect 13171 222 13229 228
rect 13171 188 13183 222
rect 13217 188 13229 222
rect 13171 182 13229 188
rect 13363 222 13421 228
rect 13363 188 13375 222
rect 13409 188 13421 222
rect 13363 182 13421 188
rect 13555 222 13613 228
rect 13555 188 13567 222
rect 13601 188 13613 222
rect 13555 182 13613 188
rect 13747 222 13805 228
rect 13747 188 13759 222
rect 13793 188 13805 222
rect 13747 182 13805 188
rect 13939 222 13997 228
rect 13939 188 13951 222
rect 13985 188 13997 222
rect 13939 182 13997 188
rect 14131 222 14189 228
rect 14131 188 14143 222
rect 14177 188 14189 222
rect 14131 182 14189 188
rect 14323 222 14381 228
rect 14323 188 14335 222
rect 14369 188 14381 222
rect 14323 182 14381 188
rect 14515 222 14573 228
rect 14515 188 14527 222
rect 14561 188 14573 222
rect 14515 182 14573 188
rect 14707 222 14765 228
rect 14707 188 14719 222
rect 14753 188 14765 222
rect 14707 182 14765 188
rect 14899 222 14957 228
rect 14899 188 14911 222
rect 14945 188 14957 222
rect 14899 182 14957 188
rect 15091 222 15149 228
rect 15091 188 15103 222
rect 15137 188 15149 222
rect 15091 182 15149 188
rect 15283 222 15341 228
rect 15283 188 15295 222
rect 15329 188 15341 222
rect 15283 182 15341 188
rect 15475 222 15533 228
rect 15475 188 15487 222
rect 15521 188 15533 222
rect 15475 182 15533 188
rect 15667 222 15725 228
rect 15667 188 15679 222
rect 15713 188 15725 222
rect 15667 182 15725 188
rect 15859 222 15917 228
rect 15859 188 15871 222
rect 15905 188 15917 222
rect 15859 182 15917 188
rect 16051 222 16109 228
rect 16051 188 16063 222
rect 16097 188 16109 222
rect 16051 182 16109 188
rect 16243 222 16301 228
rect 16243 188 16255 222
rect 16289 188 16301 222
rect 16243 182 16301 188
rect 16435 222 16493 228
rect 16435 188 16447 222
rect 16481 188 16493 222
rect 16435 182 16493 188
rect 16627 222 16685 228
rect 16627 188 16639 222
rect 16673 188 16685 222
rect 16627 182 16685 188
rect 16819 222 16877 228
rect 16819 188 16831 222
rect 16865 188 16877 222
rect 16819 182 16877 188
rect 17011 222 17069 228
rect 17011 188 17023 222
rect 17057 188 17069 222
rect 17011 182 17069 188
rect 17203 222 17261 228
rect 17203 188 17215 222
rect 17249 188 17261 222
rect 17203 182 17261 188
rect 17395 222 17453 228
rect 17395 188 17407 222
rect 17441 188 17453 222
rect 17395 182 17453 188
rect 17587 222 17645 228
rect 17587 188 17599 222
rect 17633 188 17645 222
rect 17587 182 17645 188
rect 17779 222 17837 228
rect 17779 188 17791 222
rect 17825 188 17837 222
rect 17779 182 17837 188
rect 17971 222 18029 228
rect 17971 188 17983 222
rect 18017 188 18029 222
rect 17971 182 18029 188
rect 18163 222 18221 228
rect 18163 188 18175 222
rect 18209 188 18221 222
rect 18163 182 18221 188
rect 18355 222 18413 228
rect 18355 188 18367 222
rect 18401 188 18413 222
rect 18355 182 18413 188
rect 18547 222 18605 228
rect 18547 188 18559 222
rect 18593 188 18605 222
rect 18547 182 18605 188
rect 18739 222 18797 228
rect 18739 188 18751 222
rect 18785 188 18797 222
rect 18739 182 18797 188
rect 18931 222 18989 228
rect 18931 188 18943 222
rect 18977 188 18989 222
rect 18931 182 18989 188
rect 19123 222 19181 228
rect 19123 188 19135 222
rect 19169 188 19181 222
rect 19123 182 19181 188
rect -19223 138 -19177 150
rect -19223 -138 -19217 138
rect -19183 -138 -19177 138
rect -19223 -150 -19177 -138
rect -19127 138 -19081 150
rect -19127 -138 -19121 138
rect -19087 -138 -19081 138
rect -19127 -150 -19081 -138
rect -19031 138 -18985 150
rect -19031 -138 -19025 138
rect -18991 -138 -18985 138
rect -19031 -150 -18985 -138
rect -18935 138 -18889 150
rect -18935 -138 -18929 138
rect -18895 -138 -18889 138
rect -18935 -150 -18889 -138
rect -18839 138 -18793 150
rect -18839 -138 -18833 138
rect -18799 -138 -18793 138
rect -18839 -150 -18793 -138
rect -18743 138 -18697 150
rect -18743 -138 -18737 138
rect -18703 -138 -18697 138
rect -18743 -150 -18697 -138
rect -18647 138 -18601 150
rect -18647 -138 -18641 138
rect -18607 -138 -18601 138
rect -18647 -150 -18601 -138
rect -18551 138 -18505 150
rect -18551 -138 -18545 138
rect -18511 -138 -18505 138
rect -18551 -150 -18505 -138
rect -18455 138 -18409 150
rect -18455 -138 -18449 138
rect -18415 -138 -18409 138
rect -18455 -150 -18409 -138
rect -18359 138 -18313 150
rect -18359 -138 -18353 138
rect -18319 -138 -18313 138
rect -18359 -150 -18313 -138
rect -18263 138 -18217 150
rect -18263 -138 -18257 138
rect -18223 -138 -18217 138
rect -18263 -150 -18217 -138
rect -18167 138 -18121 150
rect -18167 -138 -18161 138
rect -18127 -138 -18121 138
rect -18167 -150 -18121 -138
rect -18071 138 -18025 150
rect -18071 -138 -18065 138
rect -18031 -138 -18025 138
rect -18071 -150 -18025 -138
rect -17975 138 -17929 150
rect -17975 -138 -17969 138
rect -17935 -138 -17929 138
rect -17975 -150 -17929 -138
rect -17879 138 -17833 150
rect -17879 -138 -17873 138
rect -17839 -138 -17833 138
rect -17879 -150 -17833 -138
rect -17783 138 -17737 150
rect -17783 -138 -17777 138
rect -17743 -138 -17737 138
rect -17783 -150 -17737 -138
rect -17687 138 -17641 150
rect -17687 -138 -17681 138
rect -17647 -138 -17641 138
rect -17687 -150 -17641 -138
rect -17591 138 -17545 150
rect -17591 -138 -17585 138
rect -17551 -138 -17545 138
rect -17591 -150 -17545 -138
rect -17495 138 -17449 150
rect -17495 -138 -17489 138
rect -17455 -138 -17449 138
rect -17495 -150 -17449 -138
rect -17399 138 -17353 150
rect -17399 -138 -17393 138
rect -17359 -138 -17353 138
rect -17399 -150 -17353 -138
rect -17303 138 -17257 150
rect -17303 -138 -17297 138
rect -17263 -138 -17257 138
rect -17303 -150 -17257 -138
rect -17207 138 -17161 150
rect -17207 -138 -17201 138
rect -17167 -138 -17161 138
rect -17207 -150 -17161 -138
rect -17111 138 -17065 150
rect -17111 -138 -17105 138
rect -17071 -138 -17065 138
rect -17111 -150 -17065 -138
rect -17015 138 -16969 150
rect -17015 -138 -17009 138
rect -16975 -138 -16969 138
rect -17015 -150 -16969 -138
rect -16919 138 -16873 150
rect -16919 -138 -16913 138
rect -16879 -138 -16873 138
rect -16919 -150 -16873 -138
rect -16823 138 -16777 150
rect -16823 -138 -16817 138
rect -16783 -138 -16777 138
rect -16823 -150 -16777 -138
rect -16727 138 -16681 150
rect -16727 -138 -16721 138
rect -16687 -138 -16681 138
rect -16727 -150 -16681 -138
rect -16631 138 -16585 150
rect -16631 -138 -16625 138
rect -16591 -138 -16585 138
rect -16631 -150 -16585 -138
rect -16535 138 -16489 150
rect -16535 -138 -16529 138
rect -16495 -138 -16489 138
rect -16535 -150 -16489 -138
rect -16439 138 -16393 150
rect -16439 -138 -16433 138
rect -16399 -138 -16393 138
rect -16439 -150 -16393 -138
rect -16343 138 -16297 150
rect -16343 -138 -16337 138
rect -16303 -138 -16297 138
rect -16343 -150 -16297 -138
rect -16247 138 -16201 150
rect -16247 -138 -16241 138
rect -16207 -138 -16201 138
rect -16247 -150 -16201 -138
rect -16151 138 -16105 150
rect -16151 -138 -16145 138
rect -16111 -138 -16105 138
rect -16151 -150 -16105 -138
rect -16055 138 -16009 150
rect -16055 -138 -16049 138
rect -16015 -138 -16009 138
rect -16055 -150 -16009 -138
rect -15959 138 -15913 150
rect -15959 -138 -15953 138
rect -15919 -138 -15913 138
rect -15959 -150 -15913 -138
rect -15863 138 -15817 150
rect -15863 -138 -15857 138
rect -15823 -138 -15817 138
rect -15863 -150 -15817 -138
rect -15767 138 -15721 150
rect -15767 -138 -15761 138
rect -15727 -138 -15721 138
rect -15767 -150 -15721 -138
rect -15671 138 -15625 150
rect -15671 -138 -15665 138
rect -15631 -138 -15625 138
rect -15671 -150 -15625 -138
rect -15575 138 -15529 150
rect -15575 -138 -15569 138
rect -15535 -138 -15529 138
rect -15575 -150 -15529 -138
rect -15479 138 -15433 150
rect -15479 -138 -15473 138
rect -15439 -138 -15433 138
rect -15479 -150 -15433 -138
rect -15383 138 -15337 150
rect -15383 -138 -15377 138
rect -15343 -138 -15337 138
rect -15383 -150 -15337 -138
rect -15287 138 -15241 150
rect -15287 -138 -15281 138
rect -15247 -138 -15241 138
rect -15287 -150 -15241 -138
rect -15191 138 -15145 150
rect -15191 -138 -15185 138
rect -15151 -138 -15145 138
rect -15191 -150 -15145 -138
rect -15095 138 -15049 150
rect -15095 -138 -15089 138
rect -15055 -138 -15049 138
rect -15095 -150 -15049 -138
rect -14999 138 -14953 150
rect -14999 -138 -14993 138
rect -14959 -138 -14953 138
rect -14999 -150 -14953 -138
rect -14903 138 -14857 150
rect -14903 -138 -14897 138
rect -14863 -138 -14857 138
rect -14903 -150 -14857 -138
rect -14807 138 -14761 150
rect -14807 -138 -14801 138
rect -14767 -138 -14761 138
rect -14807 -150 -14761 -138
rect -14711 138 -14665 150
rect -14711 -138 -14705 138
rect -14671 -138 -14665 138
rect -14711 -150 -14665 -138
rect -14615 138 -14569 150
rect -14615 -138 -14609 138
rect -14575 -138 -14569 138
rect -14615 -150 -14569 -138
rect -14519 138 -14473 150
rect -14519 -138 -14513 138
rect -14479 -138 -14473 138
rect -14519 -150 -14473 -138
rect -14423 138 -14377 150
rect -14423 -138 -14417 138
rect -14383 -138 -14377 138
rect -14423 -150 -14377 -138
rect -14327 138 -14281 150
rect -14327 -138 -14321 138
rect -14287 -138 -14281 138
rect -14327 -150 -14281 -138
rect -14231 138 -14185 150
rect -14231 -138 -14225 138
rect -14191 -138 -14185 138
rect -14231 -150 -14185 -138
rect -14135 138 -14089 150
rect -14135 -138 -14129 138
rect -14095 -138 -14089 138
rect -14135 -150 -14089 -138
rect -14039 138 -13993 150
rect -14039 -138 -14033 138
rect -13999 -138 -13993 138
rect -14039 -150 -13993 -138
rect -13943 138 -13897 150
rect -13943 -138 -13937 138
rect -13903 -138 -13897 138
rect -13943 -150 -13897 -138
rect -13847 138 -13801 150
rect -13847 -138 -13841 138
rect -13807 -138 -13801 138
rect -13847 -150 -13801 -138
rect -13751 138 -13705 150
rect -13751 -138 -13745 138
rect -13711 -138 -13705 138
rect -13751 -150 -13705 -138
rect -13655 138 -13609 150
rect -13655 -138 -13649 138
rect -13615 -138 -13609 138
rect -13655 -150 -13609 -138
rect -13559 138 -13513 150
rect -13559 -138 -13553 138
rect -13519 -138 -13513 138
rect -13559 -150 -13513 -138
rect -13463 138 -13417 150
rect -13463 -138 -13457 138
rect -13423 -138 -13417 138
rect -13463 -150 -13417 -138
rect -13367 138 -13321 150
rect -13367 -138 -13361 138
rect -13327 -138 -13321 138
rect -13367 -150 -13321 -138
rect -13271 138 -13225 150
rect -13271 -138 -13265 138
rect -13231 -138 -13225 138
rect -13271 -150 -13225 -138
rect -13175 138 -13129 150
rect -13175 -138 -13169 138
rect -13135 -138 -13129 138
rect -13175 -150 -13129 -138
rect -13079 138 -13033 150
rect -13079 -138 -13073 138
rect -13039 -138 -13033 138
rect -13079 -150 -13033 -138
rect -12983 138 -12937 150
rect -12983 -138 -12977 138
rect -12943 -138 -12937 138
rect -12983 -150 -12937 -138
rect -12887 138 -12841 150
rect -12887 -138 -12881 138
rect -12847 -138 -12841 138
rect -12887 -150 -12841 -138
rect -12791 138 -12745 150
rect -12791 -138 -12785 138
rect -12751 -138 -12745 138
rect -12791 -150 -12745 -138
rect -12695 138 -12649 150
rect -12695 -138 -12689 138
rect -12655 -138 -12649 138
rect -12695 -150 -12649 -138
rect -12599 138 -12553 150
rect -12599 -138 -12593 138
rect -12559 -138 -12553 138
rect -12599 -150 -12553 -138
rect -12503 138 -12457 150
rect -12503 -138 -12497 138
rect -12463 -138 -12457 138
rect -12503 -150 -12457 -138
rect -12407 138 -12361 150
rect -12407 -138 -12401 138
rect -12367 -138 -12361 138
rect -12407 -150 -12361 -138
rect -12311 138 -12265 150
rect -12311 -138 -12305 138
rect -12271 -138 -12265 138
rect -12311 -150 -12265 -138
rect -12215 138 -12169 150
rect -12215 -138 -12209 138
rect -12175 -138 -12169 138
rect -12215 -150 -12169 -138
rect -12119 138 -12073 150
rect -12119 -138 -12113 138
rect -12079 -138 -12073 138
rect -12119 -150 -12073 -138
rect -12023 138 -11977 150
rect -12023 -138 -12017 138
rect -11983 -138 -11977 138
rect -12023 -150 -11977 -138
rect -11927 138 -11881 150
rect -11927 -138 -11921 138
rect -11887 -138 -11881 138
rect -11927 -150 -11881 -138
rect -11831 138 -11785 150
rect -11831 -138 -11825 138
rect -11791 -138 -11785 138
rect -11831 -150 -11785 -138
rect -11735 138 -11689 150
rect -11735 -138 -11729 138
rect -11695 -138 -11689 138
rect -11735 -150 -11689 -138
rect -11639 138 -11593 150
rect -11639 -138 -11633 138
rect -11599 -138 -11593 138
rect -11639 -150 -11593 -138
rect -11543 138 -11497 150
rect -11543 -138 -11537 138
rect -11503 -138 -11497 138
rect -11543 -150 -11497 -138
rect -11447 138 -11401 150
rect -11447 -138 -11441 138
rect -11407 -138 -11401 138
rect -11447 -150 -11401 -138
rect -11351 138 -11305 150
rect -11351 -138 -11345 138
rect -11311 -138 -11305 138
rect -11351 -150 -11305 -138
rect -11255 138 -11209 150
rect -11255 -138 -11249 138
rect -11215 -138 -11209 138
rect -11255 -150 -11209 -138
rect -11159 138 -11113 150
rect -11159 -138 -11153 138
rect -11119 -138 -11113 138
rect -11159 -150 -11113 -138
rect -11063 138 -11017 150
rect -11063 -138 -11057 138
rect -11023 -138 -11017 138
rect -11063 -150 -11017 -138
rect -10967 138 -10921 150
rect -10967 -138 -10961 138
rect -10927 -138 -10921 138
rect -10967 -150 -10921 -138
rect -10871 138 -10825 150
rect -10871 -138 -10865 138
rect -10831 -138 -10825 138
rect -10871 -150 -10825 -138
rect -10775 138 -10729 150
rect -10775 -138 -10769 138
rect -10735 -138 -10729 138
rect -10775 -150 -10729 -138
rect -10679 138 -10633 150
rect -10679 -138 -10673 138
rect -10639 -138 -10633 138
rect -10679 -150 -10633 -138
rect -10583 138 -10537 150
rect -10583 -138 -10577 138
rect -10543 -138 -10537 138
rect -10583 -150 -10537 -138
rect -10487 138 -10441 150
rect -10487 -138 -10481 138
rect -10447 -138 -10441 138
rect -10487 -150 -10441 -138
rect -10391 138 -10345 150
rect -10391 -138 -10385 138
rect -10351 -138 -10345 138
rect -10391 -150 -10345 -138
rect -10295 138 -10249 150
rect -10295 -138 -10289 138
rect -10255 -138 -10249 138
rect -10295 -150 -10249 -138
rect -10199 138 -10153 150
rect -10199 -138 -10193 138
rect -10159 -138 -10153 138
rect -10199 -150 -10153 -138
rect -10103 138 -10057 150
rect -10103 -138 -10097 138
rect -10063 -138 -10057 138
rect -10103 -150 -10057 -138
rect -10007 138 -9961 150
rect -10007 -138 -10001 138
rect -9967 -138 -9961 138
rect -10007 -150 -9961 -138
rect -9911 138 -9865 150
rect -9911 -138 -9905 138
rect -9871 -138 -9865 138
rect -9911 -150 -9865 -138
rect -9815 138 -9769 150
rect -9815 -138 -9809 138
rect -9775 -138 -9769 138
rect -9815 -150 -9769 -138
rect -9719 138 -9673 150
rect -9719 -138 -9713 138
rect -9679 -138 -9673 138
rect -9719 -150 -9673 -138
rect -9623 138 -9577 150
rect -9623 -138 -9617 138
rect -9583 -138 -9577 138
rect -9623 -150 -9577 -138
rect -9527 138 -9481 150
rect -9527 -138 -9521 138
rect -9487 -138 -9481 138
rect -9527 -150 -9481 -138
rect -9431 138 -9385 150
rect -9431 -138 -9425 138
rect -9391 -138 -9385 138
rect -9431 -150 -9385 -138
rect -9335 138 -9289 150
rect -9335 -138 -9329 138
rect -9295 -138 -9289 138
rect -9335 -150 -9289 -138
rect -9239 138 -9193 150
rect -9239 -138 -9233 138
rect -9199 -138 -9193 138
rect -9239 -150 -9193 -138
rect -9143 138 -9097 150
rect -9143 -138 -9137 138
rect -9103 -138 -9097 138
rect -9143 -150 -9097 -138
rect -9047 138 -9001 150
rect -9047 -138 -9041 138
rect -9007 -138 -9001 138
rect -9047 -150 -9001 -138
rect -8951 138 -8905 150
rect -8951 -138 -8945 138
rect -8911 -138 -8905 138
rect -8951 -150 -8905 -138
rect -8855 138 -8809 150
rect -8855 -138 -8849 138
rect -8815 -138 -8809 138
rect -8855 -150 -8809 -138
rect -8759 138 -8713 150
rect -8759 -138 -8753 138
rect -8719 -138 -8713 138
rect -8759 -150 -8713 -138
rect -8663 138 -8617 150
rect -8663 -138 -8657 138
rect -8623 -138 -8617 138
rect -8663 -150 -8617 -138
rect -8567 138 -8521 150
rect -8567 -138 -8561 138
rect -8527 -138 -8521 138
rect -8567 -150 -8521 -138
rect -8471 138 -8425 150
rect -8471 -138 -8465 138
rect -8431 -138 -8425 138
rect -8471 -150 -8425 -138
rect -8375 138 -8329 150
rect -8375 -138 -8369 138
rect -8335 -138 -8329 138
rect -8375 -150 -8329 -138
rect -8279 138 -8233 150
rect -8279 -138 -8273 138
rect -8239 -138 -8233 138
rect -8279 -150 -8233 -138
rect -8183 138 -8137 150
rect -8183 -138 -8177 138
rect -8143 -138 -8137 138
rect -8183 -150 -8137 -138
rect -8087 138 -8041 150
rect -8087 -138 -8081 138
rect -8047 -138 -8041 138
rect -8087 -150 -8041 -138
rect -7991 138 -7945 150
rect -7991 -138 -7985 138
rect -7951 -138 -7945 138
rect -7991 -150 -7945 -138
rect -7895 138 -7849 150
rect -7895 -138 -7889 138
rect -7855 -138 -7849 138
rect -7895 -150 -7849 -138
rect -7799 138 -7753 150
rect -7799 -138 -7793 138
rect -7759 -138 -7753 138
rect -7799 -150 -7753 -138
rect -7703 138 -7657 150
rect -7703 -138 -7697 138
rect -7663 -138 -7657 138
rect -7703 -150 -7657 -138
rect -7607 138 -7561 150
rect -7607 -138 -7601 138
rect -7567 -138 -7561 138
rect -7607 -150 -7561 -138
rect -7511 138 -7465 150
rect -7511 -138 -7505 138
rect -7471 -138 -7465 138
rect -7511 -150 -7465 -138
rect -7415 138 -7369 150
rect -7415 -138 -7409 138
rect -7375 -138 -7369 138
rect -7415 -150 -7369 -138
rect -7319 138 -7273 150
rect -7319 -138 -7313 138
rect -7279 -138 -7273 138
rect -7319 -150 -7273 -138
rect -7223 138 -7177 150
rect -7223 -138 -7217 138
rect -7183 -138 -7177 138
rect -7223 -150 -7177 -138
rect -7127 138 -7081 150
rect -7127 -138 -7121 138
rect -7087 -138 -7081 138
rect -7127 -150 -7081 -138
rect -7031 138 -6985 150
rect -7031 -138 -7025 138
rect -6991 -138 -6985 138
rect -7031 -150 -6985 -138
rect -6935 138 -6889 150
rect -6935 -138 -6929 138
rect -6895 -138 -6889 138
rect -6935 -150 -6889 -138
rect -6839 138 -6793 150
rect -6839 -138 -6833 138
rect -6799 -138 -6793 138
rect -6839 -150 -6793 -138
rect -6743 138 -6697 150
rect -6743 -138 -6737 138
rect -6703 -138 -6697 138
rect -6743 -150 -6697 -138
rect -6647 138 -6601 150
rect -6647 -138 -6641 138
rect -6607 -138 -6601 138
rect -6647 -150 -6601 -138
rect -6551 138 -6505 150
rect -6551 -138 -6545 138
rect -6511 -138 -6505 138
rect -6551 -150 -6505 -138
rect -6455 138 -6409 150
rect -6455 -138 -6449 138
rect -6415 -138 -6409 138
rect -6455 -150 -6409 -138
rect -6359 138 -6313 150
rect -6359 -138 -6353 138
rect -6319 -138 -6313 138
rect -6359 -150 -6313 -138
rect -6263 138 -6217 150
rect -6263 -138 -6257 138
rect -6223 -138 -6217 138
rect -6263 -150 -6217 -138
rect -6167 138 -6121 150
rect -6167 -138 -6161 138
rect -6127 -138 -6121 138
rect -6167 -150 -6121 -138
rect -6071 138 -6025 150
rect -6071 -138 -6065 138
rect -6031 -138 -6025 138
rect -6071 -150 -6025 -138
rect -5975 138 -5929 150
rect -5975 -138 -5969 138
rect -5935 -138 -5929 138
rect -5975 -150 -5929 -138
rect -5879 138 -5833 150
rect -5879 -138 -5873 138
rect -5839 -138 -5833 138
rect -5879 -150 -5833 -138
rect -5783 138 -5737 150
rect -5783 -138 -5777 138
rect -5743 -138 -5737 138
rect -5783 -150 -5737 -138
rect -5687 138 -5641 150
rect -5687 -138 -5681 138
rect -5647 -138 -5641 138
rect -5687 -150 -5641 -138
rect -5591 138 -5545 150
rect -5591 -138 -5585 138
rect -5551 -138 -5545 138
rect -5591 -150 -5545 -138
rect -5495 138 -5449 150
rect -5495 -138 -5489 138
rect -5455 -138 -5449 138
rect -5495 -150 -5449 -138
rect -5399 138 -5353 150
rect -5399 -138 -5393 138
rect -5359 -138 -5353 138
rect -5399 -150 -5353 -138
rect -5303 138 -5257 150
rect -5303 -138 -5297 138
rect -5263 -138 -5257 138
rect -5303 -150 -5257 -138
rect -5207 138 -5161 150
rect -5207 -138 -5201 138
rect -5167 -138 -5161 138
rect -5207 -150 -5161 -138
rect -5111 138 -5065 150
rect -5111 -138 -5105 138
rect -5071 -138 -5065 138
rect -5111 -150 -5065 -138
rect -5015 138 -4969 150
rect -5015 -138 -5009 138
rect -4975 -138 -4969 138
rect -5015 -150 -4969 -138
rect -4919 138 -4873 150
rect -4919 -138 -4913 138
rect -4879 -138 -4873 138
rect -4919 -150 -4873 -138
rect -4823 138 -4777 150
rect -4823 -138 -4817 138
rect -4783 -138 -4777 138
rect -4823 -150 -4777 -138
rect -4727 138 -4681 150
rect -4727 -138 -4721 138
rect -4687 -138 -4681 138
rect -4727 -150 -4681 -138
rect -4631 138 -4585 150
rect -4631 -138 -4625 138
rect -4591 -138 -4585 138
rect -4631 -150 -4585 -138
rect -4535 138 -4489 150
rect -4535 -138 -4529 138
rect -4495 -138 -4489 138
rect -4535 -150 -4489 -138
rect -4439 138 -4393 150
rect -4439 -138 -4433 138
rect -4399 -138 -4393 138
rect -4439 -150 -4393 -138
rect -4343 138 -4297 150
rect -4343 -138 -4337 138
rect -4303 -138 -4297 138
rect -4343 -150 -4297 -138
rect -4247 138 -4201 150
rect -4247 -138 -4241 138
rect -4207 -138 -4201 138
rect -4247 -150 -4201 -138
rect -4151 138 -4105 150
rect -4151 -138 -4145 138
rect -4111 -138 -4105 138
rect -4151 -150 -4105 -138
rect -4055 138 -4009 150
rect -4055 -138 -4049 138
rect -4015 -138 -4009 138
rect -4055 -150 -4009 -138
rect -3959 138 -3913 150
rect -3959 -138 -3953 138
rect -3919 -138 -3913 138
rect -3959 -150 -3913 -138
rect -3863 138 -3817 150
rect -3863 -138 -3857 138
rect -3823 -138 -3817 138
rect -3863 -150 -3817 -138
rect -3767 138 -3721 150
rect -3767 -138 -3761 138
rect -3727 -138 -3721 138
rect -3767 -150 -3721 -138
rect -3671 138 -3625 150
rect -3671 -138 -3665 138
rect -3631 -138 -3625 138
rect -3671 -150 -3625 -138
rect -3575 138 -3529 150
rect -3575 -138 -3569 138
rect -3535 -138 -3529 138
rect -3575 -150 -3529 -138
rect -3479 138 -3433 150
rect -3479 -138 -3473 138
rect -3439 -138 -3433 138
rect -3479 -150 -3433 -138
rect -3383 138 -3337 150
rect -3383 -138 -3377 138
rect -3343 -138 -3337 138
rect -3383 -150 -3337 -138
rect -3287 138 -3241 150
rect -3287 -138 -3281 138
rect -3247 -138 -3241 138
rect -3287 -150 -3241 -138
rect -3191 138 -3145 150
rect -3191 -138 -3185 138
rect -3151 -138 -3145 138
rect -3191 -150 -3145 -138
rect -3095 138 -3049 150
rect -3095 -138 -3089 138
rect -3055 -138 -3049 138
rect -3095 -150 -3049 -138
rect -2999 138 -2953 150
rect -2999 -138 -2993 138
rect -2959 -138 -2953 138
rect -2999 -150 -2953 -138
rect -2903 138 -2857 150
rect -2903 -138 -2897 138
rect -2863 -138 -2857 138
rect -2903 -150 -2857 -138
rect -2807 138 -2761 150
rect -2807 -138 -2801 138
rect -2767 -138 -2761 138
rect -2807 -150 -2761 -138
rect -2711 138 -2665 150
rect -2711 -138 -2705 138
rect -2671 -138 -2665 138
rect -2711 -150 -2665 -138
rect -2615 138 -2569 150
rect -2615 -138 -2609 138
rect -2575 -138 -2569 138
rect -2615 -150 -2569 -138
rect -2519 138 -2473 150
rect -2519 -138 -2513 138
rect -2479 -138 -2473 138
rect -2519 -150 -2473 -138
rect -2423 138 -2377 150
rect -2423 -138 -2417 138
rect -2383 -138 -2377 138
rect -2423 -150 -2377 -138
rect -2327 138 -2281 150
rect -2327 -138 -2321 138
rect -2287 -138 -2281 138
rect -2327 -150 -2281 -138
rect -2231 138 -2185 150
rect -2231 -138 -2225 138
rect -2191 -138 -2185 138
rect -2231 -150 -2185 -138
rect -2135 138 -2089 150
rect -2135 -138 -2129 138
rect -2095 -138 -2089 138
rect -2135 -150 -2089 -138
rect -2039 138 -1993 150
rect -2039 -138 -2033 138
rect -1999 -138 -1993 138
rect -2039 -150 -1993 -138
rect -1943 138 -1897 150
rect -1943 -138 -1937 138
rect -1903 -138 -1897 138
rect -1943 -150 -1897 -138
rect -1847 138 -1801 150
rect -1847 -138 -1841 138
rect -1807 -138 -1801 138
rect -1847 -150 -1801 -138
rect -1751 138 -1705 150
rect -1751 -138 -1745 138
rect -1711 -138 -1705 138
rect -1751 -150 -1705 -138
rect -1655 138 -1609 150
rect -1655 -138 -1649 138
rect -1615 -138 -1609 138
rect -1655 -150 -1609 -138
rect -1559 138 -1513 150
rect -1559 -138 -1553 138
rect -1519 -138 -1513 138
rect -1559 -150 -1513 -138
rect -1463 138 -1417 150
rect -1463 -138 -1457 138
rect -1423 -138 -1417 138
rect -1463 -150 -1417 -138
rect -1367 138 -1321 150
rect -1367 -138 -1361 138
rect -1327 -138 -1321 138
rect -1367 -150 -1321 -138
rect -1271 138 -1225 150
rect -1271 -138 -1265 138
rect -1231 -138 -1225 138
rect -1271 -150 -1225 -138
rect -1175 138 -1129 150
rect -1175 -138 -1169 138
rect -1135 -138 -1129 138
rect -1175 -150 -1129 -138
rect -1079 138 -1033 150
rect -1079 -138 -1073 138
rect -1039 -138 -1033 138
rect -1079 -150 -1033 -138
rect -983 138 -937 150
rect -983 -138 -977 138
rect -943 -138 -937 138
rect -983 -150 -937 -138
rect -887 138 -841 150
rect -887 -138 -881 138
rect -847 -138 -841 138
rect -887 -150 -841 -138
rect -791 138 -745 150
rect -791 -138 -785 138
rect -751 -138 -745 138
rect -791 -150 -745 -138
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
rect 745 138 791 150
rect 745 -138 751 138
rect 785 -138 791 138
rect 745 -150 791 -138
rect 841 138 887 150
rect 841 -138 847 138
rect 881 -138 887 138
rect 841 -150 887 -138
rect 937 138 983 150
rect 937 -138 943 138
rect 977 -138 983 138
rect 937 -150 983 -138
rect 1033 138 1079 150
rect 1033 -138 1039 138
rect 1073 -138 1079 138
rect 1033 -150 1079 -138
rect 1129 138 1175 150
rect 1129 -138 1135 138
rect 1169 -138 1175 138
rect 1129 -150 1175 -138
rect 1225 138 1271 150
rect 1225 -138 1231 138
rect 1265 -138 1271 138
rect 1225 -150 1271 -138
rect 1321 138 1367 150
rect 1321 -138 1327 138
rect 1361 -138 1367 138
rect 1321 -150 1367 -138
rect 1417 138 1463 150
rect 1417 -138 1423 138
rect 1457 -138 1463 138
rect 1417 -150 1463 -138
rect 1513 138 1559 150
rect 1513 -138 1519 138
rect 1553 -138 1559 138
rect 1513 -150 1559 -138
rect 1609 138 1655 150
rect 1609 -138 1615 138
rect 1649 -138 1655 138
rect 1609 -150 1655 -138
rect 1705 138 1751 150
rect 1705 -138 1711 138
rect 1745 -138 1751 138
rect 1705 -150 1751 -138
rect 1801 138 1847 150
rect 1801 -138 1807 138
rect 1841 -138 1847 138
rect 1801 -150 1847 -138
rect 1897 138 1943 150
rect 1897 -138 1903 138
rect 1937 -138 1943 138
rect 1897 -150 1943 -138
rect 1993 138 2039 150
rect 1993 -138 1999 138
rect 2033 -138 2039 138
rect 1993 -150 2039 -138
rect 2089 138 2135 150
rect 2089 -138 2095 138
rect 2129 -138 2135 138
rect 2089 -150 2135 -138
rect 2185 138 2231 150
rect 2185 -138 2191 138
rect 2225 -138 2231 138
rect 2185 -150 2231 -138
rect 2281 138 2327 150
rect 2281 -138 2287 138
rect 2321 -138 2327 138
rect 2281 -150 2327 -138
rect 2377 138 2423 150
rect 2377 -138 2383 138
rect 2417 -138 2423 138
rect 2377 -150 2423 -138
rect 2473 138 2519 150
rect 2473 -138 2479 138
rect 2513 -138 2519 138
rect 2473 -150 2519 -138
rect 2569 138 2615 150
rect 2569 -138 2575 138
rect 2609 -138 2615 138
rect 2569 -150 2615 -138
rect 2665 138 2711 150
rect 2665 -138 2671 138
rect 2705 -138 2711 138
rect 2665 -150 2711 -138
rect 2761 138 2807 150
rect 2761 -138 2767 138
rect 2801 -138 2807 138
rect 2761 -150 2807 -138
rect 2857 138 2903 150
rect 2857 -138 2863 138
rect 2897 -138 2903 138
rect 2857 -150 2903 -138
rect 2953 138 2999 150
rect 2953 -138 2959 138
rect 2993 -138 2999 138
rect 2953 -150 2999 -138
rect 3049 138 3095 150
rect 3049 -138 3055 138
rect 3089 -138 3095 138
rect 3049 -150 3095 -138
rect 3145 138 3191 150
rect 3145 -138 3151 138
rect 3185 -138 3191 138
rect 3145 -150 3191 -138
rect 3241 138 3287 150
rect 3241 -138 3247 138
rect 3281 -138 3287 138
rect 3241 -150 3287 -138
rect 3337 138 3383 150
rect 3337 -138 3343 138
rect 3377 -138 3383 138
rect 3337 -150 3383 -138
rect 3433 138 3479 150
rect 3433 -138 3439 138
rect 3473 -138 3479 138
rect 3433 -150 3479 -138
rect 3529 138 3575 150
rect 3529 -138 3535 138
rect 3569 -138 3575 138
rect 3529 -150 3575 -138
rect 3625 138 3671 150
rect 3625 -138 3631 138
rect 3665 -138 3671 138
rect 3625 -150 3671 -138
rect 3721 138 3767 150
rect 3721 -138 3727 138
rect 3761 -138 3767 138
rect 3721 -150 3767 -138
rect 3817 138 3863 150
rect 3817 -138 3823 138
rect 3857 -138 3863 138
rect 3817 -150 3863 -138
rect 3913 138 3959 150
rect 3913 -138 3919 138
rect 3953 -138 3959 138
rect 3913 -150 3959 -138
rect 4009 138 4055 150
rect 4009 -138 4015 138
rect 4049 -138 4055 138
rect 4009 -150 4055 -138
rect 4105 138 4151 150
rect 4105 -138 4111 138
rect 4145 -138 4151 138
rect 4105 -150 4151 -138
rect 4201 138 4247 150
rect 4201 -138 4207 138
rect 4241 -138 4247 138
rect 4201 -150 4247 -138
rect 4297 138 4343 150
rect 4297 -138 4303 138
rect 4337 -138 4343 138
rect 4297 -150 4343 -138
rect 4393 138 4439 150
rect 4393 -138 4399 138
rect 4433 -138 4439 138
rect 4393 -150 4439 -138
rect 4489 138 4535 150
rect 4489 -138 4495 138
rect 4529 -138 4535 138
rect 4489 -150 4535 -138
rect 4585 138 4631 150
rect 4585 -138 4591 138
rect 4625 -138 4631 138
rect 4585 -150 4631 -138
rect 4681 138 4727 150
rect 4681 -138 4687 138
rect 4721 -138 4727 138
rect 4681 -150 4727 -138
rect 4777 138 4823 150
rect 4777 -138 4783 138
rect 4817 -138 4823 138
rect 4777 -150 4823 -138
rect 4873 138 4919 150
rect 4873 -138 4879 138
rect 4913 -138 4919 138
rect 4873 -150 4919 -138
rect 4969 138 5015 150
rect 4969 -138 4975 138
rect 5009 -138 5015 138
rect 4969 -150 5015 -138
rect 5065 138 5111 150
rect 5065 -138 5071 138
rect 5105 -138 5111 138
rect 5065 -150 5111 -138
rect 5161 138 5207 150
rect 5161 -138 5167 138
rect 5201 -138 5207 138
rect 5161 -150 5207 -138
rect 5257 138 5303 150
rect 5257 -138 5263 138
rect 5297 -138 5303 138
rect 5257 -150 5303 -138
rect 5353 138 5399 150
rect 5353 -138 5359 138
rect 5393 -138 5399 138
rect 5353 -150 5399 -138
rect 5449 138 5495 150
rect 5449 -138 5455 138
rect 5489 -138 5495 138
rect 5449 -150 5495 -138
rect 5545 138 5591 150
rect 5545 -138 5551 138
rect 5585 -138 5591 138
rect 5545 -150 5591 -138
rect 5641 138 5687 150
rect 5641 -138 5647 138
rect 5681 -138 5687 138
rect 5641 -150 5687 -138
rect 5737 138 5783 150
rect 5737 -138 5743 138
rect 5777 -138 5783 138
rect 5737 -150 5783 -138
rect 5833 138 5879 150
rect 5833 -138 5839 138
rect 5873 -138 5879 138
rect 5833 -150 5879 -138
rect 5929 138 5975 150
rect 5929 -138 5935 138
rect 5969 -138 5975 138
rect 5929 -150 5975 -138
rect 6025 138 6071 150
rect 6025 -138 6031 138
rect 6065 -138 6071 138
rect 6025 -150 6071 -138
rect 6121 138 6167 150
rect 6121 -138 6127 138
rect 6161 -138 6167 138
rect 6121 -150 6167 -138
rect 6217 138 6263 150
rect 6217 -138 6223 138
rect 6257 -138 6263 138
rect 6217 -150 6263 -138
rect 6313 138 6359 150
rect 6313 -138 6319 138
rect 6353 -138 6359 138
rect 6313 -150 6359 -138
rect 6409 138 6455 150
rect 6409 -138 6415 138
rect 6449 -138 6455 138
rect 6409 -150 6455 -138
rect 6505 138 6551 150
rect 6505 -138 6511 138
rect 6545 -138 6551 138
rect 6505 -150 6551 -138
rect 6601 138 6647 150
rect 6601 -138 6607 138
rect 6641 -138 6647 138
rect 6601 -150 6647 -138
rect 6697 138 6743 150
rect 6697 -138 6703 138
rect 6737 -138 6743 138
rect 6697 -150 6743 -138
rect 6793 138 6839 150
rect 6793 -138 6799 138
rect 6833 -138 6839 138
rect 6793 -150 6839 -138
rect 6889 138 6935 150
rect 6889 -138 6895 138
rect 6929 -138 6935 138
rect 6889 -150 6935 -138
rect 6985 138 7031 150
rect 6985 -138 6991 138
rect 7025 -138 7031 138
rect 6985 -150 7031 -138
rect 7081 138 7127 150
rect 7081 -138 7087 138
rect 7121 -138 7127 138
rect 7081 -150 7127 -138
rect 7177 138 7223 150
rect 7177 -138 7183 138
rect 7217 -138 7223 138
rect 7177 -150 7223 -138
rect 7273 138 7319 150
rect 7273 -138 7279 138
rect 7313 -138 7319 138
rect 7273 -150 7319 -138
rect 7369 138 7415 150
rect 7369 -138 7375 138
rect 7409 -138 7415 138
rect 7369 -150 7415 -138
rect 7465 138 7511 150
rect 7465 -138 7471 138
rect 7505 -138 7511 138
rect 7465 -150 7511 -138
rect 7561 138 7607 150
rect 7561 -138 7567 138
rect 7601 -138 7607 138
rect 7561 -150 7607 -138
rect 7657 138 7703 150
rect 7657 -138 7663 138
rect 7697 -138 7703 138
rect 7657 -150 7703 -138
rect 7753 138 7799 150
rect 7753 -138 7759 138
rect 7793 -138 7799 138
rect 7753 -150 7799 -138
rect 7849 138 7895 150
rect 7849 -138 7855 138
rect 7889 -138 7895 138
rect 7849 -150 7895 -138
rect 7945 138 7991 150
rect 7945 -138 7951 138
rect 7985 -138 7991 138
rect 7945 -150 7991 -138
rect 8041 138 8087 150
rect 8041 -138 8047 138
rect 8081 -138 8087 138
rect 8041 -150 8087 -138
rect 8137 138 8183 150
rect 8137 -138 8143 138
rect 8177 -138 8183 138
rect 8137 -150 8183 -138
rect 8233 138 8279 150
rect 8233 -138 8239 138
rect 8273 -138 8279 138
rect 8233 -150 8279 -138
rect 8329 138 8375 150
rect 8329 -138 8335 138
rect 8369 -138 8375 138
rect 8329 -150 8375 -138
rect 8425 138 8471 150
rect 8425 -138 8431 138
rect 8465 -138 8471 138
rect 8425 -150 8471 -138
rect 8521 138 8567 150
rect 8521 -138 8527 138
rect 8561 -138 8567 138
rect 8521 -150 8567 -138
rect 8617 138 8663 150
rect 8617 -138 8623 138
rect 8657 -138 8663 138
rect 8617 -150 8663 -138
rect 8713 138 8759 150
rect 8713 -138 8719 138
rect 8753 -138 8759 138
rect 8713 -150 8759 -138
rect 8809 138 8855 150
rect 8809 -138 8815 138
rect 8849 -138 8855 138
rect 8809 -150 8855 -138
rect 8905 138 8951 150
rect 8905 -138 8911 138
rect 8945 -138 8951 138
rect 8905 -150 8951 -138
rect 9001 138 9047 150
rect 9001 -138 9007 138
rect 9041 -138 9047 138
rect 9001 -150 9047 -138
rect 9097 138 9143 150
rect 9097 -138 9103 138
rect 9137 -138 9143 138
rect 9097 -150 9143 -138
rect 9193 138 9239 150
rect 9193 -138 9199 138
rect 9233 -138 9239 138
rect 9193 -150 9239 -138
rect 9289 138 9335 150
rect 9289 -138 9295 138
rect 9329 -138 9335 138
rect 9289 -150 9335 -138
rect 9385 138 9431 150
rect 9385 -138 9391 138
rect 9425 -138 9431 138
rect 9385 -150 9431 -138
rect 9481 138 9527 150
rect 9481 -138 9487 138
rect 9521 -138 9527 138
rect 9481 -150 9527 -138
rect 9577 138 9623 150
rect 9577 -138 9583 138
rect 9617 -138 9623 138
rect 9577 -150 9623 -138
rect 9673 138 9719 150
rect 9673 -138 9679 138
rect 9713 -138 9719 138
rect 9673 -150 9719 -138
rect 9769 138 9815 150
rect 9769 -138 9775 138
rect 9809 -138 9815 138
rect 9769 -150 9815 -138
rect 9865 138 9911 150
rect 9865 -138 9871 138
rect 9905 -138 9911 138
rect 9865 -150 9911 -138
rect 9961 138 10007 150
rect 9961 -138 9967 138
rect 10001 -138 10007 138
rect 9961 -150 10007 -138
rect 10057 138 10103 150
rect 10057 -138 10063 138
rect 10097 -138 10103 138
rect 10057 -150 10103 -138
rect 10153 138 10199 150
rect 10153 -138 10159 138
rect 10193 -138 10199 138
rect 10153 -150 10199 -138
rect 10249 138 10295 150
rect 10249 -138 10255 138
rect 10289 -138 10295 138
rect 10249 -150 10295 -138
rect 10345 138 10391 150
rect 10345 -138 10351 138
rect 10385 -138 10391 138
rect 10345 -150 10391 -138
rect 10441 138 10487 150
rect 10441 -138 10447 138
rect 10481 -138 10487 138
rect 10441 -150 10487 -138
rect 10537 138 10583 150
rect 10537 -138 10543 138
rect 10577 -138 10583 138
rect 10537 -150 10583 -138
rect 10633 138 10679 150
rect 10633 -138 10639 138
rect 10673 -138 10679 138
rect 10633 -150 10679 -138
rect 10729 138 10775 150
rect 10729 -138 10735 138
rect 10769 -138 10775 138
rect 10729 -150 10775 -138
rect 10825 138 10871 150
rect 10825 -138 10831 138
rect 10865 -138 10871 138
rect 10825 -150 10871 -138
rect 10921 138 10967 150
rect 10921 -138 10927 138
rect 10961 -138 10967 138
rect 10921 -150 10967 -138
rect 11017 138 11063 150
rect 11017 -138 11023 138
rect 11057 -138 11063 138
rect 11017 -150 11063 -138
rect 11113 138 11159 150
rect 11113 -138 11119 138
rect 11153 -138 11159 138
rect 11113 -150 11159 -138
rect 11209 138 11255 150
rect 11209 -138 11215 138
rect 11249 -138 11255 138
rect 11209 -150 11255 -138
rect 11305 138 11351 150
rect 11305 -138 11311 138
rect 11345 -138 11351 138
rect 11305 -150 11351 -138
rect 11401 138 11447 150
rect 11401 -138 11407 138
rect 11441 -138 11447 138
rect 11401 -150 11447 -138
rect 11497 138 11543 150
rect 11497 -138 11503 138
rect 11537 -138 11543 138
rect 11497 -150 11543 -138
rect 11593 138 11639 150
rect 11593 -138 11599 138
rect 11633 -138 11639 138
rect 11593 -150 11639 -138
rect 11689 138 11735 150
rect 11689 -138 11695 138
rect 11729 -138 11735 138
rect 11689 -150 11735 -138
rect 11785 138 11831 150
rect 11785 -138 11791 138
rect 11825 -138 11831 138
rect 11785 -150 11831 -138
rect 11881 138 11927 150
rect 11881 -138 11887 138
rect 11921 -138 11927 138
rect 11881 -150 11927 -138
rect 11977 138 12023 150
rect 11977 -138 11983 138
rect 12017 -138 12023 138
rect 11977 -150 12023 -138
rect 12073 138 12119 150
rect 12073 -138 12079 138
rect 12113 -138 12119 138
rect 12073 -150 12119 -138
rect 12169 138 12215 150
rect 12169 -138 12175 138
rect 12209 -138 12215 138
rect 12169 -150 12215 -138
rect 12265 138 12311 150
rect 12265 -138 12271 138
rect 12305 -138 12311 138
rect 12265 -150 12311 -138
rect 12361 138 12407 150
rect 12361 -138 12367 138
rect 12401 -138 12407 138
rect 12361 -150 12407 -138
rect 12457 138 12503 150
rect 12457 -138 12463 138
rect 12497 -138 12503 138
rect 12457 -150 12503 -138
rect 12553 138 12599 150
rect 12553 -138 12559 138
rect 12593 -138 12599 138
rect 12553 -150 12599 -138
rect 12649 138 12695 150
rect 12649 -138 12655 138
rect 12689 -138 12695 138
rect 12649 -150 12695 -138
rect 12745 138 12791 150
rect 12745 -138 12751 138
rect 12785 -138 12791 138
rect 12745 -150 12791 -138
rect 12841 138 12887 150
rect 12841 -138 12847 138
rect 12881 -138 12887 138
rect 12841 -150 12887 -138
rect 12937 138 12983 150
rect 12937 -138 12943 138
rect 12977 -138 12983 138
rect 12937 -150 12983 -138
rect 13033 138 13079 150
rect 13033 -138 13039 138
rect 13073 -138 13079 138
rect 13033 -150 13079 -138
rect 13129 138 13175 150
rect 13129 -138 13135 138
rect 13169 -138 13175 138
rect 13129 -150 13175 -138
rect 13225 138 13271 150
rect 13225 -138 13231 138
rect 13265 -138 13271 138
rect 13225 -150 13271 -138
rect 13321 138 13367 150
rect 13321 -138 13327 138
rect 13361 -138 13367 138
rect 13321 -150 13367 -138
rect 13417 138 13463 150
rect 13417 -138 13423 138
rect 13457 -138 13463 138
rect 13417 -150 13463 -138
rect 13513 138 13559 150
rect 13513 -138 13519 138
rect 13553 -138 13559 138
rect 13513 -150 13559 -138
rect 13609 138 13655 150
rect 13609 -138 13615 138
rect 13649 -138 13655 138
rect 13609 -150 13655 -138
rect 13705 138 13751 150
rect 13705 -138 13711 138
rect 13745 -138 13751 138
rect 13705 -150 13751 -138
rect 13801 138 13847 150
rect 13801 -138 13807 138
rect 13841 -138 13847 138
rect 13801 -150 13847 -138
rect 13897 138 13943 150
rect 13897 -138 13903 138
rect 13937 -138 13943 138
rect 13897 -150 13943 -138
rect 13993 138 14039 150
rect 13993 -138 13999 138
rect 14033 -138 14039 138
rect 13993 -150 14039 -138
rect 14089 138 14135 150
rect 14089 -138 14095 138
rect 14129 -138 14135 138
rect 14089 -150 14135 -138
rect 14185 138 14231 150
rect 14185 -138 14191 138
rect 14225 -138 14231 138
rect 14185 -150 14231 -138
rect 14281 138 14327 150
rect 14281 -138 14287 138
rect 14321 -138 14327 138
rect 14281 -150 14327 -138
rect 14377 138 14423 150
rect 14377 -138 14383 138
rect 14417 -138 14423 138
rect 14377 -150 14423 -138
rect 14473 138 14519 150
rect 14473 -138 14479 138
rect 14513 -138 14519 138
rect 14473 -150 14519 -138
rect 14569 138 14615 150
rect 14569 -138 14575 138
rect 14609 -138 14615 138
rect 14569 -150 14615 -138
rect 14665 138 14711 150
rect 14665 -138 14671 138
rect 14705 -138 14711 138
rect 14665 -150 14711 -138
rect 14761 138 14807 150
rect 14761 -138 14767 138
rect 14801 -138 14807 138
rect 14761 -150 14807 -138
rect 14857 138 14903 150
rect 14857 -138 14863 138
rect 14897 -138 14903 138
rect 14857 -150 14903 -138
rect 14953 138 14999 150
rect 14953 -138 14959 138
rect 14993 -138 14999 138
rect 14953 -150 14999 -138
rect 15049 138 15095 150
rect 15049 -138 15055 138
rect 15089 -138 15095 138
rect 15049 -150 15095 -138
rect 15145 138 15191 150
rect 15145 -138 15151 138
rect 15185 -138 15191 138
rect 15145 -150 15191 -138
rect 15241 138 15287 150
rect 15241 -138 15247 138
rect 15281 -138 15287 138
rect 15241 -150 15287 -138
rect 15337 138 15383 150
rect 15337 -138 15343 138
rect 15377 -138 15383 138
rect 15337 -150 15383 -138
rect 15433 138 15479 150
rect 15433 -138 15439 138
rect 15473 -138 15479 138
rect 15433 -150 15479 -138
rect 15529 138 15575 150
rect 15529 -138 15535 138
rect 15569 -138 15575 138
rect 15529 -150 15575 -138
rect 15625 138 15671 150
rect 15625 -138 15631 138
rect 15665 -138 15671 138
rect 15625 -150 15671 -138
rect 15721 138 15767 150
rect 15721 -138 15727 138
rect 15761 -138 15767 138
rect 15721 -150 15767 -138
rect 15817 138 15863 150
rect 15817 -138 15823 138
rect 15857 -138 15863 138
rect 15817 -150 15863 -138
rect 15913 138 15959 150
rect 15913 -138 15919 138
rect 15953 -138 15959 138
rect 15913 -150 15959 -138
rect 16009 138 16055 150
rect 16009 -138 16015 138
rect 16049 -138 16055 138
rect 16009 -150 16055 -138
rect 16105 138 16151 150
rect 16105 -138 16111 138
rect 16145 -138 16151 138
rect 16105 -150 16151 -138
rect 16201 138 16247 150
rect 16201 -138 16207 138
rect 16241 -138 16247 138
rect 16201 -150 16247 -138
rect 16297 138 16343 150
rect 16297 -138 16303 138
rect 16337 -138 16343 138
rect 16297 -150 16343 -138
rect 16393 138 16439 150
rect 16393 -138 16399 138
rect 16433 -138 16439 138
rect 16393 -150 16439 -138
rect 16489 138 16535 150
rect 16489 -138 16495 138
rect 16529 -138 16535 138
rect 16489 -150 16535 -138
rect 16585 138 16631 150
rect 16585 -138 16591 138
rect 16625 -138 16631 138
rect 16585 -150 16631 -138
rect 16681 138 16727 150
rect 16681 -138 16687 138
rect 16721 -138 16727 138
rect 16681 -150 16727 -138
rect 16777 138 16823 150
rect 16777 -138 16783 138
rect 16817 -138 16823 138
rect 16777 -150 16823 -138
rect 16873 138 16919 150
rect 16873 -138 16879 138
rect 16913 -138 16919 138
rect 16873 -150 16919 -138
rect 16969 138 17015 150
rect 16969 -138 16975 138
rect 17009 -138 17015 138
rect 16969 -150 17015 -138
rect 17065 138 17111 150
rect 17065 -138 17071 138
rect 17105 -138 17111 138
rect 17065 -150 17111 -138
rect 17161 138 17207 150
rect 17161 -138 17167 138
rect 17201 -138 17207 138
rect 17161 -150 17207 -138
rect 17257 138 17303 150
rect 17257 -138 17263 138
rect 17297 -138 17303 138
rect 17257 -150 17303 -138
rect 17353 138 17399 150
rect 17353 -138 17359 138
rect 17393 -138 17399 138
rect 17353 -150 17399 -138
rect 17449 138 17495 150
rect 17449 -138 17455 138
rect 17489 -138 17495 138
rect 17449 -150 17495 -138
rect 17545 138 17591 150
rect 17545 -138 17551 138
rect 17585 -138 17591 138
rect 17545 -150 17591 -138
rect 17641 138 17687 150
rect 17641 -138 17647 138
rect 17681 -138 17687 138
rect 17641 -150 17687 -138
rect 17737 138 17783 150
rect 17737 -138 17743 138
rect 17777 -138 17783 138
rect 17737 -150 17783 -138
rect 17833 138 17879 150
rect 17833 -138 17839 138
rect 17873 -138 17879 138
rect 17833 -150 17879 -138
rect 17929 138 17975 150
rect 17929 -138 17935 138
rect 17969 -138 17975 138
rect 17929 -150 17975 -138
rect 18025 138 18071 150
rect 18025 -138 18031 138
rect 18065 -138 18071 138
rect 18025 -150 18071 -138
rect 18121 138 18167 150
rect 18121 -138 18127 138
rect 18161 -138 18167 138
rect 18121 -150 18167 -138
rect 18217 138 18263 150
rect 18217 -138 18223 138
rect 18257 -138 18263 138
rect 18217 -150 18263 -138
rect 18313 138 18359 150
rect 18313 -138 18319 138
rect 18353 -138 18359 138
rect 18313 -150 18359 -138
rect 18409 138 18455 150
rect 18409 -138 18415 138
rect 18449 -138 18455 138
rect 18409 -150 18455 -138
rect 18505 138 18551 150
rect 18505 -138 18511 138
rect 18545 -138 18551 138
rect 18505 -150 18551 -138
rect 18601 138 18647 150
rect 18601 -138 18607 138
rect 18641 -138 18647 138
rect 18601 -150 18647 -138
rect 18697 138 18743 150
rect 18697 -138 18703 138
rect 18737 -138 18743 138
rect 18697 -150 18743 -138
rect 18793 138 18839 150
rect 18793 -138 18799 138
rect 18833 -138 18839 138
rect 18793 -150 18839 -138
rect 18889 138 18935 150
rect 18889 -138 18895 138
rect 18929 -138 18935 138
rect 18889 -150 18935 -138
rect 18985 138 19031 150
rect 18985 -138 18991 138
rect 19025 -138 19031 138
rect 18985 -150 19031 -138
rect 19081 138 19127 150
rect 19081 -138 19087 138
rect 19121 -138 19127 138
rect 19081 -150 19127 -138
rect 19177 138 19223 150
rect 19177 -138 19183 138
rect 19217 -138 19223 138
rect 19177 -150 19223 -138
rect -19181 -188 -19123 -182
rect -19181 -222 -19169 -188
rect -19135 -222 -19123 -188
rect -19181 -228 -19123 -222
rect -18989 -188 -18931 -182
rect -18989 -222 -18977 -188
rect -18943 -222 -18931 -188
rect -18989 -228 -18931 -222
rect -18797 -188 -18739 -182
rect -18797 -222 -18785 -188
rect -18751 -222 -18739 -188
rect -18797 -228 -18739 -222
rect -18605 -188 -18547 -182
rect -18605 -222 -18593 -188
rect -18559 -222 -18547 -188
rect -18605 -228 -18547 -222
rect -18413 -188 -18355 -182
rect -18413 -222 -18401 -188
rect -18367 -222 -18355 -188
rect -18413 -228 -18355 -222
rect -18221 -188 -18163 -182
rect -18221 -222 -18209 -188
rect -18175 -222 -18163 -188
rect -18221 -228 -18163 -222
rect -18029 -188 -17971 -182
rect -18029 -222 -18017 -188
rect -17983 -222 -17971 -188
rect -18029 -228 -17971 -222
rect -17837 -188 -17779 -182
rect -17837 -222 -17825 -188
rect -17791 -222 -17779 -188
rect -17837 -228 -17779 -222
rect -17645 -188 -17587 -182
rect -17645 -222 -17633 -188
rect -17599 -222 -17587 -188
rect -17645 -228 -17587 -222
rect -17453 -188 -17395 -182
rect -17453 -222 -17441 -188
rect -17407 -222 -17395 -188
rect -17453 -228 -17395 -222
rect -17261 -188 -17203 -182
rect -17261 -222 -17249 -188
rect -17215 -222 -17203 -188
rect -17261 -228 -17203 -222
rect -17069 -188 -17011 -182
rect -17069 -222 -17057 -188
rect -17023 -222 -17011 -188
rect -17069 -228 -17011 -222
rect -16877 -188 -16819 -182
rect -16877 -222 -16865 -188
rect -16831 -222 -16819 -188
rect -16877 -228 -16819 -222
rect -16685 -188 -16627 -182
rect -16685 -222 -16673 -188
rect -16639 -222 -16627 -188
rect -16685 -228 -16627 -222
rect -16493 -188 -16435 -182
rect -16493 -222 -16481 -188
rect -16447 -222 -16435 -188
rect -16493 -228 -16435 -222
rect -16301 -188 -16243 -182
rect -16301 -222 -16289 -188
rect -16255 -222 -16243 -188
rect -16301 -228 -16243 -222
rect -16109 -188 -16051 -182
rect -16109 -222 -16097 -188
rect -16063 -222 -16051 -188
rect -16109 -228 -16051 -222
rect -15917 -188 -15859 -182
rect -15917 -222 -15905 -188
rect -15871 -222 -15859 -188
rect -15917 -228 -15859 -222
rect -15725 -188 -15667 -182
rect -15725 -222 -15713 -188
rect -15679 -222 -15667 -188
rect -15725 -228 -15667 -222
rect -15533 -188 -15475 -182
rect -15533 -222 -15521 -188
rect -15487 -222 -15475 -188
rect -15533 -228 -15475 -222
rect -15341 -188 -15283 -182
rect -15341 -222 -15329 -188
rect -15295 -222 -15283 -188
rect -15341 -228 -15283 -222
rect -15149 -188 -15091 -182
rect -15149 -222 -15137 -188
rect -15103 -222 -15091 -188
rect -15149 -228 -15091 -222
rect -14957 -188 -14899 -182
rect -14957 -222 -14945 -188
rect -14911 -222 -14899 -188
rect -14957 -228 -14899 -222
rect -14765 -188 -14707 -182
rect -14765 -222 -14753 -188
rect -14719 -222 -14707 -188
rect -14765 -228 -14707 -222
rect -14573 -188 -14515 -182
rect -14573 -222 -14561 -188
rect -14527 -222 -14515 -188
rect -14573 -228 -14515 -222
rect -14381 -188 -14323 -182
rect -14381 -222 -14369 -188
rect -14335 -222 -14323 -188
rect -14381 -228 -14323 -222
rect -14189 -188 -14131 -182
rect -14189 -222 -14177 -188
rect -14143 -222 -14131 -188
rect -14189 -228 -14131 -222
rect -13997 -188 -13939 -182
rect -13997 -222 -13985 -188
rect -13951 -222 -13939 -188
rect -13997 -228 -13939 -222
rect -13805 -188 -13747 -182
rect -13805 -222 -13793 -188
rect -13759 -222 -13747 -188
rect -13805 -228 -13747 -222
rect -13613 -188 -13555 -182
rect -13613 -222 -13601 -188
rect -13567 -222 -13555 -188
rect -13613 -228 -13555 -222
rect -13421 -188 -13363 -182
rect -13421 -222 -13409 -188
rect -13375 -222 -13363 -188
rect -13421 -228 -13363 -222
rect -13229 -188 -13171 -182
rect -13229 -222 -13217 -188
rect -13183 -222 -13171 -188
rect -13229 -228 -13171 -222
rect -13037 -188 -12979 -182
rect -13037 -222 -13025 -188
rect -12991 -222 -12979 -188
rect -13037 -228 -12979 -222
rect -12845 -188 -12787 -182
rect -12845 -222 -12833 -188
rect -12799 -222 -12787 -188
rect -12845 -228 -12787 -222
rect -12653 -188 -12595 -182
rect -12653 -222 -12641 -188
rect -12607 -222 -12595 -188
rect -12653 -228 -12595 -222
rect -12461 -188 -12403 -182
rect -12461 -222 -12449 -188
rect -12415 -222 -12403 -188
rect -12461 -228 -12403 -222
rect -12269 -188 -12211 -182
rect -12269 -222 -12257 -188
rect -12223 -222 -12211 -188
rect -12269 -228 -12211 -222
rect -12077 -188 -12019 -182
rect -12077 -222 -12065 -188
rect -12031 -222 -12019 -188
rect -12077 -228 -12019 -222
rect -11885 -188 -11827 -182
rect -11885 -222 -11873 -188
rect -11839 -222 -11827 -188
rect -11885 -228 -11827 -222
rect -11693 -188 -11635 -182
rect -11693 -222 -11681 -188
rect -11647 -222 -11635 -188
rect -11693 -228 -11635 -222
rect -11501 -188 -11443 -182
rect -11501 -222 -11489 -188
rect -11455 -222 -11443 -188
rect -11501 -228 -11443 -222
rect -11309 -188 -11251 -182
rect -11309 -222 -11297 -188
rect -11263 -222 -11251 -188
rect -11309 -228 -11251 -222
rect -11117 -188 -11059 -182
rect -11117 -222 -11105 -188
rect -11071 -222 -11059 -188
rect -11117 -228 -11059 -222
rect -10925 -188 -10867 -182
rect -10925 -222 -10913 -188
rect -10879 -222 -10867 -188
rect -10925 -228 -10867 -222
rect -10733 -188 -10675 -182
rect -10733 -222 -10721 -188
rect -10687 -222 -10675 -188
rect -10733 -228 -10675 -222
rect -10541 -188 -10483 -182
rect -10541 -222 -10529 -188
rect -10495 -222 -10483 -188
rect -10541 -228 -10483 -222
rect -10349 -188 -10291 -182
rect -10349 -222 -10337 -188
rect -10303 -222 -10291 -188
rect -10349 -228 -10291 -222
rect -10157 -188 -10099 -182
rect -10157 -222 -10145 -188
rect -10111 -222 -10099 -188
rect -10157 -228 -10099 -222
rect -9965 -188 -9907 -182
rect -9965 -222 -9953 -188
rect -9919 -222 -9907 -188
rect -9965 -228 -9907 -222
rect -9773 -188 -9715 -182
rect -9773 -222 -9761 -188
rect -9727 -222 -9715 -188
rect -9773 -228 -9715 -222
rect -9581 -188 -9523 -182
rect -9581 -222 -9569 -188
rect -9535 -222 -9523 -188
rect -9581 -228 -9523 -222
rect -9389 -188 -9331 -182
rect -9389 -222 -9377 -188
rect -9343 -222 -9331 -188
rect -9389 -228 -9331 -222
rect -9197 -188 -9139 -182
rect -9197 -222 -9185 -188
rect -9151 -222 -9139 -188
rect -9197 -228 -9139 -222
rect -9005 -188 -8947 -182
rect -9005 -222 -8993 -188
rect -8959 -222 -8947 -188
rect -9005 -228 -8947 -222
rect -8813 -188 -8755 -182
rect -8813 -222 -8801 -188
rect -8767 -222 -8755 -188
rect -8813 -228 -8755 -222
rect -8621 -188 -8563 -182
rect -8621 -222 -8609 -188
rect -8575 -222 -8563 -188
rect -8621 -228 -8563 -222
rect -8429 -188 -8371 -182
rect -8429 -222 -8417 -188
rect -8383 -222 -8371 -188
rect -8429 -228 -8371 -222
rect -8237 -188 -8179 -182
rect -8237 -222 -8225 -188
rect -8191 -222 -8179 -188
rect -8237 -228 -8179 -222
rect -8045 -188 -7987 -182
rect -8045 -222 -8033 -188
rect -7999 -222 -7987 -188
rect -8045 -228 -7987 -222
rect -7853 -188 -7795 -182
rect -7853 -222 -7841 -188
rect -7807 -222 -7795 -188
rect -7853 -228 -7795 -222
rect -7661 -188 -7603 -182
rect -7661 -222 -7649 -188
rect -7615 -222 -7603 -188
rect -7661 -228 -7603 -222
rect -7469 -188 -7411 -182
rect -7469 -222 -7457 -188
rect -7423 -222 -7411 -188
rect -7469 -228 -7411 -222
rect -7277 -188 -7219 -182
rect -7277 -222 -7265 -188
rect -7231 -222 -7219 -188
rect -7277 -228 -7219 -222
rect -7085 -188 -7027 -182
rect -7085 -222 -7073 -188
rect -7039 -222 -7027 -188
rect -7085 -228 -7027 -222
rect -6893 -188 -6835 -182
rect -6893 -222 -6881 -188
rect -6847 -222 -6835 -188
rect -6893 -228 -6835 -222
rect -6701 -188 -6643 -182
rect -6701 -222 -6689 -188
rect -6655 -222 -6643 -188
rect -6701 -228 -6643 -222
rect -6509 -188 -6451 -182
rect -6509 -222 -6497 -188
rect -6463 -222 -6451 -188
rect -6509 -228 -6451 -222
rect -6317 -188 -6259 -182
rect -6317 -222 -6305 -188
rect -6271 -222 -6259 -188
rect -6317 -228 -6259 -222
rect -6125 -188 -6067 -182
rect -6125 -222 -6113 -188
rect -6079 -222 -6067 -188
rect -6125 -228 -6067 -222
rect -5933 -188 -5875 -182
rect -5933 -222 -5921 -188
rect -5887 -222 -5875 -188
rect -5933 -228 -5875 -222
rect -5741 -188 -5683 -182
rect -5741 -222 -5729 -188
rect -5695 -222 -5683 -188
rect -5741 -228 -5683 -222
rect -5549 -188 -5491 -182
rect -5549 -222 -5537 -188
rect -5503 -222 -5491 -188
rect -5549 -228 -5491 -222
rect -5357 -188 -5299 -182
rect -5357 -222 -5345 -188
rect -5311 -222 -5299 -188
rect -5357 -228 -5299 -222
rect -5165 -188 -5107 -182
rect -5165 -222 -5153 -188
rect -5119 -222 -5107 -188
rect -5165 -228 -5107 -222
rect -4973 -188 -4915 -182
rect -4973 -222 -4961 -188
rect -4927 -222 -4915 -188
rect -4973 -228 -4915 -222
rect -4781 -188 -4723 -182
rect -4781 -222 -4769 -188
rect -4735 -222 -4723 -188
rect -4781 -228 -4723 -222
rect -4589 -188 -4531 -182
rect -4589 -222 -4577 -188
rect -4543 -222 -4531 -188
rect -4589 -228 -4531 -222
rect -4397 -188 -4339 -182
rect -4397 -222 -4385 -188
rect -4351 -222 -4339 -188
rect -4397 -228 -4339 -222
rect -4205 -188 -4147 -182
rect -4205 -222 -4193 -188
rect -4159 -222 -4147 -188
rect -4205 -228 -4147 -222
rect -4013 -188 -3955 -182
rect -4013 -222 -4001 -188
rect -3967 -222 -3955 -188
rect -4013 -228 -3955 -222
rect -3821 -188 -3763 -182
rect -3821 -222 -3809 -188
rect -3775 -222 -3763 -188
rect -3821 -228 -3763 -222
rect -3629 -188 -3571 -182
rect -3629 -222 -3617 -188
rect -3583 -222 -3571 -188
rect -3629 -228 -3571 -222
rect -3437 -188 -3379 -182
rect -3437 -222 -3425 -188
rect -3391 -222 -3379 -188
rect -3437 -228 -3379 -222
rect -3245 -188 -3187 -182
rect -3245 -222 -3233 -188
rect -3199 -222 -3187 -188
rect -3245 -228 -3187 -222
rect -3053 -188 -2995 -182
rect -3053 -222 -3041 -188
rect -3007 -222 -2995 -188
rect -3053 -228 -2995 -222
rect -2861 -188 -2803 -182
rect -2861 -222 -2849 -188
rect -2815 -222 -2803 -188
rect -2861 -228 -2803 -222
rect -2669 -188 -2611 -182
rect -2669 -222 -2657 -188
rect -2623 -222 -2611 -188
rect -2669 -228 -2611 -222
rect -2477 -188 -2419 -182
rect -2477 -222 -2465 -188
rect -2431 -222 -2419 -188
rect -2477 -228 -2419 -222
rect -2285 -188 -2227 -182
rect -2285 -222 -2273 -188
rect -2239 -222 -2227 -188
rect -2285 -228 -2227 -222
rect -2093 -188 -2035 -182
rect -2093 -222 -2081 -188
rect -2047 -222 -2035 -188
rect -2093 -228 -2035 -222
rect -1901 -188 -1843 -182
rect -1901 -222 -1889 -188
rect -1855 -222 -1843 -188
rect -1901 -228 -1843 -222
rect -1709 -188 -1651 -182
rect -1709 -222 -1697 -188
rect -1663 -222 -1651 -188
rect -1709 -228 -1651 -222
rect -1517 -188 -1459 -182
rect -1517 -222 -1505 -188
rect -1471 -222 -1459 -188
rect -1517 -228 -1459 -222
rect -1325 -188 -1267 -182
rect -1325 -222 -1313 -188
rect -1279 -222 -1267 -188
rect -1325 -228 -1267 -222
rect -1133 -188 -1075 -182
rect -1133 -222 -1121 -188
rect -1087 -222 -1075 -188
rect -1133 -228 -1075 -222
rect -941 -188 -883 -182
rect -941 -222 -929 -188
rect -895 -222 -883 -188
rect -941 -228 -883 -222
rect -749 -188 -691 -182
rect -749 -222 -737 -188
rect -703 -222 -691 -188
rect -749 -228 -691 -222
rect -557 -188 -499 -182
rect -557 -222 -545 -188
rect -511 -222 -499 -188
rect -557 -228 -499 -222
rect -365 -188 -307 -182
rect -365 -222 -353 -188
rect -319 -222 -307 -188
rect -365 -228 -307 -222
rect -173 -188 -115 -182
rect -173 -222 -161 -188
rect -127 -222 -115 -188
rect -173 -228 -115 -222
rect 19 -188 77 -182
rect 19 -222 31 -188
rect 65 -222 77 -188
rect 19 -228 77 -222
rect 211 -188 269 -182
rect 211 -222 223 -188
rect 257 -222 269 -188
rect 211 -228 269 -222
rect 403 -188 461 -182
rect 403 -222 415 -188
rect 449 -222 461 -188
rect 403 -228 461 -222
rect 595 -188 653 -182
rect 595 -222 607 -188
rect 641 -222 653 -188
rect 595 -228 653 -222
rect 787 -188 845 -182
rect 787 -222 799 -188
rect 833 -222 845 -188
rect 787 -228 845 -222
rect 979 -188 1037 -182
rect 979 -222 991 -188
rect 1025 -222 1037 -188
rect 979 -228 1037 -222
rect 1171 -188 1229 -182
rect 1171 -222 1183 -188
rect 1217 -222 1229 -188
rect 1171 -228 1229 -222
rect 1363 -188 1421 -182
rect 1363 -222 1375 -188
rect 1409 -222 1421 -188
rect 1363 -228 1421 -222
rect 1555 -188 1613 -182
rect 1555 -222 1567 -188
rect 1601 -222 1613 -188
rect 1555 -228 1613 -222
rect 1747 -188 1805 -182
rect 1747 -222 1759 -188
rect 1793 -222 1805 -188
rect 1747 -228 1805 -222
rect 1939 -188 1997 -182
rect 1939 -222 1951 -188
rect 1985 -222 1997 -188
rect 1939 -228 1997 -222
rect 2131 -188 2189 -182
rect 2131 -222 2143 -188
rect 2177 -222 2189 -188
rect 2131 -228 2189 -222
rect 2323 -188 2381 -182
rect 2323 -222 2335 -188
rect 2369 -222 2381 -188
rect 2323 -228 2381 -222
rect 2515 -188 2573 -182
rect 2515 -222 2527 -188
rect 2561 -222 2573 -188
rect 2515 -228 2573 -222
rect 2707 -188 2765 -182
rect 2707 -222 2719 -188
rect 2753 -222 2765 -188
rect 2707 -228 2765 -222
rect 2899 -188 2957 -182
rect 2899 -222 2911 -188
rect 2945 -222 2957 -188
rect 2899 -228 2957 -222
rect 3091 -188 3149 -182
rect 3091 -222 3103 -188
rect 3137 -222 3149 -188
rect 3091 -228 3149 -222
rect 3283 -188 3341 -182
rect 3283 -222 3295 -188
rect 3329 -222 3341 -188
rect 3283 -228 3341 -222
rect 3475 -188 3533 -182
rect 3475 -222 3487 -188
rect 3521 -222 3533 -188
rect 3475 -228 3533 -222
rect 3667 -188 3725 -182
rect 3667 -222 3679 -188
rect 3713 -222 3725 -188
rect 3667 -228 3725 -222
rect 3859 -188 3917 -182
rect 3859 -222 3871 -188
rect 3905 -222 3917 -188
rect 3859 -228 3917 -222
rect 4051 -188 4109 -182
rect 4051 -222 4063 -188
rect 4097 -222 4109 -188
rect 4051 -228 4109 -222
rect 4243 -188 4301 -182
rect 4243 -222 4255 -188
rect 4289 -222 4301 -188
rect 4243 -228 4301 -222
rect 4435 -188 4493 -182
rect 4435 -222 4447 -188
rect 4481 -222 4493 -188
rect 4435 -228 4493 -222
rect 4627 -188 4685 -182
rect 4627 -222 4639 -188
rect 4673 -222 4685 -188
rect 4627 -228 4685 -222
rect 4819 -188 4877 -182
rect 4819 -222 4831 -188
rect 4865 -222 4877 -188
rect 4819 -228 4877 -222
rect 5011 -188 5069 -182
rect 5011 -222 5023 -188
rect 5057 -222 5069 -188
rect 5011 -228 5069 -222
rect 5203 -188 5261 -182
rect 5203 -222 5215 -188
rect 5249 -222 5261 -188
rect 5203 -228 5261 -222
rect 5395 -188 5453 -182
rect 5395 -222 5407 -188
rect 5441 -222 5453 -188
rect 5395 -228 5453 -222
rect 5587 -188 5645 -182
rect 5587 -222 5599 -188
rect 5633 -222 5645 -188
rect 5587 -228 5645 -222
rect 5779 -188 5837 -182
rect 5779 -222 5791 -188
rect 5825 -222 5837 -188
rect 5779 -228 5837 -222
rect 5971 -188 6029 -182
rect 5971 -222 5983 -188
rect 6017 -222 6029 -188
rect 5971 -228 6029 -222
rect 6163 -188 6221 -182
rect 6163 -222 6175 -188
rect 6209 -222 6221 -188
rect 6163 -228 6221 -222
rect 6355 -188 6413 -182
rect 6355 -222 6367 -188
rect 6401 -222 6413 -188
rect 6355 -228 6413 -222
rect 6547 -188 6605 -182
rect 6547 -222 6559 -188
rect 6593 -222 6605 -188
rect 6547 -228 6605 -222
rect 6739 -188 6797 -182
rect 6739 -222 6751 -188
rect 6785 -222 6797 -188
rect 6739 -228 6797 -222
rect 6931 -188 6989 -182
rect 6931 -222 6943 -188
rect 6977 -222 6989 -188
rect 6931 -228 6989 -222
rect 7123 -188 7181 -182
rect 7123 -222 7135 -188
rect 7169 -222 7181 -188
rect 7123 -228 7181 -222
rect 7315 -188 7373 -182
rect 7315 -222 7327 -188
rect 7361 -222 7373 -188
rect 7315 -228 7373 -222
rect 7507 -188 7565 -182
rect 7507 -222 7519 -188
rect 7553 -222 7565 -188
rect 7507 -228 7565 -222
rect 7699 -188 7757 -182
rect 7699 -222 7711 -188
rect 7745 -222 7757 -188
rect 7699 -228 7757 -222
rect 7891 -188 7949 -182
rect 7891 -222 7903 -188
rect 7937 -222 7949 -188
rect 7891 -228 7949 -222
rect 8083 -188 8141 -182
rect 8083 -222 8095 -188
rect 8129 -222 8141 -188
rect 8083 -228 8141 -222
rect 8275 -188 8333 -182
rect 8275 -222 8287 -188
rect 8321 -222 8333 -188
rect 8275 -228 8333 -222
rect 8467 -188 8525 -182
rect 8467 -222 8479 -188
rect 8513 -222 8525 -188
rect 8467 -228 8525 -222
rect 8659 -188 8717 -182
rect 8659 -222 8671 -188
rect 8705 -222 8717 -188
rect 8659 -228 8717 -222
rect 8851 -188 8909 -182
rect 8851 -222 8863 -188
rect 8897 -222 8909 -188
rect 8851 -228 8909 -222
rect 9043 -188 9101 -182
rect 9043 -222 9055 -188
rect 9089 -222 9101 -188
rect 9043 -228 9101 -222
rect 9235 -188 9293 -182
rect 9235 -222 9247 -188
rect 9281 -222 9293 -188
rect 9235 -228 9293 -222
rect 9427 -188 9485 -182
rect 9427 -222 9439 -188
rect 9473 -222 9485 -188
rect 9427 -228 9485 -222
rect 9619 -188 9677 -182
rect 9619 -222 9631 -188
rect 9665 -222 9677 -188
rect 9619 -228 9677 -222
rect 9811 -188 9869 -182
rect 9811 -222 9823 -188
rect 9857 -222 9869 -188
rect 9811 -228 9869 -222
rect 10003 -188 10061 -182
rect 10003 -222 10015 -188
rect 10049 -222 10061 -188
rect 10003 -228 10061 -222
rect 10195 -188 10253 -182
rect 10195 -222 10207 -188
rect 10241 -222 10253 -188
rect 10195 -228 10253 -222
rect 10387 -188 10445 -182
rect 10387 -222 10399 -188
rect 10433 -222 10445 -188
rect 10387 -228 10445 -222
rect 10579 -188 10637 -182
rect 10579 -222 10591 -188
rect 10625 -222 10637 -188
rect 10579 -228 10637 -222
rect 10771 -188 10829 -182
rect 10771 -222 10783 -188
rect 10817 -222 10829 -188
rect 10771 -228 10829 -222
rect 10963 -188 11021 -182
rect 10963 -222 10975 -188
rect 11009 -222 11021 -188
rect 10963 -228 11021 -222
rect 11155 -188 11213 -182
rect 11155 -222 11167 -188
rect 11201 -222 11213 -188
rect 11155 -228 11213 -222
rect 11347 -188 11405 -182
rect 11347 -222 11359 -188
rect 11393 -222 11405 -188
rect 11347 -228 11405 -222
rect 11539 -188 11597 -182
rect 11539 -222 11551 -188
rect 11585 -222 11597 -188
rect 11539 -228 11597 -222
rect 11731 -188 11789 -182
rect 11731 -222 11743 -188
rect 11777 -222 11789 -188
rect 11731 -228 11789 -222
rect 11923 -188 11981 -182
rect 11923 -222 11935 -188
rect 11969 -222 11981 -188
rect 11923 -228 11981 -222
rect 12115 -188 12173 -182
rect 12115 -222 12127 -188
rect 12161 -222 12173 -188
rect 12115 -228 12173 -222
rect 12307 -188 12365 -182
rect 12307 -222 12319 -188
rect 12353 -222 12365 -188
rect 12307 -228 12365 -222
rect 12499 -188 12557 -182
rect 12499 -222 12511 -188
rect 12545 -222 12557 -188
rect 12499 -228 12557 -222
rect 12691 -188 12749 -182
rect 12691 -222 12703 -188
rect 12737 -222 12749 -188
rect 12691 -228 12749 -222
rect 12883 -188 12941 -182
rect 12883 -222 12895 -188
rect 12929 -222 12941 -188
rect 12883 -228 12941 -222
rect 13075 -188 13133 -182
rect 13075 -222 13087 -188
rect 13121 -222 13133 -188
rect 13075 -228 13133 -222
rect 13267 -188 13325 -182
rect 13267 -222 13279 -188
rect 13313 -222 13325 -188
rect 13267 -228 13325 -222
rect 13459 -188 13517 -182
rect 13459 -222 13471 -188
rect 13505 -222 13517 -188
rect 13459 -228 13517 -222
rect 13651 -188 13709 -182
rect 13651 -222 13663 -188
rect 13697 -222 13709 -188
rect 13651 -228 13709 -222
rect 13843 -188 13901 -182
rect 13843 -222 13855 -188
rect 13889 -222 13901 -188
rect 13843 -228 13901 -222
rect 14035 -188 14093 -182
rect 14035 -222 14047 -188
rect 14081 -222 14093 -188
rect 14035 -228 14093 -222
rect 14227 -188 14285 -182
rect 14227 -222 14239 -188
rect 14273 -222 14285 -188
rect 14227 -228 14285 -222
rect 14419 -188 14477 -182
rect 14419 -222 14431 -188
rect 14465 -222 14477 -188
rect 14419 -228 14477 -222
rect 14611 -188 14669 -182
rect 14611 -222 14623 -188
rect 14657 -222 14669 -188
rect 14611 -228 14669 -222
rect 14803 -188 14861 -182
rect 14803 -222 14815 -188
rect 14849 -222 14861 -188
rect 14803 -228 14861 -222
rect 14995 -188 15053 -182
rect 14995 -222 15007 -188
rect 15041 -222 15053 -188
rect 14995 -228 15053 -222
rect 15187 -188 15245 -182
rect 15187 -222 15199 -188
rect 15233 -222 15245 -188
rect 15187 -228 15245 -222
rect 15379 -188 15437 -182
rect 15379 -222 15391 -188
rect 15425 -222 15437 -188
rect 15379 -228 15437 -222
rect 15571 -188 15629 -182
rect 15571 -222 15583 -188
rect 15617 -222 15629 -188
rect 15571 -228 15629 -222
rect 15763 -188 15821 -182
rect 15763 -222 15775 -188
rect 15809 -222 15821 -188
rect 15763 -228 15821 -222
rect 15955 -188 16013 -182
rect 15955 -222 15967 -188
rect 16001 -222 16013 -188
rect 15955 -228 16013 -222
rect 16147 -188 16205 -182
rect 16147 -222 16159 -188
rect 16193 -222 16205 -188
rect 16147 -228 16205 -222
rect 16339 -188 16397 -182
rect 16339 -222 16351 -188
rect 16385 -222 16397 -188
rect 16339 -228 16397 -222
rect 16531 -188 16589 -182
rect 16531 -222 16543 -188
rect 16577 -222 16589 -188
rect 16531 -228 16589 -222
rect 16723 -188 16781 -182
rect 16723 -222 16735 -188
rect 16769 -222 16781 -188
rect 16723 -228 16781 -222
rect 16915 -188 16973 -182
rect 16915 -222 16927 -188
rect 16961 -222 16973 -188
rect 16915 -228 16973 -222
rect 17107 -188 17165 -182
rect 17107 -222 17119 -188
rect 17153 -222 17165 -188
rect 17107 -228 17165 -222
rect 17299 -188 17357 -182
rect 17299 -222 17311 -188
rect 17345 -222 17357 -188
rect 17299 -228 17357 -222
rect 17491 -188 17549 -182
rect 17491 -222 17503 -188
rect 17537 -222 17549 -188
rect 17491 -228 17549 -222
rect 17683 -188 17741 -182
rect 17683 -222 17695 -188
rect 17729 -222 17741 -188
rect 17683 -228 17741 -222
rect 17875 -188 17933 -182
rect 17875 -222 17887 -188
rect 17921 -222 17933 -188
rect 17875 -228 17933 -222
rect 18067 -188 18125 -182
rect 18067 -222 18079 -188
rect 18113 -222 18125 -188
rect 18067 -228 18125 -222
rect 18259 -188 18317 -182
rect 18259 -222 18271 -188
rect 18305 -222 18317 -188
rect 18259 -228 18317 -222
rect 18451 -188 18509 -182
rect 18451 -222 18463 -188
rect 18497 -222 18509 -188
rect 18451 -228 18509 -222
rect 18643 -188 18701 -182
rect 18643 -222 18655 -188
rect 18689 -222 18701 -188
rect 18643 -228 18701 -222
rect 18835 -188 18893 -182
rect 18835 -222 18847 -188
rect 18881 -222 18893 -188
rect 18835 -228 18893 -222
rect 19027 -188 19085 -182
rect 19027 -222 19039 -188
rect 19073 -222 19085 -188
rect 19027 -228 19085 -222
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -19314 -307 19314 307
string parameters w 1.5 l 0.150 m 1 nf 400 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
