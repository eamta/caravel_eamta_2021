magic
tech sky130A
timestamp 1624050559
<< end >>
