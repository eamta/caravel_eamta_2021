magic
tech sky130A
magscale 1 2
timestamp 1624138001
<< error_s >>
rect 169 756 182 784
rect -591 720 -580 748
rect -544 686 -533 720
rect -472 686 -463 748
rect 216 722 229 756
rect 276 722 297 784
rect 401 756 422 784
rect 665 756 686 784
rect 448 722 469 756
rect 712 722 733 756
rect 736 722 756 756
rect 772 722 793 784
rect 1189 756 1210 784
rect 1254 766 1270 772
rect 1226 756 1280 766
rect 1455 756 1476 784
rect 1520 766 1536 772
rect 1492 756 1546 766
rect 1220 746 1286 756
rect 1220 740 1257 746
rect 1236 722 1257 740
rect 1260 740 1286 746
rect 1486 746 1552 756
rect 1486 740 1523 746
rect 1260 722 1280 740
rect 1502 722 1523 740
rect 1526 740 1552 746
rect 1526 722 1546 740
rect 1562 722 1583 784
rect 1685 756 1708 784
rect 1750 766 1766 772
rect 1722 756 1776 766
rect 1716 746 1782 756
rect 1716 740 1755 746
rect 1732 722 1755 740
rect 1756 740 1782 746
rect 1756 722 1776 740
rect 1794 722 1813 784
rect 1921 756 1940 784
rect 1986 766 2002 772
rect 1958 756 2012 766
rect 1952 746 2018 756
rect 1952 740 1987 746
rect 1968 722 1987 740
rect 1992 740 2018 746
rect 1992 722 2012 740
rect 2026 722 2049 784
rect 285 604 413 625
rect 479 594 480 636
rect 540 604 598 625
rect 1330 604 1388 625
rect 1571 604 1699 625
rect 332 578 334 588
rect 364 578 366 588
rect 332 568 344 578
rect 354 568 366 578
rect 521 578 522 594
rect 1330 588 1346 594
rect 1650 588 1652 594
rect 1302 578 1356 588
rect 1608 578 1620 588
rect 1650 578 1662 588
rect 521 554 531 578
rect 332 544 366 552
rect 521 544 533 554
rect 545 544 565 578
rect 1296 568 1362 578
rect 1296 562 1322 568
rect 1312 544 1322 562
rect 1336 562 1362 568
rect 1602 568 1630 578
rect 1640 568 1668 578
rect 1602 562 1628 568
rect 1336 544 1356 562
rect 1618 554 1628 562
rect 1642 562 1668 568
rect 1642 554 1662 562
rect 1618 544 1662 554
rect 628 510 630 516
rect 586 500 598 510
rect 628 500 640 510
rect 1344 500 1346 542
rect 1636 534 1662 544
rect 1636 528 1652 534
rect 1418 510 1420 516
rect 1636 510 1652 516
rect 1376 500 1388 510
rect 1418 500 1430 510
rect 1608 500 1620 510
rect 1636 502 1662 510
rect 1650 500 1662 502
rect 580 490 608 500
rect 618 490 646 500
rect 580 484 606 490
rect 596 466 606 484
rect 620 484 646 490
rect 1370 490 1398 500
rect 1408 490 1436 500
rect 1370 484 1396 490
rect 620 466 640 484
rect 1386 476 1396 484
rect 1410 484 1436 490
rect 1602 492 1668 500
rect 1602 490 1630 492
rect 1640 490 1668 492
rect 1602 484 1628 490
rect 1410 476 1430 484
rect 1386 466 1430 476
rect 1618 476 1628 484
rect 1642 484 1668 490
rect 1642 476 1662 484
rect 1618 466 1630 476
rect 1640 466 1662 476
rect 596 450 630 460
rect 1404 456 1430 466
rect 1650 456 1662 466
rect 781 424 909 455
rect 1404 450 1420 456
rect 1650 450 1652 456
rect 2123 424 2251 455
rect 860 418 862 424
rect 2202 418 2204 424
rect 818 408 830 418
rect 860 408 872 418
rect 2160 408 2172 418
rect 2202 408 2214 418
rect 812 398 840 408
rect 850 398 878 408
rect 812 392 838 398
rect 828 384 838 392
rect 852 392 878 398
rect 2154 398 2182 408
rect 2192 398 2220 408
rect 2154 392 2180 398
rect 852 384 872 392
rect 828 374 840 384
rect 850 374 872 384
rect 2170 384 2180 392
rect 2194 392 2220 398
rect 2194 384 2214 392
rect 2170 374 2182 384
rect 2192 374 2214 384
rect 860 364 872 374
rect 2202 364 2214 374
rect 860 358 862 364
rect 2202 358 2204 364
rect 1152 350 1154 356
rect 2114 350 2118 356
rect -328 340 -294 346
rect 1110 340 1122 350
rect 1152 340 1164 350
rect 2114 340 2128 350
rect 446 306 456 340
rect 470 306 490 340
rect 1104 330 1132 340
rect 1142 330 1170 340
rect 1104 324 1130 330
rect 1120 316 1130 324
rect 1144 324 1170 330
rect 1144 316 1164 324
rect 1120 306 1132 316
rect 1142 306 1164 316
rect 1502 306 1512 340
rect 1526 306 1546 340
rect 2084 306 2094 340
rect 2104 330 2134 340
rect 2108 324 2134 330
rect 2108 316 2128 324
rect 2104 306 2128 316
rect 1152 296 1164 306
rect 2114 296 2128 306
rect 1152 290 1154 296
rect 2114 290 2118 296
rect 1064 282 1080 288
rect 1046 272 1090 282
rect 1046 262 1096 272
rect 1070 256 1096 262
rect 1070 254 1090 256
rect 1046 238 1090 254
rect 1236 254 1246 272
rect 1236 238 1248 254
rect 1260 238 1280 272
rect 1064 228 1090 238
rect 1064 222 1080 228
rect 178 188 182 216
rect 216 164 226 188
rect 240 164 260 188
rect 216 154 260 164
rect 276 154 288 216
rect 408 188 422 216
rect 674 188 686 216
rect 446 164 460 188
rect 470 164 490 188
rect 446 154 490 164
rect 712 164 724 188
rect 736 164 756 188
rect 712 154 756 164
rect 772 154 784 216
rect 1198 188 1210 216
rect 1464 188 1476 216
rect 1236 164 1248 188
rect 1260 164 1280 188
rect 1236 154 1280 164
rect 1502 164 1514 188
rect 1526 164 1546 188
rect 1502 154 1546 164
rect 1562 154 1574 216
rect 1694 188 1708 216
rect 1732 164 1746 188
rect 1756 164 1776 188
rect 1732 154 1776 164
rect 1794 154 1804 216
rect 1930 188 1940 216
rect 1968 164 1978 188
rect 1992 164 2012 188
rect 1968 154 2012 164
rect 2026 154 2040 216
rect 234 144 260 154
rect 464 144 490 154
rect 730 144 756 154
rect 1254 144 1280 154
rect 1520 144 1546 154
rect 1750 144 1776 154
rect 1986 144 2012 154
rect 234 138 250 144
rect 464 138 480 144
rect 730 138 746 144
rect 1254 138 1270 144
rect 1520 138 1536 144
rect 1750 138 1766 144
rect 1986 138 2002 144
<< metal1 >>
rect -1668 877 2296 910
rect -29 574 2003 607
rect -429 573 12 574
rect -1529 541 12 573
rect -1529 381 -1494 541
rect -434 517 -368 541
rect 1967 540 2003 574
rect -434 513 -383 517
rect -1282 493 -1212 499
rect -1282 481 -1276 493
rect -1409 447 -1276 481
rect -1282 435 -1276 447
rect -1218 481 -1212 493
rect -418 488 -383 513
rect 120 512 190 518
rect -1218 447 -518 481
rect 120 454 126 512
rect 184 454 190 512
rect 120 448 190 454
rect -1218 435 -1212 447
rect -1282 429 -1212 435
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect -552 373 -518 447
rect -552 339 -296 373
rect -49 342 223 373
rect 810 367 880 373
rect -49 266 -18 342
rect 810 309 816 367
rect 874 309 880 367
rect 810 303 880 309
rect 1967 305 2002 540
rect 2226 318 2296 324
rect 2226 305 2232 318
rect -542 235 -18 266
rect 1967 271 2232 305
rect -542 184 -511 235
rect 1967 185 2002 271
rect 2226 260 2232 271
rect 2290 260 2296 318
rect 2226 254 2296 260
rect -1668 0 2296 33
<< via1 >>
rect -1276 435 -1218 493
rect 126 454 184 512
rect -1110 352 -1052 410
rect 816 309 874 367
rect 2232 260 2290 318
<< metal2 >>
rect 120 512 190 910
rect -1282 493 -1212 498
rect -1282 435 -1276 493
rect -1218 435 -1212 493
rect -1282 429 -1212 435
rect 120 454 126 512
rect 184 454 190 512
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect 120 0 190 454
rect 810 367 880 910
rect 810 309 816 367
rect 874 309 880 367
rect 810 0 880 309
rect 2226 318 2296 324
rect 2226 260 2232 318
rect 2290 260 2296 318
rect 2226 254 2296 260
use xor_scan  xor_scan_0
timestamp 1624135929
transform 1 0 -1756 0 1 102
box 706 -102 1756 808
use dffc  dffc_0
timestamp 1624138001
transform 1 0 66 0 1 106
box -66 -106 2230 804
use and_scan  and_scan_0
timestamp 1624077215
transform 1 0 -1632 0 1 344
box -36 -344 582 566
<< labels >>
rlabel metal2 845 910 845 910 1 CLR
rlabel metal2 2296 288 2296 288 3 Dn
rlabel metal2 157 910 157 910 1 CLK
rlabel metal2 -1246 498 -1246 498 1 CE
rlabel metal2 -1081 346 -1081 346 5 Sout
rlabel metal1 260 910 260 910 1 VDD
rlabel metal1 226 0 226 0 5 VSS
rlabel metal1 15 16 15 16 5 VSS
rlabel space 15 852 15 852 5 VDD
<< end >>
