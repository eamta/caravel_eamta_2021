magic
tech sky130A
timestamp 1616018980
<< poly >>
rect 0 25 33 30
rect 0 8 8 25
rect 25 8 33 25
rect 0 3 33 8
<< polycont >>
rect 8 8 25 25
<< locali >>
rect 0 8 8 25
rect 25 8 33 25
<< viali >>
rect 8 8 25 25
<< metal1 >>
rect 2 25 31 31
rect 2 8 8 25
rect 25 8 31 25
rect 2 2 31 8
<< end >>
