magic
tech sky130A
magscale 1 2
timestamp 1615923543
<< error_p >>
rect -5870 372 -5812 378
rect -5752 372 -5694 378
rect -5634 372 -5576 378
rect -5516 372 -5458 378
rect -5398 372 -5340 378
rect -5280 372 -5222 378
rect -5162 372 -5104 378
rect -5044 372 -4986 378
rect -4926 372 -4868 378
rect -4808 372 -4750 378
rect -4690 372 -4632 378
rect -4572 372 -4514 378
rect -4454 372 -4396 378
rect -4336 372 -4278 378
rect -4218 372 -4160 378
rect -4100 372 -4042 378
rect -3982 372 -3924 378
rect -3864 372 -3806 378
rect -3746 372 -3688 378
rect -3628 372 -3570 378
rect -3510 372 -3452 378
rect -3392 372 -3334 378
rect -3274 372 -3216 378
rect -3156 372 -3098 378
rect -3038 372 -2980 378
rect -2920 372 -2862 378
rect -2802 372 -2744 378
rect -2684 372 -2626 378
rect -2566 372 -2508 378
rect -2448 372 -2390 378
rect -2330 372 -2272 378
rect -2212 372 -2154 378
rect -2094 372 -2036 378
rect -1976 372 -1918 378
rect -1858 372 -1800 378
rect -1740 372 -1682 378
rect -1622 372 -1564 378
rect -1504 372 -1446 378
rect -1386 372 -1328 378
rect -1268 372 -1210 378
rect -1150 372 -1092 378
rect -1032 372 -974 378
rect -914 372 -856 378
rect -796 372 -738 378
rect -678 372 -620 378
rect -560 372 -502 378
rect -442 372 -384 378
rect -324 372 -266 378
rect -206 372 -148 378
rect -88 372 -30 378
rect 30 372 88 378
rect 148 372 206 378
rect 266 372 324 378
rect 384 372 442 378
rect 502 372 560 378
rect 620 372 678 378
rect 738 372 796 378
rect 856 372 914 378
rect 974 372 1032 378
rect 1092 372 1150 378
rect 1210 372 1268 378
rect 1328 372 1386 378
rect 1446 372 1504 378
rect 1564 372 1622 378
rect 1682 372 1740 378
rect 1800 372 1858 378
rect 1918 372 1976 378
rect 2036 372 2094 378
rect 2154 372 2212 378
rect 2272 372 2330 378
rect 2390 372 2448 378
rect 2508 372 2566 378
rect 2626 372 2684 378
rect 2744 372 2802 378
rect 2862 372 2920 378
rect 2980 372 3038 378
rect 3098 372 3156 378
rect 3216 372 3274 378
rect 3334 372 3392 378
rect 3452 372 3510 378
rect 3570 372 3628 378
rect 3688 372 3746 378
rect 3806 372 3864 378
rect 3924 372 3982 378
rect 4042 372 4100 378
rect 4160 372 4218 378
rect 4278 372 4336 378
rect 4396 372 4454 378
rect 4514 372 4572 378
rect 4632 372 4690 378
rect 4750 372 4808 378
rect 4868 372 4926 378
rect 4986 372 5044 378
rect 5104 372 5162 378
rect 5222 372 5280 378
rect 5340 372 5398 378
rect 5458 372 5516 378
rect 5576 372 5634 378
rect 5694 372 5752 378
rect 5812 372 5870 378
rect -5870 338 -5858 372
rect -5752 338 -5740 372
rect -5634 338 -5622 372
rect -5516 338 -5504 372
rect -5398 338 -5386 372
rect -5280 338 -5268 372
rect -5162 338 -5150 372
rect -5044 338 -5032 372
rect -4926 338 -4914 372
rect -4808 338 -4796 372
rect -4690 338 -4678 372
rect -4572 338 -4560 372
rect -4454 338 -4442 372
rect -4336 338 -4324 372
rect -4218 338 -4206 372
rect -4100 338 -4088 372
rect -3982 338 -3970 372
rect -3864 338 -3852 372
rect -3746 338 -3734 372
rect -3628 338 -3616 372
rect -3510 338 -3498 372
rect -3392 338 -3380 372
rect -3274 338 -3262 372
rect -3156 338 -3144 372
rect -3038 338 -3026 372
rect -2920 338 -2908 372
rect -2802 338 -2790 372
rect -2684 338 -2672 372
rect -2566 338 -2554 372
rect -2448 338 -2436 372
rect -2330 338 -2318 372
rect -2212 338 -2200 372
rect -2094 338 -2082 372
rect -1976 338 -1964 372
rect -1858 338 -1846 372
rect -1740 338 -1728 372
rect -1622 338 -1610 372
rect -1504 338 -1492 372
rect -1386 338 -1374 372
rect -1268 338 -1256 372
rect -1150 338 -1138 372
rect -1032 338 -1020 372
rect -914 338 -902 372
rect -796 338 -784 372
rect -678 338 -666 372
rect -560 338 -548 372
rect -442 338 -430 372
rect -324 338 -312 372
rect -206 338 -194 372
rect -88 338 -76 372
rect 30 338 42 372
rect 148 338 160 372
rect 266 338 278 372
rect 384 338 396 372
rect 502 338 514 372
rect 620 338 632 372
rect 738 338 750 372
rect 856 338 868 372
rect 974 338 986 372
rect 1092 338 1104 372
rect 1210 338 1222 372
rect 1328 338 1340 372
rect 1446 338 1458 372
rect 1564 338 1576 372
rect 1682 338 1694 372
rect 1800 338 1812 372
rect 1918 338 1930 372
rect 2036 338 2048 372
rect 2154 338 2166 372
rect 2272 338 2284 372
rect 2390 338 2402 372
rect 2508 338 2520 372
rect 2626 338 2638 372
rect 2744 338 2756 372
rect 2862 338 2874 372
rect 2980 338 2992 372
rect 3098 338 3110 372
rect 3216 338 3228 372
rect 3334 338 3346 372
rect 3452 338 3464 372
rect 3570 338 3582 372
rect 3688 338 3700 372
rect 3806 338 3818 372
rect 3924 338 3936 372
rect 4042 338 4054 372
rect 4160 338 4172 372
rect 4278 338 4290 372
rect 4396 338 4408 372
rect 4514 338 4526 372
rect 4632 338 4644 372
rect 4750 338 4762 372
rect 4868 338 4880 372
rect 4986 338 4998 372
rect 5104 338 5116 372
rect 5222 338 5234 372
rect 5340 338 5352 372
rect 5458 338 5470 372
rect 5576 338 5588 372
rect 5694 338 5706 372
rect 5812 338 5824 372
rect -5870 332 -5812 338
rect -5752 332 -5694 338
rect -5634 332 -5576 338
rect -5516 332 -5458 338
rect -5398 332 -5340 338
rect -5280 332 -5222 338
rect -5162 332 -5104 338
rect -5044 332 -4986 338
rect -4926 332 -4868 338
rect -4808 332 -4750 338
rect -4690 332 -4632 338
rect -4572 332 -4514 338
rect -4454 332 -4396 338
rect -4336 332 -4278 338
rect -4218 332 -4160 338
rect -4100 332 -4042 338
rect -3982 332 -3924 338
rect -3864 332 -3806 338
rect -3746 332 -3688 338
rect -3628 332 -3570 338
rect -3510 332 -3452 338
rect -3392 332 -3334 338
rect -3274 332 -3216 338
rect -3156 332 -3098 338
rect -3038 332 -2980 338
rect -2920 332 -2862 338
rect -2802 332 -2744 338
rect -2684 332 -2626 338
rect -2566 332 -2508 338
rect -2448 332 -2390 338
rect -2330 332 -2272 338
rect -2212 332 -2154 338
rect -2094 332 -2036 338
rect -1976 332 -1918 338
rect -1858 332 -1800 338
rect -1740 332 -1682 338
rect -1622 332 -1564 338
rect -1504 332 -1446 338
rect -1386 332 -1328 338
rect -1268 332 -1210 338
rect -1150 332 -1092 338
rect -1032 332 -974 338
rect -914 332 -856 338
rect -796 332 -738 338
rect -678 332 -620 338
rect -560 332 -502 338
rect -442 332 -384 338
rect -324 332 -266 338
rect -206 332 -148 338
rect -88 332 -30 338
rect 30 332 88 338
rect 148 332 206 338
rect 266 332 324 338
rect 384 332 442 338
rect 502 332 560 338
rect 620 332 678 338
rect 738 332 796 338
rect 856 332 914 338
rect 974 332 1032 338
rect 1092 332 1150 338
rect 1210 332 1268 338
rect 1328 332 1386 338
rect 1446 332 1504 338
rect 1564 332 1622 338
rect 1682 332 1740 338
rect 1800 332 1858 338
rect 1918 332 1976 338
rect 2036 332 2094 338
rect 2154 332 2212 338
rect 2272 332 2330 338
rect 2390 332 2448 338
rect 2508 332 2566 338
rect 2626 332 2684 338
rect 2744 332 2802 338
rect 2862 332 2920 338
rect 2980 332 3038 338
rect 3098 332 3156 338
rect 3216 332 3274 338
rect 3334 332 3392 338
rect 3452 332 3510 338
rect 3570 332 3628 338
rect 3688 332 3746 338
rect 3806 332 3864 338
rect 3924 332 3982 338
rect 4042 332 4100 338
rect 4160 332 4218 338
rect 4278 332 4336 338
rect 4396 332 4454 338
rect 4514 332 4572 338
rect 4632 332 4690 338
rect 4750 332 4808 338
rect 4868 332 4926 338
rect 4986 332 5044 338
rect 5104 332 5162 338
rect 5222 332 5280 338
rect 5340 332 5398 338
rect 5458 332 5516 338
rect 5576 332 5634 338
rect 5694 332 5752 338
rect 5812 332 5870 338
rect -5870 -338 -5812 -332
rect -5752 -338 -5694 -332
rect -5634 -338 -5576 -332
rect -5516 -338 -5458 -332
rect -5398 -338 -5340 -332
rect -5280 -338 -5222 -332
rect -5162 -338 -5104 -332
rect -5044 -338 -4986 -332
rect -4926 -338 -4868 -332
rect -4808 -338 -4750 -332
rect -4690 -338 -4632 -332
rect -4572 -338 -4514 -332
rect -4454 -338 -4396 -332
rect -4336 -338 -4278 -332
rect -4218 -338 -4160 -332
rect -4100 -338 -4042 -332
rect -3982 -338 -3924 -332
rect -3864 -338 -3806 -332
rect -3746 -338 -3688 -332
rect -3628 -338 -3570 -332
rect -3510 -338 -3452 -332
rect -3392 -338 -3334 -332
rect -3274 -338 -3216 -332
rect -3156 -338 -3098 -332
rect -3038 -338 -2980 -332
rect -2920 -338 -2862 -332
rect -2802 -338 -2744 -332
rect -2684 -338 -2626 -332
rect -2566 -338 -2508 -332
rect -2448 -338 -2390 -332
rect -2330 -338 -2272 -332
rect -2212 -338 -2154 -332
rect -2094 -338 -2036 -332
rect -1976 -338 -1918 -332
rect -1858 -338 -1800 -332
rect -1740 -338 -1682 -332
rect -1622 -338 -1564 -332
rect -1504 -338 -1446 -332
rect -1386 -338 -1328 -332
rect -1268 -338 -1210 -332
rect -1150 -338 -1092 -332
rect -1032 -338 -974 -332
rect -914 -338 -856 -332
rect -796 -338 -738 -332
rect -678 -338 -620 -332
rect -560 -338 -502 -332
rect -442 -338 -384 -332
rect -324 -338 -266 -332
rect -206 -338 -148 -332
rect -88 -338 -30 -332
rect 30 -338 88 -332
rect 148 -338 206 -332
rect 266 -338 324 -332
rect 384 -338 442 -332
rect 502 -338 560 -332
rect 620 -338 678 -332
rect 738 -338 796 -332
rect 856 -338 914 -332
rect 974 -338 1032 -332
rect 1092 -338 1150 -332
rect 1210 -338 1268 -332
rect 1328 -338 1386 -332
rect 1446 -338 1504 -332
rect 1564 -338 1622 -332
rect 1682 -338 1740 -332
rect 1800 -338 1858 -332
rect 1918 -338 1976 -332
rect 2036 -338 2094 -332
rect 2154 -338 2212 -332
rect 2272 -338 2330 -332
rect 2390 -338 2448 -332
rect 2508 -338 2566 -332
rect 2626 -338 2684 -332
rect 2744 -338 2802 -332
rect 2862 -338 2920 -332
rect 2980 -338 3038 -332
rect 3098 -338 3156 -332
rect 3216 -338 3274 -332
rect 3334 -338 3392 -332
rect 3452 -338 3510 -332
rect 3570 -338 3628 -332
rect 3688 -338 3746 -332
rect 3806 -338 3864 -332
rect 3924 -338 3982 -332
rect 4042 -338 4100 -332
rect 4160 -338 4218 -332
rect 4278 -338 4336 -332
rect 4396 -338 4454 -332
rect 4514 -338 4572 -332
rect 4632 -338 4690 -332
rect 4750 -338 4808 -332
rect 4868 -338 4926 -332
rect 4986 -338 5044 -332
rect 5104 -338 5162 -332
rect 5222 -338 5280 -332
rect 5340 -338 5398 -332
rect 5458 -338 5516 -332
rect 5576 -338 5634 -332
rect 5694 -338 5752 -332
rect 5812 -338 5870 -332
rect -5870 -372 -5858 -338
rect -5752 -372 -5740 -338
rect -5634 -372 -5622 -338
rect -5516 -372 -5504 -338
rect -5398 -372 -5386 -338
rect -5280 -372 -5268 -338
rect -5162 -372 -5150 -338
rect -5044 -372 -5032 -338
rect -4926 -372 -4914 -338
rect -4808 -372 -4796 -338
rect -4690 -372 -4678 -338
rect -4572 -372 -4560 -338
rect -4454 -372 -4442 -338
rect -4336 -372 -4324 -338
rect -4218 -372 -4206 -338
rect -4100 -372 -4088 -338
rect -3982 -372 -3970 -338
rect -3864 -372 -3852 -338
rect -3746 -372 -3734 -338
rect -3628 -372 -3616 -338
rect -3510 -372 -3498 -338
rect -3392 -372 -3380 -338
rect -3274 -372 -3262 -338
rect -3156 -372 -3144 -338
rect -3038 -372 -3026 -338
rect -2920 -372 -2908 -338
rect -2802 -372 -2790 -338
rect -2684 -372 -2672 -338
rect -2566 -372 -2554 -338
rect -2448 -372 -2436 -338
rect -2330 -372 -2318 -338
rect -2212 -372 -2200 -338
rect -2094 -372 -2082 -338
rect -1976 -372 -1964 -338
rect -1858 -372 -1846 -338
rect -1740 -372 -1728 -338
rect -1622 -372 -1610 -338
rect -1504 -372 -1492 -338
rect -1386 -372 -1374 -338
rect -1268 -372 -1256 -338
rect -1150 -372 -1138 -338
rect -1032 -372 -1020 -338
rect -914 -372 -902 -338
rect -796 -372 -784 -338
rect -678 -372 -666 -338
rect -560 -372 -548 -338
rect -442 -372 -430 -338
rect -324 -372 -312 -338
rect -206 -372 -194 -338
rect -88 -372 -76 -338
rect 30 -372 42 -338
rect 148 -372 160 -338
rect 266 -372 278 -338
rect 384 -372 396 -338
rect 502 -372 514 -338
rect 620 -372 632 -338
rect 738 -372 750 -338
rect 856 -372 868 -338
rect 974 -372 986 -338
rect 1092 -372 1104 -338
rect 1210 -372 1222 -338
rect 1328 -372 1340 -338
rect 1446 -372 1458 -338
rect 1564 -372 1576 -338
rect 1682 -372 1694 -338
rect 1800 -372 1812 -338
rect 1918 -372 1930 -338
rect 2036 -372 2048 -338
rect 2154 -372 2166 -338
rect 2272 -372 2284 -338
rect 2390 -372 2402 -338
rect 2508 -372 2520 -338
rect 2626 -372 2638 -338
rect 2744 -372 2756 -338
rect 2862 -372 2874 -338
rect 2980 -372 2992 -338
rect 3098 -372 3110 -338
rect 3216 -372 3228 -338
rect 3334 -372 3346 -338
rect 3452 -372 3464 -338
rect 3570 -372 3582 -338
rect 3688 -372 3700 -338
rect 3806 -372 3818 -338
rect 3924 -372 3936 -338
rect 4042 -372 4054 -338
rect 4160 -372 4172 -338
rect 4278 -372 4290 -338
rect 4396 -372 4408 -338
rect 4514 -372 4526 -338
rect 4632 -372 4644 -338
rect 4750 -372 4762 -338
rect 4868 -372 4880 -338
rect 4986 -372 4998 -338
rect 5104 -372 5116 -338
rect 5222 -372 5234 -338
rect 5340 -372 5352 -338
rect 5458 -372 5470 -338
rect 5576 -372 5588 -338
rect 5694 -372 5706 -338
rect 5812 -372 5824 -338
rect -5870 -378 -5812 -372
rect -5752 -378 -5694 -372
rect -5634 -378 -5576 -372
rect -5516 -378 -5458 -372
rect -5398 -378 -5340 -372
rect -5280 -378 -5222 -372
rect -5162 -378 -5104 -372
rect -5044 -378 -4986 -372
rect -4926 -378 -4868 -372
rect -4808 -378 -4750 -372
rect -4690 -378 -4632 -372
rect -4572 -378 -4514 -372
rect -4454 -378 -4396 -372
rect -4336 -378 -4278 -372
rect -4218 -378 -4160 -372
rect -4100 -378 -4042 -372
rect -3982 -378 -3924 -372
rect -3864 -378 -3806 -372
rect -3746 -378 -3688 -372
rect -3628 -378 -3570 -372
rect -3510 -378 -3452 -372
rect -3392 -378 -3334 -372
rect -3274 -378 -3216 -372
rect -3156 -378 -3098 -372
rect -3038 -378 -2980 -372
rect -2920 -378 -2862 -372
rect -2802 -378 -2744 -372
rect -2684 -378 -2626 -372
rect -2566 -378 -2508 -372
rect -2448 -378 -2390 -372
rect -2330 -378 -2272 -372
rect -2212 -378 -2154 -372
rect -2094 -378 -2036 -372
rect -1976 -378 -1918 -372
rect -1858 -378 -1800 -372
rect -1740 -378 -1682 -372
rect -1622 -378 -1564 -372
rect -1504 -378 -1446 -372
rect -1386 -378 -1328 -372
rect -1268 -378 -1210 -372
rect -1150 -378 -1092 -372
rect -1032 -378 -974 -372
rect -914 -378 -856 -372
rect -796 -378 -738 -372
rect -678 -378 -620 -372
rect -560 -378 -502 -372
rect -442 -378 -384 -372
rect -324 -378 -266 -372
rect -206 -378 -148 -372
rect -88 -378 -30 -372
rect 30 -378 88 -372
rect 148 -378 206 -372
rect 266 -378 324 -372
rect 384 -378 442 -372
rect 502 -378 560 -372
rect 620 -378 678 -372
rect 738 -378 796 -372
rect 856 -378 914 -372
rect 974 -378 1032 -372
rect 1092 -378 1150 -372
rect 1210 -378 1268 -372
rect 1328 -378 1386 -372
rect 1446 -378 1504 -372
rect 1564 -378 1622 -372
rect 1682 -378 1740 -372
rect 1800 -378 1858 -372
rect 1918 -378 1976 -372
rect 2036 -378 2094 -372
rect 2154 -378 2212 -372
rect 2272 -378 2330 -372
rect 2390 -378 2448 -372
rect 2508 -378 2566 -372
rect 2626 -378 2684 -372
rect 2744 -378 2802 -372
rect 2862 -378 2920 -372
rect 2980 -378 3038 -372
rect 3098 -378 3156 -372
rect 3216 -378 3274 -372
rect 3334 -378 3392 -372
rect 3452 -378 3510 -372
rect 3570 -378 3628 -372
rect 3688 -378 3746 -372
rect 3806 -378 3864 -372
rect 3924 -378 3982 -372
rect 4042 -378 4100 -372
rect 4160 -378 4218 -372
rect 4278 -378 4336 -372
rect 4396 -378 4454 -372
rect 4514 -378 4572 -372
rect 4632 -378 4690 -372
rect 4750 -378 4808 -372
rect 4868 -378 4926 -372
rect 4986 -378 5044 -372
rect 5104 -378 5162 -372
rect 5222 -378 5280 -372
rect 5340 -378 5398 -372
rect 5458 -378 5516 -372
rect 5576 -378 5634 -372
rect 5694 -378 5752 -372
rect 5812 -378 5870 -372
<< nmos >>
rect -5871 -300 -5811 300
rect -5753 -300 -5693 300
rect -5635 -300 -5575 300
rect -5517 -300 -5457 300
rect -5399 -300 -5339 300
rect -5281 -300 -5221 300
rect -5163 -300 -5103 300
rect -5045 -300 -4985 300
rect -4927 -300 -4867 300
rect -4809 -300 -4749 300
rect -4691 -300 -4631 300
rect -4573 -300 -4513 300
rect -4455 -300 -4395 300
rect -4337 -300 -4277 300
rect -4219 -300 -4159 300
rect -4101 -300 -4041 300
rect -3983 -300 -3923 300
rect -3865 -300 -3805 300
rect -3747 -300 -3687 300
rect -3629 -300 -3569 300
rect -3511 -300 -3451 300
rect -3393 -300 -3333 300
rect -3275 -300 -3215 300
rect -3157 -300 -3097 300
rect -3039 -300 -2979 300
rect -2921 -300 -2861 300
rect -2803 -300 -2743 300
rect -2685 -300 -2625 300
rect -2567 -300 -2507 300
rect -2449 -300 -2389 300
rect -2331 -300 -2271 300
rect -2213 -300 -2153 300
rect -2095 -300 -2035 300
rect -1977 -300 -1917 300
rect -1859 -300 -1799 300
rect -1741 -300 -1681 300
rect -1623 -300 -1563 300
rect -1505 -300 -1445 300
rect -1387 -300 -1327 300
rect -1269 -300 -1209 300
rect -1151 -300 -1091 300
rect -1033 -300 -973 300
rect -915 -300 -855 300
rect -797 -300 -737 300
rect -679 -300 -619 300
rect -561 -300 -501 300
rect -443 -300 -383 300
rect -325 -300 -265 300
rect -207 -300 -147 300
rect -89 -300 -29 300
rect 29 -300 89 300
rect 147 -300 207 300
rect 265 -300 325 300
rect 383 -300 443 300
rect 501 -300 561 300
rect 619 -300 679 300
rect 737 -300 797 300
rect 855 -300 915 300
rect 973 -300 1033 300
rect 1091 -300 1151 300
rect 1209 -300 1269 300
rect 1327 -300 1387 300
rect 1445 -300 1505 300
rect 1563 -300 1623 300
rect 1681 -300 1741 300
rect 1799 -300 1859 300
rect 1917 -300 1977 300
rect 2035 -300 2095 300
rect 2153 -300 2213 300
rect 2271 -300 2331 300
rect 2389 -300 2449 300
rect 2507 -300 2567 300
rect 2625 -300 2685 300
rect 2743 -300 2803 300
rect 2861 -300 2921 300
rect 2979 -300 3039 300
rect 3097 -300 3157 300
rect 3215 -300 3275 300
rect 3333 -300 3393 300
rect 3451 -300 3511 300
rect 3569 -300 3629 300
rect 3687 -300 3747 300
rect 3805 -300 3865 300
rect 3923 -300 3983 300
rect 4041 -300 4101 300
rect 4159 -300 4219 300
rect 4277 -300 4337 300
rect 4395 -300 4455 300
rect 4513 -300 4573 300
rect 4631 -300 4691 300
rect 4749 -300 4809 300
rect 4867 -300 4927 300
rect 4985 -300 5045 300
rect 5103 -300 5163 300
rect 5221 -300 5281 300
rect 5339 -300 5399 300
rect 5457 -300 5517 300
rect 5575 -300 5635 300
rect 5693 -300 5753 300
rect 5811 -300 5871 300
<< ndiff >>
rect -5929 288 -5871 300
rect -5929 -288 -5917 288
rect -5883 -288 -5871 288
rect -5929 -300 -5871 -288
rect -5811 288 -5753 300
rect -5811 -288 -5799 288
rect -5765 -288 -5753 288
rect -5811 -300 -5753 -288
rect -5693 288 -5635 300
rect -5693 -288 -5681 288
rect -5647 -288 -5635 288
rect -5693 -300 -5635 -288
rect -5575 288 -5517 300
rect -5575 -288 -5563 288
rect -5529 -288 -5517 288
rect -5575 -300 -5517 -288
rect -5457 288 -5399 300
rect -5457 -288 -5445 288
rect -5411 -288 -5399 288
rect -5457 -300 -5399 -288
rect -5339 288 -5281 300
rect -5339 -288 -5327 288
rect -5293 -288 -5281 288
rect -5339 -300 -5281 -288
rect -5221 288 -5163 300
rect -5221 -288 -5209 288
rect -5175 -288 -5163 288
rect -5221 -300 -5163 -288
rect -5103 288 -5045 300
rect -5103 -288 -5091 288
rect -5057 -288 -5045 288
rect -5103 -300 -5045 -288
rect -4985 288 -4927 300
rect -4985 -288 -4973 288
rect -4939 -288 -4927 288
rect -4985 -300 -4927 -288
rect -4867 288 -4809 300
rect -4867 -288 -4855 288
rect -4821 -288 -4809 288
rect -4867 -300 -4809 -288
rect -4749 288 -4691 300
rect -4749 -288 -4737 288
rect -4703 -288 -4691 288
rect -4749 -300 -4691 -288
rect -4631 288 -4573 300
rect -4631 -288 -4619 288
rect -4585 -288 -4573 288
rect -4631 -300 -4573 -288
rect -4513 288 -4455 300
rect -4513 -288 -4501 288
rect -4467 -288 -4455 288
rect -4513 -300 -4455 -288
rect -4395 288 -4337 300
rect -4395 -288 -4383 288
rect -4349 -288 -4337 288
rect -4395 -300 -4337 -288
rect -4277 288 -4219 300
rect -4277 -288 -4265 288
rect -4231 -288 -4219 288
rect -4277 -300 -4219 -288
rect -4159 288 -4101 300
rect -4159 -288 -4147 288
rect -4113 -288 -4101 288
rect -4159 -300 -4101 -288
rect -4041 288 -3983 300
rect -4041 -288 -4029 288
rect -3995 -288 -3983 288
rect -4041 -300 -3983 -288
rect -3923 288 -3865 300
rect -3923 -288 -3911 288
rect -3877 -288 -3865 288
rect -3923 -300 -3865 -288
rect -3805 288 -3747 300
rect -3805 -288 -3793 288
rect -3759 -288 -3747 288
rect -3805 -300 -3747 -288
rect -3687 288 -3629 300
rect -3687 -288 -3675 288
rect -3641 -288 -3629 288
rect -3687 -300 -3629 -288
rect -3569 288 -3511 300
rect -3569 -288 -3557 288
rect -3523 -288 -3511 288
rect -3569 -300 -3511 -288
rect -3451 288 -3393 300
rect -3451 -288 -3439 288
rect -3405 -288 -3393 288
rect -3451 -300 -3393 -288
rect -3333 288 -3275 300
rect -3333 -288 -3321 288
rect -3287 -288 -3275 288
rect -3333 -300 -3275 -288
rect -3215 288 -3157 300
rect -3215 -288 -3203 288
rect -3169 -288 -3157 288
rect -3215 -300 -3157 -288
rect -3097 288 -3039 300
rect -3097 -288 -3085 288
rect -3051 -288 -3039 288
rect -3097 -300 -3039 -288
rect -2979 288 -2921 300
rect -2979 -288 -2967 288
rect -2933 -288 -2921 288
rect -2979 -300 -2921 -288
rect -2861 288 -2803 300
rect -2861 -288 -2849 288
rect -2815 -288 -2803 288
rect -2861 -300 -2803 -288
rect -2743 288 -2685 300
rect -2743 -288 -2731 288
rect -2697 -288 -2685 288
rect -2743 -300 -2685 -288
rect -2625 288 -2567 300
rect -2625 -288 -2613 288
rect -2579 -288 -2567 288
rect -2625 -300 -2567 -288
rect -2507 288 -2449 300
rect -2507 -288 -2495 288
rect -2461 -288 -2449 288
rect -2507 -300 -2449 -288
rect -2389 288 -2331 300
rect -2389 -288 -2377 288
rect -2343 -288 -2331 288
rect -2389 -300 -2331 -288
rect -2271 288 -2213 300
rect -2271 -288 -2259 288
rect -2225 -288 -2213 288
rect -2271 -300 -2213 -288
rect -2153 288 -2095 300
rect -2153 -288 -2141 288
rect -2107 -288 -2095 288
rect -2153 -300 -2095 -288
rect -2035 288 -1977 300
rect -2035 -288 -2023 288
rect -1989 -288 -1977 288
rect -2035 -300 -1977 -288
rect -1917 288 -1859 300
rect -1917 -288 -1905 288
rect -1871 -288 -1859 288
rect -1917 -300 -1859 -288
rect -1799 288 -1741 300
rect -1799 -288 -1787 288
rect -1753 -288 -1741 288
rect -1799 -300 -1741 -288
rect -1681 288 -1623 300
rect -1681 -288 -1669 288
rect -1635 -288 -1623 288
rect -1681 -300 -1623 -288
rect -1563 288 -1505 300
rect -1563 -288 -1551 288
rect -1517 -288 -1505 288
rect -1563 -300 -1505 -288
rect -1445 288 -1387 300
rect -1445 -288 -1433 288
rect -1399 -288 -1387 288
rect -1445 -300 -1387 -288
rect -1327 288 -1269 300
rect -1327 -288 -1315 288
rect -1281 -288 -1269 288
rect -1327 -300 -1269 -288
rect -1209 288 -1151 300
rect -1209 -288 -1197 288
rect -1163 -288 -1151 288
rect -1209 -300 -1151 -288
rect -1091 288 -1033 300
rect -1091 -288 -1079 288
rect -1045 -288 -1033 288
rect -1091 -300 -1033 -288
rect -973 288 -915 300
rect -973 -288 -961 288
rect -927 -288 -915 288
rect -973 -300 -915 -288
rect -855 288 -797 300
rect -855 -288 -843 288
rect -809 -288 -797 288
rect -855 -300 -797 -288
rect -737 288 -679 300
rect -737 -288 -725 288
rect -691 -288 -679 288
rect -737 -300 -679 -288
rect -619 288 -561 300
rect -619 -288 -607 288
rect -573 -288 -561 288
rect -619 -300 -561 -288
rect -501 288 -443 300
rect -501 -288 -489 288
rect -455 -288 -443 288
rect -501 -300 -443 -288
rect -383 288 -325 300
rect -383 -288 -371 288
rect -337 -288 -325 288
rect -383 -300 -325 -288
rect -265 288 -207 300
rect -265 -288 -253 288
rect -219 -288 -207 288
rect -265 -300 -207 -288
rect -147 288 -89 300
rect -147 -288 -135 288
rect -101 -288 -89 288
rect -147 -300 -89 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 89 288 147 300
rect 89 -288 101 288
rect 135 -288 147 288
rect 89 -300 147 -288
rect 207 288 265 300
rect 207 -288 219 288
rect 253 -288 265 288
rect 207 -300 265 -288
rect 325 288 383 300
rect 325 -288 337 288
rect 371 -288 383 288
rect 325 -300 383 -288
rect 443 288 501 300
rect 443 -288 455 288
rect 489 -288 501 288
rect 443 -300 501 -288
rect 561 288 619 300
rect 561 -288 573 288
rect 607 -288 619 288
rect 561 -300 619 -288
rect 679 288 737 300
rect 679 -288 691 288
rect 725 -288 737 288
rect 679 -300 737 -288
rect 797 288 855 300
rect 797 -288 809 288
rect 843 -288 855 288
rect 797 -300 855 -288
rect 915 288 973 300
rect 915 -288 927 288
rect 961 -288 973 288
rect 915 -300 973 -288
rect 1033 288 1091 300
rect 1033 -288 1045 288
rect 1079 -288 1091 288
rect 1033 -300 1091 -288
rect 1151 288 1209 300
rect 1151 -288 1163 288
rect 1197 -288 1209 288
rect 1151 -300 1209 -288
rect 1269 288 1327 300
rect 1269 -288 1281 288
rect 1315 -288 1327 288
rect 1269 -300 1327 -288
rect 1387 288 1445 300
rect 1387 -288 1399 288
rect 1433 -288 1445 288
rect 1387 -300 1445 -288
rect 1505 288 1563 300
rect 1505 -288 1517 288
rect 1551 -288 1563 288
rect 1505 -300 1563 -288
rect 1623 288 1681 300
rect 1623 -288 1635 288
rect 1669 -288 1681 288
rect 1623 -300 1681 -288
rect 1741 288 1799 300
rect 1741 -288 1753 288
rect 1787 -288 1799 288
rect 1741 -300 1799 -288
rect 1859 288 1917 300
rect 1859 -288 1871 288
rect 1905 -288 1917 288
rect 1859 -300 1917 -288
rect 1977 288 2035 300
rect 1977 -288 1989 288
rect 2023 -288 2035 288
rect 1977 -300 2035 -288
rect 2095 288 2153 300
rect 2095 -288 2107 288
rect 2141 -288 2153 288
rect 2095 -300 2153 -288
rect 2213 288 2271 300
rect 2213 -288 2225 288
rect 2259 -288 2271 288
rect 2213 -300 2271 -288
rect 2331 288 2389 300
rect 2331 -288 2343 288
rect 2377 -288 2389 288
rect 2331 -300 2389 -288
rect 2449 288 2507 300
rect 2449 -288 2461 288
rect 2495 -288 2507 288
rect 2449 -300 2507 -288
rect 2567 288 2625 300
rect 2567 -288 2579 288
rect 2613 -288 2625 288
rect 2567 -300 2625 -288
rect 2685 288 2743 300
rect 2685 -288 2697 288
rect 2731 -288 2743 288
rect 2685 -300 2743 -288
rect 2803 288 2861 300
rect 2803 -288 2815 288
rect 2849 -288 2861 288
rect 2803 -300 2861 -288
rect 2921 288 2979 300
rect 2921 -288 2933 288
rect 2967 -288 2979 288
rect 2921 -300 2979 -288
rect 3039 288 3097 300
rect 3039 -288 3051 288
rect 3085 -288 3097 288
rect 3039 -300 3097 -288
rect 3157 288 3215 300
rect 3157 -288 3169 288
rect 3203 -288 3215 288
rect 3157 -300 3215 -288
rect 3275 288 3333 300
rect 3275 -288 3287 288
rect 3321 -288 3333 288
rect 3275 -300 3333 -288
rect 3393 288 3451 300
rect 3393 -288 3405 288
rect 3439 -288 3451 288
rect 3393 -300 3451 -288
rect 3511 288 3569 300
rect 3511 -288 3523 288
rect 3557 -288 3569 288
rect 3511 -300 3569 -288
rect 3629 288 3687 300
rect 3629 -288 3641 288
rect 3675 -288 3687 288
rect 3629 -300 3687 -288
rect 3747 288 3805 300
rect 3747 -288 3759 288
rect 3793 -288 3805 288
rect 3747 -300 3805 -288
rect 3865 288 3923 300
rect 3865 -288 3877 288
rect 3911 -288 3923 288
rect 3865 -300 3923 -288
rect 3983 288 4041 300
rect 3983 -288 3995 288
rect 4029 -288 4041 288
rect 3983 -300 4041 -288
rect 4101 288 4159 300
rect 4101 -288 4113 288
rect 4147 -288 4159 288
rect 4101 -300 4159 -288
rect 4219 288 4277 300
rect 4219 -288 4231 288
rect 4265 -288 4277 288
rect 4219 -300 4277 -288
rect 4337 288 4395 300
rect 4337 -288 4349 288
rect 4383 -288 4395 288
rect 4337 -300 4395 -288
rect 4455 288 4513 300
rect 4455 -288 4467 288
rect 4501 -288 4513 288
rect 4455 -300 4513 -288
rect 4573 288 4631 300
rect 4573 -288 4585 288
rect 4619 -288 4631 288
rect 4573 -300 4631 -288
rect 4691 288 4749 300
rect 4691 -288 4703 288
rect 4737 -288 4749 288
rect 4691 -300 4749 -288
rect 4809 288 4867 300
rect 4809 -288 4821 288
rect 4855 -288 4867 288
rect 4809 -300 4867 -288
rect 4927 288 4985 300
rect 4927 -288 4939 288
rect 4973 -288 4985 288
rect 4927 -300 4985 -288
rect 5045 288 5103 300
rect 5045 -288 5057 288
rect 5091 -288 5103 288
rect 5045 -300 5103 -288
rect 5163 288 5221 300
rect 5163 -288 5175 288
rect 5209 -288 5221 288
rect 5163 -300 5221 -288
rect 5281 288 5339 300
rect 5281 -288 5293 288
rect 5327 -288 5339 288
rect 5281 -300 5339 -288
rect 5399 288 5457 300
rect 5399 -288 5411 288
rect 5445 -288 5457 288
rect 5399 -300 5457 -288
rect 5517 288 5575 300
rect 5517 -288 5529 288
rect 5563 -288 5575 288
rect 5517 -300 5575 -288
rect 5635 288 5693 300
rect 5635 -288 5647 288
rect 5681 -288 5693 288
rect 5635 -300 5693 -288
rect 5753 288 5811 300
rect 5753 -288 5765 288
rect 5799 -288 5811 288
rect 5753 -300 5811 -288
rect 5871 288 5929 300
rect 5871 -288 5883 288
rect 5917 -288 5929 288
rect 5871 -300 5929 -288
<< ndiffc >>
rect -5917 -288 -5883 288
rect -5799 -288 -5765 288
rect -5681 -288 -5647 288
rect -5563 -288 -5529 288
rect -5445 -288 -5411 288
rect -5327 -288 -5293 288
rect -5209 -288 -5175 288
rect -5091 -288 -5057 288
rect -4973 -288 -4939 288
rect -4855 -288 -4821 288
rect -4737 -288 -4703 288
rect -4619 -288 -4585 288
rect -4501 -288 -4467 288
rect -4383 -288 -4349 288
rect -4265 -288 -4231 288
rect -4147 -288 -4113 288
rect -4029 -288 -3995 288
rect -3911 -288 -3877 288
rect -3793 -288 -3759 288
rect -3675 -288 -3641 288
rect -3557 -288 -3523 288
rect -3439 -288 -3405 288
rect -3321 -288 -3287 288
rect -3203 -288 -3169 288
rect -3085 -288 -3051 288
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect 3051 -288 3085 288
rect 3169 -288 3203 288
rect 3287 -288 3321 288
rect 3405 -288 3439 288
rect 3523 -288 3557 288
rect 3641 -288 3675 288
rect 3759 -288 3793 288
rect 3877 -288 3911 288
rect 3995 -288 4029 288
rect 4113 -288 4147 288
rect 4231 -288 4265 288
rect 4349 -288 4383 288
rect 4467 -288 4501 288
rect 4585 -288 4619 288
rect 4703 -288 4737 288
rect 4821 -288 4855 288
rect 4939 -288 4973 288
rect 5057 -288 5091 288
rect 5175 -288 5209 288
rect 5293 -288 5327 288
rect 5411 -288 5445 288
rect 5529 -288 5563 288
rect 5647 -288 5681 288
rect 5765 -288 5799 288
rect 5883 -288 5917 288
<< poly >>
rect -5874 372 -5808 388
rect -5874 338 -5858 372
rect -5824 338 -5808 372
rect -5874 322 -5808 338
rect -5756 372 -5690 388
rect -5756 338 -5740 372
rect -5706 338 -5690 372
rect -5756 322 -5690 338
rect -5638 372 -5572 388
rect -5638 338 -5622 372
rect -5588 338 -5572 372
rect -5638 322 -5572 338
rect -5520 372 -5454 388
rect -5520 338 -5504 372
rect -5470 338 -5454 372
rect -5520 322 -5454 338
rect -5402 372 -5336 388
rect -5402 338 -5386 372
rect -5352 338 -5336 372
rect -5402 322 -5336 338
rect -5284 372 -5218 388
rect -5284 338 -5268 372
rect -5234 338 -5218 372
rect -5284 322 -5218 338
rect -5166 372 -5100 388
rect -5166 338 -5150 372
rect -5116 338 -5100 372
rect -5166 322 -5100 338
rect -5048 372 -4982 388
rect -5048 338 -5032 372
rect -4998 338 -4982 372
rect -5048 322 -4982 338
rect -4930 372 -4864 388
rect -4930 338 -4914 372
rect -4880 338 -4864 372
rect -4930 322 -4864 338
rect -4812 372 -4746 388
rect -4812 338 -4796 372
rect -4762 338 -4746 372
rect -4812 322 -4746 338
rect -4694 372 -4628 388
rect -4694 338 -4678 372
rect -4644 338 -4628 372
rect -4694 322 -4628 338
rect -4576 372 -4510 388
rect -4576 338 -4560 372
rect -4526 338 -4510 372
rect -4576 322 -4510 338
rect -4458 372 -4392 388
rect -4458 338 -4442 372
rect -4408 338 -4392 372
rect -4458 322 -4392 338
rect -4340 372 -4274 388
rect -4340 338 -4324 372
rect -4290 338 -4274 372
rect -4340 322 -4274 338
rect -4222 372 -4156 388
rect -4222 338 -4206 372
rect -4172 338 -4156 372
rect -4222 322 -4156 338
rect -4104 372 -4038 388
rect -4104 338 -4088 372
rect -4054 338 -4038 372
rect -4104 322 -4038 338
rect -3986 372 -3920 388
rect -3986 338 -3970 372
rect -3936 338 -3920 372
rect -3986 322 -3920 338
rect -3868 372 -3802 388
rect -3868 338 -3852 372
rect -3818 338 -3802 372
rect -3868 322 -3802 338
rect -3750 372 -3684 388
rect -3750 338 -3734 372
rect -3700 338 -3684 372
rect -3750 322 -3684 338
rect -3632 372 -3566 388
rect -3632 338 -3616 372
rect -3582 338 -3566 372
rect -3632 322 -3566 338
rect -3514 372 -3448 388
rect -3514 338 -3498 372
rect -3464 338 -3448 372
rect -3514 322 -3448 338
rect -3396 372 -3330 388
rect -3396 338 -3380 372
rect -3346 338 -3330 372
rect -3396 322 -3330 338
rect -3278 372 -3212 388
rect -3278 338 -3262 372
rect -3228 338 -3212 372
rect -3278 322 -3212 338
rect -3160 372 -3094 388
rect -3160 338 -3144 372
rect -3110 338 -3094 372
rect -3160 322 -3094 338
rect -3042 372 -2976 388
rect -3042 338 -3026 372
rect -2992 338 -2976 372
rect -3042 322 -2976 338
rect -2924 372 -2858 388
rect -2924 338 -2908 372
rect -2874 338 -2858 372
rect -2924 322 -2858 338
rect -2806 372 -2740 388
rect -2806 338 -2790 372
rect -2756 338 -2740 372
rect -2806 322 -2740 338
rect -2688 372 -2622 388
rect -2688 338 -2672 372
rect -2638 338 -2622 372
rect -2688 322 -2622 338
rect -2570 372 -2504 388
rect -2570 338 -2554 372
rect -2520 338 -2504 372
rect -2570 322 -2504 338
rect -2452 372 -2386 388
rect -2452 338 -2436 372
rect -2402 338 -2386 372
rect -2452 322 -2386 338
rect -2334 372 -2268 388
rect -2334 338 -2318 372
rect -2284 338 -2268 372
rect -2334 322 -2268 338
rect -2216 372 -2150 388
rect -2216 338 -2200 372
rect -2166 338 -2150 372
rect -2216 322 -2150 338
rect -2098 372 -2032 388
rect -2098 338 -2082 372
rect -2048 338 -2032 372
rect -2098 322 -2032 338
rect -1980 372 -1914 388
rect -1980 338 -1964 372
rect -1930 338 -1914 372
rect -1980 322 -1914 338
rect -1862 372 -1796 388
rect -1862 338 -1846 372
rect -1812 338 -1796 372
rect -1862 322 -1796 338
rect -1744 372 -1678 388
rect -1744 338 -1728 372
rect -1694 338 -1678 372
rect -1744 322 -1678 338
rect -1626 372 -1560 388
rect -1626 338 -1610 372
rect -1576 338 -1560 372
rect -1626 322 -1560 338
rect -1508 372 -1442 388
rect -1508 338 -1492 372
rect -1458 338 -1442 372
rect -1508 322 -1442 338
rect -1390 372 -1324 388
rect -1390 338 -1374 372
rect -1340 338 -1324 372
rect -1390 322 -1324 338
rect -1272 372 -1206 388
rect -1272 338 -1256 372
rect -1222 338 -1206 372
rect -1272 322 -1206 338
rect -1154 372 -1088 388
rect -1154 338 -1138 372
rect -1104 338 -1088 372
rect -1154 322 -1088 338
rect -1036 372 -970 388
rect -1036 338 -1020 372
rect -986 338 -970 372
rect -1036 322 -970 338
rect -918 372 -852 388
rect -918 338 -902 372
rect -868 338 -852 372
rect -918 322 -852 338
rect -800 372 -734 388
rect -800 338 -784 372
rect -750 338 -734 372
rect -800 322 -734 338
rect -682 372 -616 388
rect -682 338 -666 372
rect -632 338 -616 372
rect -682 322 -616 338
rect -564 372 -498 388
rect -564 338 -548 372
rect -514 338 -498 372
rect -564 322 -498 338
rect -446 372 -380 388
rect -446 338 -430 372
rect -396 338 -380 372
rect -446 322 -380 338
rect -328 372 -262 388
rect -328 338 -312 372
rect -278 338 -262 372
rect -328 322 -262 338
rect -210 372 -144 388
rect -210 338 -194 372
rect -160 338 -144 372
rect -210 322 -144 338
rect -92 372 -26 388
rect -92 338 -76 372
rect -42 338 -26 372
rect -92 322 -26 338
rect 26 372 92 388
rect 26 338 42 372
rect 76 338 92 372
rect 26 322 92 338
rect 144 372 210 388
rect 144 338 160 372
rect 194 338 210 372
rect 144 322 210 338
rect 262 372 328 388
rect 262 338 278 372
rect 312 338 328 372
rect 262 322 328 338
rect 380 372 446 388
rect 380 338 396 372
rect 430 338 446 372
rect 380 322 446 338
rect 498 372 564 388
rect 498 338 514 372
rect 548 338 564 372
rect 498 322 564 338
rect 616 372 682 388
rect 616 338 632 372
rect 666 338 682 372
rect 616 322 682 338
rect 734 372 800 388
rect 734 338 750 372
rect 784 338 800 372
rect 734 322 800 338
rect 852 372 918 388
rect 852 338 868 372
rect 902 338 918 372
rect 852 322 918 338
rect 970 372 1036 388
rect 970 338 986 372
rect 1020 338 1036 372
rect 970 322 1036 338
rect 1088 372 1154 388
rect 1088 338 1104 372
rect 1138 338 1154 372
rect 1088 322 1154 338
rect 1206 372 1272 388
rect 1206 338 1222 372
rect 1256 338 1272 372
rect 1206 322 1272 338
rect 1324 372 1390 388
rect 1324 338 1340 372
rect 1374 338 1390 372
rect 1324 322 1390 338
rect 1442 372 1508 388
rect 1442 338 1458 372
rect 1492 338 1508 372
rect 1442 322 1508 338
rect 1560 372 1626 388
rect 1560 338 1576 372
rect 1610 338 1626 372
rect 1560 322 1626 338
rect 1678 372 1744 388
rect 1678 338 1694 372
rect 1728 338 1744 372
rect 1678 322 1744 338
rect 1796 372 1862 388
rect 1796 338 1812 372
rect 1846 338 1862 372
rect 1796 322 1862 338
rect 1914 372 1980 388
rect 1914 338 1930 372
rect 1964 338 1980 372
rect 1914 322 1980 338
rect 2032 372 2098 388
rect 2032 338 2048 372
rect 2082 338 2098 372
rect 2032 322 2098 338
rect 2150 372 2216 388
rect 2150 338 2166 372
rect 2200 338 2216 372
rect 2150 322 2216 338
rect 2268 372 2334 388
rect 2268 338 2284 372
rect 2318 338 2334 372
rect 2268 322 2334 338
rect 2386 372 2452 388
rect 2386 338 2402 372
rect 2436 338 2452 372
rect 2386 322 2452 338
rect 2504 372 2570 388
rect 2504 338 2520 372
rect 2554 338 2570 372
rect 2504 322 2570 338
rect 2622 372 2688 388
rect 2622 338 2638 372
rect 2672 338 2688 372
rect 2622 322 2688 338
rect 2740 372 2806 388
rect 2740 338 2756 372
rect 2790 338 2806 372
rect 2740 322 2806 338
rect 2858 372 2924 388
rect 2858 338 2874 372
rect 2908 338 2924 372
rect 2858 322 2924 338
rect 2976 372 3042 388
rect 2976 338 2992 372
rect 3026 338 3042 372
rect 2976 322 3042 338
rect 3094 372 3160 388
rect 3094 338 3110 372
rect 3144 338 3160 372
rect 3094 322 3160 338
rect 3212 372 3278 388
rect 3212 338 3228 372
rect 3262 338 3278 372
rect 3212 322 3278 338
rect 3330 372 3396 388
rect 3330 338 3346 372
rect 3380 338 3396 372
rect 3330 322 3396 338
rect 3448 372 3514 388
rect 3448 338 3464 372
rect 3498 338 3514 372
rect 3448 322 3514 338
rect 3566 372 3632 388
rect 3566 338 3582 372
rect 3616 338 3632 372
rect 3566 322 3632 338
rect 3684 372 3750 388
rect 3684 338 3700 372
rect 3734 338 3750 372
rect 3684 322 3750 338
rect 3802 372 3868 388
rect 3802 338 3818 372
rect 3852 338 3868 372
rect 3802 322 3868 338
rect 3920 372 3986 388
rect 3920 338 3936 372
rect 3970 338 3986 372
rect 3920 322 3986 338
rect 4038 372 4104 388
rect 4038 338 4054 372
rect 4088 338 4104 372
rect 4038 322 4104 338
rect 4156 372 4222 388
rect 4156 338 4172 372
rect 4206 338 4222 372
rect 4156 322 4222 338
rect 4274 372 4340 388
rect 4274 338 4290 372
rect 4324 338 4340 372
rect 4274 322 4340 338
rect 4392 372 4458 388
rect 4392 338 4408 372
rect 4442 338 4458 372
rect 4392 322 4458 338
rect 4510 372 4576 388
rect 4510 338 4526 372
rect 4560 338 4576 372
rect 4510 322 4576 338
rect 4628 372 4694 388
rect 4628 338 4644 372
rect 4678 338 4694 372
rect 4628 322 4694 338
rect 4746 372 4812 388
rect 4746 338 4762 372
rect 4796 338 4812 372
rect 4746 322 4812 338
rect 4864 372 4930 388
rect 4864 338 4880 372
rect 4914 338 4930 372
rect 4864 322 4930 338
rect 4982 372 5048 388
rect 4982 338 4998 372
rect 5032 338 5048 372
rect 4982 322 5048 338
rect 5100 372 5166 388
rect 5100 338 5116 372
rect 5150 338 5166 372
rect 5100 322 5166 338
rect 5218 372 5284 388
rect 5218 338 5234 372
rect 5268 338 5284 372
rect 5218 322 5284 338
rect 5336 372 5402 388
rect 5336 338 5352 372
rect 5386 338 5402 372
rect 5336 322 5402 338
rect 5454 372 5520 388
rect 5454 338 5470 372
rect 5504 338 5520 372
rect 5454 322 5520 338
rect 5572 372 5638 388
rect 5572 338 5588 372
rect 5622 338 5638 372
rect 5572 322 5638 338
rect 5690 372 5756 388
rect 5690 338 5706 372
rect 5740 338 5756 372
rect 5690 322 5756 338
rect 5808 372 5874 388
rect 5808 338 5824 372
rect 5858 338 5874 372
rect 5808 322 5874 338
rect -5871 300 -5811 322
rect -5753 300 -5693 322
rect -5635 300 -5575 322
rect -5517 300 -5457 322
rect -5399 300 -5339 322
rect -5281 300 -5221 322
rect -5163 300 -5103 322
rect -5045 300 -4985 322
rect -4927 300 -4867 322
rect -4809 300 -4749 322
rect -4691 300 -4631 322
rect -4573 300 -4513 322
rect -4455 300 -4395 322
rect -4337 300 -4277 322
rect -4219 300 -4159 322
rect -4101 300 -4041 322
rect -3983 300 -3923 322
rect -3865 300 -3805 322
rect -3747 300 -3687 322
rect -3629 300 -3569 322
rect -3511 300 -3451 322
rect -3393 300 -3333 322
rect -3275 300 -3215 322
rect -3157 300 -3097 322
rect -3039 300 -2979 322
rect -2921 300 -2861 322
rect -2803 300 -2743 322
rect -2685 300 -2625 322
rect -2567 300 -2507 322
rect -2449 300 -2389 322
rect -2331 300 -2271 322
rect -2213 300 -2153 322
rect -2095 300 -2035 322
rect -1977 300 -1917 322
rect -1859 300 -1799 322
rect -1741 300 -1681 322
rect -1623 300 -1563 322
rect -1505 300 -1445 322
rect -1387 300 -1327 322
rect -1269 300 -1209 322
rect -1151 300 -1091 322
rect -1033 300 -973 322
rect -915 300 -855 322
rect -797 300 -737 322
rect -679 300 -619 322
rect -561 300 -501 322
rect -443 300 -383 322
rect -325 300 -265 322
rect -207 300 -147 322
rect -89 300 -29 322
rect 29 300 89 322
rect 147 300 207 322
rect 265 300 325 322
rect 383 300 443 322
rect 501 300 561 322
rect 619 300 679 322
rect 737 300 797 322
rect 855 300 915 322
rect 973 300 1033 322
rect 1091 300 1151 322
rect 1209 300 1269 322
rect 1327 300 1387 322
rect 1445 300 1505 322
rect 1563 300 1623 322
rect 1681 300 1741 322
rect 1799 300 1859 322
rect 1917 300 1977 322
rect 2035 300 2095 322
rect 2153 300 2213 322
rect 2271 300 2331 322
rect 2389 300 2449 322
rect 2507 300 2567 322
rect 2625 300 2685 322
rect 2743 300 2803 322
rect 2861 300 2921 322
rect 2979 300 3039 322
rect 3097 300 3157 322
rect 3215 300 3275 322
rect 3333 300 3393 322
rect 3451 300 3511 322
rect 3569 300 3629 322
rect 3687 300 3747 322
rect 3805 300 3865 322
rect 3923 300 3983 322
rect 4041 300 4101 322
rect 4159 300 4219 322
rect 4277 300 4337 322
rect 4395 300 4455 322
rect 4513 300 4573 322
rect 4631 300 4691 322
rect 4749 300 4809 322
rect 4867 300 4927 322
rect 4985 300 5045 322
rect 5103 300 5163 322
rect 5221 300 5281 322
rect 5339 300 5399 322
rect 5457 300 5517 322
rect 5575 300 5635 322
rect 5693 300 5753 322
rect 5811 300 5871 322
rect -5871 -322 -5811 -300
rect -5753 -322 -5693 -300
rect -5635 -322 -5575 -300
rect -5517 -322 -5457 -300
rect -5399 -322 -5339 -300
rect -5281 -322 -5221 -300
rect -5163 -322 -5103 -300
rect -5045 -322 -4985 -300
rect -4927 -322 -4867 -300
rect -4809 -322 -4749 -300
rect -4691 -322 -4631 -300
rect -4573 -322 -4513 -300
rect -4455 -322 -4395 -300
rect -4337 -322 -4277 -300
rect -4219 -322 -4159 -300
rect -4101 -322 -4041 -300
rect -3983 -322 -3923 -300
rect -3865 -322 -3805 -300
rect -3747 -322 -3687 -300
rect -3629 -322 -3569 -300
rect -3511 -322 -3451 -300
rect -3393 -322 -3333 -300
rect -3275 -322 -3215 -300
rect -3157 -322 -3097 -300
rect -3039 -322 -2979 -300
rect -2921 -322 -2861 -300
rect -2803 -322 -2743 -300
rect -2685 -322 -2625 -300
rect -2567 -322 -2507 -300
rect -2449 -322 -2389 -300
rect -2331 -322 -2271 -300
rect -2213 -322 -2153 -300
rect -2095 -322 -2035 -300
rect -1977 -322 -1917 -300
rect -1859 -322 -1799 -300
rect -1741 -322 -1681 -300
rect -1623 -322 -1563 -300
rect -1505 -322 -1445 -300
rect -1387 -322 -1327 -300
rect -1269 -322 -1209 -300
rect -1151 -322 -1091 -300
rect -1033 -322 -973 -300
rect -915 -322 -855 -300
rect -797 -322 -737 -300
rect -679 -322 -619 -300
rect -561 -322 -501 -300
rect -443 -322 -383 -300
rect -325 -322 -265 -300
rect -207 -322 -147 -300
rect -89 -322 -29 -300
rect 29 -322 89 -300
rect 147 -322 207 -300
rect 265 -322 325 -300
rect 383 -322 443 -300
rect 501 -322 561 -300
rect 619 -322 679 -300
rect 737 -322 797 -300
rect 855 -322 915 -300
rect 973 -322 1033 -300
rect 1091 -322 1151 -300
rect 1209 -322 1269 -300
rect 1327 -322 1387 -300
rect 1445 -322 1505 -300
rect 1563 -322 1623 -300
rect 1681 -322 1741 -300
rect 1799 -322 1859 -300
rect 1917 -322 1977 -300
rect 2035 -322 2095 -300
rect 2153 -322 2213 -300
rect 2271 -322 2331 -300
rect 2389 -322 2449 -300
rect 2507 -322 2567 -300
rect 2625 -322 2685 -300
rect 2743 -322 2803 -300
rect 2861 -322 2921 -300
rect 2979 -322 3039 -300
rect 3097 -322 3157 -300
rect 3215 -322 3275 -300
rect 3333 -322 3393 -300
rect 3451 -322 3511 -300
rect 3569 -322 3629 -300
rect 3687 -322 3747 -300
rect 3805 -322 3865 -300
rect 3923 -322 3983 -300
rect 4041 -322 4101 -300
rect 4159 -322 4219 -300
rect 4277 -322 4337 -300
rect 4395 -322 4455 -300
rect 4513 -322 4573 -300
rect 4631 -322 4691 -300
rect 4749 -322 4809 -300
rect 4867 -322 4927 -300
rect 4985 -322 5045 -300
rect 5103 -322 5163 -300
rect 5221 -322 5281 -300
rect 5339 -322 5399 -300
rect 5457 -322 5517 -300
rect 5575 -322 5635 -300
rect 5693 -322 5753 -300
rect 5811 -322 5871 -300
rect -5874 -338 -5808 -322
rect -5874 -372 -5858 -338
rect -5824 -372 -5808 -338
rect -5874 -388 -5808 -372
rect -5756 -338 -5690 -322
rect -5756 -372 -5740 -338
rect -5706 -372 -5690 -338
rect -5756 -388 -5690 -372
rect -5638 -338 -5572 -322
rect -5638 -372 -5622 -338
rect -5588 -372 -5572 -338
rect -5638 -388 -5572 -372
rect -5520 -338 -5454 -322
rect -5520 -372 -5504 -338
rect -5470 -372 -5454 -338
rect -5520 -388 -5454 -372
rect -5402 -338 -5336 -322
rect -5402 -372 -5386 -338
rect -5352 -372 -5336 -338
rect -5402 -388 -5336 -372
rect -5284 -338 -5218 -322
rect -5284 -372 -5268 -338
rect -5234 -372 -5218 -338
rect -5284 -388 -5218 -372
rect -5166 -338 -5100 -322
rect -5166 -372 -5150 -338
rect -5116 -372 -5100 -338
rect -5166 -388 -5100 -372
rect -5048 -338 -4982 -322
rect -5048 -372 -5032 -338
rect -4998 -372 -4982 -338
rect -5048 -388 -4982 -372
rect -4930 -338 -4864 -322
rect -4930 -372 -4914 -338
rect -4880 -372 -4864 -338
rect -4930 -388 -4864 -372
rect -4812 -338 -4746 -322
rect -4812 -372 -4796 -338
rect -4762 -372 -4746 -338
rect -4812 -388 -4746 -372
rect -4694 -338 -4628 -322
rect -4694 -372 -4678 -338
rect -4644 -372 -4628 -338
rect -4694 -388 -4628 -372
rect -4576 -338 -4510 -322
rect -4576 -372 -4560 -338
rect -4526 -372 -4510 -338
rect -4576 -388 -4510 -372
rect -4458 -338 -4392 -322
rect -4458 -372 -4442 -338
rect -4408 -372 -4392 -338
rect -4458 -388 -4392 -372
rect -4340 -338 -4274 -322
rect -4340 -372 -4324 -338
rect -4290 -372 -4274 -338
rect -4340 -388 -4274 -372
rect -4222 -338 -4156 -322
rect -4222 -372 -4206 -338
rect -4172 -372 -4156 -338
rect -4222 -388 -4156 -372
rect -4104 -338 -4038 -322
rect -4104 -372 -4088 -338
rect -4054 -372 -4038 -338
rect -4104 -388 -4038 -372
rect -3986 -338 -3920 -322
rect -3986 -372 -3970 -338
rect -3936 -372 -3920 -338
rect -3986 -388 -3920 -372
rect -3868 -338 -3802 -322
rect -3868 -372 -3852 -338
rect -3818 -372 -3802 -338
rect -3868 -388 -3802 -372
rect -3750 -338 -3684 -322
rect -3750 -372 -3734 -338
rect -3700 -372 -3684 -338
rect -3750 -388 -3684 -372
rect -3632 -338 -3566 -322
rect -3632 -372 -3616 -338
rect -3582 -372 -3566 -338
rect -3632 -388 -3566 -372
rect -3514 -338 -3448 -322
rect -3514 -372 -3498 -338
rect -3464 -372 -3448 -338
rect -3514 -388 -3448 -372
rect -3396 -338 -3330 -322
rect -3396 -372 -3380 -338
rect -3346 -372 -3330 -338
rect -3396 -388 -3330 -372
rect -3278 -338 -3212 -322
rect -3278 -372 -3262 -338
rect -3228 -372 -3212 -338
rect -3278 -388 -3212 -372
rect -3160 -338 -3094 -322
rect -3160 -372 -3144 -338
rect -3110 -372 -3094 -338
rect -3160 -388 -3094 -372
rect -3042 -338 -2976 -322
rect -3042 -372 -3026 -338
rect -2992 -372 -2976 -338
rect -3042 -388 -2976 -372
rect -2924 -338 -2858 -322
rect -2924 -372 -2908 -338
rect -2874 -372 -2858 -338
rect -2924 -388 -2858 -372
rect -2806 -338 -2740 -322
rect -2806 -372 -2790 -338
rect -2756 -372 -2740 -338
rect -2806 -388 -2740 -372
rect -2688 -338 -2622 -322
rect -2688 -372 -2672 -338
rect -2638 -372 -2622 -338
rect -2688 -388 -2622 -372
rect -2570 -338 -2504 -322
rect -2570 -372 -2554 -338
rect -2520 -372 -2504 -338
rect -2570 -388 -2504 -372
rect -2452 -338 -2386 -322
rect -2452 -372 -2436 -338
rect -2402 -372 -2386 -338
rect -2452 -388 -2386 -372
rect -2334 -338 -2268 -322
rect -2334 -372 -2318 -338
rect -2284 -372 -2268 -338
rect -2334 -388 -2268 -372
rect -2216 -338 -2150 -322
rect -2216 -372 -2200 -338
rect -2166 -372 -2150 -338
rect -2216 -388 -2150 -372
rect -2098 -338 -2032 -322
rect -2098 -372 -2082 -338
rect -2048 -372 -2032 -338
rect -2098 -388 -2032 -372
rect -1980 -338 -1914 -322
rect -1980 -372 -1964 -338
rect -1930 -372 -1914 -338
rect -1980 -388 -1914 -372
rect -1862 -338 -1796 -322
rect -1862 -372 -1846 -338
rect -1812 -372 -1796 -338
rect -1862 -388 -1796 -372
rect -1744 -338 -1678 -322
rect -1744 -372 -1728 -338
rect -1694 -372 -1678 -338
rect -1744 -388 -1678 -372
rect -1626 -338 -1560 -322
rect -1626 -372 -1610 -338
rect -1576 -372 -1560 -338
rect -1626 -388 -1560 -372
rect -1508 -338 -1442 -322
rect -1508 -372 -1492 -338
rect -1458 -372 -1442 -338
rect -1508 -388 -1442 -372
rect -1390 -338 -1324 -322
rect -1390 -372 -1374 -338
rect -1340 -372 -1324 -338
rect -1390 -388 -1324 -372
rect -1272 -338 -1206 -322
rect -1272 -372 -1256 -338
rect -1222 -372 -1206 -338
rect -1272 -388 -1206 -372
rect -1154 -338 -1088 -322
rect -1154 -372 -1138 -338
rect -1104 -372 -1088 -338
rect -1154 -388 -1088 -372
rect -1036 -338 -970 -322
rect -1036 -372 -1020 -338
rect -986 -372 -970 -338
rect -1036 -388 -970 -372
rect -918 -338 -852 -322
rect -918 -372 -902 -338
rect -868 -372 -852 -338
rect -918 -388 -852 -372
rect -800 -338 -734 -322
rect -800 -372 -784 -338
rect -750 -372 -734 -338
rect -800 -388 -734 -372
rect -682 -338 -616 -322
rect -682 -372 -666 -338
rect -632 -372 -616 -338
rect -682 -388 -616 -372
rect -564 -338 -498 -322
rect -564 -372 -548 -338
rect -514 -372 -498 -338
rect -564 -388 -498 -372
rect -446 -338 -380 -322
rect -446 -372 -430 -338
rect -396 -372 -380 -338
rect -446 -388 -380 -372
rect -328 -338 -262 -322
rect -328 -372 -312 -338
rect -278 -372 -262 -338
rect -328 -388 -262 -372
rect -210 -338 -144 -322
rect -210 -372 -194 -338
rect -160 -372 -144 -338
rect -210 -388 -144 -372
rect -92 -338 -26 -322
rect -92 -372 -76 -338
rect -42 -372 -26 -338
rect -92 -388 -26 -372
rect 26 -338 92 -322
rect 26 -372 42 -338
rect 76 -372 92 -338
rect 26 -388 92 -372
rect 144 -338 210 -322
rect 144 -372 160 -338
rect 194 -372 210 -338
rect 144 -388 210 -372
rect 262 -338 328 -322
rect 262 -372 278 -338
rect 312 -372 328 -338
rect 262 -388 328 -372
rect 380 -338 446 -322
rect 380 -372 396 -338
rect 430 -372 446 -338
rect 380 -388 446 -372
rect 498 -338 564 -322
rect 498 -372 514 -338
rect 548 -372 564 -338
rect 498 -388 564 -372
rect 616 -338 682 -322
rect 616 -372 632 -338
rect 666 -372 682 -338
rect 616 -388 682 -372
rect 734 -338 800 -322
rect 734 -372 750 -338
rect 784 -372 800 -338
rect 734 -388 800 -372
rect 852 -338 918 -322
rect 852 -372 868 -338
rect 902 -372 918 -338
rect 852 -388 918 -372
rect 970 -338 1036 -322
rect 970 -372 986 -338
rect 1020 -372 1036 -338
rect 970 -388 1036 -372
rect 1088 -338 1154 -322
rect 1088 -372 1104 -338
rect 1138 -372 1154 -338
rect 1088 -388 1154 -372
rect 1206 -338 1272 -322
rect 1206 -372 1222 -338
rect 1256 -372 1272 -338
rect 1206 -388 1272 -372
rect 1324 -338 1390 -322
rect 1324 -372 1340 -338
rect 1374 -372 1390 -338
rect 1324 -388 1390 -372
rect 1442 -338 1508 -322
rect 1442 -372 1458 -338
rect 1492 -372 1508 -338
rect 1442 -388 1508 -372
rect 1560 -338 1626 -322
rect 1560 -372 1576 -338
rect 1610 -372 1626 -338
rect 1560 -388 1626 -372
rect 1678 -338 1744 -322
rect 1678 -372 1694 -338
rect 1728 -372 1744 -338
rect 1678 -388 1744 -372
rect 1796 -338 1862 -322
rect 1796 -372 1812 -338
rect 1846 -372 1862 -338
rect 1796 -388 1862 -372
rect 1914 -338 1980 -322
rect 1914 -372 1930 -338
rect 1964 -372 1980 -338
rect 1914 -388 1980 -372
rect 2032 -338 2098 -322
rect 2032 -372 2048 -338
rect 2082 -372 2098 -338
rect 2032 -388 2098 -372
rect 2150 -338 2216 -322
rect 2150 -372 2166 -338
rect 2200 -372 2216 -338
rect 2150 -388 2216 -372
rect 2268 -338 2334 -322
rect 2268 -372 2284 -338
rect 2318 -372 2334 -338
rect 2268 -388 2334 -372
rect 2386 -338 2452 -322
rect 2386 -372 2402 -338
rect 2436 -372 2452 -338
rect 2386 -388 2452 -372
rect 2504 -338 2570 -322
rect 2504 -372 2520 -338
rect 2554 -372 2570 -338
rect 2504 -388 2570 -372
rect 2622 -338 2688 -322
rect 2622 -372 2638 -338
rect 2672 -372 2688 -338
rect 2622 -388 2688 -372
rect 2740 -338 2806 -322
rect 2740 -372 2756 -338
rect 2790 -372 2806 -338
rect 2740 -388 2806 -372
rect 2858 -338 2924 -322
rect 2858 -372 2874 -338
rect 2908 -372 2924 -338
rect 2858 -388 2924 -372
rect 2976 -338 3042 -322
rect 2976 -372 2992 -338
rect 3026 -372 3042 -338
rect 2976 -388 3042 -372
rect 3094 -338 3160 -322
rect 3094 -372 3110 -338
rect 3144 -372 3160 -338
rect 3094 -388 3160 -372
rect 3212 -338 3278 -322
rect 3212 -372 3228 -338
rect 3262 -372 3278 -338
rect 3212 -388 3278 -372
rect 3330 -338 3396 -322
rect 3330 -372 3346 -338
rect 3380 -372 3396 -338
rect 3330 -388 3396 -372
rect 3448 -338 3514 -322
rect 3448 -372 3464 -338
rect 3498 -372 3514 -338
rect 3448 -388 3514 -372
rect 3566 -338 3632 -322
rect 3566 -372 3582 -338
rect 3616 -372 3632 -338
rect 3566 -388 3632 -372
rect 3684 -338 3750 -322
rect 3684 -372 3700 -338
rect 3734 -372 3750 -338
rect 3684 -388 3750 -372
rect 3802 -338 3868 -322
rect 3802 -372 3818 -338
rect 3852 -372 3868 -338
rect 3802 -388 3868 -372
rect 3920 -338 3986 -322
rect 3920 -372 3936 -338
rect 3970 -372 3986 -338
rect 3920 -388 3986 -372
rect 4038 -338 4104 -322
rect 4038 -372 4054 -338
rect 4088 -372 4104 -338
rect 4038 -388 4104 -372
rect 4156 -338 4222 -322
rect 4156 -372 4172 -338
rect 4206 -372 4222 -338
rect 4156 -388 4222 -372
rect 4274 -338 4340 -322
rect 4274 -372 4290 -338
rect 4324 -372 4340 -338
rect 4274 -388 4340 -372
rect 4392 -338 4458 -322
rect 4392 -372 4408 -338
rect 4442 -372 4458 -338
rect 4392 -388 4458 -372
rect 4510 -338 4576 -322
rect 4510 -372 4526 -338
rect 4560 -372 4576 -338
rect 4510 -388 4576 -372
rect 4628 -338 4694 -322
rect 4628 -372 4644 -338
rect 4678 -372 4694 -338
rect 4628 -388 4694 -372
rect 4746 -338 4812 -322
rect 4746 -372 4762 -338
rect 4796 -372 4812 -338
rect 4746 -388 4812 -372
rect 4864 -338 4930 -322
rect 4864 -372 4880 -338
rect 4914 -372 4930 -338
rect 4864 -388 4930 -372
rect 4982 -338 5048 -322
rect 4982 -372 4998 -338
rect 5032 -372 5048 -338
rect 4982 -388 5048 -372
rect 5100 -338 5166 -322
rect 5100 -372 5116 -338
rect 5150 -372 5166 -338
rect 5100 -388 5166 -372
rect 5218 -338 5284 -322
rect 5218 -372 5234 -338
rect 5268 -372 5284 -338
rect 5218 -388 5284 -372
rect 5336 -338 5402 -322
rect 5336 -372 5352 -338
rect 5386 -372 5402 -338
rect 5336 -388 5402 -372
rect 5454 -338 5520 -322
rect 5454 -372 5470 -338
rect 5504 -372 5520 -338
rect 5454 -388 5520 -372
rect 5572 -338 5638 -322
rect 5572 -372 5588 -338
rect 5622 -372 5638 -338
rect 5572 -388 5638 -372
rect 5690 -338 5756 -322
rect 5690 -372 5706 -338
rect 5740 -372 5756 -338
rect 5690 -388 5756 -372
rect 5808 -338 5874 -322
rect 5808 -372 5824 -338
rect 5858 -372 5874 -338
rect 5808 -388 5874 -372
<< polycont >>
rect -5858 338 -5824 372
rect -5740 338 -5706 372
rect -5622 338 -5588 372
rect -5504 338 -5470 372
rect -5386 338 -5352 372
rect -5268 338 -5234 372
rect -5150 338 -5116 372
rect -5032 338 -4998 372
rect -4914 338 -4880 372
rect -4796 338 -4762 372
rect -4678 338 -4644 372
rect -4560 338 -4526 372
rect -4442 338 -4408 372
rect -4324 338 -4290 372
rect -4206 338 -4172 372
rect -4088 338 -4054 372
rect -3970 338 -3936 372
rect -3852 338 -3818 372
rect -3734 338 -3700 372
rect -3616 338 -3582 372
rect -3498 338 -3464 372
rect -3380 338 -3346 372
rect -3262 338 -3228 372
rect -3144 338 -3110 372
rect -3026 338 -2992 372
rect -2908 338 -2874 372
rect -2790 338 -2756 372
rect -2672 338 -2638 372
rect -2554 338 -2520 372
rect -2436 338 -2402 372
rect -2318 338 -2284 372
rect -2200 338 -2166 372
rect -2082 338 -2048 372
rect -1964 338 -1930 372
rect -1846 338 -1812 372
rect -1728 338 -1694 372
rect -1610 338 -1576 372
rect -1492 338 -1458 372
rect -1374 338 -1340 372
rect -1256 338 -1222 372
rect -1138 338 -1104 372
rect -1020 338 -986 372
rect -902 338 -868 372
rect -784 338 -750 372
rect -666 338 -632 372
rect -548 338 -514 372
rect -430 338 -396 372
rect -312 338 -278 372
rect -194 338 -160 372
rect -76 338 -42 372
rect 42 338 76 372
rect 160 338 194 372
rect 278 338 312 372
rect 396 338 430 372
rect 514 338 548 372
rect 632 338 666 372
rect 750 338 784 372
rect 868 338 902 372
rect 986 338 1020 372
rect 1104 338 1138 372
rect 1222 338 1256 372
rect 1340 338 1374 372
rect 1458 338 1492 372
rect 1576 338 1610 372
rect 1694 338 1728 372
rect 1812 338 1846 372
rect 1930 338 1964 372
rect 2048 338 2082 372
rect 2166 338 2200 372
rect 2284 338 2318 372
rect 2402 338 2436 372
rect 2520 338 2554 372
rect 2638 338 2672 372
rect 2756 338 2790 372
rect 2874 338 2908 372
rect 2992 338 3026 372
rect 3110 338 3144 372
rect 3228 338 3262 372
rect 3346 338 3380 372
rect 3464 338 3498 372
rect 3582 338 3616 372
rect 3700 338 3734 372
rect 3818 338 3852 372
rect 3936 338 3970 372
rect 4054 338 4088 372
rect 4172 338 4206 372
rect 4290 338 4324 372
rect 4408 338 4442 372
rect 4526 338 4560 372
rect 4644 338 4678 372
rect 4762 338 4796 372
rect 4880 338 4914 372
rect 4998 338 5032 372
rect 5116 338 5150 372
rect 5234 338 5268 372
rect 5352 338 5386 372
rect 5470 338 5504 372
rect 5588 338 5622 372
rect 5706 338 5740 372
rect 5824 338 5858 372
rect -5858 -372 -5824 -338
rect -5740 -372 -5706 -338
rect -5622 -372 -5588 -338
rect -5504 -372 -5470 -338
rect -5386 -372 -5352 -338
rect -5268 -372 -5234 -338
rect -5150 -372 -5116 -338
rect -5032 -372 -4998 -338
rect -4914 -372 -4880 -338
rect -4796 -372 -4762 -338
rect -4678 -372 -4644 -338
rect -4560 -372 -4526 -338
rect -4442 -372 -4408 -338
rect -4324 -372 -4290 -338
rect -4206 -372 -4172 -338
rect -4088 -372 -4054 -338
rect -3970 -372 -3936 -338
rect -3852 -372 -3818 -338
rect -3734 -372 -3700 -338
rect -3616 -372 -3582 -338
rect -3498 -372 -3464 -338
rect -3380 -372 -3346 -338
rect -3262 -372 -3228 -338
rect -3144 -372 -3110 -338
rect -3026 -372 -2992 -338
rect -2908 -372 -2874 -338
rect -2790 -372 -2756 -338
rect -2672 -372 -2638 -338
rect -2554 -372 -2520 -338
rect -2436 -372 -2402 -338
rect -2318 -372 -2284 -338
rect -2200 -372 -2166 -338
rect -2082 -372 -2048 -338
rect -1964 -372 -1930 -338
rect -1846 -372 -1812 -338
rect -1728 -372 -1694 -338
rect -1610 -372 -1576 -338
rect -1492 -372 -1458 -338
rect -1374 -372 -1340 -338
rect -1256 -372 -1222 -338
rect -1138 -372 -1104 -338
rect -1020 -372 -986 -338
rect -902 -372 -868 -338
rect -784 -372 -750 -338
rect -666 -372 -632 -338
rect -548 -372 -514 -338
rect -430 -372 -396 -338
rect -312 -372 -278 -338
rect -194 -372 -160 -338
rect -76 -372 -42 -338
rect 42 -372 76 -338
rect 160 -372 194 -338
rect 278 -372 312 -338
rect 396 -372 430 -338
rect 514 -372 548 -338
rect 632 -372 666 -338
rect 750 -372 784 -338
rect 868 -372 902 -338
rect 986 -372 1020 -338
rect 1104 -372 1138 -338
rect 1222 -372 1256 -338
rect 1340 -372 1374 -338
rect 1458 -372 1492 -338
rect 1576 -372 1610 -338
rect 1694 -372 1728 -338
rect 1812 -372 1846 -338
rect 1930 -372 1964 -338
rect 2048 -372 2082 -338
rect 2166 -372 2200 -338
rect 2284 -372 2318 -338
rect 2402 -372 2436 -338
rect 2520 -372 2554 -338
rect 2638 -372 2672 -338
rect 2756 -372 2790 -338
rect 2874 -372 2908 -338
rect 2992 -372 3026 -338
rect 3110 -372 3144 -338
rect 3228 -372 3262 -338
rect 3346 -372 3380 -338
rect 3464 -372 3498 -338
rect 3582 -372 3616 -338
rect 3700 -372 3734 -338
rect 3818 -372 3852 -338
rect 3936 -372 3970 -338
rect 4054 -372 4088 -338
rect 4172 -372 4206 -338
rect 4290 -372 4324 -338
rect 4408 -372 4442 -338
rect 4526 -372 4560 -338
rect 4644 -372 4678 -338
rect 4762 -372 4796 -338
rect 4880 -372 4914 -338
rect 4998 -372 5032 -338
rect 5116 -372 5150 -338
rect 5234 -372 5268 -338
rect 5352 -372 5386 -338
rect 5470 -372 5504 -338
rect 5588 -372 5622 -338
rect 5706 -372 5740 -338
rect 5824 -372 5858 -338
<< locali >>
rect -5874 338 -5858 372
rect -5824 338 -5808 372
rect -5756 338 -5740 372
rect -5706 338 -5690 372
rect -5638 338 -5622 372
rect -5588 338 -5572 372
rect -5520 338 -5504 372
rect -5470 338 -5454 372
rect -5402 338 -5386 372
rect -5352 338 -5336 372
rect -5284 338 -5268 372
rect -5234 338 -5218 372
rect -5166 338 -5150 372
rect -5116 338 -5100 372
rect -5048 338 -5032 372
rect -4998 338 -4982 372
rect -4930 338 -4914 372
rect -4880 338 -4864 372
rect -4812 338 -4796 372
rect -4762 338 -4746 372
rect -4694 338 -4678 372
rect -4644 338 -4628 372
rect -4576 338 -4560 372
rect -4526 338 -4510 372
rect -4458 338 -4442 372
rect -4408 338 -4392 372
rect -4340 338 -4324 372
rect -4290 338 -4274 372
rect -4222 338 -4206 372
rect -4172 338 -4156 372
rect -4104 338 -4088 372
rect -4054 338 -4038 372
rect -3986 338 -3970 372
rect -3936 338 -3920 372
rect -3868 338 -3852 372
rect -3818 338 -3802 372
rect -3750 338 -3734 372
rect -3700 338 -3684 372
rect -3632 338 -3616 372
rect -3582 338 -3566 372
rect -3514 338 -3498 372
rect -3464 338 -3448 372
rect -3396 338 -3380 372
rect -3346 338 -3330 372
rect -3278 338 -3262 372
rect -3228 338 -3212 372
rect -3160 338 -3144 372
rect -3110 338 -3094 372
rect -3042 338 -3026 372
rect -2992 338 -2976 372
rect -2924 338 -2908 372
rect -2874 338 -2858 372
rect -2806 338 -2790 372
rect -2756 338 -2740 372
rect -2688 338 -2672 372
rect -2638 338 -2622 372
rect -2570 338 -2554 372
rect -2520 338 -2504 372
rect -2452 338 -2436 372
rect -2402 338 -2386 372
rect -2334 338 -2318 372
rect -2284 338 -2268 372
rect -2216 338 -2200 372
rect -2166 338 -2150 372
rect -2098 338 -2082 372
rect -2048 338 -2032 372
rect -1980 338 -1964 372
rect -1930 338 -1914 372
rect -1862 338 -1846 372
rect -1812 338 -1796 372
rect -1744 338 -1728 372
rect -1694 338 -1678 372
rect -1626 338 -1610 372
rect -1576 338 -1560 372
rect -1508 338 -1492 372
rect -1458 338 -1442 372
rect -1390 338 -1374 372
rect -1340 338 -1324 372
rect -1272 338 -1256 372
rect -1222 338 -1206 372
rect -1154 338 -1138 372
rect -1104 338 -1088 372
rect -1036 338 -1020 372
rect -986 338 -970 372
rect -918 338 -902 372
rect -868 338 -852 372
rect -800 338 -784 372
rect -750 338 -734 372
rect -682 338 -666 372
rect -632 338 -616 372
rect -564 338 -548 372
rect -514 338 -498 372
rect -446 338 -430 372
rect -396 338 -380 372
rect -328 338 -312 372
rect -278 338 -262 372
rect -210 338 -194 372
rect -160 338 -144 372
rect -92 338 -76 372
rect -42 338 -26 372
rect 26 338 42 372
rect 76 338 92 372
rect 144 338 160 372
rect 194 338 210 372
rect 262 338 278 372
rect 312 338 328 372
rect 380 338 396 372
rect 430 338 446 372
rect 498 338 514 372
rect 548 338 564 372
rect 616 338 632 372
rect 666 338 682 372
rect 734 338 750 372
rect 784 338 800 372
rect 852 338 868 372
rect 902 338 918 372
rect 970 338 986 372
rect 1020 338 1036 372
rect 1088 338 1104 372
rect 1138 338 1154 372
rect 1206 338 1222 372
rect 1256 338 1272 372
rect 1324 338 1340 372
rect 1374 338 1390 372
rect 1442 338 1458 372
rect 1492 338 1508 372
rect 1560 338 1576 372
rect 1610 338 1626 372
rect 1678 338 1694 372
rect 1728 338 1744 372
rect 1796 338 1812 372
rect 1846 338 1862 372
rect 1914 338 1930 372
rect 1964 338 1980 372
rect 2032 338 2048 372
rect 2082 338 2098 372
rect 2150 338 2166 372
rect 2200 338 2216 372
rect 2268 338 2284 372
rect 2318 338 2334 372
rect 2386 338 2402 372
rect 2436 338 2452 372
rect 2504 338 2520 372
rect 2554 338 2570 372
rect 2622 338 2638 372
rect 2672 338 2688 372
rect 2740 338 2756 372
rect 2790 338 2806 372
rect 2858 338 2874 372
rect 2908 338 2924 372
rect 2976 338 2992 372
rect 3026 338 3042 372
rect 3094 338 3110 372
rect 3144 338 3160 372
rect 3212 338 3228 372
rect 3262 338 3278 372
rect 3330 338 3346 372
rect 3380 338 3396 372
rect 3448 338 3464 372
rect 3498 338 3514 372
rect 3566 338 3582 372
rect 3616 338 3632 372
rect 3684 338 3700 372
rect 3734 338 3750 372
rect 3802 338 3818 372
rect 3852 338 3868 372
rect 3920 338 3936 372
rect 3970 338 3986 372
rect 4038 338 4054 372
rect 4088 338 4104 372
rect 4156 338 4172 372
rect 4206 338 4222 372
rect 4274 338 4290 372
rect 4324 338 4340 372
rect 4392 338 4408 372
rect 4442 338 4458 372
rect 4510 338 4526 372
rect 4560 338 4576 372
rect 4628 338 4644 372
rect 4678 338 4694 372
rect 4746 338 4762 372
rect 4796 338 4812 372
rect 4864 338 4880 372
rect 4914 338 4930 372
rect 4982 338 4998 372
rect 5032 338 5048 372
rect 5100 338 5116 372
rect 5150 338 5166 372
rect 5218 338 5234 372
rect 5268 338 5284 372
rect 5336 338 5352 372
rect 5386 338 5402 372
rect 5454 338 5470 372
rect 5504 338 5520 372
rect 5572 338 5588 372
rect 5622 338 5638 372
rect 5690 338 5706 372
rect 5740 338 5756 372
rect 5808 338 5824 372
rect 5858 338 5874 372
rect -5917 288 -5883 304
rect -5917 -304 -5883 -288
rect -5799 288 -5765 304
rect -5799 -304 -5765 -288
rect -5681 288 -5647 304
rect -5681 -304 -5647 -288
rect -5563 288 -5529 304
rect -5563 -304 -5529 -288
rect -5445 288 -5411 304
rect -5445 -304 -5411 -288
rect -5327 288 -5293 304
rect -5327 -304 -5293 -288
rect -5209 288 -5175 304
rect -5209 -304 -5175 -288
rect -5091 288 -5057 304
rect -5091 -304 -5057 -288
rect -4973 288 -4939 304
rect -4973 -304 -4939 -288
rect -4855 288 -4821 304
rect -4855 -304 -4821 -288
rect -4737 288 -4703 304
rect -4737 -304 -4703 -288
rect -4619 288 -4585 304
rect -4619 -304 -4585 -288
rect -4501 288 -4467 304
rect -4501 -304 -4467 -288
rect -4383 288 -4349 304
rect -4383 -304 -4349 -288
rect -4265 288 -4231 304
rect -4265 -304 -4231 -288
rect -4147 288 -4113 304
rect -4147 -304 -4113 -288
rect -4029 288 -3995 304
rect -4029 -304 -3995 -288
rect -3911 288 -3877 304
rect -3911 -304 -3877 -288
rect -3793 288 -3759 304
rect -3793 -304 -3759 -288
rect -3675 288 -3641 304
rect -3675 -304 -3641 -288
rect -3557 288 -3523 304
rect -3557 -304 -3523 -288
rect -3439 288 -3405 304
rect -3439 -304 -3405 -288
rect -3321 288 -3287 304
rect -3321 -304 -3287 -288
rect -3203 288 -3169 304
rect -3203 -304 -3169 -288
rect -3085 288 -3051 304
rect -3085 -304 -3051 -288
rect -2967 288 -2933 304
rect -2967 -304 -2933 -288
rect -2849 288 -2815 304
rect -2849 -304 -2815 -288
rect -2731 288 -2697 304
rect -2731 -304 -2697 -288
rect -2613 288 -2579 304
rect -2613 -304 -2579 -288
rect -2495 288 -2461 304
rect -2495 -304 -2461 -288
rect -2377 288 -2343 304
rect -2377 -304 -2343 -288
rect -2259 288 -2225 304
rect -2259 -304 -2225 -288
rect -2141 288 -2107 304
rect -2141 -304 -2107 -288
rect -2023 288 -1989 304
rect -2023 -304 -1989 -288
rect -1905 288 -1871 304
rect -1905 -304 -1871 -288
rect -1787 288 -1753 304
rect -1787 -304 -1753 -288
rect -1669 288 -1635 304
rect -1669 -304 -1635 -288
rect -1551 288 -1517 304
rect -1551 -304 -1517 -288
rect -1433 288 -1399 304
rect -1433 -304 -1399 -288
rect -1315 288 -1281 304
rect -1315 -304 -1281 -288
rect -1197 288 -1163 304
rect -1197 -304 -1163 -288
rect -1079 288 -1045 304
rect -1079 -304 -1045 -288
rect -961 288 -927 304
rect -961 -304 -927 -288
rect -843 288 -809 304
rect -843 -304 -809 -288
rect -725 288 -691 304
rect -725 -304 -691 -288
rect -607 288 -573 304
rect -607 -304 -573 -288
rect -489 288 -455 304
rect -489 -304 -455 -288
rect -371 288 -337 304
rect -371 -304 -337 -288
rect -253 288 -219 304
rect -253 -304 -219 -288
rect -135 288 -101 304
rect -135 -304 -101 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 101 288 135 304
rect 101 -304 135 -288
rect 219 288 253 304
rect 219 -304 253 -288
rect 337 288 371 304
rect 337 -304 371 -288
rect 455 288 489 304
rect 455 -304 489 -288
rect 573 288 607 304
rect 573 -304 607 -288
rect 691 288 725 304
rect 691 -304 725 -288
rect 809 288 843 304
rect 809 -304 843 -288
rect 927 288 961 304
rect 927 -304 961 -288
rect 1045 288 1079 304
rect 1045 -304 1079 -288
rect 1163 288 1197 304
rect 1163 -304 1197 -288
rect 1281 288 1315 304
rect 1281 -304 1315 -288
rect 1399 288 1433 304
rect 1399 -304 1433 -288
rect 1517 288 1551 304
rect 1517 -304 1551 -288
rect 1635 288 1669 304
rect 1635 -304 1669 -288
rect 1753 288 1787 304
rect 1753 -304 1787 -288
rect 1871 288 1905 304
rect 1871 -304 1905 -288
rect 1989 288 2023 304
rect 1989 -304 2023 -288
rect 2107 288 2141 304
rect 2107 -304 2141 -288
rect 2225 288 2259 304
rect 2225 -304 2259 -288
rect 2343 288 2377 304
rect 2343 -304 2377 -288
rect 2461 288 2495 304
rect 2461 -304 2495 -288
rect 2579 288 2613 304
rect 2579 -304 2613 -288
rect 2697 288 2731 304
rect 2697 -304 2731 -288
rect 2815 288 2849 304
rect 2815 -304 2849 -288
rect 2933 288 2967 304
rect 2933 -304 2967 -288
rect 3051 288 3085 304
rect 3051 -304 3085 -288
rect 3169 288 3203 304
rect 3169 -304 3203 -288
rect 3287 288 3321 304
rect 3287 -304 3321 -288
rect 3405 288 3439 304
rect 3405 -304 3439 -288
rect 3523 288 3557 304
rect 3523 -304 3557 -288
rect 3641 288 3675 304
rect 3641 -304 3675 -288
rect 3759 288 3793 304
rect 3759 -304 3793 -288
rect 3877 288 3911 304
rect 3877 -304 3911 -288
rect 3995 288 4029 304
rect 3995 -304 4029 -288
rect 4113 288 4147 304
rect 4113 -304 4147 -288
rect 4231 288 4265 304
rect 4231 -304 4265 -288
rect 4349 288 4383 304
rect 4349 -304 4383 -288
rect 4467 288 4501 304
rect 4467 -304 4501 -288
rect 4585 288 4619 304
rect 4585 -304 4619 -288
rect 4703 288 4737 304
rect 4703 -304 4737 -288
rect 4821 288 4855 304
rect 4821 -304 4855 -288
rect 4939 288 4973 304
rect 4939 -304 4973 -288
rect 5057 288 5091 304
rect 5057 -304 5091 -288
rect 5175 288 5209 304
rect 5175 -304 5209 -288
rect 5293 288 5327 304
rect 5293 -304 5327 -288
rect 5411 288 5445 304
rect 5411 -304 5445 -288
rect 5529 288 5563 304
rect 5529 -304 5563 -288
rect 5647 288 5681 304
rect 5647 -304 5681 -288
rect 5765 288 5799 304
rect 5765 -304 5799 -288
rect 5883 288 5917 304
rect 5883 -304 5917 -288
rect -5874 -372 -5858 -338
rect -5824 -372 -5808 -338
rect -5756 -372 -5740 -338
rect -5706 -372 -5690 -338
rect -5638 -372 -5622 -338
rect -5588 -372 -5572 -338
rect -5520 -372 -5504 -338
rect -5470 -372 -5454 -338
rect -5402 -372 -5386 -338
rect -5352 -372 -5336 -338
rect -5284 -372 -5268 -338
rect -5234 -372 -5218 -338
rect -5166 -372 -5150 -338
rect -5116 -372 -5100 -338
rect -5048 -372 -5032 -338
rect -4998 -372 -4982 -338
rect -4930 -372 -4914 -338
rect -4880 -372 -4864 -338
rect -4812 -372 -4796 -338
rect -4762 -372 -4746 -338
rect -4694 -372 -4678 -338
rect -4644 -372 -4628 -338
rect -4576 -372 -4560 -338
rect -4526 -372 -4510 -338
rect -4458 -372 -4442 -338
rect -4408 -372 -4392 -338
rect -4340 -372 -4324 -338
rect -4290 -372 -4274 -338
rect -4222 -372 -4206 -338
rect -4172 -372 -4156 -338
rect -4104 -372 -4088 -338
rect -4054 -372 -4038 -338
rect -3986 -372 -3970 -338
rect -3936 -372 -3920 -338
rect -3868 -372 -3852 -338
rect -3818 -372 -3802 -338
rect -3750 -372 -3734 -338
rect -3700 -372 -3684 -338
rect -3632 -372 -3616 -338
rect -3582 -372 -3566 -338
rect -3514 -372 -3498 -338
rect -3464 -372 -3448 -338
rect -3396 -372 -3380 -338
rect -3346 -372 -3330 -338
rect -3278 -372 -3262 -338
rect -3228 -372 -3212 -338
rect -3160 -372 -3144 -338
rect -3110 -372 -3094 -338
rect -3042 -372 -3026 -338
rect -2992 -372 -2976 -338
rect -2924 -372 -2908 -338
rect -2874 -372 -2858 -338
rect -2806 -372 -2790 -338
rect -2756 -372 -2740 -338
rect -2688 -372 -2672 -338
rect -2638 -372 -2622 -338
rect -2570 -372 -2554 -338
rect -2520 -372 -2504 -338
rect -2452 -372 -2436 -338
rect -2402 -372 -2386 -338
rect -2334 -372 -2318 -338
rect -2284 -372 -2268 -338
rect -2216 -372 -2200 -338
rect -2166 -372 -2150 -338
rect -2098 -372 -2082 -338
rect -2048 -372 -2032 -338
rect -1980 -372 -1964 -338
rect -1930 -372 -1914 -338
rect -1862 -372 -1846 -338
rect -1812 -372 -1796 -338
rect -1744 -372 -1728 -338
rect -1694 -372 -1678 -338
rect -1626 -372 -1610 -338
rect -1576 -372 -1560 -338
rect -1508 -372 -1492 -338
rect -1458 -372 -1442 -338
rect -1390 -372 -1374 -338
rect -1340 -372 -1324 -338
rect -1272 -372 -1256 -338
rect -1222 -372 -1206 -338
rect -1154 -372 -1138 -338
rect -1104 -372 -1088 -338
rect -1036 -372 -1020 -338
rect -986 -372 -970 -338
rect -918 -372 -902 -338
rect -868 -372 -852 -338
rect -800 -372 -784 -338
rect -750 -372 -734 -338
rect -682 -372 -666 -338
rect -632 -372 -616 -338
rect -564 -372 -548 -338
rect -514 -372 -498 -338
rect -446 -372 -430 -338
rect -396 -372 -380 -338
rect -328 -372 -312 -338
rect -278 -372 -262 -338
rect -210 -372 -194 -338
rect -160 -372 -144 -338
rect -92 -372 -76 -338
rect -42 -372 -26 -338
rect 26 -372 42 -338
rect 76 -372 92 -338
rect 144 -372 160 -338
rect 194 -372 210 -338
rect 262 -372 278 -338
rect 312 -372 328 -338
rect 380 -372 396 -338
rect 430 -372 446 -338
rect 498 -372 514 -338
rect 548 -372 564 -338
rect 616 -372 632 -338
rect 666 -372 682 -338
rect 734 -372 750 -338
rect 784 -372 800 -338
rect 852 -372 868 -338
rect 902 -372 918 -338
rect 970 -372 986 -338
rect 1020 -372 1036 -338
rect 1088 -372 1104 -338
rect 1138 -372 1154 -338
rect 1206 -372 1222 -338
rect 1256 -372 1272 -338
rect 1324 -372 1340 -338
rect 1374 -372 1390 -338
rect 1442 -372 1458 -338
rect 1492 -372 1508 -338
rect 1560 -372 1576 -338
rect 1610 -372 1626 -338
rect 1678 -372 1694 -338
rect 1728 -372 1744 -338
rect 1796 -372 1812 -338
rect 1846 -372 1862 -338
rect 1914 -372 1930 -338
rect 1964 -372 1980 -338
rect 2032 -372 2048 -338
rect 2082 -372 2098 -338
rect 2150 -372 2166 -338
rect 2200 -372 2216 -338
rect 2268 -372 2284 -338
rect 2318 -372 2334 -338
rect 2386 -372 2402 -338
rect 2436 -372 2452 -338
rect 2504 -372 2520 -338
rect 2554 -372 2570 -338
rect 2622 -372 2638 -338
rect 2672 -372 2688 -338
rect 2740 -372 2756 -338
rect 2790 -372 2806 -338
rect 2858 -372 2874 -338
rect 2908 -372 2924 -338
rect 2976 -372 2992 -338
rect 3026 -372 3042 -338
rect 3094 -372 3110 -338
rect 3144 -372 3160 -338
rect 3212 -372 3228 -338
rect 3262 -372 3278 -338
rect 3330 -372 3346 -338
rect 3380 -372 3396 -338
rect 3448 -372 3464 -338
rect 3498 -372 3514 -338
rect 3566 -372 3582 -338
rect 3616 -372 3632 -338
rect 3684 -372 3700 -338
rect 3734 -372 3750 -338
rect 3802 -372 3818 -338
rect 3852 -372 3868 -338
rect 3920 -372 3936 -338
rect 3970 -372 3986 -338
rect 4038 -372 4054 -338
rect 4088 -372 4104 -338
rect 4156 -372 4172 -338
rect 4206 -372 4222 -338
rect 4274 -372 4290 -338
rect 4324 -372 4340 -338
rect 4392 -372 4408 -338
rect 4442 -372 4458 -338
rect 4510 -372 4526 -338
rect 4560 -372 4576 -338
rect 4628 -372 4644 -338
rect 4678 -372 4694 -338
rect 4746 -372 4762 -338
rect 4796 -372 4812 -338
rect 4864 -372 4880 -338
rect 4914 -372 4930 -338
rect 4982 -372 4998 -338
rect 5032 -372 5048 -338
rect 5100 -372 5116 -338
rect 5150 -372 5166 -338
rect 5218 -372 5234 -338
rect 5268 -372 5284 -338
rect 5336 -372 5352 -338
rect 5386 -372 5402 -338
rect 5454 -372 5470 -338
rect 5504 -372 5520 -338
rect 5572 -372 5588 -338
rect 5622 -372 5638 -338
rect 5690 -372 5706 -338
rect 5740 -372 5756 -338
rect 5808 -372 5824 -338
rect 5858 -372 5874 -338
<< viali >>
rect -5858 338 -5824 372
rect -5740 338 -5706 372
rect -5622 338 -5588 372
rect -5504 338 -5470 372
rect -5386 338 -5352 372
rect -5268 338 -5234 372
rect -5150 338 -5116 372
rect -5032 338 -4998 372
rect -4914 338 -4880 372
rect -4796 338 -4762 372
rect -4678 338 -4644 372
rect -4560 338 -4526 372
rect -4442 338 -4408 372
rect -4324 338 -4290 372
rect -4206 338 -4172 372
rect -4088 338 -4054 372
rect -3970 338 -3936 372
rect -3852 338 -3818 372
rect -3734 338 -3700 372
rect -3616 338 -3582 372
rect -3498 338 -3464 372
rect -3380 338 -3346 372
rect -3262 338 -3228 372
rect -3144 338 -3110 372
rect -3026 338 -2992 372
rect -2908 338 -2874 372
rect -2790 338 -2756 372
rect -2672 338 -2638 372
rect -2554 338 -2520 372
rect -2436 338 -2402 372
rect -2318 338 -2284 372
rect -2200 338 -2166 372
rect -2082 338 -2048 372
rect -1964 338 -1930 372
rect -1846 338 -1812 372
rect -1728 338 -1694 372
rect -1610 338 -1576 372
rect -1492 338 -1458 372
rect -1374 338 -1340 372
rect -1256 338 -1222 372
rect -1138 338 -1104 372
rect -1020 338 -986 372
rect -902 338 -868 372
rect -784 338 -750 372
rect -666 338 -632 372
rect -548 338 -514 372
rect -430 338 -396 372
rect -312 338 -278 372
rect -194 338 -160 372
rect -76 338 -42 372
rect 42 338 76 372
rect 160 338 194 372
rect 278 338 312 372
rect 396 338 430 372
rect 514 338 548 372
rect 632 338 666 372
rect 750 338 784 372
rect 868 338 902 372
rect 986 338 1020 372
rect 1104 338 1138 372
rect 1222 338 1256 372
rect 1340 338 1374 372
rect 1458 338 1492 372
rect 1576 338 1610 372
rect 1694 338 1728 372
rect 1812 338 1846 372
rect 1930 338 1964 372
rect 2048 338 2082 372
rect 2166 338 2200 372
rect 2284 338 2318 372
rect 2402 338 2436 372
rect 2520 338 2554 372
rect 2638 338 2672 372
rect 2756 338 2790 372
rect 2874 338 2908 372
rect 2992 338 3026 372
rect 3110 338 3144 372
rect 3228 338 3262 372
rect 3346 338 3380 372
rect 3464 338 3498 372
rect 3582 338 3616 372
rect 3700 338 3734 372
rect 3818 338 3852 372
rect 3936 338 3970 372
rect 4054 338 4088 372
rect 4172 338 4206 372
rect 4290 338 4324 372
rect 4408 338 4442 372
rect 4526 338 4560 372
rect 4644 338 4678 372
rect 4762 338 4796 372
rect 4880 338 4914 372
rect 4998 338 5032 372
rect 5116 338 5150 372
rect 5234 338 5268 372
rect 5352 338 5386 372
rect 5470 338 5504 372
rect 5588 338 5622 372
rect 5706 338 5740 372
rect 5824 338 5858 372
rect -5917 -288 -5883 288
rect -5799 -288 -5765 288
rect -5681 -288 -5647 288
rect -5563 -288 -5529 288
rect -5445 -288 -5411 288
rect -5327 -288 -5293 288
rect -5209 -288 -5175 288
rect -5091 -288 -5057 288
rect -4973 -288 -4939 288
rect -4855 -288 -4821 288
rect -4737 -288 -4703 288
rect -4619 -288 -4585 288
rect -4501 -288 -4467 288
rect -4383 -288 -4349 288
rect -4265 -288 -4231 288
rect -4147 -288 -4113 288
rect -4029 -288 -3995 288
rect -3911 -288 -3877 288
rect -3793 -288 -3759 288
rect -3675 -288 -3641 288
rect -3557 -288 -3523 288
rect -3439 -288 -3405 288
rect -3321 -288 -3287 288
rect -3203 -288 -3169 288
rect -3085 -288 -3051 288
rect -2967 -288 -2933 288
rect -2849 -288 -2815 288
rect -2731 -288 -2697 288
rect -2613 -288 -2579 288
rect -2495 -288 -2461 288
rect -2377 -288 -2343 288
rect -2259 -288 -2225 288
rect -2141 -288 -2107 288
rect -2023 -288 -1989 288
rect -1905 -288 -1871 288
rect -1787 -288 -1753 288
rect -1669 -288 -1635 288
rect -1551 -288 -1517 288
rect -1433 -288 -1399 288
rect -1315 -288 -1281 288
rect -1197 -288 -1163 288
rect -1079 -288 -1045 288
rect -961 -288 -927 288
rect -843 -288 -809 288
rect -725 -288 -691 288
rect -607 -288 -573 288
rect -489 -288 -455 288
rect -371 -288 -337 288
rect -253 -288 -219 288
rect -135 -288 -101 288
rect -17 -288 17 288
rect 101 -288 135 288
rect 219 -288 253 288
rect 337 -288 371 288
rect 455 -288 489 288
rect 573 -288 607 288
rect 691 -288 725 288
rect 809 -288 843 288
rect 927 -288 961 288
rect 1045 -288 1079 288
rect 1163 -288 1197 288
rect 1281 -288 1315 288
rect 1399 -288 1433 288
rect 1517 -288 1551 288
rect 1635 -288 1669 288
rect 1753 -288 1787 288
rect 1871 -288 1905 288
rect 1989 -288 2023 288
rect 2107 -288 2141 288
rect 2225 -288 2259 288
rect 2343 -288 2377 288
rect 2461 -288 2495 288
rect 2579 -288 2613 288
rect 2697 -288 2731 288
rect 2815 -288 2849 288
rect 2933 -288 2967 288
rect 3051 -288 3085 288
rect 3169 -288 3203 288
rect 3287 -288 3321 288
rect 3405 -288 3439 288
rect 3523 -288 3557 288
rect 3641 -288 3675 288
rect 3759 -288 3793 288
rect 3877 -288 3911 288
rect 3995 -288 4029 288
rect 4113 -288 4147 288
rect 4231 -288 4265 288
rect 4349 -288 4383 288
rect 4467 -288 4501 288
rect 4585 -288 4619 288
rect 4703 -288 4737 288
rect 4821 -288 4855 288
rect 4939 -288 4973 288
rect 5057 -288 5091 288
rect 5175 -288 5209 288
rect 5293 -288 5327 288
rect 5411 -288 5445 288
rect 5529 -288 5563 288
rect 5647 -288 5681 288
rect 5765 -288 5799 288
rect 5883 -288 5917 288
rect -5858 -372 -5824 -338
rect -5740 -372 -5706 -338
rect -5622 -372 -5588 -338
rect -5504 -372 -5470 -338
rect -5386 -372 -5352 -338
rect -5268 -372 -5234 -338
rect -5150 -372 -5116 -338
rect -5032 -372 -4998 -338
rect -4914 -372 -4880 -338
rect -4796 -372 -4762 -338
rect -4678 -372 -4644 -338
rect -4560 -372 -4526 -338
rect -4442 -372 -4408 -338
rect -4324 -372 -4290 -338
rect -4206 -372 -4172 -338
rect -4088 -372 -4054 -338
rect -3970 -372 -3936 -338
rect -3852 -372 -3818 -338
rect -3734 -372 -3700 -338
rect -3616 -372 -3582 -338
rect -3498 -372 -3464 -338
rect -3380 -372 -3346 -338
rect -3262 -372 -3228 -338
rect -3144 -372 -3110 -338
rect -3026 -372 -2992 -338
rect -2908 -372 -2874 -338
rect -2790 -372 -2756 -338
rect -2672 -372 -2638 -338
rect -2554 -372 -2520 -338
rect -2436 -372 -2402 -338
rect -2318 -372 -2284 -338
rect -2200 -372 -2166 -338
rect -2082 -372 -2048 -338
rect -1964 -372 -1930 -338
rect -1846 -372 -1812 -338
rect -1728 -372 -1694 -338
rect -1610 -372 -1576 -338
rect -1492 -372 -1458 -338
rect -1374 -372 -1340 -338
rect -1256 -372 -1222 -338
rect -1138 -372 -1104 -338
rect -1020 -372 -986 -338
rect -902 -372 -868 -338
rect -784 -372 -750 -338
rect -666 -372 -632 -338
rect -548 -372 -514 -338
rect -430 -372 -396 -338
rect -312 -372 -278 -338
rect -194 -372 -160 -338
rect -76 -372 -42 -338
rect 42 -372 76 -338
rect 160 -372 194 -338
rect 278 -372 312 -338
rect 396 -372 430 -338
rect 514 -372 548 -338
rect 632 -372 666 -338
rect 750 -372 784 -338
rect 868 -372 902 -338
rect 986 -372 1020 -338
rect 1104 -372 1138 -338
rect 1222 -372 1256 -338
rect 1340 -372 1374 -338
rect 1458 -372 1492 -338
rect 1576 -372 1610 -338
rect 1694 -372 1728 -338
rect 1812 -372 1846 -338
rect 1930 -372 1964 -338
rect 2048 -372 2082 -338
rect 2166 -372 2200 -338
rect 2284 -372 2318 -338
rect 2402 -372 2436 -338
rect 2520 -372 2554 -338
rect 2638 -372 2672 -338
rect 2756 -372 2790 -338
rect 2874 -372 2908 -338
rect 2992 -372 3026 -338
rect 3110 -372 3144 -338
rect 3228 -372 3262 -338
rect 3346 -372 3380 -338
rect 3464 -372 3498 -338
rect 3582 -372 3616 -338
rect 3700 -372 3734 -338
rect 3818 -372 3852 -338
rect 3936 -372 3970 -338
rect 4054 -372 4088 -338
rect 4172 -372 4206 -338
rect 4290 -372 4324 -338
rect 4408 -372 4442 -338
rect 4526 -372 4560 -338
rect 4644 -372 4678 -338
rect 4762 -372 4796 -338
rect 4880 -372 4914 -338
rect 4998 -372 5032 -338
rect 5116 -372 5150 -338
rect 5234 -372 5268 -338
rect 5352 -372 5386 -338
rect 5470 -372 5504 -338
rect 5588 -372 5622 -338
rect 5706 -372 5740 -338
rect 5824 -372 5858 -338
<< metal1 >>
rect -5870 372 -5812 378
rect -5870 338 -5858 372
rect -5824 338 -5812 372
rect -5870 332 -5812 338
rect -5752 372 -5694 378
rect -5752 338 -5740 372
rect -5706 338 -5694 372
rect -5752 332 -5694 338
rect -5634 372 -5576 378
rect -5634 338 -5622 372
rect -5588 338 -5576 372
rect -5634 332 -5576 338
rect -5516 372 -5458 378
rect -5516 338 -5504 372
rect -5470 338 -5458 372
rect -5516 332 -5458 338
rect -5398 372 -5340 378
rect -5398 338 -5386 372
rect -5352 338 -5340 372
rect -5398 332 -5340 338
rect -5280 372 -5222 378
rect -5280 338 -5268 372
rect -5234 338 -5222 372
rect -5280 332 -5222 338
rect -5162 372 -5104 378
rect -5162 338 -5150 372
rect -5116 338 -5104 372
rect -5162 332 -5104 338
rect -5044 372 -4986 378
rect -5044 338 -5032 372
rect -4998 338 -4986 372
rect -5044 332 -4986 338
rect -4926 372 -4868 378
rect -4926 338 -4914 372
rect -4880 338 -4868 372
rect -4926 332 -4868 338
rect -4808 372 -4750 378
rect -4808 338 -4796 372
rect -4762 338 -4750 372
rect -4808 332 -4750 338
rect -4690 372 -4632 378
rect -4690 338 -4678 372
rect -4644 338 -4632 372
rect -4690 332 -4632 338
rect -4572 372 -4514 378
rect -4572 338 -4560 372
rect -4526 338 -4514 372
rect -4572 332 -4514 338
rect -4454 372 -4396 378
rect -4454 338 -4442 372
rect -4408 338 -4396 372
rect -4454 332 -4396 338
rect -4336 372 -4278 378
rect -4336 338 -4324 372
rect -4290 338 -4278 372
rect -4336 332 -4278 338
rect -4218 372 -4160 378
rect -4218 338 -4206 372
rect -4172 338 -4160 372
rect -4218 332 -4160 338
rect -4100 372 -4042 378
rect -4100 338 -4088 372
rect -4054 338 -4042 372
rect -4100 332 -4042 338
rect -3982 372 -3924 378
rect -3982 338 -3970 372
rect -3936 338 -3924 372
rect -3982 332 -3924 338
rect -3864 372 -3806 378
rect -3864 338 -3852 372
rect -3818 338 -3806 372
rect -3864 332 -3806 338
rect -3746 372 -3688 378
rect -3746 338 -3734 372
rect -3700 338 -3688 372
rect -3746 332 -3688 338
rect -3628 372 -3570 378
rect -3628 338 -3616 372
rect -3582 338 -3570 372
rect -3628 332 -3570 338
rect -3510 372 -3452 378
rect -3510 338 -3498 372
rect -3464 338 -3452 372
rect -3510 332 -3452 338
rect -3392 372 -3334 378
rect -3392 338 -3380 372
rect -3346 338 -3334 372
rect -3392 332 -3334 338
rect -3274 372 -3216 378
rect -3274 338 -3262 372
rect -3228 338 -3216 372
rect -3274 332 -3216 338
rect -3156 372 -3098 378
rect -3156 338 -3144 372
rect -3110 338 -3098 372
rect -3156 332 -3098 338
rect -3038 372 -2980 378
rect -3038 338 -3026 372
rect -2992 338 -2980 372
rect -3038 332 -2980 338
rect -2920 372 -2862 378
rect -2920 338 -2908 372
rect -2874 338 -2862 372
rect -2920 332 -2862 338
rect -2802 372 -2744 378
rect -2802 338 -2790 372
rect -2756 338 -2744 372
rect -2802 332 -2744 338
rect -2684 372 -2626 378
rect -2684 338 -2672 372
rect -2638 338 -2626 372
rect -2684 332 -2626 338
rect -2566 372 -2508 378
rect -2566 338 -2554 372
rect -2520 338 -2508 372
rect -2566 332 -2508 338
rect -2448 372 -2390 378
rect -2448 338 -2436 372
rect -2402 338 -2390 372
rect -2448 332 -2390 338
rect -2330 372 -2272 378
rect -2330 338 -2318 372
rect -2284 338 -2272 372
rect -2330 332 -2272 338
rect -2212 372 -2154 378
rect -2212 338 -2200 372
rect -2166 338 -2154 372
rect -2212 332 -2154 338
rect -2094 372 -2036 378
rect -2094 338 -2082 372
rect -2048 338 -2036 372
rect -2094 332 -2036 338
rect -1976 372 -1918 378
rect -1976 338 -1964 372
rect -1930 338 -1918 372
rect -1976 332 -1918 338
rect -1858 372 -1800 378
rect -1858 338 -1846 372
rect -1812 338 -1800 372
rect -1858 332 -1800 338
rect -1740 372 -1682 378
rect -1740 338 -1728 372
rect -1694 338 -1682 372
rect -1740 332 -1682 338
rect -1622 372 -1564 378
rect -1622 338 -1610 372
rect -1576 338 -1564 372
rect -1622 332 -1564 338
rect -1504 372 -1446 378
rect -1504 338 -1492 372
rect -1458 338 -1446 372
rect -1504 332 -1446 338
rect -1386 372 -1328 378
rect -1386 338 -1374 372
rect -1340 338 -1328 372
rect -1386 332 -1328 338
rect -1268 372 -1210 378
rect -1268 338 -1256 372
rect -1222 338 -1210 372
rect -1268 332 -1210 338
rect -1150 372 -1092 378
rect -1150 338 -1138 372
rect -1104 338 -1092 372
rect -1150 332 -1092 338
rect -1032 372 -974 378
rect -1032 338 -1020 372
rect -986 338 -974 372
rect -1032 332 -974 338
rect -914 372 -856 378
rect -914 338 -902 372
rect -868 338 -856 372
rect -914 332 -856 338
rect -796 372 -738 378
rect -796 338 -784 372
rect -750 338 -738 372
rect -796 332 -738 338
rect -678 372 -620 378
rect -678 338 -666 372
rect -632 338 -620 372
rect -678 332 -620 338
rect -560 372 -502 378
rect -560 338 -548 372
rect -514 338 -502 372
rect -560 332 -502 338
rect -442 372 -384 378
rect -442 338 -430 372
rect -396 338 -384 372
rect -442 332 -384 338
rect -324 372 -266 378
rect -324 338 -312 372
rect -278 338 -266 372
rect -324 332 -266 338
rect -206 372 -148 378
rect -206 338 -194 372
rect -160 338 -148 372
rect -206 332 -148 338
rect -88 372 -30 378
rect -88 338 -76 372
rect -42 338 -30 372
rect -88 332 -30 338
rect 30 372 88 378
rect 30 338 42 372
rect 76 338 88 372
rect 30 332 88 338
rect 148 372 206 378
rect 148 338 160 372
rect 194 338 206 372
rect 148 332 206 338
rect 266 372 324 378
rect 266 338 278 372
rect 312 338 324 372
rect 266 332 324 338
rect 384 372 442 378
rect 384 338 396 372
rect 430 338 442 372
rect 384 332 442 338
rect 502 372 560 378
rect 502 338 514 372
rect 548 338 560 372
rect 502 332 560 338
rect 620 372 678 378
rect 620 338 632 372
rect 666 338 678 372
rect 620 332 678 338
rect 738 372 796 378
rect 738 338 750 372
rect 784 338 796 372
rect 738 332 796 338
rect 856 372 914 378
rect 856 338 868 372
rect 902 338 914 372
rect 856 332 914 338
rect 974 372 1032 378
rect 974 338 986 372
rect 1020 338 1032 372
rect 974 332 1032 338
rect 1092 372 1150 378
rect 1092 338 1104 372
rect 1138 338 1150 372
rect 1092 332 1150 338
rect 1210 372 1268 378
rect 1210 338 1222 372
rect 1256 338 1268 372
rect 1210 332 1268 338
rect 1328 372 1386 378
rect 1328 338 1340 372
rect 1374 338 1386 372
rect 1328 332 1386 338
rect 1446 372 1504 378
rect 1446 338 1458 372
rect 1492 338 1504 372
rect 1446 332 1504 338
rect 1564 372 1622 378
rect 1564 338 1576 372
rect 1610 338 1622 372
rect 1564 332 1622 338
rect 1682 372 1740 378
rect 1682 338 1694 372
rect 1728 338 1740 372
rect 1682 332 1740 338
rect 1800 372 1858 378
rect 1800 338 1812 372
rect 1846 338 1858 372
rect 1800 332 1858 338
rect 1918 372 1976 378
rect 1918 338 1930 372
rect 1964 338 1976 372
rect 1918 332 1976 338
rect 2036 372 2094 378
rect 2036 338 2048 372
rect 2082 338 2094 372
rect 2036 332 2094 338
rect 2154 372 2212 378
rect 2154 338 2166 372
rect 2200 338 2212 372
rect 2154 332 2212 338
rect 2272 372 2330 378
rect 2272 338 2284 372
rect 2318 338 2330 372
rect 2272 332 2330 338
rect 2390 372 2448 378
rect 2390 338 2402 372
rect 2436 338 2448 372
rect 2390 332 2448 338
rect 2508 372 2566 378
rect 2508 338 2520 372
rect 2554 338 2566 372
rect 2508 332 2566 338
rect 2626 372 2684 378
rect 2626 338 2638 372
rect 2672 338 2684 372
rect 2626 332 2684 338
rect 2744 372 2802 378
rect 2744 338 2756 372
rect 2790 338 2802 372
rect 2744 332 2802 338
rect 2862 372 2920 378
rect 2862 338 2874 372
rect 2908 338 2920 372
rect 2862 332 2920 338
rect 2980 372 3038 378
rect 2980 338 2992 372
rect 3026 338 3038 372
rect 2980 332 3038 338
rect 3098 372 3156 378
rect 3098 338 3110 372
rect 3144 338 3156 372
rect 3098 332 3156 338
rect 3216 372 3274 378
rect 3216 338 3228 372
rect 3262 338 3274 372
rect 3216 332 3274 338
rect 3334 372 3392 378
rect 3334 338 3346 372
rect 3380 338 3392 372
rect 3334 332 3392 338
rect 3452 372 3510 378
rect 3452 338 3464 372
rect 3498 338 3510 372
rect 3452 332 3510 338
rect 3570 372 3628 378
rect 3570 338 3582 372
rect 3616 338 3628 372
rect 3570 332 3628 338
rect 3688 372 3746 378
rect 3688 338 3700 372
rect 3734 338 3746 372
rect 3688 332 3746 338
rect 3806 372 3864 378
rect 3806 338 3818 372
rect 3852 338 3864 372
rect 3806 332 3864 338
rect 3924 372 3982 378
rect 3924 338 3936 372
rect 3970 338 3982 372
rect 3924 332 3982 338
rect 4042 372 4100 378
rect 4042 338 4054 372
rect 4088 338 4100 372
rect 4042 332 4100 338
rect 4160 372 4218 378
rect 4160 338 4172 372
rect 4206 338 4218 372
rect 4160 332 4218 338
rect 4278 372 4336 378
rect 4278 338 4290 372
rect 4324 338 4336 372
rect 4278 332 4336 338
rect 4396 372 4454 378
rect 4396 338 4408 372
rect 4442 338 4454 372
rect 4396 332 4454 338
rect 4514 372 4572 378
rect 4514 338 4526 372
rect 4560 338 4572 372
rect 4514 332 4572 338
rect 4632 372 4690 378
rect 4632 338 4644 372
rect 4678 338 4690 372
rect 4632 332 4690 338
rect 4750 372 4808 378
rect 4750 338 4762 372
rect 4796 338 4808 372
rect 4750 332 4808 338
rect 4868 372 4926 378
rect 4868 338 4880 372
rect 4914 338 4926 372
rect 4868 332 4926 338
rect 4986 372 5044 378
rect 4986 338 4998 372
rect 5032 338 5044 372
rect 4986 332 5044 338
rect 5104 372 5162 378
rect 5104 338 5116 372
rect 5150 338 5162 372
rect 5104 332 5162 338
rect 5222 372 5280 378
rect 5222 338 5234 372
rect 5268 338 5280 372
rect 5222 332 5280 338
rect 5340 372 5398 378
rect 5340 338 5352 372
rect 5386 338 5398 372
rect 5340 332 5398 338
rect 5458 372 5516 378
rect 5458 338 5470 372
rect 5504 338 5516 372
rect 5458 332 5516 338
rect 5576 372 5634 378
rect 5576 338 5588 372
rect 5622 338 5634 372
rect 5576 332 5634 338
rect 5694 372 5752 378
rect 5694 338 5706 372
rect 5740 338 5752 372
rect 5694 332 5752 338
rect 5812 372 5870 378
rect 5812 338 5824 372
rect 5858 338 5870 372
rect 5812 332 5870 338
rect -5923 288 -5877 300
rect -5923 -288 -5917 288
rect -5883 -288 -5877 288
rect -5923 -300 -5877 -288
rect -5805 288 -5759 300
rect -5805 -288 -5799 288
rect -5765 -288 -5759 288
rect -5805 -300 -5759 -288
rect -5687 288 -5641 300
rect -5687 -288 -5681 288
rect -5647 -288 -5641 288
rect -5687 -300 -5641 -288
rect -5569 288 -5523 300
rect -5569 -288 -5563 288
rect -5529 -288 -5523 288
rect -5569 -300 -5523 -288
rect -5451 288 -5405 300
rect -5451 -288 -5445 288
rect -5411 -288 -5405 288
rect -5451 -300 -5405 -288
rect -5333 288 -5287 300
rect -5333 -288 -5327 288
rect -5293 -288 -5287 288
rect -5333 -300 -5287 -288
rect -5215 288 -5169 300
rect -5215 -288 -5209 288
rect -5175 -288 -5169 288
rect -5215 -300 -5169 -288
rect -5097 288 -5051 300
rect -5097 -288 -5091 288
rect -5057 -288 -5051 288
rect -5097 -300 -5051 -288
rect -4979 288 -4933 300
rect -4979 -288 -4973 288
rect -4939 -288 -4933 288
rect -4979 -300 -4933 -288
rect -4861 288 -4815 300
rect -4861 -288 -4855 288
rect -4821 -288 -4815 288
rect -4861 -300 -4815 -288
rect -4743 288 -4697 300
rect -4743 -288 -4737 288
rect -4703 -288 -4697 288
rect -4743 -300 -4697 -288
rect -4625 288 -4579 300
rect -4625 -288 -4619 288
rect -4585 -288 -4579 288
rect -4625 -300 -4579 -288
rect -4507 288 -4461 300
rect -4507 -288 -4501 288
rect -4467 -288 -4461 288
rect -4507 -300 -4461 -288
rect -4389 288 -4343 300
rect -4389 -288 -4383 288
rect -4349 -288 -4343 288
rect -4389 -300 -4343 -288
rect -4271 288 -4225 300
rect -4271 -288 -4265 288
rect -4231 -288 -4225 288
rect -4271 -300 -4225 -288
rect -4153 288 -4107 300
rect -4153 -288 -4147 288
rect -4113 -288 -4107 288
rect -4153 -300 -4107 -288
rect -4035 288 -3989 300
rect -4035 -288 -4029 288
rect -3995 -288 -3989 288
rect -4035 -300 -3989 -288
rect -3917 288 -3871 300
rect -3917 -288 -3911 288
rect -3877 -288 -3871 288
rect -3917 -300 -3871 -288
rect -3799 288 -3753 300
rect -3799 -288 -3793 288
rect -3759 -288 -3753 288
rect -3799 -300 -3753 -288
rect -3681 288 -3635 300
rect -3681 -288 -3675 288
rect -3641 -288 -3635 288
rect -3681 -300 -3635 -288
rect -3563 288 -3517 300
rect -3563 -288 -3557 288
rect -3523 -288 -3517 288
rect -3563 -300 -3517 -288
rect -3445 288 -3399 300
rect -3445 -288 -3439 288
rect -3405 -288 -3399 288
rect -3445 -300 -3399 -288
rect -3327 288 -3281 300
rect -3327 -288 -3321 288
rect -3287 -288 -3281 288
rect -3327 -300 -3281 -288
rect -3209 288 -3163 300
rect -3209 -288 -3203 288
rect -3169 -288 -3163 288
rect -3209 -300 -3163 -288
rect -3091 288 -3045 300
rect -3091 -288 -3085 288
rect -3051 -288 -3045 288
rect -3091 -300 -3045 -288
rect -2973 288 -2927 300
rect -2973 -288 -2967 288
rect -2933 -288 -2927 288
rect -2973 -300 -2927 -288
rect -2855 288 -2809 300
rect -2855 -288 -2849 288
rect -2815 -288 -2809 288
rect -2855 -300 -2809 -288
rect -2737 288 -2691 300
rect -2737 -288 -2731 288
rect -2697 -288 -2691 288
rect -2737 -300 -2691 -288
rect -2619 288 -2573 300
rect -2619 -288 -2613 288
rect -2579 -288 -2573 288
rect -2619 -300 -2573 -288
rect -2501 288 -2455 300
rect -2501 -288 -2495 288
rect -2461 -288 -2455 288
rect -2501 -300 -2455 -288
rect -2383 288 -2337 300
rect -2383 -288 -2377 288
rect -2343 -288 -2337 288
rect -2383 -300 -2337 -288
rect -2265 288 -2219 300
rect -2265 -288 -2259 288
rect -2225 -288 -2219 288
rect -2265 -300 -2219 -288
rect -2147 288 -2101 300
rect -2147 -288 -2141 288
rect -2107 -288 -2101 288
rect -2147 -300 -2101 -288
rect -2029 288 -1983 300
rect -2029 -288 -2023 288
rect -1989 -288 -1983 288
rect -2029 -300 -1983 -288
rect -1911 288 -1865 300
rect -1911 -288 -1905 288
rect -1871 -288 -1865 288
rect -1911 -300 -1865 -288
rect -1793 288 -1747 300
rect -1793 -288 -1787 288
rect -1753 -288 -1747 288
rect -1793 -300 -1747 -288
rect -1675 288 -1629 300
rect -1675 -288 -1669 288
rect -1635 -288 -1629 288
rect -1675 -300 -1629 -288
rect -1557 288 -1511 300
rect -1557 -288 -1551 288
rect -1517 -288 -1511 288
rect -1557 -300 -1511 -288
rect -1439 288 -1393 300
rect -1439 -288 -1433 288
rect -1399 -288 -1393 288
rect -1439 -300 -1393 -288
rect -1321 288 -1275 300
rect -1321 -288 -1315 288
rect -1281 -288 -1275 288
rect -1321 -300 -1275 -288
rect -1203 288 -1157 300
rect -1203 -288 -1197 288
rect -1163 -288 -1157 288
rect -1203 -300 -1157 -288
rect -1085 288 -1039 300
rect -1085 -288 -1079 288
rect -1045 -288 -1039 288
rect -1085 -300 -1039 -288
rect -967 288 -921 300
rect -967 -288 -961 288
rect -927 -288 -921 288
rect -967 -300 -921 -288
rect -849 288 -803 300
rect -849 -288 -843 288
rect -809 -288 -803 288
rect -849 -300 -803 -288
rect -731 288 -685 300
rect -731 -288 -725 288
rect -691 -288 -685 288
rect -731 -300 -685 -288
rect -613 288 -567 300
rect -613 -288 -607 288
rect -573 -288 -567 288
rect -613 -300 -567 -288
rect -495 288 -449 300
rect -495 -288 -489 288
rect -455 -288 -449 288
rect -495 -300 -449 -288
rect -377 288 -331 300
rect -377 -288 -371 288
rect -337 -288 -331 288
rect -377 -300 -331 -288
rect -259 288 -213 300
rect -259 -288 -253 288
rect -219 -288 -213 288
rect -259 -300 -213 -288
rect -141 288 -95 300
rect -141 -288 -135 288
rect -101 -288 -95 288
rect -141 -300 -95 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 95 288 141 300
rect 95 -288 101 288
rect 135 -288 141 288
rect 95 -300 141 -288
rect 213 288 259 300
rect 213 -288 219 288
rect 253 -288 259 288
rect 213 -300 259 -288
rect 331 288 377 300
rect 331 -288 337 288
rect 371 -288 377 288
rect 331 -300 377 -288
rect 449 288 495 300
rect 449 -288 455 288
rect 489 -288 495 288
rect 449 -300 495 -288
rect 567 288 613 300
rect 567 -288 573 288
rect 607 -288 613 288
rect 567 -300 613 -288
rect 685 288 731 300
rect 685 -288 691 288
rect 725 -288 731 288
rect 685 -300 731 -288
rect 803 288 849 300
rect 803 -288 809 288
rect 843 -288 849 288
rect 803 -300 849 -288
rect 921 288 967 300
rect 921 -288 927 288
rect 961 -288 967 288
rect 921 -300 967 -288
rect 1039 288 1085 300
rect 1039 -288 1045 288
rect 1079 -288 1085 288
rect 1039 -300 1085 -288
rect 1157 288 1203 300
rect 1157 -288 1163 288
rect 1197 -288 1203 288
rect 1157 -300 1203 -288
rect 1275 288 1321 300
rect 1275 -288 1281 288
rect 1315 -288 1321 288
rect 1275 -300 1321 -288
rect 1393 288 1439 300
rect 1393 -288 1399 288
rect 1433 -288 1439 288
rect 1393 -300 1439 -288
rect 1511 288 1557 300
rect 1511 -288 1517 288
rect 1551 -288 1557 288
rect 1511 -300 1557 -288
rect 1629 288 1675 300
rect 1629 -288 1635 288
rect 1669 -288 1675 288
rect 1629 -300 1675 -288
rect 1747 288 1793 300
rect 1747 -288 1753 288
rect 1787 -288 1793 288
rect 1747 -300 1793 -288
rect 1865 288 1911 300
rect 1865 -288 1871 288
rect 1905 -288 1911 288
rect 1865 -300 1911 -288
rect 1983 288 2029 300
rect 1983 -288 1989 288
rect 2023 -288 2029 288
rect 1983 -300 2029 -288
rect 2101 288 2147 300
rect 2101 -288 2107 288
rect 2141 -288 2147 288
rect 2101 -300 2147 -288
rect 2219 288 2265 300
rect 2219 -288 2225 288
rect 2259 -288 2265 288
rect 2219 -300 2265 -288
rect 2337 288 2383 300
rect 2337 -288 2343 288
rect 2377 -288 2383 288
rect 2337 -300 2383 -288
rect 2455 288 2501 300
rect 2455 -288 2461 288
rect 2495 -288 2501 288
rect 2455 -300 2501 -288
rect 2573 288 2619 300
rect 2573 -288 2579 288
rect 2613 -288 2619 288
rect 2573 -300 2619 -288
rect 2691 288 2737 300
rect 2691 -288 2697 288
rect 2731 -288 2737 288
rect 2691 -300 2737 -288
rect 2809 288 2855 300
rect 2809 -288 2815 288
rect 2849 -288 2855 288
rect 2809 -300 2855 -288
rect 2927 288 2973 300
rect 2927 -288 2933 288
rect 2967 -288 2973 288
rect 2927 -300 2973 -288
rect 3045 288 3091 300
rect 3045 -288 3051 288
rect 3085 -288 3091 288
rect 3045 -300 3091 -288
rect 3163 288 3209 300
rect 3163 -288 3169 288
rect 3203 -288 3209 288
rect 3163 -300 3209 -288
rect 3281 288 3327 300
rect 3281 -288 3287 288
rect 3321 -288 3327 288
rect 3281 -300 3327 -288
rect 3399 288 3445 300
rect 3399 -288 3405 288
rect 3439 -288 3445 288
rect 3399 -300 3445 -288
rect 3517 288 3563 300
rect 3517 -288 3523 288
rect 3557 -288 3563 288
rect 3517 -300 3563 -288
rect 3635 288 3681 300
rect 3635 -288 3641 288
rect 3675 -288 3681 288
rect 3635 -300 3681 -288
rect 3753 288 3799 300
rect 3753 -288 3759 288
rect 3793 -288 3799 288
rect 3753 -300 3799 -288
rect 3871 288 3917 300
rect 3871 -288 3877 288
rect 3911 -288 3917 288
rect 3871 -300 3917 -288
rect 3989 288 4035 300
rect 3989 -288 3995 288
rect 4029 -288 4035 288
rect 3989 -300 4035 -288
rect 4107 288 4153 300
rect 4107 -288 4113 288
rect 4147 -288 4153 288
rect 4107 -300 4153 -288
rect 4225 288 4271 300
rect 4225 -288 4231 288
rect 4265 -288 4271 288
rect 4225 -300 4271 -288
rect 4343 288 4389 300
rect 4343 -288 4349 288
rect 4383 -288 4389 288
rect 4343 -300 4389 -288
rect 4461 288 4507 300
rect 4461 -288 4467 288
rect 4501 -288 4507 288
rect 4461 -300 4507 -288
rect 4579 288 4625 300
rect 4579 -288 4585 288
rect 4619 -288 4625 288
rect 4579 -300 4625 -288
rect 4697 288 4743 300
rect 4697 -288 4703 288
rect 4737 -288 4743 288
rect 4697 -300 4743 -288
rect 4815 288 4861 300
rect 4815 -288 4821 288
rect 4855 -288 4861 288
rect 4815 -300 4861 -288
rect 4933 288 4979 300
rect 4933 -288 4939 288
rect 4973 -288 4979 288
rect 4933 -300 4979 -288
rect 5051 288 5097 300
rect 5051 -288 5057 288
rect 5091 -288 5097 288
rect 5051 -300 5097 -288
rect 5169 288 5215 300
rect 5169 -288 5175 288
rect 5209 -288 5215 288
rect 5169 -300 5215 -288
rect 5287 288 5333 300
rect 5287 -288 5293 288
rect 5327 -288 5333 288
rect 5287 -300 5333 -288
rect 5405 288 5451 300
rect 5405 -288 5411 288
rect 5445 -288 5451 288
rect 5405 -300 5451 -288
rect 5523 288 5569 300
rect 5523 -288 5529 288
rect 5563 -288 5569 288
rect 5523 -300 5569 -288
rect 5641 288 5687 300
rect 5641 -288 5647 288
rect 5681 -288 5687 288
rect 5641 -300 5687 -288
rect 5759 288 5805 300
rect 5759 -288 5765 288
rect 5799 -288 5805 288
rect 5759 -300 5805 -288
rect 5877 288 5923 300
rect 5877 -288 5883 288
rect 5917 -288 5923 288
rect 5877 -300 5923 -288
rect -5870 -338 -5812 -332
rect -5870 -372 -5858 -338
rect -5824 -372 -5812 -338
rect -5870 -378 -5812 -372
rect -5752 -338 -5694 -332
rect -5752 -372 -5740 -338
rect -5706 -372 -5694 -338
rect -5752 -378 -5694 -372
rect -5634 -338 -5576 -332
rect -5634 -372 -5622 -338
rect -5588 -372 -5576 -338
rect -5634 -378 -5576 -372
rect -5516 -338 -5458 -332
rect -5516 -372 -5504 -338
rect -5470 -372 -5458 -338
rect -5516 -378 -5458 -372
rect -5398 -338 -5340 -332
rect -5398 -372 -5386 -338
rect -5352 -372 -5340 -338
rect -5398 -378 -5340 -372
rect -5280 -338 -5222 -332
rect -5280 -372 -5268 -338
rect -5234 -372 -5222 -338
rect -5280 -378 -5222 -372
rect -5162 -338 -5104 -332
rect -5162 -372 -5150 -338
rect -5116 -372 -5104 -338
rect -5162 -378 -5104 -372
rect -5044 -338 -4986 -332
rect -5044 -372 -5032 -338
rect -4998 -372 -4986 -338
rect -5044 -378 -4986 -372
rect -4926 -338 -4868 -332
rect -4926 -372 -4914 -338
rect -4880 -372 -4868 -338
rect -4926 -378 -4868 -372
rect -4808 -338 -4750 -332
rect -4808 -372 -4796 -338
rect -4762 -372 -4750 -338
rect -4808 -378 -4750 -372
rect -4690 -338 -4632 -332
rect -4690 -372 -4678 -338
rect -4644 -372 -4632 -338
rect -4690 -378 -4632 -372
rect -4572 -338 -4514 -332
rect -4572 -372 -4560 -338
rect -4526 -372 -4514 -338
rect -4572 -378 -4514 -372
rect -4454 -338 -4396 -332
rect -4454 -372 -4442 -338
rect -4408 -372 -4396 -338
rect -4454 -378 -4396 -372
rect -4336 -338 -4278 -332
rect -4336 -372 -4324 -338
rect -4290 -372 -4278 -338
rect -4336 -378 -4278 -372
rect -4218 -338 -4160 -332
rect -4218 -372 -4206 -338
rect -4172 -372 -4160 -338
rect -4218 -378 -4160 -372
rect -4100 -338 -4042 -332
rect -4100 -372 -4088 -338
rect -4054 -372 -4042 -338
rect -4100 -378 -4042 -372
rect -3982 -338 -3924 -332
rect -3982 -372 -3970 -338
rect -3936 -372 -3924 -338
rect -3982 -378 -3924 -372
rect -3864 -338 -3806 -332
rect -3864 -372 -3852 -338
rect -3818 -372 -3806 -338
rect -3864 -378 -3806 -372
rect -3746 -338 -3688 -332
rect -3746 -372 -3734 -338
rect -3700 -372 -3688 -338
rect -3746 -378 -3688 -372
rect -3628 -338 -3570 -332
rect -3628 -372 -3616 -338
rect -3582 -372 -3570 -338
rect -3628 -378 -3570 -372
rect -3510 -338 -3452 -332
rect -3510 -372 -3498 -338
rect -3464 -372 -3452 -338
rect -3510 -378 -3452 -372
rect -3392 -338 -3334 -332
rect -3392 -372 -3380 -338
rect -3346 -372 -3334 -338
rect -3392 -378 -3334 -372
rect -3274 -338 -3216 -332
rect -3274 -372 -3262 -338
rect -3228 -372 -3216 -338
rect -3274 -378 -3216 -372
rect -3156 -338 -3098 -332
rect -3156 -372 -3144 -338
rect -3110 -372 -3098 -338
rect -3156 -378 -3098 -372
rect -3038 -338 -2980 -332
rect -3038 -372 -3026 -338
rect -2992 -372 -2980 -338
rect -3038 -378 -2980 -372
rect -2920 -338 -2862 -332
rect -2920 -372 -2908 -338
rect -2874 -372 -2862 -338
rect -2920 -378 -2862 -372
rect -2802 -338 -2744 -332
rect -2802 -372 -2790 -338
rect -2756 -372 -2744 -338
rect -2802 -378 -2744 -372
rect -2684 -338 -2626 -332
rect -2684 -372 -2672 -338
rect -2638 -372 -2626 -338
rect -2684 -378 -2626 -372
rect -2566 -338 -2508 -332
rect -2566 -372 -2554 -338
rect -2520 -372 -2508 -338
rect -2566 -378 -2508 -372
rect -2448 -338 -2390 -332
rect -2448 -372 -2436 -338
rect -2402 -372 -2390 -338
rect -2448 -378 -2390 -372
rect -2330 -338 -2272 -332
rect -2330 -372 -2318 -338
rect -2284 -372 -2272 -338
rect -2330 -378 -2272 -372
rect -2212 -338 -2154 -332
rect -2212 -372 -2200 -338
rect -2166 -372 -2154 -338
rect -2212 -378 -2154 -372
rect -2094 -338 -2036 -332
rect -2094 -372 -2082 -338
rect -2048 -372 -2036 -338
rect -2094 -378 -2036 -372
rect -1976 -338 -1918 -332
rect -1976 -372 -1964 -338
rect -1930 -372 -1918 -338
rect -1976 -378 -1918 -372
rect -1858 -338 -1800 -332
rect -1858 -372 -1846 -338
rect -1812 -372 -1800 -338
rect -1858 -378 -1800 -372
rect -1740 -338 -1682 -332
rect -1740 -372 -1728 -338
rect -1694 -372 -1682 -338
rect -1740 -378 -1682 -372
rect -1622 -338 -1564 -332
rect -1622 -372 -1610 -338
rect -1576 -372 -1564 -338
rect -1622 -378 -1564 -372
rect -1504 -338 -1446 -332
rect -1504 -372 -1492 -338
rect -1458 -372 -1446 -338
rect -1504 -378 -1446 -372
rect -1386 -338 -1328 -332
rect -1386 -372 -1374 -338
rect -1340 -372 -1328 -338
rect -1386 -378 -1328 -372
rect -1268 -338 -1210 -332
rect -1268 -372 -1256 -338
rect -1222 -372 -1210 -338
rect -1268 -378 -1210 -372
rect -1150 -338 -1092 -332
rect -1150 -372 -1138 -338
rect -1104 -372 -1092 -338
rect -1150 -378 -1092 -372
rect -1032 -338 -974 -332
rect -1032 -372 -1020 -338
rect -986 -372 -974 -338
rect -1032 -378 -974 -372
rect -914 -338 -856 -332
rect -914 -372 -902 -338
rect -868 -372 -856 -338
rect -914 -378 -856 -372
rect -796 -338 -738 -332
rect -796 -372 -784 -338
rect -750 -372 -738 -338
rect -796 -378 -738 -372
rect -678 -338 -620 -332
rect -678 -372 -666 -338
rect -632 -372 -620 -338
rect -678 -378 -620 -372
rect -560 -338 -502 -332
rect -560 -372 -548 -338
rect -514 -372 -502 -338
rect -560 -378 -502 -372
rect -442 -338 -384 -332
rect -442 -372 -430 -338
rect -396 -372 -384 -338
rect -442 -378 -384 -372
rect -324 -338 -266 -332
rect -324 -372 -312 -338
rect -278 -372 -266 -338
rect -324 -378 -266 -372
rect -206 -338 -148 -332
rect -206 -372 -194 -338
rect -160 -372 -148 -338
rect -206 -378 -148 -372
rect -88 -338 -30 -332
rect -88 -372 -76 -338
rect -42 -372 -30 -338
rect -88 -378 -30 -372
rect 30 -338 88 -332
rect 30 -372 42 -338
rect 76 -372 88 -338
rect 30 -378 88 -372
rect 148 -338 206 -332
rect 148 -372 160 -338
rect 194 -372 206 -338
rect 148 -378 206 -372
rect 266 -338 324 -332
rect 266 -372 278 -338
rect 312 -372 324 -338
rect 266 -378 324 -372
rect 384 -338 442 -332
rect 384 -372 396 -338
rect 430 -372 442 -338
rect 384 -378 442 -372
rect 502 -338 560 -332
rect 502 -372 514 -338
rect 548 -372 560 -338
rect 502 -378 560 -372
rect 620 -338 678 -332
rect 620 -372 632 -338
rect 666 -372 678 -338
rect 620 -378 678 -372
rect 738 -338 796 -332
rect 738 -372 750 -338
rect 784 -372 796 -338
rect 738 -378 796 -372
rect 856 -338 914 -332
rect 856 -372 868 -338
rect 902 -372 914 -338
rect 856 -378 914 -372
rect 974 -338 1032 -332
rect 974 -372 986 -338
rect 1020 -372 1032 -338
rect 974 -378 1032 -372
rect 1092 -338 1150 -332
rect 1092 -372 1104 -338
rect 1138 -372 1150 -338
rect 1092 -378 1150 -372
rect 1210 -338 1268 -332
rect 1210 -372 1222 -338
rect 1256 -372 1268 -338
rect 1210 -378 1268 -372
rect 1328 -338 1386 -332
rect 1328 -372 1340 -338
rect 1374 -372 1386 -338
rect 1328 -378 1386 -372
rect 1446 -338 1504 -332
rect 1446 -372 1458 -338
rect 1492 -372 1504 -338
rect 1446 -378 1504 -372
rect 1564 -338 1622 -332
rect 1564 -372 1576 -338
rect 1610 -372 1622 -338
rect 1564 -378 1622 -372
rect 1682 -338 1740 -332
rect 1682 -372 1694 -338
rect 1728 -372 1740 -338
rect 1682 -378 1740 -372
rect 1800 -338 1858 -332
rect 1800 -372 1812 -338
rect 1846 -372 1858 -338
rect 1800 -378 1858 -372
rect 1918 -338 1976 -332
rect 1918 -372 1930 -338
rect 1964 -372 1976 -338
rect 1918 -378 1976 -372
rect 2036 -338 2094 -332
rect 2036 -372 2048 -338
rect 2082 -372 2094 -338
rect 2036 -378 2094 -372
rect 2154 -338 2212 -332
rect 2154 -372 2166 -338
rect 2200 -372 2212 -338
rect 2154 -378 2212 -372
rect 2272 -338 2330 -332
rect 2272 -372 2284 -338
rect 2318 -372 2330 -338
rect 2272 -378 2330 -372
rect 2390 -338 2448 -332
rect 2390 -372 2402 -338
rect 2436 -372 2448 -338
rect 2390 -378 2448 -372
rect 2508 -338 2566 -332
rect 2508 -372 2520 -338
rect 2554 -372 2566 -338
rect 2508 -378 2566 -372
rect 2626 -338 2684 -332
rect 2626 -372 2638 -338
rect 2672 -372 2684 -338
rect 2626 -378 2684 -372
rect 2744 -338 2802 -332
rect 2744 -372 2756 -338
rect 2790 -372 2802 -338
rect 2744 -378 2802 -372
rect 2862 -338 2920 -332
rect 2862 -372 2874 -338
rect 2908 -372 2920 -338
rect 2862 -378 2920 -372
rect 2980 -338 3038 -332
rect 2980 -372 2992 -338
rect 3026 -372 3038 -338
rect 2980 -378 3038 -372
rect 3098 -338 3156 -332
rect 3098 -372 3110 -338
rect 3144 -372 3156 -338
rect 3098 -378 3156 -372
rect 3216 -338 3274 -332
rect 3216 -372 3228 -338
rect 3262 -372 3274 -338
rect 3216 -378 3274 -372
rect 3334 -338 3392 -332
rect 3334 -372 3346 -338
rect 3380 -372 3392 -338
rect 3334 -378 3392 -372
rect 3452 -338 3510 -332
rect 3452 -372 3464 -338
rect 3498 -372 3510 -338
rect 3452 -378 3510 -372
rect 3570 -338 3628 -332
rect 3570 -372 3582 -338
rect 3616 -372 3628 -338
rect 3570 -378 3628 -372
rect 3688 -338 3746 -332
rect 3688 -372 3700 -338
rect 3734 -372 3746 -338
rect 3688 -378 3746 -372
rect 3806 -338 3864 -332
rect 3806 -372 3818 -338
rect 3852 -372 3864 -338
rect 3806 -378 3864 -372
rect 3924 -338 3982 -332
rect 3924 -372 3936 -338
rect 3970 -372 3982 -338
rect 3924 -378 3982 -372
rect 4042 -338 4100 -332
rect 4042 -372 4054 -338
rect 4088 -372 4100 -338
rect 4042 -378 4100 -372
rect 4160 -338 4218 -332
rect 4160 -372 4172 -338
rect 4206 -372 4218 -338
rect 4160 -378 4218 -372
rect 4278 -338 4336 -332
rect 4278 -372 4290 -338
rect 4324 -372 4336 -338
rect 4278 -378 4336 -372
rect 4396 -338 4454 -332
rect 4396 -372 4408 -338
rect 4442 -372 4454 -338
rect 4396 -378 4454 -372
rect 4514 -338 4572 -332
rect 4514 -372 4526 -338
rect 4560 -372 4572 -338
rect 4514 -378 4572 -372
rect 4632 -338 4690 -332
rect 4632 -372 4644 -338
rect 4678 -372 4690 -338
rect 4632 -378 4690 -372
rect 4750 -338 4808 -332
rect 4750 -372 4762 -338
rect 4796 -372 4808 -338
rect 4750 -378 4808 -372
rect 4868 -338 4926 -332
rect 4868 -372 4880 -338
rect 4914 -372 4926 -338
rect 4868 -378 4926 -372
rect 4986 -338 5044 -332
rect 4986 -372 4998 -338
rect 5032 -372 5044 -338
rect 4986 -378 5044 -372
rect 5104 -338 5162 -332
rect 5104 -372 5116 -338
rect 5150 -372 5162 -338
rect 5104 -378 5162 -372
rect 5222 -338 5280 -332
rect 5222 -372 5234 -338
rect 5268 -372 5280 -338
rect 5222 -378 5280 -372
rect 5340 -338 5398 -332
rect 5340 -372 5352 -338
rect 5386 -372 5398 -338
rect 5340 -378 5398 -372
rect 5458 -338 5516 -332
rect 5458 -372 5470 -338
rect 5504 -372 5516 -338
rect 5458 -378 5516 -372
rect 5576 -338 5634 -332
rect 5576 -372 5588 -338
rect 5622 -372 5634 -338
rect 5576 -378 5634 -372
rect 5694 -338 5752 -332
rect 5694 -372 5706 -338
rect 5740 -372 5752 -338
rect 5694 -378 5752 -372
rect 5812 -338 5870 -332
rect 5812 -372 5824 -338
rect 5858 -372 5870 -338
rect 5812 -378 5870 -372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 3 l 0.3 m 1 nf 100 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
