**.subckt tb_and
x1 vdd vin2 out vin1 vss and
V1 vss GND 0
V2 vdd vss 1.8
V3 vin1 vss PULSE(0 {vin1} 1ps 1ps 1ps 50ns 100ns) DC{vin1} 
V4 vin2 vss PULSE(0 {vin2} 1ps 1ps 1ps 25ns 50ns) DC{vin2} 
C1 out vss 1p m=1
**** begin user architecture code



*Circuits Params

.param vin1 = 1.8
.param vin2 = 1.8
.options TEMP = 27.0

*include

.lib /home/eamta/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT

*signals to SAVE

.save all  @M.x1.xm1.msky130_fd_pr__nfet_01v8[id]  @M.x1.xm1.msky130_fd_pr__nfet_01v8[gm]  @M.x1.xm2.msky130_fd_pr__nfet_01v8[id]  @M.x1.xm2.msky130_fd_pr__nfet_01v8[gm]  @M.x1.xm3.msky130_fd_pr__nfet_01v8[id]  @M.x1.xm3.msky130_fd_pr__nfet_01v8[gm]  @M.x1.xm4.msky130_fd_pr__pfet_01v8[id]  @M.x1.xm4.msky130_fd_pr__pfet_01v8[gm]  @M.x1.xm5.msky130_fd_pr__pfet_01v8[id]  @M.x1.xm5.msky130_fd_pr__pfet_01v8[gm]  @M.x1.xm6.msky130_fd_pr__pfet_01v8[id]  @M.x1.xm6.msky130_fd_pr__pfet_01v8[gm]


*simulation

.control
  tran 0.1n 0.5us
  setplot tran1
  plot v(out) v(vin1) v(vin2)
  write tb_and_tran.raw


  reset
  dc v3 0 1.8 0.01
  setplot dc1
  plot v(out) v(vin1) v(vin2)
  write tb_and_dc.raw

  reset
  op

  set filetype= ASCII

  write tb_and.raw
  print all


.endc






**** end user architecture code
**.ends

* expanding   symbol:  /home/eamta/eamta2021/sch/and/and.sym # of pins=5
* sym_path: /home/eamta/eamta2021/sch/and/and.sym
* sch_path: /home/eamta/eamta2021/sch/and/and.sch
.subckt and  vdd vb out va vss
*.opin out
*.ipin va
*.ipin vb
*.ipin vdd
*.ipin vss
XM1 net1 va vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net2 vb net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 out net2 vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net2 va vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net2 vb vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out net2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
