magic
tech sky130A
magscale 1 2
timestamp 1616037006
<< metal3 >>
rect -2550 2472 2549 2500
rect -2550 -2472 2465 2472
rect 2529 -2472 2549 2472
rect -2550 -2500 2549 -2472
<< via3 >>
rect 2465 -2472 2529 2472
<< mimcap >>
rect -2450 2360 2350 2400
rect -2450 -2360 -2410 2360
rect 2310 -2360 2350 2360
rect -2450 -2400 2350 -2360
<< mimcapcontact >>
rect -2410 -2360 2310 2360
<< metal4 >>
rect 2449 2472 2545 2488
rect -2411 2360 2311 2361
rect -2411 -2360 -2410 2360
rect 2310 -2360 2311 2360
rect -2411 -2361 2311 -2360
rect 2449 -2472 2465 2472
rect 2529 -2472 2545 2472
rect 2449 -2488 2545 -2472
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -2550 -2500 2450 2500
string parameters w 24 l 24 val 592.32 carea 1.00 cperi 0.17 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
