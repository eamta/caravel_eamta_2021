magic
tech sky130A
magscale 1 2
timestamp 1616092564
<< error_p >>
rect -6867 -411 -6795 -405
rect -6729 -411 -6657 -405
rect -6591 -411 -6519 -405
rect -6453 -411 -6381 -405
rect -6315 -411 -6243 -405
rect -6177 -411 -6105 -405
rect -6039 -411 -5967 -405
rect -5901 -411 -5829 -405
rect -5763 -411 -5691 -405
rect -5625 -411 -5553 -405
rect -5487 -411 -5415 -405
rect -5349 -411 -5277 -405
rect -5211 -411 -5139 -405
rect -5073 -411 -5001 -405
rect -4935 -411 -4863 -405
rect -4797 -411 -4725 -405
rect -4659 -411 -4587 -405
rect -4521 -411 -4449 -405
rect -4383 -411 -4311 -405
rect -4245 -411 -4173 -405
rect -4107 -411 -4035 -405
rect -3969 -411 -3897 -405
rect -3831 -411 -3759 -405
rect -3693 -411 -3621 -405
rect -3555 -411 -3483 -405
rect -3417 -411 -3345 -405
rect -3279 -411 -3207 -405
rect -3141 -411 -3069 -405
rect -3003 -411 -2931 -405
rect -2865 -411 -2793 -405
rect -2727 -411 -2655 -405
rect -2589 -411 -2517 -405
rect -2451 -411 -2379 -405
rect -2313 -411 -2241 -405
rect -2175 -411 -2103 -405
rect -2037 -411 -1965 -405
rect -1899 -411 -1827 -405
rect -1761 -411 -1689 -405
rect -1623 -411 -1551 -405
rect -1485 -411 -1413 -405
rect -1347 -411 -1275 -405
rect -1209 -411 -1137 -405
rect -1071 -411 -999 -405
rect -933 -411 -861 -405
rect -795 -411 -723 -405
rect -657 -411 -585 -405
rect -519 -411 -447 -405
rect -381 -411 -309 -405
rect -243 -411 -171 -405
rect -105 -411 -33 -405
rect 33 -411 105 -405
rect 171 -411 243 -405
rect 309 -411 381 -405
rect 447 -411 519 -405
rect 585 -411 657 -405
rect 723 -411 795 -405
rect 861 -411 933 -405
rect 999 -411 1071 -405
rect 1137 -411 1209 -405
rect 1275 -411 1347 -405
rect 1413 -411 1485 -405
rect 1551 -411 1623 -405
rect 1689 -411 1761 -405
rect 1827 -411 1899 -405
rect 1965 -411 2037 -405
rect 2103 -411 2175 -405
rect 2241 -411 2313 -405
rect 2379 -411 2451 -405
rect 2517 -411 2589 -405
rect 2655 -411 2727 -405
rect 2793 -411 2865 -405
rect 2931 -411 3003 -405
rect 3069 -411 3141 -405
rect 3207 -411 3279 -405
rect 3345 -411 3417 -405
rect 3483 -411 3555 -405
rect 3621 -411 3693 -405
rect 3759 -411 3831 -405
rect 3897 -411 3969 -405
rect 4035 -411 4107 -405
rect 4173 -411 4245 -405
rect 4311 -411 4383 -405
rect 4449 -411 4521 -405
rect 4587 -411 4659 -405
rect 4725 -411 4797 -405
rect 4863 -411 4935 -405
rect 5001 -411 5073 -405
rect 5139 -411 5211 -405
rect 5277 -411 5349 -405
rect 5415 -411 5487 -405
rect 5553 -411 5625 -405
rect 5691 -411 5763 -405
rect 5829 -411 5901 -405
rect 5967 -411 6039 -405
rect 6105 -411 6177 -405
rect 6243 -411 6315 -405
rect 6381 -411 6453 -405
rect 6519 -411 6591 -405
rect 6657 -411 6729 -405
rect 6795 -411 6867 -405
rect -6867 -445 -6855 -411
rect -6729 -445 -6717 -411
rect -6591 -445 -6579 -411
rect -6453 -445 -6441 -411
rect -6315 -445 -6303 -411
rect -6177 -445 -6165 -411
rect -6039 -445 -6027 -411
rect -5901 -445 -5889 -411
rect -5763 -445 -5751 -411
rect -5625 -445 -5613 -411
rect -5487 -445 -5475 -411
rect -5349 -445 -5337 -411
rect -5211 -445 -5199 -411
rect -5073 -445 -5061 -411
rect -4935 -445 -4923 -411
rect -4797 -445 -4785 -411
rect -4659 -445 -4647 -411
rect -4521 -445 -4509 -411
rect -4383 -445 -4371 -411
rect -4245 -445 -4233 -411
rect -4107 -445 -4095 -411
rect -3969 -445 -3957 -411
rect -3831 -445 -3819 -411
rect -3693 -445 -3681 -411
rect -3555 -445 -3543 -411
rect -3417 -445 -3405 -411
rect -3279 -445 -3267 -411
rect -3141 -445 -3129 -411
rect -3003 -445 -2991 -411
rect -2865 -445 -2853 -411
rect -2727 -445 -2715 -411
rect -2589 -445 -2577 -411
rect -2451 -445 -2439 -411
rect -2313 -445 -2301 -411
rect -2175 -445 -2163 -411
rect -2037 -445 -2025 -411
rect -1899 -445 -1887 -411
rect -1761 -445 -1749 -411
rect -1623 -445 -1611 -411
rect -1485 -445 -1473 -411
rect -1347 -445 -1335 -411
rect -1209 -445 -1197 -411
rect -1071 -445 -1059 -411
rect -933 -445 -921 -411
rect -795 -445 -783 -411
rect -657 -445 -645 -411
rect -519 -445 -507 -411
rect -381 -445 -369 -411
rect -243 -445 -231 -411
rect -105 -445 -93 -411
rect 33 -445 45 -411
rect 171 -445 183 -411
rect 309 -445 321 -411
rect 447 -445 459 -411
rect 585 -445 597 -411
rect 723 -445 735 -411
rect 861 -445 873 -411
rect 999 -445 1011 -411
rect 1137 -445 1149 -411
rect 1275 -445 1287 -411
rect 1413 -445 1425 -411
rect 1551 -445 1563 -411
rect 1689 -445 1701 -411
rect 1827 -445 1839 -411
rect 1965 -445 1977 -411
rect 2103 -445 2115 -411
rect 2241 -445 2253 -411
rect 2379 -445 2391 -411
rect 2517 -445 2529 -411
rect 2655 -445 2667 -411
rect 2793 -445 2805 -411
rect 2931 -445 2943 -411
rect 3069 -445 3081 -411
rect 3207 -445 3219 -411
rect 3345 -445 3357 -411
rect 3483 -445 3495 -411
rect 3621 -445 3633 -411
rect 3759 -445 3771 -411
rect 3897 -445 3909 -411
rect 4035 -445 4047 -411
rect 4173 -445 4185 -411
rect 4311 -445 4323 -411
rect 4449 -445 4461 -411
rect 4587 -445 4599 -411
rect 4725 -445 4737 -411
rect 4863 -445 4875 -411
rect 5001 -445 5013 -411
rect 5139 -445 5151 -411
rect 5277 -445 5289 -411
rect 5415 -445 5427 -411
rect 5553 -445 5565 -411
rect 5691 -445 5703 -411
rect 5829 -445 5841 -411
rect 5967 -445 5979 -411
rect 6105 -445 6117 -411
rect 6243 -445 6255 -411
rect 6381 -445 6393 -411
rect 6519 -445 6531 -411
rect 6657 -445 6669 -411
rect 6795 -445 6807 -411
rect -6867 -451 -6795 -445
rect -6729 -451 -6657 -445
rect -6591 -451 -6519 -445
rect -6453 -451 -6381 -445
rect -6315 -451 -6243 -445
rect -6177 -451 -6105 -445
rect -6039 -451 -5967 -445
rect -5901 -451 -5829 -445
rect -5763 -451 -5691 -445
rect -5625 -451 -5553 -445
rect -5487 -451 -5415 -445
rect -5349 -451 -5277 -445
rect -5211 -451 -5139 -445
rect -5073 -451 -5001 -445
rect -4935 -451 -4863 -445
rect -4797 -451 -4725 -445
rect -4659 -451 -4587 -445
rect -4521 -451 -4449 -445
rect -4383 -451 -4311 -445
rect -4245 -451 -4173 -445
rect -4107 -451 -4035 -445
rect -3969 -451 -3897 -445
rect -3831 -451 -3759 -445
rect -3693 -451 -3621 -445
rect -3555 -451 -3483 -445
rect -3417 -451 -3345 -445
rect -3279 -451 -3207 -445
rect -3141 -451 -3069 -445
rect -3003 -451 -2931 -445
rect -2865 -451 -2793 -445
rect -2727 -451 -2655 -445
rect -2589 -451 -2517 -445
rect -2451 -451 -2379 -445
rect -2313 -451 -2241 -445
rect -2175 -451 -2103 -445
rect -2037 -451 -1965 -445
rect -1899 -451 -1827 -445
rect -1761 -451 -1689 -445
rect -1623 -451 -1551 -445
rect -1485 -451 -1413 -445
rect -1347 -451 -1275 -445
rect -1209 -451 -1137 -445
rect -1071 -451 -999 -445
rect -933 -451 -861 -445
rect -795 -451 -723 -445
rect -657 -451 -585 -445
rect -519 -451 -447 -445
rect -381 -451 -309 -445
rect -243 -451 -171 -445
rect -105 -451 -33 -445
rect 33 -451 105 -445
rect 171 -451 243 -445
rect 309 -451 381 -445
rect 447 -451 519 -445
rect 585 -451 657 -445
rect 723 -451 795 -445
rect 861 -451 933 -445
rect 999 -451 1071 -445
rect 1137 -451 1209 -445
rect 1275 -451 1347 -445
rect 1413 -451 1485 -445
rect 1551 -451 1623 -445
rect 1689 -451 1761 -445
rect 1827 -451 1899 -445
rect 1965 -451 2037 -445
rect 2103 -451 2175 -445
rect 2241 -451 2313 -445
rect 2379 -451 2451 -445
rect 2517 -451 2589 -445
rect 2655 -451 2727 -445
rect 2793 -451 2865 -445
rect 2931 -451 3003 -445
rect 3069 -451 3141 -445
rect 3207 -451 3279 -445
rect 3345 -451 3417 -445
rect 3483 -451 3555 -445
rect 3621 -451 3693 -445
rect 3759 -451 3831 -445
rect 3897 -451 3969 -445
rect 4035 -451 4107 -445
rect 4173 -451 4245 -445
rect 4311 -451 4383 -445
rect 4449 -451 4521 -445
rect 4587 -451 4659 -445
rect 4725 -451 4797 -445
rect 4863 -451 4935 -445
rect 5001 -451 5073 -445
rect 5139 -451 5211 -445
rect 5277 -451 5349 -445
rect 5415 -451 5487 -445
rect 5553 -451 5625 -445
rect 5691 -451 5763 -445
rect 5829 -451 5901 -445
rect 5967 -451 6039 -445
rect 6105 -451 6177 -445
rect 6243 -451 6315 -445
rect 6381 -451 6453 -445
rect 6519 -451 6591 -445
rect 6657 -451 6729 -445
rect 6795 -451 6867 -445
<< nwell >>
rect -6965 -464 6965 498
<< pmoslvt >>
rect -6871 -364 -6791 436
rect -6733 -364 -6653 436
rect -6595 -364 -6515 436
rect -6457 -364 -6377 436
rect -6319 -364 -6239 436
rect -6181 -364 -6101 436
rect -6043 -364 -5963 436
rect -5905 -364 -5825 436
rect -5767 -364 -5687 436
rect -5629 -364 -5549 436
rect -5491 -364 -5411 436
rect -5353 -364 -5273 436
rect -5215 -364 -5135 436
rect -5077 -364 -4997 436
rect -4939 -364 -4859 436
rect -4801 -364 -4721 436
rect -4663 -364 -4583 436
rect -4525 -364 -4445 436
rect -4387 -364 -4307 436
rect -4249 -364 -4169 436
rect -4111 -364 -4031 436
rect -3973 -364 -3893 436
rect -3835 -364 -3755 436
rect -3697 -364 -3617 436
rect -3559 -364 -3479 436
rect -3421 -364 -3341 436
rect -3283 -364 -3203 436
rect -3145 -364 -3065 436
rect -3007 -364 -2927 436
rect -2869 -364 -2789 436
rect -2731 -364 -2651 436
rect -2593 -364 -2513 436
rect -2455 -364 -2375 436
rect -2317 -364 -2237 436
rect -2179 -364 -2099 436
rect -2041 -364 -1961 436
rect -1903 -364 -1823 436
rect -1765 -364 -1685 436
rect -1627 -364 -1547 436
rect -1489 -364 -1409 436
rect -1351 -364 -1271 436
rect -1213 -364 -1133 436
rect -1075 -364 -995 436
rect -937 -364 -857 436
rect -799 -364 -719 436
rect -661 -364 -581 436
rect -523 -364 -443 436
rect -385 -364 -305 436
rect -247 -364 -167 436
rect -109 -364 -29 436
rect 29 -364 109 436
rect 167 -364 247 436
rect 305 -364 385 436
rect 443 -364 523 436
rect 581 -364 661 436
rect 719 -364 799 436
rect 857 -364 937 436
rect 995 -364 1075 436
rect 1133 -364 1213 436
rect 1271 -364 1351 436
rect 1409 -364 1489 436
rect 1547 -364 1627 436
rect 1685 -364 1765 436
rect 1823 -364 1903 436
rect 1961 -364 2041 436
rect 2099 -364 2179 436
rect 2237 -364 2317 436
rect 2375 -364 2455 436
rect 2513 -364 2593 436
rect 2651 -364 2731 436
rect 2789 -364 2869 436
rect 2927 -364 3007 436
rect 3065 -364 3145 436
rect 3203 -364 3283 436
rect 3341 -364 3421 436
rect 3479 -364 3559 436
rect 3617 -364 3697 436
rect 3755 -364 3835 436
rect 3893 -364 3973 436
rect 4031 -364 4111 436
rect 4169 -364 4249 436
rect 4307 -364 4387 436
rect 4445 -364 4525 436
rect 4583 -364 4663 436
rect 4721 -364 4801 436
rect 4859 -364 4939 436
rect 4997 -364 5077 436
rect 5135 -364 5215 436
rect 5273 -364 5353 436
rect 5411 -364 5491 436
rect 5549 -364 5629 436
rect 5687 -364 5767 436
rect 5825 -364 5905 436
rect 5963 -364 6043 436
rect 6101 -364 6181 436
rect 6239 -364 6319 436
rect 6377 -364 6457 436
rect 6515 -364 6595 436
rect 6653 -364 6733 436
rect 6791 -364 6871 436
<< pdiff >>
rect -6929 424 -6871 436
rect -6929 -352 -6917 424
rect -6883 -352 -6871 424
rect -6929 -364 -6871 -352
rect -6791 424 -6733 436
rect -6791 -352 -6779 424
rect -6745 -352 -6733 424
rect -6791 -364 -6733 -352
rect -6653 424 -6595 436
rect -6653 -352 -6641 424
rect -6607 -352 -6595 424
rect -6653 -364 -6595 -352
rect -6515 424 -6457 436
rect -6515 -352 -6503 424
rect -6469 -352 -6457 424
rect -6515 -364 -6457 -352
rect -6377 424 -6319 436
rect -6377 -352 -6365 424
rect -6331 -352 -6319 424
rect -6377 -364 -6319 -352
rect -6239 424 -6181 436
rect -6239 -352 -6227 424
rect -6193 -352 -6181 424
rect -6239 -364 -6181 -352
rect -6101 424 -6043 436
rect -6101 -352 -6089 424
rect -6055 -352 -6043 424
rect -6101 -364 -6043 -352
rect -5963 424 -5905 436
rect -5963 -352 -5951 424
rect -5917 -352 -5905 424
rect -5963 -364 -5905 -352
rect -5825 424 -5767 436
rect -5825 -352 -5813 424
rect -5779 -352 -5767 424
rect -5825 -364 -5767 -352
rect -5687 424 -5629 436
rect -5687 -352 -5675 424
rect -5641 -352 -5629 424
rect -5687 -364 -5629 -352
rect -5549 424 -5491 436
rect -5549 -352 -5537 424
rect -5503 -352 -5491 424
rect -5549 -364 -5491 -352
rect -5411 424 -5353 436
rect -5411 -352 -5399 424
rect -5365 -352 -5353 424
rect -5411 -364 -5353 -352
rect -5273 424 -5215 436
rect -5273 -352 -5261 424
rect -5227 -352 -5215 424
rect -5273 -364 -5215 -352
rect -5135 424 -5077 436
rect -5135 -352 -5123 424
rect -5089 -352 -5077 424
rect -5135 -364 -5077 -352
rect -4997 424 -4939 436
rect -4997 -352 -4985 424
rect -4951 -352 -4939 424
rect -4997 -364 -4939 -352
rect -4859 424 -4801 436
rect -4859 -352 -4847 424
rect -4813 -352 -4801 424
rect -4859 -364 -4801 -352
rect -4721 424 -4663 436
rect -4721 -352 -4709 424
rect -4675 -352 -4663 424
rect -4721 -364 -4663 -352
rect -4583 424 -4525 436
rect -4583 -352 -4571 424
rect -4537 -352 -4525 424
rect -4583 -364 -4525 -352
rect -4445 424 -4387 436
rect -4445 -352 -4433 424
rect -4399 -352 -4387 424
rect -4445 -364 -4387 -352
rect -4307 424 -4249 436
rect -4307 -352 -4295 424
rect -4261 -352 -4249 424
rect -4307 -364 -4249 -352
rect -4169 424 -4111 436
rect -4169 -352 -4157 424
rect -4123 -352 -4111 424
rect -4169 -364 -4111 -352
rect -4031 424 -3973 436
rect -4031 -352 -4019 424
rect -3985 -352 -3973 424
rect -4031 -364 -3973 -352
rect -3893 424 -3835 436
rect -3893 -352 -3881 424
rect -3847 -352 -3835 424
rect -3893 -364 -3835 -352
rect -3755 424 -3697 436
rect -3755 -352 -3743 424
rect -3709 -352 -3697 424
rect -3755 -364 -3697 -352
rect -3617 424 -3559 436
rect -3617 -352 -3605 424
rect -3571 -352 -3559 424
rect -3617 -364 -3559 -352
rect -3479 424 -3421 436
rect -3479 -352 -3467 424
rect -3433 -352 -3421 424
rect -3479 -364 -3421 -352
rect -3341 424 -3283 436
rect -3341 -352 -3329 424
rect -3295 -352 -3283 424
rect -3341 -364 -3283 -352
rect -3203 424 -3145 436
rect -3203 -352 -3191 424
rect -3157 -352 -3145 424
rect -3203 -364 -3145 -352
rect -3065 424 -3007 436
rect -3065 -352 -3053 424
rect -3019 -352 -3007 424
rect -3065 -364 -3007 -352
rect -2927 424 -2869 436
rect -2927 -352 -2915 424
rect -2881 -352 -2869 424
rect -2927 -364 -2869 -352
rect -2789 424 -2731 436
rect -2789 -352 -2777 424
rect -2743 -352 -2731 424
rect -2789 -364 -2731 -352
rect -2651 424 -2593 436
rect -2651 -352 -2639 424
rect -2605 -352 -2593 424
rect -2651 -364 -2593 -352
rect -2513 424 -2455 436
rect -2513 -352 -2501 424
rect -2467 -352 -2455 424
rect -2513 -364 -2455 -352
rect -2375 424 -2317 436
rect -2375 -352 -2363 424
rect -2329 -352 -2317 424
rect -2375 -364 -2317 -352
rect -2237 424 -2179 436
rect -2237 -352 -2225 424
rect -2191 -352 -2179 424
rect -2237 -364 -2179 -352
rect -2099 424 -2041 436
rect -2099 -352 -2087 424
rect -2053 -352 -2041 424
rect -2099 -364 -2041 -352
rect -1961 424 -1903 436
rect -1961 -352 -1949 424
rect -1915 -352 -1903 424
rect -1961 -364 -1903 -352
rect -1823 424 -1765 436
rect -1823 -352 -1811 424
rect -1777 -352 -1765 424
rect -1823 -364 -1765 -352
rect -1685 424 -1627 436
rect -1685 -352 -1673 424
rect -1639 -352 -1627 424
rect -1685 -364 -1627 -352
rect -1547 424 -1489 436
rect -1547 -352 -1535 424
rect -1501 -352 -1489 424
rect -1547 -364 -1489 -352
rect -1409 424 -1351 436
rect -1409 -352 -1397 424
rect -1363 -352 -1351 424
rect -1409 -364 -1351 -352
rect -1271 424 -1213 436
rect -1271 -352 -1259 424
rect -1225 -352 -1213 424
rect -1271 -364 -1213 -352
rect -1133 424 -1075 436
rect -1133 -352 -1121 424
rect -1087 -352 -1075 424
rect -1133 -364 -1075 -352
rect -995 424 -937 436
rect -995 -352 -983 424
rect -949 -352 -937 424
rect -995 -364 -937 -352
rect -857 424 -799 436
rect -857 -352 -845 424
rect -811 -352 -799 424
rect -857 -364 -799 -352
rect -719 424 -661 436
rect -719 -352 -707 424
rect -673 -352 -661 424
rect -719 -364 -661 -352
rect -581 424 -523 436
rect -581 -352 -569 424
rect -535 -352 -523 424
rect -581 -364 -523 -352
rect -443 424 -385 436
rect -443 -352 -431 424
rect -397 -352 -385 424
rect -443 -364 -385 -352
rect -305 424 -247 436
rect -305 -352 -293 424
rect -259 -352 -247 424
rect -305 -364 -247 -352
rect -167 424 -109 436
rect -167 -352 -155 424
rect -121 -352 -109 424
rect -167 -364 -109 -352
rect -29 424 29 436
rect -29 -352 -17 424
rect 17 -352 29 424
rect -29 -364 29 -352
rect 109 424 167 436
rect 109 -352 121 424
rect 155 -352 167 424
rect 109 -364 167 -352
rect 247 424 305 436
rect 247 -352 259 424
rect 293 -352 305 424
rect 247 -364 305 -352
rect 385 424 443 436
rect 385 -352 397 424
rect 431 -352 443 424
rect 385 -364 443 -352
rect 523 424 581 436
rect 523 -352 535 424
rect 569 -352 581 424
rect 523 -364 581 -352
rect 661 424 719 436
rect 661 -352 673 424
rect 707 -352 719 424
rect 661 -364 719 -352
rect 799 424 857 436
rect 799 -352 811 424
rect 845 -352 857 424
rect 799 -364 857 -352
rect 937 424 995 436
rect 937 -352 949 424
rect 983 -352 995 424
rect 937 -364 995 -352
rect 1075 424 1133 436
rect 1075 -352 1087 424
rect 1121 -352 1133 424
rect 1075 -364 1133 -352
rect 1213 424 1271 436
rect 1213 -352 1225 424
rect 1259 -352 1271 424
rect 1213 -364 1271 -352
rect 1351 424 1409 436
rect 1351 -352 1363 424
rect 1397 -352 1409 424
rect 1351 -364 1409 -352
rect 1489 424 1547 436
rect 1489 -352 1501 424
rect 1535 -352 1547 424
rect 1489 -364 1547 -352
rect 1627 424 1685 436
rect 1627 -352 1639 424
rect 1673 -352 1685 424
rect 1627 -364 1685 -352
rect 1765 424 1823 436
rect 1765 -352 1777 424
rect 1811 -352 1823 424
rect 1765 -364 1823 -352
rect 1903 424 1961 436
rect 1903 -352 1915 424
rect 1949 -352 1961 424
rect 1903 -364 1961 -352
rect 2041 424 2099 436
rect 2041 -352 2053 424
rect 2087 -352 2099 424
rect 2041 -364 2099 -352
rect 2179 424 2237 436
rect 2179 -352 2191 424
rect 2225 -352 2237 424
rect 2179 -364 2237 -352
rect 2317 424 2375 436
rect 2317 -352 2329 424
rect 2363 -352 2375 424
rect 2317 -364 2375 -352
rect 2455 424 2513 436
rect 2455 -352 2467 424
rect 2501 -352 2513 424
rect 2455 -364 2513 -352
rect 2593 424 2651 436
rect 2593 -352 2605 424
rect 2639 -352 2651 424
rect 2593 -364 2651 -352
rect 2731 424 2789 436
rect 2731 -352 2743 424
rect 2777 -352 2789 424
rect 2731 -364 2789 -352
rect 2869 424 2927 436
rect 2869 -352 2881 424
rect 2915 -352 2927 424
rect 2869 -364 2927 -352
rect 3007 424 3065 436
rect 3007 -352 3019 424
rect 3053 -352 3065 424
rect 3007 -364 3065 -352
rect 3145 424 3203 436
rect 3145 -352 3157 424
rect 3191 -352 3203 424
rect 3145 -364 3203 -352
rect 3283 424 3341 436
rect 3283 -352 3295 424
rect 3329 -352 3341 424
rect 3283 -364 3341 -352
rect 3421 424 3479 436
rect 3421 -352 3433 424
rect 3467 -352 3479 424
rect 3421 -364 3479 -352
rect 3559 424 3617 436
rect 3559 -352 3571 424
rect 3605 -352 3617 424
rect 3559 -364 3617 -352
rect 3697 424 3755 436
rect 3697 -352 3709 424
rect 3743 -352 3755 424
rect 3697 -364 3755 -352
rect 3835 424 3893 436
rect 3835 -352 3847 424
rect 3881 -352 3893 424
rect 3835 -364 3893 -352
rect 3973 424 4031 436
rect 3973 -352 3985 424
rect 4019 -352 4031 424
rect 3973 -364 4031 -352
rect 4111 424 4169 436
rect 4111 -352 4123 424
rect 4157 -352 4169 424
rect 4111 -364 4169 -352
rect 4249 424 4307 436
rect 4249 -352 4261 424
rect 4295 -352 4307 424
rect 4249 -364 4307 -352
rect 4387 424 4445 436
rect 4387 -352 4399 424
rect 4433 -352 4445 424
rect 4387 -364 4445 -352
rect 4525 424 4583 436
rect 4525 -352 4537 424
rect 4571 -352 4583 424
rect 4525 -364 4583 -352
rect 4663 424 4721 436
rect 4663 -352 4675 424
rect 4709 -352 4721 424
rect 4663 -364 4721 -352
rect 4801 424 4859 436
rect 4801 -352 4813 424
rect 4847 -352 4859 424
rect 4801 -364 4859 -352
rect 4939 424 4997 436
rect 4939 -352 4951 424
rect 4985 -352 4997 424
rect 4939 -364 4997 -352
rect 5077 424 5135 436
rect 5077 -352 5089 424
rect 5123 -352 5135 424
rect 5077 -364 5135 -352
rect 5215 424 5273 436
rect 5215 -352 5227 424
rect 5261 -352 5273 424
rect 5215 -364 5273 -352
rect 5353 424 5411 436
rect 5353 -352 5365 424
rect 5399 -352 5411 424
rect 5353 -364 5411 -352
rect 5491 424 5549 436
rect 5491 -352 5503 424
rect 5537 -352 5549 424
rect 5491 -364 5549 -352
rect 5629 424 5687 436
rect 5629 -352 5641 424
rect 5675 -352 5687 424
rect 5629 -364 5687 -352
rect 5767 424 5825 436
rect 5767 -352 5779 424
rect 5813 -352 5825 424
rect 5767 -364 5825 -352
rect 5905 424 5963 436
rect 5905 -352 5917 424
rect 5951 -352 5963 424
rect 5905 -364 5963 -352
rect 6043 424 6101 436
rect 6043 -352 6055 424
rect 6089 -352 6101 424
rect 6043 -364 6101 -352
rect 6181 424 6239 436
rect 6181 -352 6193 424
rect 6227 -352 6239 424
rect 6181 -364 6239 -352
rect 6319 424 6377 436
rect 6319 -352 6331 424
rect 6365 -352 6377 424
rect 6319 -364 6377 -352
rect 6457 424 6515 436
rect 6457 -352 6469 424
rect 6503 -352 6515 424
rect 6457 -364 6515 -352
rect 6595 424 6653 436
rect 6595 -352 6607 424
rect 6641 -352 6653 424
rect 6595 -364 6653 -352
rect 6733 424 6791 436
rect 6733 -352 6745 424
rect 6779 -352 6791 424
rect 6733 -364 6791 -352
rect 6871 424 6929 436
rect 6871 -352 6883 424
rect 6917 -352 6929 424
rect 6871 -364 6929 -352
<< pdiffc >>
rect -6917 -352 -6883 424
rect -6779 -352 -6745 424
rect -6641 -352 -6607 424
rect -6503 -352 -6469 424
rect -6365 -352 -6331 424
rect -6227 -352 -6193 424
rect -6089 -352 -6055 424
rect -5951 -352 -5917 424
rect -5813 -352 -5779 424
rect -5675 -352 -5641 424
rect -5537 -352 -5503 424
rect -5399 -352 -5365 424
rect -5261 -352 -5227 424
rect -5123 -352 -5089 424
rect -4985 -352 -4951 424
rect -4847 -352 -4813 424
rect -4709 -352 -4675 424
rect -4571 -352 -4537 424
rect -4433 -352 -4399 424
rect -4295 -352 -4261 424
rect -4157 -352 -4123 424
rect -4019 -352 -3985 424
rect -3881 -352 -3847 424
rect -3743 -352 -3709 424
rect -3605 -352 -3571 424
rect -3467 -352 -3433 424
rect -3329 -352 -3295 424
rect -3191 -352 -3157 424
rect -3053 -352 -3019 424
rect -2915 -352 -2881 424
rect -2777 -352 -2743 424
rect -2639 -352 -2605 424
rect -2501 -352 -2467 424
rect -2363 -352 -2329 424
rect -2225 -352 -2191 424
rect -2087 -352 -2053 424
rect -1949 -352 -1915 424
rect -1811 -352 -1777 424
rect -1673 -352 -1639 424
rect -1535 -352 -1501 424
rect -1397 -352 -1363 424
rect -1259 -352 -1225 424
rect -1121 -352 -1087 424
rect -983 -352 -949 424
rect -845 -352 -811 424
rect -707 -352 -673 424
rect -569 -352 -535 424
rect -431 -352 -397 424
rect -293 -352 -259 424
rect -155 -352 -121 424
rect -17 -352 17 424
rect 121 -352 155 424
rect 259 -352 293 424
rect 397 -352 431 424
rect 535 -352 569 424
rect 673 -352 707 424
rect 811 -352 845 424
rect 949 -352 983 424
rect 1087 -352 1121 424
rect 1225 -352 1259 424
rect 1363 -352 1397 424
rect 1501 -352 1535 424
rect 1639 -352 1673 424
rect 1777 -352 1811 424
rect 1915 -352 1949 424
rect 2053 -352 2087 424
rect 2191 -352 2225 424
rect 2329 -352 2363 424
rect 2467 -352 2501 424
rect 2605 -352 2639 424
rect 2743 -352 2777 424
rect 2881 -352 2915 424
rect 3019 -352 3053 424
rect 3157 -352 3191 424
rect 3295 -352 3329 424
rect 3433 -352 3467 424
rect 3571 -352 3605 424
rect 3709 -352 3743 424
rect 3847 -352 3881 424
rect 3985 -352 4019 424
rect 4123 -352 4157 424
rect 4261 -352 4295 424
rect 4399 -352 4433 424
rect 4537 -352 4571 424
rect 4675 -352 4709 424
rect 4813 -352 4847 424
rect 4951 -352 4985 424
rect 5089 -352 5123 424
rect 5227 -352 5261 424
rect 5365 -352 5399 424
rect 5503 -352 5537 424
rect 5641 -352 5675 424
rect 5779 -352 5813 424
rect 5917 -352 5951 424
rect 6055 -352 6089 424
rect 6193 -352 6227 424
rect 6331 -352 6365 424
rect 6469 -352 6503 424
rect 6607 -352 6641 424
rect 6745 -352 6779 424
rect 6883 -352 6917 424
<< poly >>
rect -6871 436 -6791 462
rect -6733 436 -6653 462
rect -6595 436 -6515 462
rect -6457 436 -6377 462
rect -6319 436 -6239 462
rect -6181 436 -6101 462
rect -6043 436 -5963 462
rect -5905 436 -5825 462
rect -5767 436 -5687 462
rect -5629 436 -5549 462
rect -5491 436 -5411 462
rect -5353 436 -5273 462
rect -5215 436 -5135 462
rect -5077 436 -4997 462
rect -4939 436 -4859 462
rect -4801 436 -4721 462
rect -4663 436 -4583 462
rect -4525 436 -4445 462
rect -4387 436 -4307 462
rect -4249 436 -4169 462
rect -4111 436 -4031 462
rect -3973 436 -3893 462
rect -3835 436 -3755 462
rect -3697 436 -3617 462
rect -3559 436 -3479 462
rect -3421 436 -3341 462
rect -3283 436 -3203 462
rect -3145 436 -3065 462
rect -3007 436 -2927 462
rect -2869 436 -2789 462
rect -2731 436 -2651 462
rect -2593 436 -2513 462
rect -2455 436 -2375 462
rect -2317 436 -2237 462
rect -2179 436 -2099 462
rect -2041 436 -1961 462
rect -1903 436 -1823 462
rect -1765 436 -1685 462
rect -1627 436 -1547 462
rect -1489 436 -1409 462
rect -1351 436 -1271 462
rect -1213 436 -1133 462
rect -1075 436 -995 462
rect -937 436 -857 462
rect -799 436 -719 462
rect -661 436 -581 462
rect -523 436 -443 462
rect -385 436 -305 462
rect -247 436 -167 462
rect -109 436 -29 462
rect 29 436 109 462
rect 167 436 247 462
rect 305 436 385 462
rect 443 436 523 462
rect 581 436 661 462
rect 719 436 799 462
rect 857 436 937 462
rect 995 436 1075 462
rect 1133 436 1213 462
rect 1271 436 1351 462
rect 1409 436 1489 462
rect 1547 436 1627 462
rect 1685 436 1765 462
rect 1823 436 1903 462
rect 1961 436 2041 462
rect 2099 436 2179 462
rect 2237 436 2317 462
rect 2375 436 2455 462
rect 2513 436 2593 462
rect 2651 436 2731 462
rect 2789 436 2869 462
rect 2927 436 3007 462
rect 3065 436 3145 462
rect 3203 436 3283 462
rect 3341 436 3421 462
rect 3479 436 3559 462
rect 3617 436 3697 462
rect 3755 436 3835 462
rect 3893 436 3973 462
rect 4031 436 4111 462
rect 4169 436 4249 462
rect 4307 436 4387 462
rect 4445 436 4525 462
rect 4583 436 4663 462
rect 4721 436 4801 462
rect 4859 436 4939 462
rect 4997 436 5077 462
rect 5135 436 5215 462
rect 5273 436 5353 462
rect 5411 436 5491 462
rect 5549 436 5629 462
rect 5687 436 5767 462
rect 5825 436 5905 462
rect 5963 436 6043 462
rect 6101 436 6181 462
rect 6239 436 6319 462
rect 6377 436 6457 462
rect 6515 436 6595 462
rect 6653 436 6733 462
rect 6791 436 6871 462
rect -6871 -411 -6791 -364
rect -6871 -445 -6855 -411
rect -6807 -445 -6791 -411
rect -6871 -461 -6791 -445
rect -6733 -411 -6653 -364
rect -6733 -445 -6717 -411
rect -6669 -445 -6653 -411
rect -6733 -461 -6653 -445
rect -6595 -411 -6515 -364
rect -6595 -445 -6579 -411
rect -6531 -445 -6515 -411
rect -6595 -461 -6515 -445
rect -6457 -411 -6377 -364
rect -6457 -445 -6441 -411
rect -6393 -445 -6377 -411
rect -6457 -461 -6377 -445
rect -6319 -411 -6239 -364
rect -6319 -445 -6303 -411
rect -6255 -445 -6239 -411
rect -6319 -461 -6239 -445
rect -6181 -411 -6101 -364
rect -6181 -445 -6165 -411
rect -6117 -445 -6101 -411
rect -6181 -461 -6101 -445
rect -6043 -411 -5963 -364
rect -6043 -445 -6027 -411
rect -5979 -445 -5963 -411
rect -6043 -461 -5963 -445
rect -5905 -411 -5825 -364
rect -5905 -445 -5889 -411
rect -5841 -445 -5825 -411
rect -5905 -461 -5825 -445
rect -5767 -411 -5687 -364
rect -5767 -445 -5751 -411
rect -5703 -445 -5687 -411
rect -5767 -461 -5687 -445
rect -5629 -411 -5549 -364
rect -5629 -445 -5613 -411
rect -5565 -445 -5549 -411
rect -5629 -461 -5549 -445
rect -5491 -411 -5411 -364
rect -5491 -445 -5475 -411
rect -5427 -445 -5411 -411
rect -5491 -461 -5411 -445
rect -5353 -411 -5273 -364
rect -5353 -445 -5337 -411
rect -5289 -445 -5273 -411
rect -5353 -461 -5273 -445
rect -5215 -411 -5135 -364
rect -5215 -445 -5199 -411
rect -5151 -445 -5135 -411
rect -5215 -461 -5135 -445
rect -5077 -411 -4997 -364
rect -5077 -445 -5061 -411
rect -5013 -445 -4997 -411
rect -5077 -461 -4997 -445
rect -4939 -411 -4859 -364
rect -4939 -445 -4923 -411
rect -4875 -445 -4859 -411
rect -4939 -461 -4859 -445
rect -4801 -411 -4721 -364
rect -4801 -445 -4785 -411
rect -4737 -445 -4721 -411
rect -4801 -461 -4721 -445
rect -4663 -411 -4583 -364
rect -4663 -445 -4647 -411
rect -4599 -445 -4583 -411
rect -4663 -461 -4583 -445
rect -4525 -411 -4445 -364
rect -4525 -445 -4509 -411
rect -4461 -445 -4445 -411
rect -4525 -461 -4445 -445
rect -4387 -411 -4307 -364
rect -4387 -445 -4371 -411
rect -4323 -445 -4307 -411
rect -4387 -461 -4307 -445
rect -4249 -411 -4169 -364
rect -4249 -445 -4233 -411
rect -4185 -445 -4169 -411
rect -4249 -461 -4169 -445
rect -4111 -411 -4031 -364
rect -4111 -445 -4095 -411
rect -4047 -445 -4031 -411
rect -4111 -461 -4031 -445
rect -3973 -411 -3893 -364
rect -3973 -445 -3957 -411
rect -3909 -445 -3893 -411
rect -3973 -461 -3893 -445
rect -3835 -411 -3755 -364
rect -3835 -445 -3819 -411
rect -3771 -445 -3755 -411
rect -3835 -461 -3755 -445
rect -3697 -411 -3617 -364
rect -3697 -445 -3681 -411
rect -3633 -445 -3617 -411
rect -3697 -461 -3617 -445
rect -3559 -411 -3479 -364
rect -3559 -445 -3543 -411
rect -3495 -445 -3479 -411
rect -3559 -461 -3479 -445
rect -3421 -411 -3341 -364
rect -3421 -445 -3405 -411
rect -3357 -445 -3341 -411
rect -3421 -461 -3341 -445
rect -3283 -411 -3203 -364
rect -3283 -445 -3267 -411
rect -3219 -445 -3203 -411
rect -3283 -461 -3203 -445
rect -3145 -411 -3065 -364
rect -3145 -445 -3129 -411
rect -3081 -445 -3065 -411
rect -3145 -461 -3065 -445
rect -3007 -411 -2927 -364
rect -3007 -445 -2991 -411
rect -2943 -445 -2927 -411
rect -3007 -461 -2927 -445
rect -2869 -411 -2789 -364
rect -2869 -445 -2853 -411
rect -2805 -445 -2789 -411
rect -2869 -461 -2789 -445
rect -2731 -411 -2651 -364
rect -2731 -445 -2715 -411
rect -2667 -445 -2651 -411
rect -2731 -461 -2651 -445
rect -2593 -411 -2513 -364
rect -2593 -445 -2577 -411
rect -2529 -445 -2513 -411
rect -2593 -461 -2513 -445
rect -2455 -411 -2375 -364
rect -2455 -445 -2439 -411
rect -2391 -445 -2375 -411
rect -2455 -461 -2375 -445
rect -2317 -411 -2237 -364
rect -2317 -445 -2301 -411
rect -2253 -445 -2237 -411
rect -2317 -461 -2237 -445
rect -2179 -411 -2099 -364
rect -2179 -445 -2163 -411
rect -2115 -445 -2099 -411
rect -2179 -461 -2099 -445
rect -2041 -411 -1961 -364
rect -2041 -445 -2025 -411
rect -1977 -445 -1961 -411
rect -2041 -461 -1961 -445
rect -1903 -411 -1823 -364
rect -1903 -445 -1887 -411
rect -1839 -445 -1823 -411
rect -1903 -461 -1823 -445
rect -1765 -411 -1685 -364
rect -1765 -445 -1749 -411
rect -1701 -445 -1685 -411
rect -1765 -461 -1685 -445
rect -1627 -411 -1547 -364
rect -1627 -445 -1611 -411
rect -1563 -445 -1547 -411
rect -1627 -461 -1547 -445
rect -1489 -411 -1409 -364
rect -1489 -445 -1473 -411
rect -1425 -445 -1409 -411
rect -1489 -461 -1409 -445
rect -1351 -411 -1271 -364
rect -1351 -445 -1335 -411
rect -1287 -445 -1271 -411
rect -1351 -461 -1271 -445
rect -1213 -411 -1133 -364
rect -1213 -445 -1197 -411
rect -1149 -445 -1133 -411
rect -1213 -461 -1133 -445
rect -1075 -411 -995 -364
rect -1075 -445 -1059 -411
rect -1011 -445 -995 -411
rect -1075 -461 -995 -445
rect -937 -411 -857 -364
rect -937 -445 -921 -411
rect -873 -445 -857 -411
rect -937 -461 -857 -445
rect -799 -411 -719 -364
rect -799 -445 -783 -411
rect -735 -445 -719 -411
rect -799 -461 -719 -445
rect -661 -411 -581 -364
rect -661 -445 -645 -411
rect -597 -445 -581 -411
rect -661 -461 -581 -445
rect -523 -411 -443 -364
rect -523 -445 -507 -411
rect -459 -445 -443 -411
rect -523 -461 -443 -445
rect -385 -411 -305 -364
rect -385 -445 -369 -411
rect -321 -445 -305 -411
rect -385 -461 -305 -445
rect -247 -411 -167 -364
rect -247 -445 -231 -411
rect -183 -445 -167 -411
rect -247 -461 -167 -445
rect -109 -411 -29 -364
rect -109 -445 -93 -411
rect -45 -445 -29 -411
rect -109 -461 -29 -445
rect 29 -411 109 -364
rect 29 -445 45 -411
rect 93 -445 109 -411
rect 29 -461 109 -445
rect 167 -411 247 -364
rect 167 -445 183 -411
rect 231 -445 247 -411
rect 167 -461 247 -445
rect 305 -411 385 -364
rect 305 -445 321 -411
rect 369 -445 385 -411
rect 305 -461 385 -445
rect 443 -411 523 -364
rect 443 -445 459 -411
rect 507 -445 523 -411
rect 443 -461 523 -445
rect 581 -411 661 -364
rect 581 -445 597 -411
rect 645 -445 661 -411
rect 581 -461 661 -445
rect 719 -411 799 -364
rect 719 -445 735 -411
rect 783 -445 799 -411
rect 719 -461 799 -445
rect 857 -411 937 -364
rect 857 -445 873 -411
rect 921 -445 937 -411
rect 857 -461 937 -445
rect 995 -411 1075 -364
rect 995 -445 1011 -411
rect 1059 -445 1075 -411
rect 995 -461 1075 -445
rect 1133 -411 1213 -364
rect 1133 -445 1149 -411
rect 1197 -445 1213 -411
rect 1133 -461 1213 -445
rect 1271 -411 1351 -364
rect 1271 -445 1287 -411
rect 1335 -445 1351 -411
rect 1271 -461 1351 -445
rect 1409 -411 1489 -364
rect 1409 -445 1425 -411
rect 1473 -445 1489 -411
rect 1409 -461 1489 -445
rect 1547 -411 1627 -364
rect 1547 -445 1563 -411
rect 1611 -445 1627 -411
rect 1547 -461 1627 -445
rect 1685 -411 1765 -364
rect 1685 -445 1701 -411
rect 1749 -445 1765 -411
rect 1685 -461 1765 -445
rect 1823 -411 1903 -364
rect 1823 -445 1839 -411
rect 1887 -445 1903 -411
rect 1823 -461 1903 -445
rect 1961 -411 2041 -364
rect 1961 -445 1977 -411
rect 2025 -445 2041 -411
rect 1961 -461 2041 -445
rect 2099 -411 2179 -364
rect 2099 -445 2115 -411
rect 2163 -445 2179 -411
rect 2099 -461 2179 -445
rect 2237 -411 2317 -364
rect 2237 -445 2253 -411
rect 2301 -445 2317 -411
rect 2237 -461 2317 -445
rect 2375 -411 2455 -364
rect 2375 -445 2391 -411
rect 2439 -445 2455 -411
rect 2375 -461 2455 -445
rect 2513 -411 2593 -364
rect 2513 -445 2529 -411
rect 2577 -445 2593 -411
rect 2513 -461 2593 -445
rect 2651 -411 2731 -364
rect 2651 -445 2667 -411
rect 2715 -445 2731 -411
rect 2651 -461 2731 -445
rect 2789 -411 2869 -364
rect 2789 -445 2805 -411
rect 2853 -445 2869 -411
rect 2789 -461 2869 -445
rect 2927 -411 3007 -364
rect 2927 -445 2943 -411
rect 2991 -445 3007 -411
rect 2927 -461 3007 -445
rect 3065 -411 3145 -364
rect 3065 -445 3081 -411
rect 3129 -445 3145 -411
rect 3065 -461 3145 -445
rect 3203 -411 3283 -364
rect 3203 -445 3219 -411
rect 3267 -445 3283 -411
rect 3203 -461 3283 -445
rect 3341 -411 3421 -364
rect 3341 -445 3357 -411
rect 3405 -445 3421 -411
rect 3341 -461 3421 -445
rect 3479 -411 3559 -364
rect 3479 -445 3495 -411
rect 3543 -445 3559 -411
rect 3479 -461 3559 -445
rect 3617 -411 3697 -364
rect 3617 -445 3633 -411
rect 3681 -445 3697 -411
rect 3617 -461 3697 -445
rect 3755 -411 3835 -364
rect 3755 -445 3771 -411
rect 3819 -445 3835 -411
rect 3755 -461 3835 -445
rect 3893 -411 3973 -364
rect 3893 -445 3909 -411
rect 3957 -445 3973 -411
rect 3893 -461 3973 -445
rect 4031 -411 4111 -364
rect 4031 -445 4047 -411
rect 4095 -445 4111 -411
rect 4031 -461 4111 -445
rect 4169 -411 4249 -364
rect 4169 -445 4185 -411
rect 4233 -445 4249 -411
rect 4169 -461 4249 -445
rect 4307 -411 4387 -364
rect 4307 -445 4323 -411
rect 4371 -445 4387 -411
rect 4307 -461 4387 -445
rect 4445 -411 4525 -364
rect 4445 -445 4461 -411
rect 4509 -445 4525 -411
rect 4445 -461 4525 -445
rect 4583 -411 4663 -364
rect 4583 -445 4599 -411
rect 4647 -445 4663 -411
rect 4583 -461 4663 -445
rect 4721 -411 4801 -364
rect 4721 -445 4737 -411
rect 4785 -445 4801 -411
rect 4721 -461 4801 -445
rect 4859 -411 4939 -364
rect 4859 -445 4875 -411
rect 4923 -445 4939 -411
rect 4859 -461 4939 -445
rect 4997 -411 5077 -364
rect 4997 -445 5013 -411
rect 5061 -445 5077 -411
rect 4997 -461 5077 -445
rect 5135 -411 5215 -364
rect 5135 -445 5151 -411
rect 5199 -445 5215 -411
rect 5135 -461 5215 -445
rect 5273 -411 5353 -364
rect 5273 -445 5289 -411
rect 5337 -445 5353 -411
rect 5273 -461 5353 -445
rect 5411 -411 5491 -364
rect 5411 -445 5427 -411
rect 5475 -445 5491 -411
rect 5411 -461 5491 -445
rect 5549 -411 5629 -364
rect 5549 -445 5565 -411
rect 5613 -445 5629 -411
rect 5549 -461 5629 -445
rect 5687 -411 5767 -364
rect 5687 -445 5703 -411
rect 5751 -445 5767 -411
rect 5687 -461 5767 -445
rect 5825 -411 5905 -364
rect 5825 -445 5841 -411
rect 5889 -445 5905 -411
rect 5825 -461 5905 -445
rect 5963 -411 6043 -364
rect 5963 -445 5979 -411
rect 6027 -445 6043 -411
rect 5963 -461 6043 -445
rect 6101 -411 6181 -364
rect 6101 -445 6117 -411
rect 6165 -445 6181 -411
rect 6101 -461 6181 -445
rect 6239 -411 6319 -364
rect 6239 -445 6255 -411
rect 6303 -445 6319 -411
rect 6239 -461 6319 -445
rect 6377 -411 6457 -364
rect 6377 -445 6393 -411
rect 6441 -445 6457 -411
rect 6377 -461 6457 -445
rect 6515 -411 6595 -364
rect 6515 -445 6531 -411
rect 6579 -445 6595 -411
rect 6515 -461 6595 -445
rect 6653 -411 6733 -364
rect 6653 -445 6669 -411
rect 6717 -445 6733 -411
rect 6653 -461 6733 -445
rect 6791 -411 6871 -364
rect 6791 -445 6807 -411
rect 6855 -445 6871 -411
rect 6791 -461 6871 -445
<< polycont >>
rect -6855 -445 -6807 -411
rect -6717 -445 -6669 -411
rect -6579 -445 -6531 -411
rect -6441 -445 -6393 -411
rect -6303 -445 -6255 -411
rect -6165 -445 -6117 -411
rect -6027 -445 -5979 -411
rect -5889 -445 -5841 -411
rect -5751 -445 -5703 -411
rect -5613 -445 -5565 -411
rect -5475 -445 -5427 -411
rect -5337 -445 -5289 -411
rect -5199 -445 -5151 -411
rect -5061 -445 -5013 -411
rect -4923 -445 -4875 -411
rect -4785 -445 -4737 -411
rect -4647 -445 -4599 -411
rect -4509 -445 -4461 -411
rect -4371 -445 -4323 -411
rect -4233 -445 -4185 -411
rect -4095 -445 -4047 -411
rect -3957 -445 -3909 -411
rect -3819 -445 -3771 -411
rect -3681 -445 -3633 -411
rect -3543 -445 -3495 -411
rect -3405 -445 -3357 -411
rect -3267 -445 -3219 -411
rect -3129 -445 -3081 -411
rect -2991 -445 -2943 -411
rect -2853 -445 -2805 -411
rect -2715 -445 -2667 -411
rect -2577 -445 -2529 -411
rect -2439 -445 -2391 -411
rect -2301 -445 -2253 -411
rect -2163 -445 -2115 -411
rect -2025 -445 -1977 -411
rect -1887 -445 -1839 -411
rect -1749 -445 -1701 -411
rect -1611 -445 -1563 -411
rect -1473 -445 -1425 -411
rect -1335 -445 -1287 -411
rect -1197 -445 -1149 -411
rect -1059 -445 -1011 -411
rect -921 -445 -873 -411
rect -783 -445 -735 -411
rect -645 -445 -597 -411
rect -507 -445 -459 -411
rect -369 -445 -321 -411
rect -231 -445 -183 -411
rect -93 -445 -45 -411
rect 45 -445 93 -411
rect 183 -445 231 -411
rect 321 -445 369 -411
rect 459 -445 507 -411
rect 597 -445 645 -411
rect 735 -445 783 -411
rect 873 -445 921 -411
rect 1011 -445 1059 -411
rect 1149 -445 1197 -411
rect 1287 -445 1335 -411
rect 1425 -445 1473 -411
rect 1563 -445 1611 -411
rect 1701 -445 1749 -411
rect 1839 -445 1887 -411
rect 1977 -445 2025 -411
rect 2115 -445 2163 -411
rect 2253 -445 2301 -411
rect 2391 -445 2439 -411
rect 2529 -445 2577 -411
rect 2667 -445 2715 -411
rect 2805 -445 2853 -411
rect 2943 -445 2991 -411
rect 3081 -445 3129 -411
rect 3219 -445 3267 -411
rect 3357 -445 3405 -411
rect 3495 -445 3543 -411
rect 3633 -445 3681 -411
rect 3771 -445 3819 -411
rect 3909 -445 3957 -411
rect 4047 -445 4095 -411
rect 4185 -445 4233 -411
rect 4323 -445 4371 -411
rect 4461 -445 4509 -411
rect 4599 -445 4647 -411
rect 4737 -445 4785 -411
rect 4875 -445 4923 -411
rect 5013 -445 5061 -411
rect 5151 -445 5199 -411
rect 5289 -445 5337 -411
rect 5427 -445 5475 -411
rect 5565 -445 5613 -411
rect 5703 -445 5751 -411
rect 5841 -445 5889 -411
rect 5979 -445 6027 -411
rect 6117 -445 6165 -411
rect 6255 -445 6303 -411
rect 6393 -445 6441 -411
rect 6531 -445 6579 -411
rect 6669 -445 6717 -411
rect 6807 -445 6855 -411
<< locali >>
rect -6917 424 -6883 440
rect -6917 -368 -6883 -352
rect -6779 424 -6745 440
rect -6779 -368 -6745 -352
rect -6641 424 -6607 440
rect -6641 -368 -6607 -352
rect -6503 424 -6469 440
rect -6503 -368 -6469 -352
rect -6365 424 -6331 440
rect -6365 -368 -6331 -352
rect -6227 424 -6193 440
rect -6227 -368 -6193 -352
rect -6089 424 -6055 440
rect -6089 -368 -6055 -352
rect -5951 424 -5917 440
rect -5951 -368 -5917 -352
rect -5813 424 -5779 440
rect -5813 -368 -5779 -352
rect -5675 424 -5641 440
rect -5675 -368 -5641 -352
rect -5537 424 -5503 440
rect -5537 -368 -5503 -352
rect -5399 424 -5365 440
rect -5399 -368 -5365 -352
rect -5261 424 -5227 440
rect -5261 -368 -5227 -352
rect -5123 424 -5089 440
rect -5123 -368 -5089 -352
rect -4985 424 -4951 440
rect -4985 -368 -4951 -352
rect -4847 424 -4813 440
rect -4847 -368 -4813 -352
rect -4709 424 -4675 440
rect -4709 -368 -4675 -352
rect -4571 424 -4537 440
rect -4571 -368 -4537 -352
rect -4433 424 -4399 440
rect -4433 -368 -4399 -352
rect -4295 424 -4261 440
rect -4295 -368 -4261 -352
rect -4157 424 -4123 440
rect -4157 -368 -4123 -352
rect -4019 424 -3985 440
rect -4019 -368 -3985 -352
rect -3881 424 -3847 440
rect -3881 -368 -3847 -352
rect -3743 424 -3709 440
rect -3743 -368 -3709 -352
rect -3605 424 -3571 440
rect -3605 -368 -3571 -352
rect -3467 424 -3433 440
rect -3467 -368 -3433 -352
rect -3329 424 -3295 440
rect -3329 -368 -3295 -352
rect -3191 424 -3157 440
rect -3191 -368 -3157 -352
rect -3053 424 -3019 440
rect -3053 -368 -3019 -352
rect -2915 424 -2881 440
rect -2915 -368 -2881 -352
rect -2777 424 -2743 440
rect -2777 -368 -2743 -352
rect -2639 424 -2605 440
rect -2639 -368 -2605 -352
rect -2501 424 -2467 440
rect -2501 -368 -2467 -352
rect -2363 424 -2329 440
rect -2363 -368 -2329 -352
rect -2225 424 -2191 440
rect -2225 -368 -2191 -352
rect -2087 424 -2053 440
rect -2087 -368 -2053 -352
rect -1949 424 -1915 440
rect -1949 -368 -1915 -352
rect -1811 424 -1777 440
rect -1811 -368 -1777 -352
rect -1673 424 -1639 440
rect -1673 -368 -1639 -352
rect -1535 424 -1501 440
rect -1535 -368 -1501 -352
rect -1397 424 -1363 440
rect -1397 -368 -1363 -352
rect -1259 424 -1225 440
rect -1259 -368 -1225 -352
rect -1121 424 -1087 440
rect -1121 -368 -1087 -352
rect -983 424 -949 440
rect -983 -368 -949 -352
rect -845 424 -811 440
rect -845 -368 -811 -352
rect -707 424 -673 440
rect -707 -368 -673 -352
rect -569 424 -535 440
rect -569 -368 -535 -352
rect -431 424 -397 440
rect -431 -368 -397 -352
rect -293 424 -259 440
rect -293 -368 -259 -352
rect -155 424 -121 440
rect -155 -368 -121 -352
rect -17 424 17 440
rect -17 -368 17 -352
rect 121 424 155 440
rect 121 -368 155 -352
rect 259 424 293 440
rect 259 -368 293 -352
rect 397 424 431 440
rect 397 -368 431 -352
rect 535 424 569 440
rect 535 -368 569 -352
rect 673 424 707 440
rect 673 -368 707 -352
rect 811 424 845 440
rect 811 -368 845 -352
rect 949 424 983 440
rect 949 -368 983 -352
rect 1087 424 1121 440
rect 1087 -368 1121 -352
rect 1225 424 1259 440
rect 1225 -368 1259 -352
rect 1363 424 1397 440
rect 1363 -368 1397 -352
rect 1501 424 1535 440
rect 1501 -368 1535 -352
rect 1639 424 1673 440
rect 1639 -368 1673 -352
rect 1777 424 1811 440
rect 1777 -368 1811 -352
rect 1915 424 1949 440
rect 1915 -368 1949 -352
rect 2053 424 2087 440
rect 2053 -368 2087 -352
rect 2191 424 2225 440
rect 2191 -368 2225 -352
rect 2329 424 2363 440
rect 2329 -368 2363 -352
rect 2467 424 2501 440
rect 2467 -368 2501 -352
rect 2605 424 2639 440
rect 2605 -368 2639 -352
rect 2743 424 2777 440
rect 2743 -368 2777 -352
rect 2881 424 2915 440
rect 2881 -368 2915 -352
rect 3019 424 3053 440
rect 3019 -368 3053 -352
rect 3157 424 3191 440
rect 3157 -368 3191 -352
rect 3295 424 3329 440
rect 3295 -368 3329 -352
rect 3433 424 3467 440
rect 3433 -368 3467 -352
rect 3571 424 3605 440
rect 3571 -368 3605 -352
rect 3709 424 3743 440
rect 3709 -368 3743 -352
rect 3847 424 3881 440
rect 3847 -368 3881 -352
rect 3985 424 4019 440
rect 3985 -368 4019 -352
rect 4123 424 4157 440
rect 4123 -368 4157 -352
rect 4261 424 4295 440
rect 4261 -368 4295 -352
rect 4399 424 4433 440
rect 4399 -368 4433 -352
rect 4537 424 4571 440
rect 4537 -368 4571 -352
rect 4675 424 4709 440
rect 4675 -368 4709 -352
rect 4813 424 4847 440
rect 4813 -368 4847 -352
rect 4951 424 4985 440
rect 4951 -368 4985 -352
rect 5089 424 5123 440
rect 5089 -368 5123 -352
rect 5227 424 5261 440
rect 5227 -368 5261 -352
rect 5365 424 5399 440
rect 5365 -368 5399 -352
rect 5503 424 5537 440
rect 5503 -368 5537 -352
rect 5641 424 5675 440
rect 5641 -368 5675 -352
rect 5779 424 5813 440
rect 5779 -368 5813 -352
rect 5917 424 5951 440
rect 5917 -368 5951 -352
rect 6055 424 6089 440
rect 6055 -368 6089 -352
rect 6193 424 6227 440
rect 6193 -368 6227 -352
rect 6331 424 6365 440
rect 6331 -368 6365 -352
rect 6469 424 6503 440
rect 6469 -368 6503 -352
rect 6607 424 6641 440
rect 6607 -368 6641 -352
rect 6745 424 6779 440
rect 6745 -368 6779 -352
rect 6883 424 6917 440
rect 6883 -368 6917 -352
rect -6871 -445 -6855 -411
rect -6807 -445 -6791 -411
rect -6733 -445 -6717 -411
rect -6669 -445 -6653 -411
rect -6595 -445 -6579 -411
rect -6531 -445 -6515 -411
rect -6457 -445 -6441 -411
rect -6393 -445 -6377 -411
rect -6319 -445 -6303 -411
rect -6255 -445 -6239 -411
rect -6181 -445 -6165 -411
rect -6117 -445 -6101 -411
rect -6043 -445 -6027 -411
rect -5979 -445 -5963 -411
rect -5905 -445 -5889 -411
rect -5841 -445 -5825 -411
rect -5767 -445 -5751 -411
rect -5703 -445 -5687 -411
rect -5629 -445 -5613 -411
rect -5565 -445 -5549 -411
rect -5491 -445 -5475 -411
rect -5427 -445 -5411 -411
rect -5353 -445 -5337 -411
rect -5289 -445 -5273 -411
rect -5215 -445 -5199 -411
rect -5151 -445 -5135 -411
rect -5077 -445 -5061 -411
rect -5013 -445 -4997 -411
rect -4939 -445 -4923 -411
rect -4875 -445 -4859 -411
rect -4801 -445 -4785 -411
rect -4737 -445 -4721 -411
rect -4663 -445 -4647 -411
rect -4599 -445 -4583 -411
rect -4525 -445 -4509 -411
rect -4461 -445 -4445 -411
rect -4387 -445 -4371 -411
rect -4323 -445 -4307 -411
rect -4249 -445 -4233 -411
rect -4185 -445 -4169 -411
rect -4111 -445 -4095 -411
rect -4047 -445 -4031 -411
rect -3973 -445 -3957 -411
rect -3909 -445 -3893 -411
rect -3835 -445 -3819 -411
rect -3771 -445 -3755 -411
rect -3697 -445 -3681 -411
rect -3633 -445 -3617 -411
rect -3559 -445 -3543 -411
rect -3495 -445 -3479 -411
rect -3421 -445 -3405 -411
rect -3357 -445 -3341 -411
rect -3283 -445 -3267 -411
rect -3219 -445 -3203 -411
rect -3145 -445 -3129 -411
rect -3081 -445 -3065 -411
rect -3007 -445 -2991 -411
rect -2943 -445 -2927 -411
rect -2869 -445 -2853 -411
rect -2805 -445 -2789 -411
rect -2731 -445 -2715 -411
rect -2667 -445 -2651 -411
rect -2593 -445 -2577 -411
rect -2529 -445 -2513 -411
rect -2455 -445 -2439 -411
rect -2391 -445 -2375 -411
rect -2317 -445 -2301 -411
rect -2253 -445 -2237 -411
rect -2179 -445 -2163 -411
rect -2115 -445 -2099 -411
rect -2041 -445 -2025 -411
rect -1977 -445 -1961 -411
rect -1903 -445 -1887 -411
rect -1839 -445 -1823 -411
rect -1765 -445 -1749 -411
rect -1701 -445 -1685 -411
rect -1627 -445 -1611 -411
rect -1563 -445 -1547 -411
rect -1489 -445 -1473 -411
rect -1425 -445 -1409 -411
rect -1351 -445 -1335 -411
rect -1287 -445 -1271 -411
rect -1213 -445 -1197 -411
rect -1149 -445 -1133 -411
rect -1075 -445 -1059 -411
rect -1011 -445 -995 -411
rect -937 -445 -921 -411
rect -873 -445 -857 -411
rect -799 -445 -783 -411
rect -735 -445 -719 -411
rect -661 -445 -645 -411
rect -597 -445 -581 -411
rect -523 -445 -507 -411
rect -459 -445 -443 -411
rect -385 -445 -369 -411
rect -321 -445 -305 -411
rect -247 -445 -231 -411
rect -183 -445 -167 -411
rect -109 -445 -93 -411
rect -45 -445 -29 -411
rect 29 -445 45 -411
rect 93 -445 109 -411
rect 167 -445 183 -411
rect 231 -445 247 -411
rect 305 -445 321 -411
rect 369 -445 385 -411
rect 443 -445 459 -411
rect 507 -445 523 -411
rect 581 -445 597 -411
rect 645 -445 661 -411
rect 719 -445 735 -411
rect 783 -445 799 -411
rect 857 -445 873 -411
rect 921 -445 937 -411
rect 995 -445 1011 -411
rect 1059 -445 1075 -411
rect 1133 -445 1149 -411
rect 1197 -445 1213 -411
rect 1271 -445 1287 -411
rect 1335 -445 1351 -411
rect 1409 -445 1425 -411
rect 1473 -445 1489 -411
rect 1547 -445 1563 -411
rect 1611 -445 1627 -411
rect 1685 -445 1701 -411
rect 1749 -445 1765 -411
rect 1823 -445 1839 -411
rect 1887 -445 1903 -411
rect 1961 -445 1977 -411
rect 2025 -445 2041 -411
rect 2099 -445 2115 -411
rect 2163 -445 2179 -411
rect 2237 -445 2253 -411
rect 2301 -445 2317 -411
rect 2375 -445 2391 -411
rect 2439 -445 2455 -411
rect 2513 -445 2529 -411
rect 2577 -445 2593 -411
rect 2651 -445 2667 -411
rect 2715 -445 2731 -411
rect 2789 -445 2805 -411
rect 2853 -445 2869 -411
rect 2927 -445 2943 -411
rect 2991 -445 3007 -411
rect 3065 -445 3081 -411
rect 3129 -445 3145 -411
rect 3203 -445 3219 -411
rect 3267 -445 3283 -411
rect 3341 -445 3357 -411
rect 3405 -445 3421 -411
rect 3479 -445 3495 -411
rect 3543 -445 3559 -411
rect 3617 -445 3633 -411
rect 3681 -445 3697 -411
rect 3755 -445 3771 -411
rect 3819 -445 3835 -411
rect 3893 -445 3909 -411
rect 3957 -445 3973 -411
rect 4031 -445 4047 -411
rect 4095 -445 4111 -411
rect 4169 -445 4185 -411
rect 4233 -445 4249 -411
rect 4307 -445 4323 -411
rect 4371 -445 4387 -411
rect 4445 -445 4461 -411
rect 4509 -445 4525 -411
rect 4583 -445 4599 -411
rect 4647 -445 4663 -411
rect 4721 -445 4737 -411
rect 4785 -445 4801 -411
rect 4859 -445 4875 -411
rect 4923 -445 4939 -411
rect 4997 -445 5013 -411
rect 5061 -445 5077 -411
rect 5135 -445 5151 -411
rect 5199 -445 5215 -411
rect 5273 -445 5289 -411
rect 5337 -445 5353 -411
rect 5411 -445 5427 -411
rect 5475 -445 5491 -411
rect 5549 -445 5565 -411
rect 5613 -445 5629 -411
rect 5687 -445 5703 -411
rect 5751 -445 5767 -411
rect 5825 -445 5841 -411
rect 5889 -445 5905 -411
rect 5963 -445 5979 -411
rect 6027 -445 6043 -411
rect 6101 -445 6117 -411
rect 6165 -445 6181 -411
rect 6239 -445 6255 -411
rect 6303 -445 6319 -411
rect 6377 -445 6393 -411
rect 6441 -445 6457 -411
rect 6515 -445 6531 -411
rect 6579 -445 6595 -411
rect 6653 -445 6669 -411
rect 6717 -445 6733 -411
rect 6791 -445 6807 -411
rect 6855 -445 6871 -411
<< viali >>
rect -6917 -352 -6883 424
rect -6779 -352 -6745 424
rect -6641 -352 -6607 424
rect -6503 -352 -6469 424
rect -6365 -352 -6331 424
rect -6227 -352 -6193 424
rect -6089 -352 -6055 424
rect -5951 -352 -5917 424
rect -5813 -352 -5779 424
rect -5675 -352 -5641 424
rect -5537 -352 -5503 424
rect -5399 -352 -5365 424
rect -5261 -352 -5227 424
rect -5123 -352 -5089 424
rect -4985 -352 -4951 424
rect -4847 -352 -4813 424
rect -4709 -352 -4675 424
rect -4571 -352 -4537 424
rect -4433 -352 -4399 424
rect -4295 -352 -4261 424
rect -4157 -352 -4123 424
rect -4019 -352 -3985 424
rect -3881 -352 -3847 424
rect -3743 -352 -3709 424
rect -3605 -352 -3571 424
rect -3467 -352 -3433 424
rect -3329 -352 -3295 424
rect -3191 -352 -3157 424
rect -3053 -352 -3019 424
rect -2915 -352 -2881 424
rect -2777 -352 -2743 424
rect -2639 -352 -2605 424
rect -2501 -352 -2467 424
rect -2363 -352 -2329 424
rect -2225 -352 -2191 424
rect -2087 -352 -2053 424
rect -1949 -352 -1915 424
rect -1811 -352 -1777 424
rect -1673 -352 -1639 424
rect -1535 -352 -1501 424
rect -1397 -352 -1363 424
rect -1259 -352 -1225 424
rect -1121 -352 -1087 424
rect -983 -352 -949 424
rect -845 -352 -811 424
rect -707 -352 -673 424
rect -569 -352 -535 424
rect -431 -352 -397 424
rect -293 -352 -259 424
rect -155 -352 -121 424
rect -17 -352 17 424
rect 121 -352 155 424
rect 259 -352 293 424
rect 397 -352 431 424
rect 535 -352 569 424
rect 673 -352 707 424
rect 811 -352 845 424
rect 949 -352 983 424
rect 1087 -352 1121 424
rect 1225 -352 1259 424
rect 1363 -352 1397 424
rect 1501 -352 1535 424
rect 1639 -352 1673 424
rect 1777 -352 1811 424
rect 1915 -352 1949 424
rect 2053 -352 2087 424
rect 2191 -352 2225 424
rect 2329 -352 2363 424
rect 2467 -352 2501 424
rect 2605 -352 2639 424
rect 2743 -352 2777 424
rect 2881 -352 2915 424
rect 3019 -352 3053 424
rect 3157 -352 3191 424
rect 3295 -352 3329 424
rect 3433 -352 3467 424
rect 3571 -352 3605 424
rect 3709 -352 3743 424
rect 3847 -352 3881 424
rect 3985 -352 4019 424
rect 4123 -352 4157 424
rect 4261 -352 4295 424
rect 4399 -352 4433 424
rect 4537 -352 4571 424
rect 4675 -352 4709 424
rect 4813 -352 4847 424
rect 4951 -352 4985 424
rect 5089 -352 5123 424
rect 5227 -352 5261 424
rect 5365 -352 5399 424
rect 5503 -352 5537 424
rect 5641 -352 5675 424
rect 5779 -352 5813 424
rect 5917 -352 5951 424
rect 6055 -352 6089 424
rect 6193 -352 6227 424
rect 6331 -352 6365 424
rect 6469 -352 6503 424
rect 6607 -352 6641 424
rect 6745 -352 6779 424
rect 6883 -352 6917 424
rect -6855 -445 -6807 -411
rect -6717 -445 -6669 -411
rect -6579 -445 -6531 -411
rect -6441 -445 -6393 -411
rect -6303 -445 -6255 -411
rect -6165 -445 -6117 -411
rect -6027 -445 -5979 -411
rect -5889 -445 -5841 -411
rect -5751 -445 -5703 -411
rect -5613 -445 -5565 -411
rect -5475 -445 -5427 -411
rect -5337 -445 -5289 -411
rect -5199 -445 -5151 -411
rect -5061 -445 -5013 -411
rect -4923 -445 -4875 -411
rect -4785 -445 -4737 -411
rect -4647 -445 -4599 -411
rect -4509 -445 -4461 -411
rect -4371 -445 -4323 -411
rect -4233 -445 -4185 -411
rect -4095 -445 -4047 -411
rect -3957 -445 -3909 -411
rect -3819 -445 -3771 -411
rect -3681 -445 -3633 -411
rect -3543 -445 -3495 -411
rect -3405 -445 -3357 -411
rect -3267 -445 -3219 -411
rect -3129 -445 -3081 -411
rect -2991 -445 -2943 -411
rect -2853 -445 -2805 -411
rect -2715 -445 -2667 -411
rect -2577 -445 -2529 -411
rect -2439 -445 -2391 -411
rect -2301 -445 -2253 -411
rect -2163 -445 -2115 -411
rect -2025 -445 -1977 -411
rect -1887 -445 -1839 -411
rect -1749 -445 -1701 -411
rect -1611 -445 -1563 -411
rect -1473 -445 -1425 -411
rect -1335 -445 -1287 -411
rect -1197 -445 -1149 -411
rect -1059 -445 -1011 -411
rect -921 -445 -873 -411
rect -783 -445 -735 -411
rect -645 -445 -597 -411
rect -507 -445 -459 -411
rect -369 -445 -321 -411
rect -231 -445 -183 -411
rect -93 -445 -45 -411
rect 45 -445 93 -411
rect 183 -445 231 -411
rect 321 -445 369 -411
rect 459 -445 507 -411
rect 597 -445 645 -411
rect 735 -445 783 -411
rect 873 -445 921 -411
rect 1011 -445 1059 -411
rect 1149 -445 1197 -411
rect 1287 -445 1335 -411
rect 1425 -445 1473 -411
rect 1563 -445 1611 -411
rect 1701 -445 1749 -411
rect 1839 -445 1887 -411
rect 1977 -445 2025 -411
rect 2115 -445 2163 -411
rect 2253 -445 2301 -411
rect 2391 -445 2439 -411
rect 2529 -445 2577 -411
rect 2667 -445 2715 -411
rect 2805 -445 2853 -411
rect 2943 -445 2991 -411
rect 3081 -445 3129 -411
rect 3219 -445 3267 -411
rect 3357 -445 3405 -411
rect 3495 -445 3543 -411
rect 3633 -445 3681 -411
rect 3771 -445 3819 -411
rect 3909 -445 3957 -411
rect 4047 -445 4095 -411
rect 4185 -445 4233 -411
rect 4323 -445 4371 -411
rect 4461 -445 4509 -411
rect 4599 -445 4647 -411
rect 4737 -445 4785 -411
rect 4875 -445 4923 -411
rect 5013 -445 5061 -411
rect 5151 -445 5199 -411
rect 5289 -445 5337 -411
rect 5427 -445 5475 -411
rect 5565 -445 5613 -411
rect 5703 -445 5751 -411
rect 5841 -445 5889 -411
rect 5979 -445 6027 -411
rect 6117 -445 6165 -411
rect 6255 -445 6303 -411
rect 6393 -445 6441 -411
rect 6531 -445 6579 -411
rect 6669 -445 6717 -411
rect 6807 -445 6855 -411
<< metal1 >>
rect -6923 424 -6877 436
rect -6923 -352 -6917 424
rect -6883 -352 -6877 424
rect -6923 -364 -6877 -352
rect -6785 424 -6739 436
rect -6785 -352 -6779 424
rect -6745 -352 -6739 424
rect -6785 -364 -6739 -352
rect -6647 424 -6601 436
rect -6647 -352 -6641 424
rect -6607 -352 -6601 424
rect -6647 -364 -6601 -352
rect -6509 424 -6463 436
rect -6509 -352 -6503 424
rect -6469 -352 -6463 424
rect -6509 -364 -6463 -352
rect -6371 424 -6325 436
rect -6371 -352 -6365 424
rect -6331 -352 -6325 424
rect -6371 -364 -6325 -352
rect -6233 424 -6187 436
rect -6233 -352 -6227 424
rect -6193 -352 -6187 424
rect -6233 -364 -6187 -352
rect -6095 424 -6049 436
rect -6095 -352 -6089 424
rect -6055 -352 -6049 424
rect -6095 -364 -6049 -352
rect -5957 424 -5911 436
rect -5957 -352 -5951 424
rect -5917 -352 -5911 424
rect -5957 -364 -5911 -352
rect -5819 424 -5773 436
rect -5819 -352 -5813 424
rect -5779 -352 -5773 424
rect -5819 -364 -5773 -352
rect -5681 424 -5635 436
rect -5681 -352 -5675 424
rect -5641 -352 -5635 424
rect -5681 -364 -5635 -352
rect -5543 424 -5497 436
rect -5543 -352 -5537 424
rect -5503 -352 -5497 424
rect -5543 -364 -5497 -352
rect -5405 424 -5359 436
rect -5405 -352 -5399 424
rect -5365 -352 -5359 424
rect -5405 -364 -5359 -352
rect -5267 424 -5221 436
rect -5267 -352 -5261 424
rect -5227 -352 -5221 424
rect -5267 -364 -5221 -352
rect -5129 424 -5083 436
rect -5129 -352 -5123 424
rect -5089 -352 -5083 424
rect -5129 -364 -5083 -352
rect -4991 424 -4945 436
rect -4991 -352 -4985 424
rect -4951 -352 -4945 424
rect -4991 -364 -4945 -352
rect -4853 424 -4807 436
rect -4853 -352 -4847 424
rect -4813 -352 -4807 424
rect -4853 -364 -4807 -352
rect -4715 424 -4669 436
rect -4715 -352 -4709 424
rect -4675 -352 -4669 424
rect -4715 -364 -4669 -352
rect -4577 424 -4531 436
rect -4577 -352 -4571 424
rect -4537 -352 -4531 424
rect -4577 -364 -4531 -352
rect -4439 424 -4393 436
rect -4439 -352 -4433 424
rect -4399 -352 -4393 424
rect -4439 -364 -4393 -352
rect -4301 424 -4255 436
rect -4301 -352 -4295 424
rect -4261 -352 -4255 424
rect -4301 -364 -4255 -352
rect -4163 424 -4117 436
rect -4163 -352 -4157 424
rect -4123 -352 -4117 424
rect -4163 -364 -4117 -352
rect -4025 424 -3979 436
rect -4025 -352 -4019 424
rect -3985 -352 -3979 424
rect -4025 -364 -3979 -352
rect -3887 424 -3841 436
rect -3887 -352 -3881 424
rect -3847 -352 -3841 424
rect -3887 -364 -3841 -352
rect -3749 424 -3703 436
rect -3749 -352 -3743 424
rect -3709 -352 -3703 424
rect -3749 -364 -3703 -352
rect -3611 424 -3565 436
rect -3611 -352 -3605 424
rect -3571 -352 -3565 424
rect -3611 -364 -3565 -352
rect -3473 424 -3427 436
rect -3473 -352 -3467 424
rect -3433 -352 -3427 424
rect -3473 -364 -3427 -352
rect -3335 424 -3289 436
rect -3335 -352 -3329 424
rect -3295 -352 -3289 424
rect -3335 -364 -3289 -352
rect -3197 424 -3151 436
rect -3197 -352 -3191 424
rect -3157 -352 -3151 424
rect -3197 -364 -3151 -352
rect -3059 424 -3013 436
rect -3059 -352 -3053 424
rect -3019 -352 -3013 424
rect -3059 -364 -3013 -352
rect -2921 424 -2875 436
rect -2921 -352 -2915 424
rect -2881 -352 -2875 424
rect -2921 -364 -2875 -352
rect -2783 424 -2737 436
rect -2783 -352 -2777 424
rect -2743 -352 -2737 424
rect -2783 -364 -2737 -352
rect -2645 424 -2599 436
rect -2645 -352 -2639 424
rect -2605 -352 -2599 424
rect -2645 -364 -2599 -352
rect -2507 424 -2461 436
rect -2507 -352 -2501 424
rect -2467 -352 -2461 424
rect -2507 -364 -2461 -352
rect -2369 424 -2323 436
rect -2369 -352 -2363 424
rect -2329 -352 -2323 424
rect -2369 -364 -2323 -352
rect -2231 424 -2185 436
rect -2231 -352 -2225 424
rect -2191 -352 -2185 424
rect -2231 -364 -2185 -352
rect -2093 424 -2047 436
rect -2093 -352 -2087 424
rect -2053 -352 -2047 424
rect -2093 -364 -2047 -352
rect -1955 424 -1909 436
rect -1955 -352 -1949 424
rect -1915 -352 -1909 424
rect -1955 -364 -1909 -352
rect -1817 424 -1771 436
rect -1817 -352 -1811 424
rect -1777 -352 -1771 424
rect -1817 -364 -1771 -352
rect -1679 424 -1633 436
rect -1679 -352 -1673 424
rect -1639 -352 -1633 424
rect -1679 -364 -1633 -352
rect -1541 424 -1495 436
rect -1541 -352 -1535 424
rect -1501 -352 -1495 424
rect -1541 -364 -1495 -352
rect -1403 424 -1357 436
rect -1403 -352 -1397 424
rect -1363 -352 -1357 424
rect -1403 -364 -1357 -352
rect -1265 424 -1219 436
rect -1265 -352 -1259 424
rect -1225 -352 -1219 424
rect -1265 -364 -1219 -352
rect -1127 424 -1081 436
rect -1127 -352 -1121 424
rect -1087 -352 -1081 424
rect -1127 -364 -1081 -352
rect -989 424 -943 436
rect -989 -352 -983 424
rect -949 -352 -943 424
rect -989 -364 -943 -352
rect -851 424 -805 436
rect -851 -352 -845 424
rect -811 -352 -805 424
rect -851 -364 -805 -352
rect -713 424 -667 436
rect -713 -352 -707 424
rect -673 -352 -667 424
rect -713 -364 -667 -352
rect -575 424 -529 436
rect -575 -352 -569 424
rect -535 -352 -529 424
rect -575 -364 -529 -352
rect -437 424 -391 436
rect -437 -352 -431 424
rect -397 -352 -391 424
rect -437 -364 -391 -352
rect -299 424 -253 436
rect -299 -352 -293 424
rect -259 -352 -253 424
rect -299 -364 -253 -352
rect -161 424 -115 436
rect -161 -352 -155 424
rect -121 -352 -115 424
rect -161 -364 -115 -352
rect -23 424 23 436
rect -23 -352 -17 424
rect 17 -352 23 424
rect -23 -364 23 -352
rect 115 424 161 436
rect 115 -352 121 424
rect 155 -352 161 424
rect 115 -364 161 -352
rect 253 424 299 436
rect 253 -352 259 424
rect 293 -352 299 424
rect 253 -364 299 -352
rect 391 424 437 436
rect 391 -352 397 424
rect 431 -352 437 424
rect 391 -364 437 -352
rect 529 424 575 436
rect 529 -352 535 424
rect 569 -352 575 424
rect 529 -364 575 -352
rect 667 424 713 436
rect 667 -352 673 424
rect 707 -352 713 424
rect 667 -364 713 -352
rect 805 424 851 436
rect 805 -352 811 424
rect 845 -352 851 424
rect 805 -364 851 -352
rect 943 424 989 436
rect 943 -352 949 424
rect 983 -352 989 424
rect 943 -364 989 -352
rect 1081 424 1127 436
rect 1081 -352 1087 424
rect 1121 -352 1127 424
rect 1081 -364 1127 -352
rect 1219 424 1265 436
rect 1219 -352 1225 424
rect 1259 -352 1265 424
rect 1219 -364 1265 -352
rect 1357 424 1403 436
rect 1357 -352 1363 424
rect 1397 -352 1403 424
rect 1357 -364 1403 -352
rect 1495 424 1541 436
rect 1495 -352 1501 424
rect 1535 -352 1541 424
rect 1495 -364 1541 -352
rect 1633 424 1679 436
rect 1633 -352 1639 424
rect 1673 -352 1679 424
rect 1633 -364 1679 -352
rect 1771 424 1817 436
rect 1771 -352 1777 424
rect 1811 -352 1817 424
rect 1771 -364 1817 -352
rect 1909 424 1955 436
rect 1909 -352 1915 424
rect 1949 -352 1955 424
rect 1909 -364 1955 -352
rect 2047 424 2093 436
rect 2047 -352 2053 424
rect 2087 -352 2093 424
rect 2047 -364 2093 -352
rect 2185 424 2231 436
rect 2185 -352 2191 424
rect 2225 -352 2231 424
rect 2185 -364 2231 -352
rect 2323 424 2369 436
rect 2323 -352 2329 424
rect 2363 -352 2369 424
rect 2323 -364 2369 -352
rect 2461 424 2507 436
rect 2461 -352 2467 424
rect 2501 -352 2507 424
rect 2461 -364 2507 -352
rect 2599 424 2645 436
rect 2599 -352 2605 424
rect 2639 -352 2645 424
rect 2599 -364 2645 -352
rect 2737 424 2783 436
rect 2737 -352 2743 424
rect 2777 -352 2783 424
rect 2737 -364 2783 -352
rect 2875 424 2921 436
rect 2875 -352 2881 424
rect 2915 -352 2921 424
rect 2875 -364 2921 -352
rect 3013 424 3059 436
rect 3013 -352 3019 424
rect 3053 -352 3059 424
rect 3013 -364 3059 -352
rect 3151 424 3197 436
rect 3151 -352 3157 424
rect 3191 -352 3197 424
rect 3151 -364 3197 -352
rect 3289 424 3335 436
rect 3289 -352 3295 424
rect 3329 -352 3335 424
rect 3289 -364 3335 -352
rect 3427 424 3473 436
rect 3427 -352 3433 424
rect 3467 -352 3473 424
rect 3427 -364 3473 -352
rect 3565 424 3611 436
rect 3565 -352 3571 424
rect 3605 -352 3611 424
rect 3565 -364 3611 -352
rect 3703 424 3749 436
rect 3703 -352 3709 424
rect 3743 -352 3749 424
rect 3703 -364 3749 -352
rect 3841 424 3887 436
rect 3841 -352 3847 424
rect 3881 -352 3887 424
rect 3841 -364 3887 -352
rect 3979 424 4025 436
rect 3979 -352 3985 424
rect 4019 -352 4025 424
rect 3979 -364 4025 -352
rect 4117 424 4163 436
rect 4117 -352 4123 424
rect 4157 -352 4163 424
rect 4117 -364 4163 -352
rect 4255 424 4301 436
rect 4255 -352 4261 424
rect 4295 -352 4301 424
rect 4255 -364 4301 -352
rect 4393 424 4439 436
rect 4393 -352 4399 424
rect 4433 -352 4439 424
rect 4393 -364 4439 -352
rect 4531 424 4577 436
rect 4531 -352 4537 424
rect 4571 -352 4577 424
rect 4531 -364 4577 -352
rect 4669 424 4715 436
rect 4669 -352 4675 424
rect 4709 -352 4715 424
rect 4669 -364 4715 -352
rect 4807 424 4853 436
rect 4807 -352 4813 424
rect 4847 -352 4853 424
rect 4807 -364 4853 -352
rect 4945 424 4991 436
rect 4945 -352 4951 424
rect 4985 -352 4991 424
rect 4945 -364 4991 -352
rect 5083 424 5129 436
rect 5083 -352 5089 424
rect 5123 -352 5129 424
rect 5083 -364 5129 -352
rect 5221 424 5267 436
rect 5221 -352 5227 424
rect 5261 -352 5267 424
rect 5221 -364 5267 -352
rect 5359 424 5405 436
rect 5359 -352 5365 424
rect 5399 -352 5405 424
rect 5359 -364 5405 -352
rect 5497 424 5543 436
rect 5497 -352 5503 424
rect 5537 -352 5543 424
rect 5497 -364 5543 -352
rect 5635 424 5681 436
rect 5635 -352 5641 424
rect 5675 -352 5681 424
rect 5635 -364 5681 -352
rect 5773 424 5819 436
rect 5773 -352 5779 424
rect 5813 -352 5819 424
rect 5773 -364 5819 -352
rect 5911 424 5957 436
rect 5911 -352 5917 424
rect 5951 -352 5957 424
rect 5911 -364 5957 -352
rect 6049 424 6095 436
rect 6049 -352 6055 424
rect 6089 -352 6095 424
rect 6049 -364 6095 -352
rect 6187 424 6233 436
rect 6187 -352 6193 424
rect 6227 -352 6233 424
rect 6187 -364 6233 -352
rect 6325 424 6371 436
rect 6325 -352 6331 424
rect 6365 -352 6371 424
rect 6325 -364 6371 -352
rect 6463 424 6509 436
rect 6463 -352 6469 424
rect 6503 -352 6509 424
rect 6463 -364 6509 -352
rect 6601 424 6647 436
rect 6601 -352 6607 424
rect 6641 -352 6647 424
rect 6601 -364 6647 -352
rect 6739 424 6785 436
rect 6739 -352 6745 424
rect 6779 -352 6785 424
rect 6739 -364 6785 -352
rect 6877 424 6923 436
rect 6877 -352 6883 424
rect 6917 -352 6923 424
rect 6877 -364 6923 -352
rect -6867 -411 -6795 -405
rect -6867 -445 -6855 -411
rect -6807 -445 -6795 -411
rect -6867 -451 -6795 -445
rect -6729 -411 -6657 -405
rect -6729 -445 -6717 -411
rect -6669 -445 -6657 -411
rect -6729 -451 -6657 -445
rect -6591 -411 -6519 -405
rect -6591 -445 -6579 -411
rect -6531 -445 -6519 -411
rect -6591 -451 -6519 -445
rect -6453 -411 -6381 -405
rect -6453 -445 -6441 -411
rect -6393 -445 -6381 -411
rect -6453 -451 -6381 -445
rect -6315 -411 -6243 -405
rect -6315 -445 -6303 -411
rect -6255 -445 -6243 -411
rect -6315 -451 -6243 -445
rect -6177 -411 -6105 -405
rect -6177 -445 -6165 -411
rect -6117 -445 -6105 -411
rect -6177 -451 -6105 -445
rect -6039 -411 -5967 -405
rect -6039 -445 -6027 -411
rect -5979 -445 -5967 -411
rect -6039 -451 -5967 -445
rect -5901 -411 -5829 -405
rect -5901 -445 -5889 -411
rect -5841 -445 -5829 -411
rect -5901 -451 -5829 -445
rect -5763 -411 -5691 -405
rect -5763 -445 -5751 -411
rect -5703 -445 -5691 -411
rect -5763 -451 -5691 -445
rect -5625 -411 -5553 -405
rect -5625 -445 -5613 -411
rect -5565 -445 -5553 -411
rect -5625 -451 -5553 -445
rect -5487 -411 -5415 -405
rect -5487 -445 -5475 -411
rect -5427 -445 -5415 -411
rect -5487 -451 -5415 -445
rect -5349 -411 -5277 -405
rect -5349 -445 -5337 -411
rect -5289 -445 -5277 -411
rect -5349 -451 -5277 -445
rect -5211 -411 -5139 -405
rect -5211 -445 -5199 -411
rect -5151 -445 -5139 -411
rect -5211 -451 -5139 -445
rect -5073 -411 -5001 -405
rect -5073 -445 -5061 -411
rect -5013 -445 -5001 -411
rect -5073 -451 -5001 -445
rect -4935 -411 -4863 -405
rect -4935 -445 -4923 -411
rect -4875 -445 -4863 -411
rect -4935 -451 -4863 -445
rect -4797 -411 -4725 -405
rect -4797 -445 -4785 -411
rect -4737 -445 -4725 -411
rect -4797 -451 -4725 -445
rect -4659 -411 -4587 -405
rect -4659 -445 -4647 -411
rect -4599 -445 -4587 -411
rect -4659 -451 -4587 -445
rect -4521 -411 -4449 -405
rect -4521 -445 -4509 -411
rect -4461 -445 -4449 -411
rect -4521 -451 -4449 -445
rect -4383 -411 -4311 -405
rect -4383 -445 -4371 -411
rect -4323 -445 -4311 -411
rect -4383 -451 -4311 -445
rect -4245 -411 -4173 -405
rect -4245 -445 -4233 -411
rect -4185 -445 -4173 -411
rect -4245 -451 -4173 -445
rect -4107 -411 -4035 -405
rect -4107 -445 -4095 -411
rect -4047 -445 -4035 -411
rect -4107 -451 -4035 -445
rect -3969 -411 -3897 -405
rect -3969 -445 -3957 -411
rect -3909 -445 -3897 -411
rect -3969 -451 -3897 -445
rect -3831 -411 -3759 -405
rect -3831 -445 -3819 -411
rect -3771 -445 -3759 -411
rect -3831 -451 -3759 -445
rect -3693 -411 -3621 -405
rect -3693 -445 -3681 -411
rect -3633 -445 -3621 -411
rect -3693 -451 -3621 -445
rect -3555 -411 -3483 -405
rect -3555 -445 -3543 -411
rect -3495 -445 -3483 -411
rect -3555 -451 -3483 -445
rect -3417 -411 -3345 -405
rect -3417 -445 -3405 -411
rect -3357 -445 -3345 -411
rect -3417 -451 -3345 -445
rect -3279 -411 -3207 -405
rect -3279 -445 -3267 -411
rect -3219 -445 -3207 -411
rect -3279 -451 -3207 -445
rect -3141 -411 -3069 -405
rect -3141 -445 -3129 -411
rect -3081 -445 -3069 -411
rect -3141 -451 -3069 -445
rect -3003 -411 -2931 -405
rect -3003 -445 -2991 -411
rect -2943 -445 -2931 -411
rect -3003 -451 -2931 -445
rect -2865 -411 -2793 -405
rect -2865 -445 -2853 -411
rect -2805 -445 -2793 -411
rect -2865 -451 -2793 -445
rect -2727 -411 -2655 -405
rect -2727 -445 -2715 -411
rect -2667 -445 -2655 -411
rect -2727 -451 -2655 -445
rect -2589 -411 -2517 -405
rect -2589 -445 -2577 -411
rect -2529 -445 -2517 -411
rect -2589 -451 -2517 -445
rect -2451 -411 -2379 -405
rect -2451 -445 -2439 -411
rect -2391 -445 -2379 -411
rect -2451 -451 -2379 -445
rect -2313 -411 -2241 -405
rect -2313 -445 -2301 -411
rect -2253 -445 -2241 -411
rect -2313 -451 -2241 -445
rect -2175 -411 -2103 -405
rect -2175 -445 -2163 -411
rect -2115 -445 -2103 -411
rect -2175 -451 -2103 -445
rect -2037 -411 -1965 -405
rect -2037 -445 -2025 -411
rect -1977 -445 -1965 -411
rect -2037 -451 -1965 -445
rect -1899 -411 -1827 -405
rect -1899 -445 -1887 -411
rect -1839 -445 -1827 -411
rect -1899 -451 -1827 -445
rect -1761 -411 -1689 -405
rect -1761 -445 -1749 -411
rect -1701 -445 -1689 -411
rect -1761 -451 -1689 -445
rect -1623 -411 -1551 -405
rect -1623 -445 -1611 -411
rect -1563 -445 -1551 -411
rect -1623 -451 -1551 -445
rect -1485 -411 -1413 -405
rect -1485 -445 -1473 -411
rect -1425 -445 -1413 -411
rect -1485 -451 -1413 -445
rect -1347 -411 -1275 -405
rect -1347 -445 -1335 -411
rect -1287 -445 -1275 -411
rect -1347 -451 -1275 -445
rect -1209 -411 -1137 -405
rect -1209 -445 -1197 -411
rect -1149 -445 -1137 -411
rect -1209 -451 -1137 -445
rect -1071 -411 -999 -405
rect -1071 -445 -1059 -411
rect -1011 -445 -999 -411
rect -1071 -451 -999 -445
rect -933 -411 -861 -405
rect -933 -445 -921 -411
rect -873 -445 -861 -411
rect -933 -451 -861 -445
rect -795 -411 -723 -405
rect -795 -445 -783 -411
rect -735 -445 -723 -411
rect -795 -451 -723 -445
rect -657 -411 -585 -405
rect -657 -445 -645 -411
rect -597 -445 -585 -411
rect -657 -451 -585 -445
rect -519 -411 -447 -405
rect -519 -445 -507 -411
rect -459 -445 -447 -411
rect -519 -451 -447 -445
rect -381 -411 -309 -405
rect -381 -445 -369 -411
rect -321 -445 -309 -411
rect -381 -451 -309 -445
rect -243 -411 -171 -405
rect -243 -445 -231 -411
rect -183 -445 -171 -411
rect -243 -451 -171 -445
rect -105 -411 -33 -405
rect -105 -445 -93 -411
rect -45 -445 -33 -411
rect -105 -451 -33 -445
rect 33 -411 105 -405
rect 33 -445 45 -411
rect 93 -445 105 -411
rect 33 -451 105 -445
rect 171 -411 243 -405
rect 171 -445 183 -411
rect 231 -445 243 -411
rect 171 -451 243 -445
rect 309 -411 381 -405
rect 309 -445 321 -411
rect 369 -445 381 -411
rect 309 -451 381 -445
rect 447 -411 519 -405
rect 447 -445 459 -411
rect 507 -445 519 -411
rect 447 -451 519 -445
rect 585 -411 657 -405
rect 585 -445 597 -411
rect 645 -445 657 -411
rect 585 -451 657 -445
rect 723 -411 795 -405
rect 723 -445 735 -411
rect 783 -445 795 -411
rect 723 -451 795 -445
rect 861 -411 933 -405
rect 861 -445 873 -411
rect 921 -445 933 -411
rect 861 -451 933 -445
rect 999 -411 1071 -405
rect 999 -445 1011 -411
rect 1059 -445 1071 -411
rect 999 -451 1071 -445
rect 1137 -411 1209 -405
rect 1137 -445 1149 -411
rect 1197 -445 1209 -411
rect 1137 -451 1209 -445
rect 1275 -411 1347 -405
rect 1275 -445 1287 -411
rect 1335 -445 1347 -411
rect 1275 -451 1347 -445
rect 1413 -411 1485 -405
rect 1413 -445 1425 -411
rect 1473 -445 1485 -411
rect 1413 -451 1485 -445
rect 1551 -411 1623 -405
rect 1551 -445 1563 -411
rect 1611 -445 1623 -411
rect 1551 -451 1623 -445
rect 1689 -411 1761 -405
rect 1689 -445 1701 -411
rect 1749 -445 1761 -411
rect 1689 -451 1761 -445
rect 1827 -411 1899 -405
rect 1827 -445 1839 -411
rect 1887 -445 1899 -411
rect 1827 -451 1899 -445
rect 1965 -411 2037 -405
rect 1965 -445 1977 -411
rect 2025 -445 2037 -411
rect 1965 -451 2037 -445
rect 2103 -411 2175 -405
rect 2103 -445 2115 -411
rect 2163 -445 2175 -411
rect 2103 -451 2175 -445
rect 2241 -411 2313 -405
rect 2241 -445 2253 -411
rect 2301 -445 2313 -411
rect 2241 -451 2313 -445
rect 2379 -411 2451 -405
rect 2379 -445 2391 -411
rect 2439 -445 2451 -411
rect 2379 -451 2451 -445
rect 2517 -411 2589 -405
rect 2517 -445 2529 -411
rect 2577 -445 2589 -411
rect 2517 -451 2589 -445
rect 2655 -411 2727 -405
rect 2655 -445 2667 -411
rect 2715 -445 2727 -411
rect 2655 -451 2727 -445
rect 2793 -411 2865 -405
rect 2793 -445 2805 -411
rect 2853 -445 2865 -411
rect 2793 -451 2865 -445
rect 2931 -411 3003 -405
rect 2931 -445 2943 -411
rect 2991 -445 3003 -411
rect 2931 -451 3003 -445
rect 3069 -411 3141 -405
rect 3069 -445 3081 -411
rect 3129 -445 3141 -411
rect 3069 -451 3141 -445
rect 3207 -411 3279 -405
rect 3207 -445 3219 -411
rect 3267 -445 3279 -411
rect 3207 -451 3279 -445
rect 3345 -411 3417 -405
rect 3345 -445 3357 -411
rect 3405 -445 3417 -411
rect 3345 -451 3417 -445
rect 3483 -411 3555 -405
rect 3483 -445 3495 -411
rect 3543 -445 3555 -411
rect 3483 -451 3555 -445
rect 3621 -411 3693 -405
rect 3621 -445 3633 -411
rect 3681 -445 3693 -411
rect 3621 -451 3693 -445
rect 3759 -411 3831 -405
rect 3759 -445 3771 -411
rect 3819 -445 3831 -411
rect 3759 -451 3831 -445
rect 3897 -411 3969 -405
rect 3897 -445 3909 -411
rect 3957 -445 3969 -411
rect 3897 -451 3969 -445
rect 4035 -411 4107 -405
rect 4035 -445 4047 -411
rect 4095 -445 4107 -411
rect 4035 -451 4107 -445
rect 4173 -411 4245 -405
rect 4173 -445 4185 -411
rect 4233 -445 4245 -411
rect 4173 -451 4245 -445
rect 4311 -411 4383 -405
rect 4311 -445 4323 -411
rect 4371 -445 4383 -411
rect 4311 -451 4383 -445
rect 4449 -411 4521 -405
rect 4449 -445 4461 -411
rect 4509 -445 4521 -411
rect 4449 -451 4521 -445
rect 4587 -411 4659 -405
rect 4587 -445 4599 -411
rect 4647 -445 4659 -411
rect 4587 -451 4659 -445
rect 4725 -411 4797 -405
rect 4725 -445 4737 -411
rect 4785 -445 4797 -411
rect 4725 -451 4797 -445
rect 4863 -411 4935 -405
rect 4863 -445 4875 -411
rect 4923 -445 4935 -411
rect 4863 -451 4935 -445
rect 5001 -411 5073 -405
rect 5001 -445 5013 -411
rect 5061 -445 5073 -411
rect 5001 -451 5073 -445
rect 5139 -411 5211 -405
rect 5139 -445 5151 -411
rect 5199 -445 5211 -411
rect 5139 -451 5211 -445
rect 5277 -411 5349 -405
rect 5277 -445 5289 -411
rect 5337 -445 5349 -411
rect 5277 -451 5349 -445
rect 5415 -411 5487 -405
rect 5415 -445 5427 -411
rect 5475 -445 5487 -411
rect 5415 -451 5487 -445
rect 5553 -411 5625 -405
rect 5553 -445 5565 -411
rect 5613 -445 5625 -411
rect 5553 -451 5625 -445
rect 5691 -411 5763 -405
rect 5691 -445 5703 -411
rect 5751 -445 5763 -411
rect 5691 -451 5763 -445
rect 5829 -411 5901 -405
rect 5829 -445 5841 -411
rect 5889 -445 5901 -411
rect 5829 -451 5901 -445
rect 5967 -411 6039 -405
rect 5967 -445 5979 -411
rect 6027 -445 6039 -411
rect 5967 -451 6039 -445
rect 6105 -411 6177 -405
rect 6105 -445 6117 -411
rect 6165 -445 6177 -411
rect 6105 -451 6177 -445
rect 6243 -411 6315 -405
rect 6243 -445 6255 -411
rect 6303 -445 6315 -411
rect 6243 -451 6315 -445
rect 6381 -411 6453 -405
rect 6381 -445 6393 -411
rect 6441 -445 6453 -411
rect 6381 -451 6453 -445
rect 6519 -411 6591 -405
rect 6519 -445 6531 -411
rect 6579 -445 6591 -411
rect 6519 -451 6591 -445
rect 6657 -411 6729 -405
rect 6657 -445 6669 -411
rect 6717 -445 6729 -411
rect 6657 -451 6729 -445
rect 6795 -411 6867 -405
rect 6795 -445 6807 -411
rect 6855 -445 6867 -411
rect 6795 -451 6867 -445
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 4 l 0.4 m 1 nf 100 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
