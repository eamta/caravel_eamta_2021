magic
tech sky130A
magscale 1 2
timestamp 1616876989
<< pwell >>
rect -4967 -360 4967 360
<< nmos >>
rect -4767 -150 -4737 150
rect -4671 -150 -4641 150
rect -4575 -150 -4545 150
rect -4479 -150 -4449 150
rect -4383 -150 -4353 150
rect -4287 -150 -4257 150
rect -4191 -150 -4161 150
rect -4095 -150 -4065 150
rect -3999 -150 -3969 150
rect -3903 -150 -3873 150
rect -3807 -150 -3777 150
rect -3711 -150 -3681 150
rect -3615 -150 -3585 150
rect -3519 -150 -3489 150
rect -3423 -150 -3393 150
rect -3327 -150 -3297 150
rect -3231 -150 -3201 150
rect -3135 -150 -3105 150
rect -3039 -150 -3009 150
rect -2943 -150 -2913 150
rect -2847 -150 -2817 150
rect -2751 -150 -2721 150
rect -2655 -150 -2625 150
rect -2559 -150 -2529 150
rect -2463 -150 -2433 150
rect -2367 -150 -2337 150
rect -2271 -150 -2241 150
rect -2175 -150 -2145 150
rect -2079 -150 -2049 150
rect -1983 -150 -1953 150
rect -1887 -150 -1857 150
rect -1791 -150 -1761 150
rect -1695 -150 -1665 150
rect -1599 -150 -1569 150
rect -1503 -150 -1473 150
rect -1407 -150 -1377 150
rect -1311 -150 -1281 150
rect -1215 -150 -1185 150
rect -1119 -150 -1089 150
rect -1023 -150 -993 150
rect -927 -150 -897 150
rect -831 -150 -801 150
rect -735 -150 -705 150
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
rect 705 -150 735 150
rect 801 -150 831 150
rect 897 -150 927 150
rect 993 -150 1023 150
rect 1089 -150 1119 150
rect 1185 -150 1215 150
rect 1281 -150 1311 150
rect 1377 -150 1407 150
rect 1473 -150 1503 150
rect 1569 -150 1599 150
rect 1665 -150 1695 150
rect 1761 -150 1791 150
rect 1857 -150 1887 150
rect 1953 -150 1983 150
rect 2049 -150 2079 150
rect 2145 -150 2175 150
rect 2241 -150 2271 150
rect 2337 -150 2367 150
rect 2433 -150 2463 150
rect 2529 -150 2559 150
rect 2625 -150 2655 150
rect 2721 -150 2751 150
rect 2817 -150 2847 150
rect 2913 -150 2943 150
rect 3009 -150 3039 150
rect 3105 -150 3135 150
rect 3201 -150 3231 150
rect 3297 -150 3327 150
rect 3393 -150 3423 150
rect 3489 -150 3519 150
rect 3585 -150 3615 150
rect 3681 -150 3711 150
rect 3777 -150 3807 150
rect 3873 -150 3903 150
rect 3969 -150 3999 150
rect 4065 -150 4095 150
rect 4161 -150 4191 150
rect 4257 -150 4287 150
rect 4353 -150 4383 150
rect 4449 -150 4479 150
rect 4545 -150 4575 150
rect 4641 -150 4671 150
rect 4737 -150 4767 150
<< ndiff >>
rect -4829 138 -4767 150
rect -4829 -138 -4817 138
rect -4783 -138 -4767 138
rect -4829 -150 -4767 -138
rect -4737 138 -4671 150
rect -4737 -138 -4721 138
rect -4687 -138 -4671 138
rect -4737 -150 -4671 -138
rect -4641 138 -4575 150
rect -4641 -138 -4625 138
rect -4591 -138 -4575 138
rect -4641 -150 -4575 -138
rect -4545 138 -4479 150
rect -4545 -138 -4529 138
rect -4495 -138 -4479 138
rect -4545 -150 -4479 -138
rect -4449 138 -4383 150
rect -4449 -138 -4433 138
rect -4399 -138 -4383 138
rect -4449 -150 -4383 -138
rect -4353 138 -4287 150
rect -4353 -138 -4337 138
rect -4303 -138 -4287 138
rect -4353 -150 -4287 -138
rect -4257 138 -4191 150
rect -4257 -138 -4241 138
rect -4207 -138 -4191 138
rect -4257 -150 -4191 -138
rect -4161 138 -4095 150
rect -4161 -138 -4145 138
rect -4111 -138 -4095 138
rect -4161 -150 -4095 -138
rect -4065 138 -3999 150
rect -4065 -138 -4049 138
rect -4015 -138 -3999 138
rect -4065 -150 -3999 -138
rect -3969 138 -3903 150
rect -3969 -138 -3953 138
rect -3919 -138 -3903 138
rect -3969 -150 -3903 -138
rect -3873 138 -3807 150
rect -3873 -138 -3857 138
rect -3823 -138 -3807 138
rect -3873 -150 -3807 -138
rect -3777 138 -3711 150
rect -3777 -138 -3761 138
rect -3727 -138 -3711 138
rect -3777 -150 -3711 -138
rect -3681 138 -3615 150
rect -3681 -138 -3665 138
rect -3631 -138 -3615 138
rect -3681 -150 -3615 -138
rect -3585 138 -3519 150
rect -3585 -138 -3569 138
rect -3535 -138 -3519 138
rect -3585 -150 -3519 -138
rect -3489 138 -3423 150
rect -3489 -138 -3473 138
rect -3439 -138 -3423 138
rect -3489 -150 -3423 -138
rect -3393 138 -3327 150
rect -3393 -138 -3377 138
rect -3343 -138 -3327 138
rect -3393 -150 -3327 -138
rect -3297 138 -3231 150
rect -3297 -138 -3281 138
rect -3247 -138 -3231 138
rect -3297 -150 -3231 -138
rect -3201 138 -3135 150
rect -3201 -138 -3185 138
rect -3151 -138 -3135 138
rect -3201 -150 -3135 -138
rect -3105 138 -3039 150
rect -3105 -138 -3089 138
rect -3055 -138 -3039 138
rect -3105 -150 -3039 -138
rect -3009 138 -2943 150
rect -3009 -138 -2993 138
rect -2959 -138 -2943 138
rect -3009 -150 -2943 -138
rect -2913 138 -2847 150
rect -2913 -138 -2897 138
rect -2863 -138 -2847 138
rect -2913 -150 -2847 -138
rect -2817 138 -2751 150
rect -2817 -138 -2801 138
rect -2767 -138 -2751 138
rect -2817 -150 -2751 -138
rect -2721 138 -2655 150
rect -2721 -138 -2705 138
rect -2671 -138 -2655 138
rect -2721 -150 -2655 -138
rect -2625 138 -2559 150
rect -2625 -138 -2609 138
rect -2575 -138 -2559 138
rect -2625 -150 -2559 -138
rect -2529 138 -2463 150
rect -2529 -138 -2513 138
rect -2479 -138 -2463 138
rect -2529 -150 -2463 -138
rect -2433 138 -2367 150
rect -2433 -138 -2417 138
rect -2383 -138 -2367 138
rect -2433 -150 -2367 -138
rect -2337 138 -2271 150
rect -2337 -138 -2321 138
rect -2287 -138 -2271 138
rect -2337 -150 -2271 -138
rect -2241 138 -2175 150
rect -2241 -138 -2225 138
rect -2191 -138 -2175 138
rect -2241 -150 -2175 -138
rect -2145 138 -2079 150
rect -2145 -138 -2129 138
rect -2095 -138 -2079 138
rect -2145 -150 -2079 -138
rect -2049 138 -1983 150
rect -2049 -138 -2033 138
rect -1999 -138 -1983 138
rect -2049 -150 -1983 -138
rect -1953 138 -1887 150
rect -1953 -138 -1937 138
rect -1903 -138 -1887 138
rect -1953 -150 -1887 -138
rect -1857 138 -1791 150
rect -1857 -138 -1841 138
rect -1807 -138 -1791 138
rect -1857 -150 -1791 -138
rect -1761 138 -1695 150
rect -1761 -138 -1745 138
rect -1711 -138 -1695 138
rect -1761 -150 -1695 -138
rect -1665 138 -1599 150
rect -1665 -138 -1649 138
rect -1615 -138 -1599 138
rect -1665 -150 -1599 -138
rect -1569 138 -1503 150
rect -1569 -138 -1553 138
rect -1519 -138 -1503 138
rect -1569 -150 -1503 -138
rect -1473 138 -1407 150
rect -1473 -138 -1457 138
rect -1423 -138 -1407 138
rect -1473 -150 -1407 -138
rect -1377 138 -1311 150
rect -1377 -138 -1361 138
rect -1327 -138 -1311 138
rect -1377 -150 -1311 -138
rect -1281 138 -1215 150
rect -1281 -138 -1265 138
rect -1231 -138 -1215 138
rect -1281 -150 -1215 -138
rect -1185 138 -1119 150
rect -1185 -138 -1169 138
rect -1135 -138 -1119 138
rect -1185 -150 -1119 -138
rect -1089 138 -1023 150
rect -1089 -138 -1073 138
rect -1039 -138 -1023 138
rect -1089 -150 -1023 -138
rect -993 138 -927 150
rect -993 -138 -977 138
rect -943 -138 -927 138
rect -993 -150 -927 -138
rect -897 138 -831 150
rect -897 -138 -881 138
rect -847 -138 -831 138
rect -897 -150 -831 -138
rect -801 138 -735 150
rect -801 -138 -785 138
rect -751 -138 -735 138
rect -801 -150 -735 -138
rect -705 138 -639 150
rect -705 -138 -689 138
rect -655 -138 -639 138
rect -705 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 705 150
rect 639 -138 655 138
rect 689 -138 705 138
rect 639 -150 705 -138
rect 735 138 801 150
rect 735 -138 751 138
rect 785 -138 801 138
rect 735 -150 801 -138
rect 831 138 897 150
rect 831 -138 847 138
rect 881 -138 897 138
rect 831 -150 897 -138
rect 927 138 993 150
rect 927 -138 943 138
rect 977 -138 993 138
rect 927 -150 993 -138
rect 1023 138 1089 150
rect 1023 -138 1039 138
rect 1073 -138 1089 138
rect 1023 -150 1089 -138
rect 1119 138 1185 150
rect 1119 -138 1135 138
rect 1169 -138 1185 138
rect 1119 -150 1185 -138
rect 1215 138 1281 150
rect 1215 -138 1231 138
rect 1265 -138 1281 138
rect 1215 -150 1281 -138
rect 1311 138 1377 150
rect 1311 -138 1327 138
rect 1361 -138 1377 138
rect 1311 -150 1377 -138
rect 1407 138 1473 150
rect 1407 -138 1423 138
rect 1457 -138 1473 138
rect 1407 -150 1473 -138
rect 1503 138 1569 150
rect 1503 -138 1519 138
rect 1553 -138 1569 138
rect 1503 -150 1569 -138
rect 1599 138 1665 150
rect 1599 -138 1615 138
rect 1649 -138 1665 138
rect 1599 -150 1665 -138
rect 1695 138 1761 150
rect 1695 -138 1711 138
rect 1745 -138 1761 138
rect 1695 -150 1761 -138
rect 1791 138 1857 150
rect 1791 -138 1807 138
rect 1841 -138 1857 138
rect 1791 -150 1857 -138
rect 1887 138 1953 150
rect 1887 -138 1903 138
rect 1937 -138 1953 138
rect 1887 -150 1953 -138
rect 1983 138 2049 150
rect 1983 -138 1999 138
rect 2033 -138 2049 138
rect 1983 -150 2049 -138
rect 2079 138 2145 150
rect 2079 -138 2095 138
rect 2129 -138 2145 138
rect 2079 -150 2145 -138
rect 2175 138 2241 150
rect 2175 -138 2191 138
rect 2225 -138 2241 138
rect 2175 -150 2241 -138
rect 2271 138 2337 150
rect 2271 -138 2287 138
rect 2321 -138 2337 138
rect 2271 -150 2337 -138
rect 2367 138 2433 150
rect 2367 -138 2383 138
rect 2417 -138 2433 138
rect 2367 -150 2433 -138
rect 2463 138 2529 150
rect 2463 -138 2479 138
rect 2513 -138 2529 138
rect 2463 -150 2529 -138
rect 2559 138 2625 150
rect 2559 -138 2575 138
rect 2609 -138 2625 138
rect 2559 -150 2625 -138
rect 2655 138 2721 150
rect 2655 -138 2671 138
rect 2705 -138 2721 138
rect 2655 -150 2721 -138
rect 2751 138 2817 150
rect 2751 -138 2767 138
rect 2801 -138 2817 138
rect 2751 -150 2817 -138
rect 2847 138 2913 150
rect 2847 -138 2863 138
rect 2897 -138 2913 138
rect 2847 -150 2913 -138
rect 2943 138 3009 150
rect 2943 -138 2959 138
rect 2993 -138 3009 138
rect 2943 -150 3009 -138
rect 3039 138 3105 150
rect 3039 -138 3055 138
rect 3089 -138 3105 138
rect 3039 -150 3105 -138
rect 3135 138 3201 150
rect 3135 -138 3151 138
rect 3185 -138 3201 138
rect 3135 -150 3201 -138
rect 3231 138 3297 150
rect 3231 -138 3247 138
rect 3281 -138 3297 138
rect 3231 -150 3297 -138
rect 3327 138 3393 150
rect 3327 -138 3343 138
rect 3377 -138 3393 138
rect 3327 -150 3393 -138
rect 3423 138 3489 150
rect 3423 -138 3439 138
rect 3473 -138 3489 138
rect 3423 -150 3489 -138
rect 3519 138 3585 150
rect 3519 -138 3535 138
rect 3569 -138 3585 138
rect 3519 -150 3585 -138
rect 3615 138 3681 150
rect 3615 -138 3631 138
rect 3665 -138 3681 138
rect 3615 -150 3681 -138
rect 3711 138 3777 150
rect 3711 -138 3727 138
rect 3761 -138 3777 138
rect 3711 -150 3777 -138
rect 3807 138 3873 150
rect 3807 -138 3823 138
rect 3857 -138 3873 138
rect 3807 -150 3873 -138
rect 3903 138 3969 150
rect 3903 -138 3919 138
rect 3953 -138 3969 138
rect 3903 -150 3969 -138
rect 3999 138 4065 150
rect 3999 -138 4015 138
rect 4049 -138 4065 138
rect 3999 -150 4065 -138
rect 4095 138 4161 150
rect 4095 -138 4111 138
rect 4145 -138 4161 138
rect 4095 -150 4161 -138
rect 4191 138 4257 150
rect 4191 -138 4207 138
rect 4241 -138 4257 138
rect 4191 -150 4257 -138
rect 4287 138 4353 150
rect 4287 -138 4303 138
rect 4337 -138 4353 138
rect 4287 -150 4353 -138
rect 4383 138 4449 150
rect 4383 -138 4399 138
rect 4433 -138 4449 138
rect 4383 -150 4449 -138
rect 4479 138 4545 150
rect 4479 -138 4495 138
rect 4529 -138 4545 138
rect 4479 -150 4545 -138
rect 4575 138 4641 150
rect 4575 -138 4591 138
rect 4625 -138 4641 138
rect 4575 -150 4641 -138
rect 4671 138 4737 150
rect 4671 -138 4687 138
rect 4721 -138 4737 138
rect 4671 -150 4737 -138
rect 4767 138 4829 150
rect 4767 -138 4783 138
rect 4817 -138 4829 138
rect 4767 -150 4829 -138
<< ndiffc >>
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
<< psubdiff >>
rect -4931 290 -4835 324
rect 4835 290 4931 324
rect -4931 228 -4897 290
rect 4897 228 4931 290
rect -4931 -290 -4897 -228
rect 4897 -290 4931 -228
rect -4931 -324 -4835 -290
rect 4835 -324 4931 -290
<< psubdiffcont >>
rect -4835 290 4835 324
rect -4931 -228 -4897 228
rect 4897 -228 4931 228
rect -4835 -324 4835 -290
<< poly >>
rect -4767 232 4767 242
rect -4767 191 -4721 232
rect 4719 191 4767 232
rect -4767 176 4767 191
rect -4767 150 -4737 176
rect -4671 150 -4641 176
rect -4575 150 -4545 176
rect -4479 150 -4449 176
rect -4383 150 -4353 176
rect -4287 150 -4257 176
rect -4191 150 -4161 176
rect -4095 150 -4065 176
rect -3999 150 -3969 176
rect -3903 150 -3873 176
rect -3807 150 -3777 176
rect -3711 150 -3681 176
rect -3615 150 -3585 176
rect -3519 150 -3489 176
rect -3423 150 -3393 176
rect -3327 150 -3297 176
rect -3231 150 -3201 176
rect -3135 150 -3105 176
rect -3039 150 -3009 176
rect -2943 150 -2913 176
rect -2847 150 -2817 176
rect -2751 150 -2721 176
rect -2655 150 -2625 176
rect -2559 150 -2529 176
rect -2463 150 -2433 176
rect -2367 150 -2337 176
rect -2271 150 -2241 176
rect -2175 150 -2145 176
rect -2079 150 -2049 176
rect -1983 150 -1953 176
rect -1887 150 -1857 176
rect -1791 150 -1761 176
rect -1695 150 -1665 176
rect -1599 150 -1569 176
rect -1503 150 -1473 176
rect -1407 150 -1377 176
rect -1311 150 -1281 176
rect -1215 150 -1185 176
rect -1119 150 -1089 176
rect -1023 150 -993 176
rect -927 150 -897 176
rect -831 150 -801 176
rect -735 150 -705 176
rect -639 150 -609 176
rect -543 150 -513 176
rect -447 150 -417 176
rect -351 150 -321 176
rect -255 150 -225 176
rect -159 150 -129 176
rect -63 150 -33 176
rect 33 150 63 176
rect 129 150 159 176
rect 225 150 255 176
rect 321 150 351 176
rect 417 150 447 176
rect 513 150 543 176
rect 609 150 639 176
rect 705 150 735 176
rect 801 150 831 176
rect 897 150 927 176
rect 993 150 1023 176
rect 1089 150 1119 176
rect 1185 150 1215 176
rect 1281 150 1311 176
rect 1377 150 1407 176
rect 1473 150 1503 176
rect 1569 150 1599 176
rect 1665 150 1695 176
rect 1761 150 1791 176
rect 1857 150 1887 176
rect 1953 150 1983 176
rect 2049 150 2079 176
rect 2145 150 2175 176
rect 2241 150 2271 176
rect 2337 150 2367 176
rect 2433 150 2463 176
rect 2529 150 2559 176
rect 2625 150 2655 176
rect 2721 150 2751 176
rect 2817 150 2847 176
rect 2913 150 2943 176
rect 3009 150 3039 176
rect 3105 150 3135 176
rect 3201 150 3231 176
rect 3297 150 3327 176
rect 3393 150 3423 176
rect 3489 150 3519 176
rect 3585 150 3615 176
rect 3681 150 3711 176
rect 3777 150 3807 176
rect 3873 150 3903 176
rect 3969 150 3999 176
rect 4065 150 4095 176
rect 4161 150 4191 176
rect 4257 150 4287 176
rect 4353 150 4383 176
rect 4449 150 4479 176
rect 4545 150 4575 176
rect 4641 150 4671 176
rect 4737 150 4767 176
rect -4767 -176 -4737 -150
rect -4671 -176 -4641 -150
rect -4575 -176 -4545 -150
rect -4479 -176 -4449 -150
rect -4383 -176 -4353 -150
rect -4287 -176 -4257 -150
rect -4191 -176 -4161 -150
rect -4095 -176 -4065 -150
rect -3999 -176 -3969 -150
rect -3903 -176 -3873 -150
rect -3807 -176 -3777 -150
rect -3711 -176 -3681 -150
rect -3615 -176 -3585 -150
rect -3519 -176 -3489 -150
rect -3423 -176 -3393 -150
rect -3327 -176 -3297 -150
rect -3231 -176 -3201 -150
rect -3135 -176 -3105 -150
rect -3039 -176 -3009 -150
rect -2943 -176 -2913 -150
rect -2847 -176 -2817 -150
rect -2751 -176 -2721 -150
rect -2655 -176 -2625 -150
rect -2559 -176 -2529 -150
rect -2463 -176 -2433 -150
rect -2367 -176 -2337 -150
rect -2271 -176 -2241 -150
rect -2175 -176 -2145 -150
rect -2079 -176 -2049 -150
rect -1983 -176 -1953 -150
rect -1887 -176 -1857 -150
rect -1791 -176 -1761 -150
rect -1695 -176 -1665 -150
rect -1599 -176 -1569 -150
rect -1503 -176 -1473 -150
rect -1407 -176 -1377 -150
rect -1311 -176 -1281 -150
rect -1215 -176 -1185 -150
rect -1119 -176 -1089 -150
rect -1023 -176 -993 -150
rect -927 -176 -897 -150
rect -831 -176 -801 -150
rect -735 -176 -705 -150
rect -639 -176 -609 -150
rect -543 -176 -513 -150
rect -447 -176 -417 -150
rect -351 -176 -321 -150
rect -255 -176 -225 -150
rect -159 -176 -129 -150
rect -63 -176 -33 -150
rect 33 -176 63 -150
rect 129 -176 159 -150
rect 225 -176 255 -150
rect 321 -176 351 -150
rect 417 -176 447 -150
rect 513 -176 543 -150
rect 609 -176 639 -150
rect 705 -176 735 -150
rect 801 -176 831 -150
rect 897 -176 927 -150
rect 993 -176 1023 -150
rect 1089 -176 1119 -150
rect 1185 -176 1215 -150
rect 1281 -176 1311 -150
rect 1377 -176 1407 -150
rect 1473 -176 1503 -150
rect 1569 -176 1599 -150
rect 1665 -176 1695 -150
rect 1761 -176 1791 -150
rect 1857 -176 1887 -150
rect 1953 -176 1983 -150
rect 2049 -176 2079 -150
rect 2145 -176 2175 -150
rect 2241 -176 2271 -150
rect 2337 -176 2367 -150
rect 2433 -176 2463 -150
rect 2529 -176 2559 -150
rect 2625 -176 2655 -150
rect 2721 -176 2751 -150
rect 2817 -176 2847 -150
rect 2913 -176 2943 -150
rect 3009 -176 3039 -150
rect 3105 -176 3135 -150
rect 3201 -176 3231 -150
rect 3297 -176 3327 -150
rect 3393 -176 3423 -150
rect 3489 -176 3519 -150
rect 3585 -176 3615 -150
rect 3681 -176 3711 -150
rect 3777 -176 3807 -150
rect 3873 -176 3903 -150
rect 3969 -176 3999 -150
rect 4065 -176 4095 -150
rect 4161 -176 4191 -150
rect 4257 -176 4287 -150
rect 4353 -176 4383 -150
rect 4449 -176 4479 -150
rect 4545 -176 4575 -150
rect 4641 -176 4671 -150
rect 4737 -176 4767 -150
<< polycont >>
rect -4721 191 4719 232
<< locali >>
rect -4931 290 -4835 324
rect 4835 290 4931 324
rect -4931 228 -4897 290
rect 4897 228 4931 290
rect -4817 138 -4783 154
rect -4817 -154 -4783 -138
rect -4721 138 -4687 154
rect -4721 -154 -4687 -138
rect -4625 138 -4591 154
rect -4625 -154 -4591 -138
rect -4529 138 -4495 154
rect -4529 -154 -4495 -138
rect -4433 138 -4399 154
rect -4433 -154 -4399 -138
rect -4337 138 -4303 154
rect -4337 -154 -4303 -138
rect -4241 138 -4207 154
rect -4241 -154 -4207 -138
rect -4145 138 -4111 154
rect -4145 -154 -4111 -138
rect -4049 138 -4015 154
rect -4049 -154 -4015 -138
rect -3953 138 -3919 154
rect -3953 -154 -3919 -138
rect -3857 138 -3823 154
rect -3857 -154 -3823 -138
rect -3761 138 -3727 154
rect -3761 -154 -3727 -138
rect -3665 138 -3631 154
rect -3665 -154 -3631 -138
rect -3569 138 -3535 154
rect -3569 -154 -3535 -138
rect -3473 138 -3439 154
rect -3473 -154 -3439 -138
rect -3377 138 -3343 154
rect -3377 -154 -3343 -138
rect -3281 138 -3247 154
rect -3281 -154 -3247 -138
rect -3185 138 -3151 154
rect -3185 -154 -3151 -138
rect -3089 138 -3055 154
rect -3089 -154 -3055 -138
rect -2993 138 -2959 154
rect -2993 -154 -2959 -138
rect -2897 138 -2863 154
rect -2897 -154 -2863 -138
rect -2801 138 -2767 154
rect -2801 -154 -2767 -138
rect -2705 138 -2671 154
rect -2705 -154 -2671 -138
rect -2609 138 -2575 154
rect -2609 -154 -2575 -138
rect -2513 138 -2479 154
rect -2513 -154 -2479 -138
rect -2417 138 -2383 154
rect -2417 -154 -2383 -138
rect -2321 138 -2287 154
rect -2321 -154 -2287 -138
rect -2225 138 -2191 154
rect -2225 -154 -2191 -138
rect -2129 138 -2095 154
rect -2129 -154 -2095 -138
rect -2033 138 -1999 154
rect -2033 -154 -1999 -138
rect -1937 138 -1903 154
rect -1937 -154 -1903 -138
rect -1841 138 -1807 154
rect -1841 -154 -1807 -138
rect -1745 138 -1711 154
rect -1745 -154 -1711 -138
rect -1649 138 -1615 154
rect -1649 -154 -1615 -138
rect -1553 138 -1519 154
rect -1553 -154 -1519 -138
rect -1457 138 -1423 154
rect -1457 -154 -1423 -138
rect -1361 138 -1327 154
rect -1361 -154 -1327 -138
rect -1265 138 -1231 154
rect -1265 -154 -1231 -138
rect -1169 138 -1135 154
rect -1169 -154 -1135 -138
rect -1073 138 -1039 154
rect -1073 -154 -1039 -138
rect -977 138 -943 154
rect -977 -154 -943 -138
rect -881 138 -847 154
rect -881 -154 -847 -138
rect -785 138 -751 154
rect -785 -154 -751 -138
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect 751 138 785 154
rect 751 -154 785 -138
rect 847 138 881 154
rect 847 -154 881 -138
rect 943 138 977 154
rect 943 -154 977 -138
rect 1039 138 1073 154
rect 1039 -154 1073 -138
rect 1135 138 1169 154
rect 1135 -154 1169 -138
rect 1231 138 1265 154
rect 1231 -154 1265 -138
rect 1327 138 1361 154
rect 1327 -154 1361 -138
rect 1423 138 1457 154
rect 1423 -154 1457 -138
rect 1519 138 1553 154
rect 1519 -154 1553 -138
rect 1615 138 1649 154
rect 1615 -154 1649 -138
rect 1711 138 1745 154
rect 1711 -154 1745 -138
rect 1807 138 1841 154
rect 1807 -154 1841 -138
rect 1903 138 1937 154
rect 1903 -154 1937 -138
rect 1999 138 2033 154
rect 1999 -154 2033 -138
rect 2095 138 2129 154
rect 2095 -154 2129 -138
rect 2191 138 2225 154
rect 2191 -154 2225 -138
rect 2287 138 2321 154
rect 2287 -154 2321 -138
rect 2383 138 2417 154
rect 2383 -154 2417 -138
rect 2479 138 2513 154
rect 2479 -154 2513 -138
rect 2575 138 2609 154
rect 2575 -154 2609 -138
rect 2671 138 2705 154
rect 2671 -154 2705 -138
rect 2767 138 2801 154
rect 2767 -154 2801 -138
rect 2863 138 2897 154
rect 2863 -154 2897 -138
rect 2959 138 2993 154
rect 2959 -154 2993 -138
rect 3055 138 3089 154
rect 3055 -154 3089 -138
rect 3151 138 3185 154
rect 3151 -154 3185 -138
rect 3247 138 3281 154
rect 3247 -154 3281 -138
rect 3343 138 3377 154
rect 3343 -154 3377 -138
rect 3439 138 3473 154
rect 3439 -154 3473 -138
rect 3535 138 3569 154
rect 3535 -154 3569 -138
rect 3631 138 3665 154
rect 3631 -154 3665 -138
rect 3727 138 3761 154
rect 3727 -154 3761 -138
rect 3823 138 3857 154
rect 3823 -154 3857 -138
rect 3919 138 3953 154
rect 3919 -154 3953 -138
rect 4015 138 4049 154
rect 4015 -154 4049 -138
rect 4111 138 4145 154
rect 4111 -154 4145 -138
rect 4207 138 4241 154
rect 4207 -154 4241 -138
rect 4303 138 4337 154
rect 4303 -154 4337 -138
rect 4399 138 4433 154
rect 4399 -154 4433 -138
rect 4495 138 4529 154
rect 4495 -154 4529 -138
rect 4591 138 4625 154
rect 4591 -154 4625 -138
rect 4687 138 4721 154
rect 4687 -154 4721 -138
rect 4783 138 4817 154
rect 4783 -154 4817 -138
rect -4931 -290 -4897 -228
rect 4897 -290 4931 -228
rect -4931 -324 -4835 -290
rect 4835 -324 4931 -290
<< viali >>
rect -4737 191 -4721 232
rect -4721 191 4719 232
rect 4719 191 4738 232
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
rect -4835 -324 4835 -290
<< metal1 >>
rect -4749 232 4750 238
rect -4749 191 -4737 232
rect 4738 191 4750 232
rect -4749 185 4750 191
rect -4842 -153 -4832 155
rect -4768 -153 -4758 155
rect -4727 138 -4681 150
rect -4727 -138 -4721 138
rect -4687 -138 -4681 138
rect -4727 -201 -4681 -138
rect -4650 -154 -4640 154
rect -4576 -154 -4566 154
rect -4535 138 -4489 150
rect -4535 -138 -4529 138
rect -4495 -138 -4489 138
rect -4535 -201 -4489 -138
rect -4458 -154 -4448 154
rect -4384 -154 -4374 154
rect -4343 138 -4297 150
rect -4343 -138 -4337 138
rect -4303 -138 -4297 138
rect -4343 -201 -4297 -138
rect -4266 -154 -4256 154
rect -4192 -154 -4182 154
rect -4151 138 -4105 150
rect -4151 -138 -4145 138
rect -4111 -138 -4105 138
rect -4151 -201 -4105 -138
rect -4074 -154 -4064 154
rect -4000 -154 -3990 154
rect -3959 138 -3913 150
rect -3959 -138 -3953 138
rect -3919 -138 -3913 138
rect -3959 -201 -3913 -138
rect -3882 -154 -3872 154
rect -3808 -154 -3798 154
rect -3767 138 -3721 150
rect -3767 -138 -3761 138
rect -3727 -138 -3721 138
rect -3767 -201 -3721 -138
rect -3690 -154 -3680 154
rect -3616 -154 -3606 154
rect -3575 138 -3529 150
rect -3575 -138 -3569 138
rect -3535 -138 -3529 138
rect -3575 -201 -3529 -138
rect -3498 -154 -3488 154
rect -3424 -154 -3414 154
rect -3383 138 -3337 150
rect -3383 -138 -3377 138
rect -3343 -138 -3337 138
rect -3383 -201 -3337 -138
rect -3306 -154 -3296 154
rect -3232 -154 -3222 154
rect -3191 138 -3145 150
rect -3191 -138 -3185 138
rect -3151 -138 -3145 138
rect -3191 -201 -3145 -138
rect -3114 -154 -3104 154
rect -3040 -154 -3030 154
rect -2999 138 -2953 150
rect -2999 -138 -2993 138
rect -2959 -138 -2953 138
rect -2999 -201 -2953 -138
rect -2922 -154 -2912 154
rect -2848 -154 -2838 154
rect -2807 138 -2761 150
rect -2807 -138 -2801 138
rect -2767 -138 -2761 138
rect -2807 -201 -2761 -138
rect -2730 -154 -2720 154
rect -2656 -154 -2646 154
rect -2615 138 -2569 150
rect -2615 -138 -2609 138
rect -2575 -138 -2569 138
rect -2615 -201 -2569 -138
rect -2538 -154 -2528 154
rect -2464 -154 -2454 154
rect -2423 138 -2377 150
rect -2423 -138 -2417 138
rect -2383 -138 -2377 138
rect -2423 -201 -2377 -138
rect -2346 -154 -2336 154
rect -2272 -154 -2262 154
rect -2231 138 -2185 150
rect -2231 -138 -2225 138
rect -2191 -138 -2185 138
rect -2231 -201 -2185 -138
rect -2154 -154 -2144 154
rect -2080 -154 -2070 154
rect -2039 138 -1993 150
rect -2039 -138 -2033 138
rect -1999 -138 -1993 138
rect -2039 -201 -1993 -138
rect -1962 -154 -1952 154
rect -1888 -154 -1878 154
rect -1847 138 -1801 150
rect -1847 -138 -1841 138
rect -1807 -138 -1801 138
rect -1847 -201 -1801 -138
rect -1770 -154 -1760 154
rect -1696 -154 -1686 154
rect -1655 138 -1609 150
rect -1655 -138 -1649 138
rect -1615 -138 -1609 138
rect -1655 -201 -1609 -138
rect -1578 -154 -1568 154
rect -1504 -154 -1494 154
rect -1463 138 -1417 150
rect -1463 -138 -1457 138
rect -1423 -138 -1417 138
rect -1463 -201 -1417 -138
rect -1386 -154 -1376 154
rect -1312 -154 -1302 154
rect -1271 138 -1225 150
rect -1271 -138 -1265 138
rect -1231 -138 -1225 138
rect -1271 -201 -1225 -138
rect -1194 -154 -1184 154
rect -1120 -154 -1110 154
rect -1079 138 -1033 150
rect -1079 -138 -1073 138
rect -1039 -138 -1033 138
rect -1079 -201 -1033 -138
rect -1002 -154 -992 154
rect -928 -154 -918 154
rect -887 138 -841 150
rect -887 -138 -881 138
rect -847 -138 -841 138
rect -887 -201 -841 -138
rect -810 -154 -800 154
rect -736 -154 -726 154
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -201 -649 -138
rect -618 -154 -608 154
rect -544 -154 -534 154
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -201 -457 -138
rect -426 -154 -416 154
rect -352 -154 -342 154
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -201 -265 -138
rect -234 -154 -224 154
rect -160 -154 -150 154
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -201 -73 -138
rect -42 -154 -32 154
rect 32 -154 42 154
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -201 119 -138
rect 150 -154 160 154
rect 224 -154 234 154
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -201 311 -138
rect 342 -154 352 154
rect 416 -154 426 154
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -201 503 -138
rect 534 -154 544 154
rect 608 -154 618 154
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -201 695 -138
rect 726 -154 736 154
rect 800 -154 810 154
rect 841 138 887 150
rect 841 -138 847 138
rect 881 -138 887 138
rect 841 -201 887 -138
rect 918 -154 928 154
rect 992 -154 1002 154
rect 1033 138 1079 150
rect 1033 -138 1039 138
rect 1073 -138 1079 138
rect 1033 -201 1079 -138
rect 1110 -154 1120 154
rect 1184 -154 1194 154
rect 1225 138 1271 150
rect 1225 -138 1231 138
rect 1265 -138 1271 138
rect 1225 -201 1271 -138
rect 1302 -154 1312 154
rect 1376 -154 1386 154
rect 1417 138 1463 150
rect 1417 -138 1423 138
rect 1457 -138 1463 138
rect 1417 -201 1463 -138
rect 1494 -154 1504 154
rect 1568 -154 1578 154
rect 1609 138 1655 150
rect 1609 -138 1615 138
rect 1649 -138 1655 138
rect 1609 -201 1655 -138
rect 1686 -154 1696 154
rect 1760 -154 1770 154
rect 1801 138 1847 150
rect 1801 -138 1807 138
rect 1841 -138 1847 138
rect 1801 -201 1847 -138
rect 1878 -154 1888 154
rect 1952 -154 1962 154
rect 1993 138 2039 150
rect 1993 -138 1999 138
rect 2033 -138 2039 138
rect 1993 -201 2039 -138
rect 2070 -154 2080 154
rect 2144 -154 2154 154
rect 2185 138 2231 150
rect 2185 -138 2191 138
rect 2225 -138 2231 138
rect 2185 -201 2231 -138
rect 2262 -154 2272 154
rect 2336 -154 2346 154
rect 2377 138 2423 150
rect 2377 -138 2383 138
rect 2417 -138 2423 138
rect 2377 -201 2423 -138
rect 2454 -154 2464 154
rect 2528 -154 2538 154
rect 2569 138 2615 150
rect 2569 -138 2575 138
rect 2609 -138 2615 138
rect 2569 -201 2615 -138
rect 2646 -154 2656 154
rect 2720 -154 2730 154
rect 2761 138 2807 150
rect 2761 -138 2767 138
rect 2801 -138 2807 138
rect 2761 -201 2807 -138
rect 2838 -154 2848 154
rect 2912 -154 2922 154
rect 2953 138 2999 150
rect 2953 -138 2959 138
rect 2993 -138 2999 138
rect 2953 -201 2999 -138
rect 3030 -154 3040 154
rect 3104 -154 3114 154
rect 3145 138 3191 150
rect 3145 -138 3151 138
rect 3185 -138 3191 138
rect 3145 -201 3191 -138
rect 3222 -154 3232 154
rect 3296 -154 3306 154
rect 3337 138 3383 150
rect 3337 -138 3343 138
rect 3377 -138 3383 138
rect 3337 -201 3383 -138
rect 3414 -154 3424 154
rect 3488 -154 3498 154
rect 3529 138 3575 150
rect 3529 -138 3535 138
rect 3569 -138 3575 138
rect 3529 -201 3575 -138
rect 3606 -154 3616 154
rect 3680 -154 3690 154
rect 3721 138 3767 150
rect 3721 -138 3727 138
rect 3761 -138 3767 138
rect 3721 -201 3767 -138
rect 3798 -154 3808 154
rect 3872 -154 3882 154
rect 3913 138 3959 150
rect 3913 -138 3919 138
rect 3953 -138 3959 138
rect 3913 -201 3959 -138
rect 3990 -154 4000 154
rect 4064 -154 4074 154
rect 4105 138 4151 150
rect 4105 -138 4111 138
rect 4145 -138 4151 138
rect 4105 -201 4151 -138
rect 4182 -154 4192 154
rect 4256 -154 4266 154
rect 4297 138 4343 150
rect 4297 -138 4303 138
rect 4337 -138 4343 138
rect 4297 -201 4343 -138
rect 4374 -154 4384 154
rect 4448 -154 4458 154
rect 4489 138 4535 150
rect 4489 -138 4495 138
rect 4529 -138 4535 138
rect 4489 -201 4535 -138
rect 4566 -154 4576 154
rect 4640 -154 4650 154
rect 4681 138 4727 150
rect 4681 -138 4687 138
rect 4721 -138 4727 138
rect 4681 -201 4727 -138
rect 4758 -154 4768 154
rect 4832 -154 4842 154
rect -4847 -290 4847 -201
rect -4847 -324 -4835 -290
rect 4835 -324 4847 -290
rect -4847 -330 4847 -324
<< via1 >>
rect -4832 138 -4768 155
rect -4832 -138 -4817 138
rect -4817 -138 -4783 138
rect -4783 -138 -4768 138
rect -4832 -153 -4768 -138
rect -4640 138 -4576 154
rect -4640 -138 -4625 138
rect -4625 -138 -4591 138
rect -4591 -138 -4576 138
rect -4640 -154 -4576 -138
rect -4448 138 -4384 154
rect -4448 -138 -4433 138
rect -4433 -138 -4399 138
rect -4399 -138 -4384 138
rect -4448 -154 -4384 -138
rect -4256 138 -4192 154
rect -4256 -138 -4241 138
rect -4241 -138 -4207 138
rect -4207 -138 -4192 138
rect -4256 -154 -4192 -138
rect -4064 138 -4000 154
rect -4064 -138 -4049 138
rect -4049 -138 -4015 138
rect -4015 -138 -4000 138
rect -4064 -154 -4000 -138
rect -3872 138 -3808 154
rect -3872 -138 -3857 138
rect -3857 -138 -3823 138
rect -3823 -138 -3808 138
rect -3872 -154 -3808 -138
rect -3680 138 -3616 154
rect -3680 -138 -3665 138
rect -3665 -138 -3631 138
rect -3631 -138 -3616 138
rect -3680 -154 -3616 -138
rect -3488 138 -3424 154
rect -3488 -138 -3473 138
rect -3473 -138 -3439 138
rect -3439 -138 -3424 138
rect -3488 -154 -3424 -138
rect -3296 138 -3232 154
rect -3296 -138 -3281 138
rect -3281 -138 -3247 138
rect -3247 -138 -3232 138
rect -3296 -154 -3232 -138
rect -3104 138 -3040 154
rect -3104 -138 -3089 138
rect -3089 -138 -3055 138
rect -3055 -138 -3040 138
rect -3104 -154 -3040 -138
rect -2912 138 -2848 154
rect -2912 -138 -2897 138
rect -2897 -138 -2863 138
rect -2863 -138 -2848 138
rect -2912 -154 -2848 -138
rect -2720 138 -2656 154
rect -2720 -138 -2705 138
rect -2705 -138 -2671 138
rect -2671 -138 -2656 138
rect -2720 -154 -2656 -138
rect -2528 138 -2464 154
rect -2528 -138 -2513 138
rect -2513 -138 -2479 138
rect -2479 -138 -2464 138
rect -2528 -154 -2464 -138
rect -2336 138 -2272 154
rect -2336 -138 -2321 138
rect -2321 -138 -2287 138
rect -2287 -138 -2272 138
rect -2336 -154 -2272 -138
rect -2144 138 -2080 154
rect -2144 -138 -2129 138
rect -2129 -138 -2095 138
rect -2095 -138 -2080 138
rect -2144 -154 -2080 -138
rect -1952 138 -1888 154
rect -1952 -138 -1937 138
rect -1937 -138 -1903 138
rect -1903 -138 -1888 138
rect -1952 -154 -1888 -138
rect -1760 138 -1696 154
rect -1760 -138 -1745 138
rect -1745 -138 -1711 138
rect -1711 -138 -1696 138
rect -1760 -154 -1696 -138
rect -1568 138 -1504 154
rect -1568 -138 -1553 138
rect -1553 -138 -1519 138
rect -1519 -138 -1504 138
rect -1568 -154 -1504 -138
rect -1376 138 -1312 154
rect -1376 -138 -1361 138
rect -1361 -138 -1327 138
rect -1327 -138 -1312 138
rect -1376 -154 -1312 -138
rect -1184 138 -1120 154
rect -1184 -138 -1169 138
rect -1169 -138 -1135 138
rect -1135 -138 -1120 138
rect -1184 -154 -1120 -138
rect -992 138 -928 154
rect -992 -138 -977 138
rect -977 -138 -943 138
rect -943 -138 -928 138
rect -992 -154 -928 -138
rect -800 138 -736 154
rect -800 -138 -785 138
rect -785 -138 -751 138
rect -751 -138 -736 138
rect -800 -154 -736 -138
rect -608 138 -544 154
rect -608 -138 -593 138
rect -593 -138 -559 138
rect -559 -138 -544 138
rect -608 -154 -544 -138
rect -416 138 -352 154
rect -416 -138 -401 138
rect -401 -138 -367 138
rect -367 -138 -352 138
rect -416 -154 -352 -138
rect -224 138 -160 154
rect -224 -138 -209 138
rect -209 -138 -175 138
rect -175 -138 -160 138
rect -224 -154 -160 -138
rect -32 138 32 154
rect -32 -138 -17 138
rect -17 -138 17 138
rect 17 -138 32 138
rect -32 -154 32 -138
rect 160 138 224 154
rect 160 -138 175 138
rect 175 -138 209 138
rect 209 -138 224 138
rect 160 -154 224 -138
rect 352 138 416 154
rect 352 -138 367 138
rect 367 -138 401 138
rect 401 -138 416 138
rect 352 -154 416 -138
rect 544 138 608 154
rect 544 -138 559 138
rect 559 -138 593 138
rect 593 -138 608 138
rect 544 -154 608 -138
rect 736 138 800 154
rect 736 -138 751 138
rect 751 -138 785 138
rect 785 -138 800 138
rect 736 -154 800 -138
rect 928 138 992 154
rect 928 -138 943 138
rect 943 -138 977 138
rect 977 -138 992 138
rect 928 -154 992 -138
rect 1120 138 1184 154
rect 1120 -138 1135 138
rect 1135 -138 1169 138
rect 1169 -138 1184 138
rect 1120 -154 1184 -138
rect 1312 138 1376 154
rect 1312 -138 1327 138
rect 1327 -138 1361 138
rect 1361 -138 1376 138
rect 1312 -154 1376 -138
rect 1504 138 1568 154
rect 1504 -138 1519 138
rect 1519 -138 1553 138
rect 1553 -138 1568 138
rect 1504 -154 1568 -138
rect 1696 138 1760 154
rect 1696 -138 1711 138
rect 1711 -138 1745 138
rect 1745 -138 1760 138
rect 1696 -154 1760 -138
rect 1888 138 1952 154
rect 1888 -138 1903 138
rect 1903 -138 1937 138
rect 1937 -138 1952 138
rect 1888 -154 1952 -138
rect 2080 138 2144 154
rect 2080 -138 2095 138
rect 2095 -138 2129 138
rect 2129 -138 2144 138
rect 2080 -154 2144 -138
rect 2272 138 2336 154
rect 2272 -138 2287 138
rect 2287 -138 2321 138
rect 2321 -138 2336 138
rect 2272 -154 2336 -138
rect 2464 138 2528 154
rect 2464 -138 2479 138
rect 2479 -138 2513 138
rect 2513 -138 2528 138
rect 2464 -154 2528 -138
rect 2656 138 2720 154
rect 2656 -138 2671 138
rect 2671 -138 2705 138
rect 2705 -138 2720 138
rect 2656 -154 2720 -138
rect 2848 138 2912 154
rect 2848 -138 2863 138
rect 2863 -138 2897 138
rect 2897 -138 2912 138
rect 2848 -154 2912 -138
rect 3040 138 3104 154
rect 3040 -138 3055 138
rect 3055 -138 3089 138
rect 3089 -138 3104 138
rect 3040 -154 3104 -138
rect 3232 138 3296 154
rect 3232 -138 3247 138
rect 3247 -138 3281 138
rect 3281 -138 3296 138
rect 3232 -154 3296 -138
rect 3424 138 3488 154
rect 3424 -138 3439 138
rect 3439 -138 3473 138
rect 3473 -138 3488 138
rect 3424 -154 3488 -138
rect 3616 138 3680 154
rect 3616 -138 3631 138
rect 3631 -138 3665 138
rect 3665 -138 3680 138
rect 3616 -154 3680 -138
rect 3808 138 3872 154
rect 3808 -138 3823 138
rect 3823 -138 3857 138
rect 3857 -138 3872 138
rect 3808 -154 3872 -138
rect 4000 138 4064 154
rect 4000 -138 4015 138
rect 4015 -138 4049 138
rect 4049 -138 4064 138
rect 4000 -154 4064 -138
rect 4192 138 4256 154
rect 4192 -138 4207 138
rect 4207 -138 4241 138
rect 4241 -138 4256 138
rect 4192 -154 4256 -138
rect 4384 138 4448 154
rect 4384 -138 4399 138
rect 4399 -138 4433 138
rect 4433 -138 4448 138
rect 4384 -154 4448 -138
rect 4576 138 4640 154
rect 4576 -138 4591 138
rect 4591 -138 4625 138
rect 4625 -138 4640 138
rect 4576 -154 4640 -138
rect 4768 138 4832 154
rect 4768 -138 4783 138
rect 4783 -138 4817 138
rect 4817 -138 4832 138
rect 4768 -154 4832 -138
<< metal2 >>
rect -4832 155 -4768 165
rect -4832 -163 -4768 -153
rect -4640 154 -4576 164
rect -4640 -164 -4576 -154
rect -4448 154 -4384 164
rect -4448 -164 -4384 -154
rect -4256 154 -4192 164
rect -4256 -164 -4192 -154
rect -4064 154 -4000 164
rect -4064 -164 -4000 -154
rect -3872 154 -3808 164
rect -3872 -164 -3808 -154
rect -3680 154 -3616 164
rect -3680 -164 -3616 -154
rect -3488 154 -3424 164
rect -3488 -164 -3424 -154
rect -3296 154 -3232 164
rect -3296 -164 -3232 -154
rect -3104 154 -3040 164
rect -3104 -164 -3040 -154
rect -2912 154 -2848 164
rect -2912 -164 -2848 -154
rect -2720 154 -2656 164
rect -2720 -164 -2656 -154
rect -2528 154 -2464 164
rect -2528 -164 -2464 -154
rect -2336 154 -2272 164
rect -2336 -164 -2272 -154
rect -2144 154 -2080 164
rect -2144 -164 -2080 -154
rect -1952 154 -1888 164
rect -1952 -164 -1888 -154
rect -1760 154 -1696 164
rect -1760 -164 -1696 -154
rect -1568 154 -1504 164
rect -1568 -164 -1504 -154
rect -1376 154 -1312 164
rect -1376 -164 -1312 -154
rect -1184 154 -1120 164
rect -1184 -164 -1120 -154
rect -992 154 -928 164
rect -992 -164 -928 -154
rect -800 154 -736 164
rect -800 -164 -736 -154
rect -608 154 -544 164
rect -608 -164 -544 -154
rect -416 154 -352 164
rect -416 -164 -352 -154
rect -224 154 -160 164
rect -224 -164 -160 -154
rect -32 154 32 164
rect -32 -164 32 -154
rect 160 154 224 164
rect 160 -164 224 -154
rect 352 154 416 164
rect 352 -164 416 -154
rect 544 154 608 164
rect 544 -164 608 -154
rect 736 154 800 164
rect 736 -164 800 -154
rect 928 154 992 164
rect 928 -164 992 -154
rect 1120 154 1184 164
rect 1120 -164 1184 -154
rect 1312 154 1376 164
rect 1312 -164 1376 -154
rect 1504 154 1568 164
rect 1504 -164 1568 -154
rect 1696 154 1760 164
rect 1696 -164 1760 -154
rect 1888 154 1952 164
rect 1888 -164 1952 -154
rect 2080 154 2144 164
rect 2080 -164 2144 -154
rect 2272 154 2336 164
rect 2272 -164 2336 -154
rect 2464 154 2528 164
rect 2464 -164 2528 -154
rect 2656 154 2720 164
rect 2656 -164 2720 -154
rect 2848 154 2912 164
rect 2848 -164 2912 -154
rect 3040 154 3104 164
rect 3040 -164 3104 -154
rect 3232 154 3296 164
rect 3232 -164 3296 -154
rect 3424 154 3488 164
rect 3424 -164 3488 -154
rect 3616 154 3680 164
rect 3616 -164 3680 -154
rect 3808 154 3872 164
rect 3808 -164 3872 -154
rect 4000 154 4064 164
rect 4000 -164 4064 -154
rect 4192 154 4256 164
rect 4192 -164 4256 -154
rect 4384 154 4448 164
rect 4384 -164 4448 -154
rect 4576 154 4640 164
rect 4576 -164 4640 -154
rect 4768 154 4832 164
rect 4768 -164 4832 -154
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -4914 -307 4914 307
string parameters w 1.5 l 0.150 m 1 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
