magic
tech sky130A
magscale 1 2
timestamp 1624077215
<< error_p >>
rect 1165 618 1176 646
rect 1212 584 1223 618
rect 1284 584 1293 646
rect 1020 380 1024 414
rect 1130 308 1132 342
rect 904 238 908 272
rect 1462 244 1464 272
rect 1430 238 1464 244
rect 1174 90 1176 128
rect 1212 54 1214 90
<< nwell >>
rect 706 430 1756 808
<< nmos >>
rect 800 28 830 118
rect 1000 26 1030 206
rect 1088 26 1118 206
rect 1342 26 1372 206
rect 1430 26 1460 206
rect 1632 28 1662 118
<< pmos >>
rect 800 466 830 646
rect 1000 466 1030 646
rect 1088 466 1118 646
rect 1342 466 1372 646
rect 1430 466 1460 646
rect 1632 466 1662 646
<< ndiff >>
rect 742 88 800 118
rect 742 54 754 88
rect 788 54 800 88
rect 742 28 800 54
rect 830 88 888 118
rect 830 54 842 88
rect 876 54 888 88
rect 830 28 888 54
rect 942 88 1000 206
rect 942 54 954 88
rect 988 54 1000 88
rect 942 26 1000 54
rect 1030 88 1088 206
rect 1030 54 1042 88
rect 1076 54 1088 88
rect 1030 26 1088 54
rect 1118 88 1176 206
rect 1118 54 1130 88
rect 1164 54 1176 88
rect 1118 26 1176 54
rect 1284 88 1342 206
rect 1284 54 1296 88
rect 1330 54 1342 88
rect 1284 26 1342 54
rect 1372 26 1430 206
rect 1460 88 1518 206
rect 1460 54 1472 88
rect 1506 54 1518 88
rect 1460 26 1518 54
rect 1574 88 1632 118
rect 1574 54 1586 88
rect 1620 54 1632 88
rect 1574 28 1632 54
rect 1662 88 1720 118
rect 1662 54 1674 88
rect 1708 54 1720 88
rect 1662 28 1720 54
<< pdiff >>
rect 742 618 800 646
rect 742 584 754 618
rect 788 584 800 618
rect 742 466 800 584
rect 830 618 888 646
rect 830 584 842 618
rect 876 584 888 618
rect 830 466 888 584
rect 942 618 1000 646
rect 942 584 954 618
rect 988 584 1000 618
rect 942 466 1000 584
rect 1030 618 1088 646
rect 1030 584 1042 618
rect 1076 584 1088 618
rect 1030 466 1088 584
rect 1118 618 1176 646
rect 1118 584 1130 618
rect 1164 584 1176 618
rect 1118 466 1176 584
rect 1284 618 1342 646
rect 1284 584 1296 618
rect 1330 584 1342 618
rect 1284 466 1342 584
rect 1372 618 1430 646
rect 1372 584 1384 618
rect 1418 584 1430 618
rect 1372 466 1430 584
rect 1460 618 1518 646
rect 1460 584 1472 618
rect 1506 584 1518 618
rect 1460 466 1518 584
rect 1574 618 1632 646
rect 1574 584 1586 618
rect 1620 584 1632 618
rect 1574 466 1632 584
rect 1662 618 1720 646
rect 1662 584 1674 618
rect 1708 584 1720 618
rect 1662 466 1720 584
<< ndiffc >>
rect 754 54 788 88
rect 842 54 876 88
rect 954 54 988 88
rect 1042 54 1076 88
rect 1130 54 1164 88
rect 1296 54 1330 88
rect 1472 54 1506 88
rect 1586 54 1620 88
rect 1674 54 1708 88
<< pdiffc >>
rect 754 584 788 618
rect 842 584 876 618
rect 954 584 988 618
rect 1042 584 1076 618
rect 1130 584 1164 618
rect 1296 584 1330 618
rect 1384 584 1418 618
rect 1472 584 1506 618
rect 1586 584 1620 618
rect 1674 584 1708 618
<< psubdiff >>
rect 762 -64 786 -30
rect 1678 -64 1702 -30
<< nsubdiff >>
rect 762 736 786 770
rect 1676 736 1700 770
<< psubdiffcont >>
rect 786 -64 1678 -30
<< nsubdiffcont >>
rect 786 736 1676 770
<< poly >>
rect 800 646 830 672
rect 1000 646 1030 672
rect 1088 646 1118 672
rect 1342 646 1372 672
rect 1430 646 1460 672
rect 1632 646 1662 672
rect 1196 618 1262 632
rect 1196 584 1212 618
rect 1246 584 1262 618
rect 1196 566 1262 584
rect 800 288 830 466
rect 1000 430 1030 466
rect 970 414 1038 430
rect 970 380 990 414
rect 1020 380 1038 414
rect 970 364 1038 380
rect 800 272 922 288
rect 800 238 874 272
rect 904 238 922 272
rect 800 222 922 238
rect 800 118 830 222
rect 1000 206 1030 364
rect 1088 358 1118 466
rect 1080 342 1146 358
rect 1080 308 1098 342
rect 1130 308 1146 342
rect 1080 292 1146 308
rect 1088 206 1118 292
rect 800 2 830 28
rect 1212 104 1246 566
rect 1342 430 1372 466
rect 1322 414 1388 430
rect 1322 380 1338 414
rect 1372 380 1388 414
rect 1322 364 1388 380
rect 1342 206 1372 364
rect 1430 288 1460 466
rect 1632 430 1662 466
rect 1566 414 1662 430
rect 1566 380 1582 414
rect 1616 380 1662 414
rect 1566 364 1662 380
rect 1414 272 1478 288
rect 1414 238 1430 272
rect 1462 238 1478 272
rect 1414 222 1478 238
rect 1430 206 1460 222
rect 1196 90 1262 104
rect 1196 54 1212 90
rect 1246 54 1262 90
rect 1196 38 1262 54
rect 1632 118 1662 364
rect 1000 0 1030 26
rect 1088 0 1118 26
rect 1342 0 1372 26
rect 1430 0 1460 26
rect 1632 2 1662 28
<< polycont >>
rect 1212 584 1246 618
rect 990 380 1020 414
rect 874 238 904 272
rect 1098 308 1130 342
rect 1338 380 1372 414
rect 1582 380 1616 414
rect 1430 238 1462 272
rect 1212 54 1246 90
<< locali >>
rect 754 736 786 770
rect 1676 736 1692 770
rect 754 618 788 634
rect 754 414 788 584
rect 842 618 876 736
rect 842 568 876 584
rect 954 618 988 634
rect 954 534 988 584
rect 1042 618 1076 736
rect 1212 668 1506 702
rect 1042 568 1076 584
rect 1130 618 1164 634
rect 1130 534 1164 584
rect 1212 618 1246 668
rect 1212 568 1246 584
rect 1296 618 1330 668
rect 1296 568 1330 584
rect 1384 618 1418 634
rect 1384 534 1418 584
rect 1472 618 1506 668
rect 1472 568 1506 584
rect 1586 618 1620 736
rect 1586 568 1620 584
rect 1674 618 1708 634
rect 954 500 1418 534
rect 754 380 990 414
rect 1020 380 1040 414
rect 1322 380 1338 414
rect 1372 380 1582 414
rect 1616 380 1632 414
rect 754 88 788 380
rect 1674 342 1708 584
rect 1080 308 1098 342
rect 1130 308 1708 342
rect 854 238 874 272
rect 904 238 1428 272
rect 1462 238 1478 272
rect 754 38 788 54
rect 842 88 876 104
rect 842 -30 876 54
rect 954 88 988 104
rect 954 -30 988 54
rect 1042 88 1088 104
rect 1076 54 1088 88
rect 1042 38 1088 54
rect 1130 90 1330 104
rect 1130 88 1212 90
rect 1164 54 1212 88
rect 1246 88 1330 90
rect 1246 54 1296 88
rect 1130 38 1330 54
rect 1472 88 1506 104
rect 1472 -30 1506 54
rect 1586 88 1620 104
rect 1586 -30 1620 54
rect 1674 88 1708 308
rect 1674 38 1708 54
rect 754 -64 786 -30
rect 1678 -64 1694 -30
<< viali >>
rect 786 736 1676 770
rect 1338 380 1372 414
rect 1428 238 1430 272
rect 1430 238 1462 272
rect 1212 54 1246 90
rect 786 -64 1676 -30
<< metal1 >>
rect 706 770 1756 808
rect 706 736 786 770
rect 1676 736 1756 770
rect 706 698 1756 736
rect 1322 414 1388 430
rect 1322 380 1338 414
rect 1372 380 1388 414
rect 1322 364 1388 380
rect 1414 272 1478 288
rect 1414 238 1428 272
rect 1462 238 1478 272
rect 1414 222 1478 238
rect 1196 90 1262 104
rect 1196 54 1212 90
rect 1246 54 1262 90
rect 1196 38 1262 54
rect 706 -30 1756 8
rect 706 -64 786 -30
rect 1676 -64 1756 -30
rect 706 -102 1756 -64
<< labels >>
rlabel metal1 1196 38 1262 54 5 Z
rlabel metal1 1228 808 1228 808 1 VDD
rlabel metal1 1228 -102 1228 -102 5 VSS
rlabel metal1 1446 222 1446 222 5 B
rlabel metal1 1322 364 1388 380 5 A
<< end >>
