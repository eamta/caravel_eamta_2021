magic
tech sky130A
timestamp 1624067212
<< nwell >>
rect 1848 1107 1859 1156
rect 1819 38 1831 87
rect 1826 -1135 1838 -1080
<< poly >>
rect 3 1173 13 1185
rect 39 1173 49 1185
rect 1847 1173 1858 1185
rect 1847 1172 1857 1173
rect 1847 -1031 1857 -1009
<< metal1 >>
rect -60 1084 110 1185
rect 1848 1107 1859 1156
rect -60 137 40 1084
rect 1886 701 1986 1185
rect 1867 638 1986 701
rect 1858 588 1986 638
rect 1867 520 1986 588
rect -60 -88 130 137
rect 1819 38 1831 87
rect -60 -1035 40 -88
rect 1886 -472 1986 520
rect 1869 -529 1986 -472
rect 1857 -580 1986 -529
rect 1869 -653 1986 -580
rect -60 -1173 111 -1035
rect 1826 -1135 1838 -1080
rect 1886 -1173 1986 -653
<< metal2 >>
rect 1551 779 1579 807
rect 1551 414 1579 442
rect 1551 -394 1579 -366
rect 1551 -759 1579 -731
use c2b  c2b_1
timestamp 1624067212
transform 1 0 79 0 1 -575
box -79 -598 1793 587
use c2b  c2b_0
timestamp 1624067212
transform 1 0 79 0 1 598
box -79 -598 1793 587
<< labels >>
rlabel poly 3 1173 13 1185 1 clr
rlabel poly 39 1173 49 1185 1 clk
rlabel poly 1847 1172 1857 1184 1 ce
rlabel metal2 1551 779 1579 807 1 b0
rlabel metal2 1551 414 1579 442 1 b1
rlabel metal2 1551 -394 1579 -366 1 b2
rlabel metal2 1551 -759 1579 -731 1 b3
rlabel metal1 -48 1151 -14 1174 1 vdd
rlabel metal1 1906 1136 1964 1172 1 vss
rlabel poly 1847 -1031 1857 -1009 1 out
<< end >>
