**.subckt tb_inverter
x1 vdd out vin vss inverter
V1 vss GND 0
V2 vdd vss 1.8
V3 vin vss PULSE(0 {Vin} 1ps 1ps 1ps 50ns 100ns) DC{Vin} 
x2 vdd outb out vss inverter
C1 outb vss 1p m=1
**** begin user architecture code



* Parametros del circuito
.param Vin = 1.8
.options TEMP = 27.0

* Include
.lib /home/eamta/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT

* Signals to SAVE
.save all  @M.X1.XM1.msky130_fd_pr__nfet_01v8[id] @M.X1.XM1.msky130_fd_pr__nfet_01v8[gm]  @M.X1.XM2.msky130_fd_pr__pfet_01v8[id] @M.X1.XM2.msky130_fd_pr__pfet_01v8[gm]

*simulation
.control
  tran 0.1n 300ns
  setplot tran1
  plot v(out) v(vin)
  write tb_inverter_tran.raw

  reset
  dc V3 0 1.8 0.01
  setplot dc1
  plot v(out) v(vin)
  write tb_inverter_dc.raw

.endc



**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
* sym_path: /home/eamta/caravel_eamta_2021/track_vlsi/ledesma/sch/inverter.sym
* sch_path: /home/eamta/caravel_eamta_2021/track_vlsi/ledesma/sch/inverter.sch
.subckt inverter  vdd out in vss
*.opin out
*.ipin in
*.ipin vdd
*.ipin vss
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
