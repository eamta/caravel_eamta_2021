magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -1181 999 -1123 1005
rect -989 999 -931 1005
rect -797 999 -739 1005
rect -605 999 -547 1005
rect -413 999 -355 1005
rect -221 999 -163 1005
rect -29 999 29 1005
rect 163 999 221 1005
rect 355 999 413 1005
rect 547 999 605 1005
rect 739 999 797 1005
rect 931 999 989 1005
rect 1123 999 1181 1005
rect -1181 965 -1169 999
rect -989 965 -977 999
rect -797 965 -785 999
rect -605 965 -593 999
rect -413 965 -401 999
rect -221 965 -209 999
rect -29 965 -17 999
rect 163 965 175 999
rect 355 965 367 999
rect 547 965 559 999
rect 739 965 751 999
rect 931 965 943 999
rect 1123 965 1135 999
rect -1181 959 -1123 965
rect -989 959 -931 965
rect -797 959 -739 965
rect -605 959 -547 965
rect -413 959 -355 965
rect -221 959 -163 965
rect -29 959 29 965
rect 163 959 221 965
rect 355 959 413 965
rect 547 959 605 965
rect 739 959 797 965
rect 931 959 989 965
rect 1123 959 1181 965
rect -1085 589 -1027 595
rect -893 589 -835 595
rect -701 589 -643 595
rect -509 589 -451 595
rect -317 589 -259 595
rect -125 589 -67 595
rect 67 589 125 595
rect 259 589 317 595
rect 451 589 509 595
rect 643 589 701 595
rect 835 589 893 595
rect 1027 589 1085 595
rect -1085 555 -1073 589
rect -893 555 -881 589
rect -701 555 -689 589
rect -509 555 -497 589
rect -317 555 -305 589
rect -125 555 -113 589
rect 67 555 79 589
rect 259 555 271 589
rect 451 555 463 589
rect 643 555 655 589
rect 835 555 847 589
rect 1027 555 1039 589
rect -1085 549 -1027 555
rect -893 549 -835 555
rect -701 549 -643 555
rect -509 549 -451 555
rect -317 549 -259 555
rect -125 549 -67 555
rect 67 549 125 555
rect 259 549 317 555
rect 451 549 509 555
rect 643 549 701 555
rect 835 549 893 555
rect 1027 549 1085 555
rect -1085 481 -1027 487
rect -893 481 -835 487
rect -701 481 -643 487
rect -509 481 -451 487
rect -317 481 -259 487
rect -125 481 -67 487
rect 67 481 125 487
rect 259 481 317 487
rect 451 481 509 487
rect 643 481 701 487
rect 835 481 893 487
rect 1027 481 1085 487
rect -1085 447 -1073 481
rect -893 447 -881 481
rect -701 447 -689 481
rect -509 447 -497 481
rect -317 447 -305 481
rect -125 447 -113 481
rect 67 447 79 481
rect 259 447 271 481
rect 451 447 463 481
rect 643 447 655 481
rect 835 447 847 481
rect 1027 447 1039 481
rect -1085 441 -1027 447
rect -893 441 -835 447
rect -701 441 -643 447
rect -509 441 -451 447
rect -317 441 -259 447
rect -125 441 -67 447
rect 67 441 125 447
rect 259 441 317 447
rect 451 441 509 447
rect 643 441 701 447
rect 835 441 893 447
rect 1027 441 1085 447
rect -1181 71 -1123 77
rect -989 71 -931 77
rect -797 71 -739 77
rect -605 71 -547 77
rect -413 71 -355 77
rect -221 71 -163 77
rect -29 71 29 77
rect 163 71 221 77
rect 355 71 413 77
rect 547 71 605 77
rect 739 71 797 77
rect 931 71 989 77
rect 1123 71 1181 77
rect -1181 37 -1169 71
rect -989 37 -977 71
rect -797 37 -785 71
rect -605 37 -593 71
rect -413 37 -401 71
rect -221 37 -209 71
rect -29 37 -17 71
rect 163 37 175 71
rect 355 37 367 71
rect 547 37 559 71
rect 739 37 751 71
rect 931 37 943 71
rect 1123 37 1135 71
rect -1181 31 -1123 37
rect -989 31 -931 37
rect -797 31 -739 37
rect -605 31 -547 37
rect -413 31 -355 37
rect -221 31 -163 37
rect -29 31 29 37
rect 163 31 221 37
rect 355 31 413 37
rect 547 31 605 37
rect 739 31 797 37
rect 931 31 989 37
rect 1123 31 1181 37
rect -1181 -37 -1123 -31
rect -989 -37 -931 -31
rect -797 -37 -739 -31
rect -605 -37 -547 -31
rect -413 -37 -355 -31
rect -221 -37 -163 -31
rect -29 -37 29 -31
rect 163 -37 221 -31
rect 355 -37 413 -31
rect 547 -37 605 -31
rect 739 -37 797 -31
rect 931 -37 989 -31
rect 1123 -37 1181 -31
rect -1181 -71 -1169 -37
rect -989 -71 -977 -37
rect -797 -71 -785 -37
rect -605 -71 -593 -37
rect -413 -71 -401 -37
rect -221 -71 -209 -37
rect -29 -71 -17 -37
rect 163 -71 175 -37
rect 355 -71 367 -37
rect 547 -71 559 -37
rect 739 -71 751 -37
rect 931 -71 943 -37
rect 1123 -71 1135 -37
rect -1181 -77 -1123 -71
rect -989 -77 -931 -71
rect -797 -77 -739 -71
rect -605 -77 -547 -71
rect -413 -77 -355 -71
rect -221 -77 -163 -71
rect -29 -77 29 -71
rect 163 -77 221 -71
rect 355 -77 413 -71
rect 547 -77 605 -71
rect 739 -77 797 -71
rect 931 -77 989 -71
rect 1123 -77 1181 -71
rect -1085 -447 -1027 -441
rect -893 -447 -835 -441
rect -701 -447 -643 -441
rect -509 -447 -451 -441
rect -317 -447 -259 -441
rect -125 -447 -67 -441
rect 67 -447 125 -441
rect 259 -447 317 -441
rect 451 -447 509 -441
rect 643 -447 701 -441
rect 835 -447 893 -441
rect 1027 -447 1085 -441
rect -1085 -481 -1073 -447
rect -893 -481 -881 -447
rect -701 -481 -689 -447
rect -509 -481 -497 -447
rect -317 -481 -305 -447
rect -125 -481 -113 -447
rect 67 -481 79 -447
rect 259 -481 271 -447
rect 451 -481 463 -447
rect 643 -481 655 -447
rect 835 -481 847 -447
rect 1027 -481 1039 -447
rect -1085 -487 -1027 -481
rect -893 -487 -835 -481
rect -701 -487 -643 -481
rect -509 -487 -451 -481
rect -317 -487 -259 -481
rect -125 -487 -67 -481
rect 67 -487 125 -481
rect 259 -487 317 -481
rect 451 -487 509 -481
rect 643 -487 701 -481
rect 835 -487 893 -481
rect 1027 -487 1085 -481
rect -1085 -555 -1027 -549
rect -893 -555 -835 -549
rect -701 -555 -643 -549
rect -509 -555 -451 -549
rect -317 -555 -259 -549
rect -125 -555 -67 -549
rect 67 -555 125 -549
rect 259 -555 317 -549
rect 451 -555 509 -549
rect 643 -555 701 -549
rect 835 -555 893 -549
rect 1027 -555 1085 -549
rect -1085 -589 -1073 -555
rect -893 -589 -881 -555
rect -701 -589 -689 -555
rect -509 -589 -497 -555
rect -317 -589 -305 -555
rect -125 -589 -113 -555
rect 67 -589 79 -555
rect 259 -589 271 -555
rect 451 -589 463 -555
rect 643 -589 655 -555
rect 835 -589 847 -555
rect 1027 -589 1039 -555
rect -1085 -595 -1027 -589
rect -893 -595 -835 -589
rect -701 -595 -643 -589
rect -509 -595 -451 -589
rect -317 -595 -259 -589
rect -125 -595 -67 -589
rect 67 -595 125 -589
rect 259 -595 317 -589
rect 451 -595 509 -589
rect 643 -595 701 -589
rect 835 -595 893 -589
rect 1027 -595 1085 -589
rect -1181 -965 -1123 -959
rect -989 -965 -931 -959
rect -797 -965 -739 -959
rect -605 -965 -547 -959
rect -413 -965 -355 -959
rect -221 -965 -163 -959
rect -29 -965 29 -959
rect 163 -965 221 -959
rect 355 -965 413 -959
rect 547 -965 605 -959
rect 739 -965 797 -959
rect 931 -965 989 -959
rect 1123 -965 1181 -959
rect -1181 -999 -1169 -965
rect -989 -999 -977 -965
rect -797 -999 -785 -965
rect -605 -999 -593 -965
rect -413 -999 -401 -965
rect -221 -999 -209 -965
rect -29 -999 -17 -965
rect 163 -999 175 -965
rect 355 -999 367 -965
rect 547 -999 559 -965
rect 739 -999 751 -965
rect 931 -999 943 -965
rect 1123 -999 1135 -965
rect -1181 -1005 -1123 -999
rect -989 -1005 -931 -999
rect -797 -1005 -739 -999
rect -605 -1005 -547 -999
rect -413 -1005 -355 -999
rect -221 -1005 -163 -999
rect -29 -1005 29 -999
rect 163 -1005 221 -999
rect 355 -1005 413 -999
rect 547 -1005 605 -999
rect 739 -1005 797 -999
rect 931 -1005 989 -999
rect 1123 -1005 1181 -999
<< pwell >>
rect -1367 -1137 1367 1137
<< nmos >>
rect -1167 627 -1137 927
rect -1071 627 -1041 927
rect -975 627 -945 927
rect -879 627 -849 927
rect -783 627 -753 927
rect -687 627 -657 927
rect -591 627 -561 927
rect -495 627 -465 927
rect -399 627 -369 927
rect -303 627 -273 927
rect -207 627 -177 927
rect -111 627 -81 927
rect -15 627 15 927
rect 81 627 111 927
rect 177 627 207 927
rect 273 627 303 927
rect 369 627 399 927
rect 465 627 495 927
rect 561 627 591 927
rect 657 627 687 927
rect 753 627 783 927
rect 849 627 879 927
rect 945 627 975 927
rect 1041 627 1071 927
rect 1137 627 1167 927
rect -1167 109 -1137 409
rect -1071 109 -1041 409
rect -975 109 -945 409
rect -879 109 -849 409
rect -783 109 -753 409
rect -687 109 -657 409
rect -591 109 -561 409
rect -495 109 -465 409
rect -399 109 -369 409
rect -303 109 -273 409
rect -207 109 -177 409
rect -111 109 -81 409
rect -15 109 15 409
rect 81 109 111 409
rect 177 109 207 409
rect 273 109 303 409
rect 369 109 399 409
rect 465 109 495 409
rect 561 109 591 409
rect 657 109 687 409
rect 753 109 783 409
rect 849 109 879 409
rect 945 109 975 409
rect 1041 109 1071 409
rect 1137 109 1167 409
rect -1167 -409 -1137 -109
rect -1071 -409 -1041 -109
rect -975 -409 -945 -109
rect -879 -409 -849 -109
rect -783 -409 -753 -109
rect -687 -409 -657 -109
rect -591 -409 -561 -109
rect -495 -409 -465 -109
rect -399 -409 -369 -109
rect -303 -409 -273 -109
rect -207 -409 -177 -109
rect -111 -409 -81 -109
rect -15 -409 15 -109
rect 81 -409 111 -109
rect 177 -409 207 -109
rect 273 -409 303 -109
rect 369 -409 399 -109
rect 465 -409 495 -109
rect 561 -409 591 -109
rect 657 -409 687 -109
rect 753 -409 783 -109
rect 849 -409 879 -109
rect 945 -409 975 -109
rect 1041 -409 1071 -109
rect 1137 -409 1167 -109
rect -1167 -927 -1137 -627
rect -1071 -927 -1041 -627
rect -975 -927 -945 -627
rect -879 -927 -849 -627
rect -783 -927 -753 -627
rect -687 -927 -657 -627
rect -591 -927 -561 -627
rect -495 -927 -465 -627
rect -399 -927 -369 -627
rect -303 -927 -273 -627
rect -207 -927 -177 -627
rect -111 -927 -81 -627
rect -15 -927 15 -627
rect 81 -927 111 -627
rect 177 -927 207 -627
rect 273 -927 303 -627
rect 369 -927 399 -627
rect 465 -927 495 -627
rect 561 -927 591 -627
rect 657 -927 687 -627
rect 753 -927 783 -627
rect 849 -927 879 -627
rect 945 -927 975 -627
rect 1041 -927 1071 -627
rect 1137 -927 1167 -627
<< ndiff >>
rect -1229 915 -1167 927
rect -1229 639 -1217 915
rect -1183 639 -1167 915
rect -1229 627 -1167 639
rect -1137 915 -1071 927
rect -1137 639 -1121 915
rect -1087 639 -1071 915
rect -1137 627 -1071 639
rect -1041 915 -975 927
rect -1041 639 -1025 915
rect -991 639 -975 915
rect -1041 627 -975 639
rect -945 915 -879 927
rect -945 639 -929 915
rect -895 639 -879 915
rect -945 627 -879 639
rect -849 915 -783 927
rect -849 639 -833 915
rect -799 639 -783 915
rect -849 627 -783 639
rect -753 915 -687 927
rect -753 639 -737 915
rect -703 639 -687 915
rect -753 627 -687 639
rect -657 915 -591 927
rect -657 639 -641 915
rect -607 639 -591 915
rect -657 627 -591 639
rect -561 915 -495 927
rect -561 639 -545 915
rect -511 639 -495 915
rect -561 627 -495 639
rect -465 915 -399 927
rect -465 639 -449 915
rect -415 639 -399 915
rect -465 627 -399 639
rect -369 915 -303 927
rect -369 639 -353 915
rect -319 639 -303 915
rect -369 627 -303 639
rect -273 915 -207 927
rect -273 639 -257 915
rect -223 639 -207 915
rect -273 627 -207 639
rect -177 915 -111 927
rect -177 639 -161 915
rect -127 639 -111 915
rect -177 627 -111 639
rect -81 915 -15 927
rect -81 639 -65 915
rect -31 639 -15 915
rect -81 627 -15 639
rect 15 915 81 927
rect 15 639 31 915
rect 65 639 81 915
rect 15 627 81 639
rect 111 915 177 927
rect 111 639 127 915
rect 161 639 177 915
rect 111 627 177 639
rect 207 915 273 927
rect 207 639 223 915
rect 257 639 273 915
rect 207 627 273 639
rect 303 915 369 927
rect 303 639 319 915
rect 353 639 369 915
rect 303 627 369 639
rect 399 915 465 927
rect 399 639 415 915
rect 449 639 465 915
rect 399 627 465 639
rect 495 915 561 927
rect 495 639 511 915
rect 545 639 561 915
rect 495 627 561 639
rect 591 915 657 927
rect 591 639 607 915
rect 641 639 657 915
rect 591 627 657 639
rect 687 915 753 927
rect 687 639 703 915
rect 737 639 753 915
rect 687 627 753 639
rect 783 915 849 927
rect 783 639 799 915
rect 833 639 849 915
rect 783 627 849 639
rect 879 915 945 927
rect 879 639 895 915
rect 929 639 945 915
rect 879 627 945 639
rect 975 915 1041 927
rect 975 639 991 915
rect 1025 639 1041 915
rect 975 627 1041 639
rect 1071 915 1137 927
rect 1071 639 1087 915
rect 1121 639 1137 915
rect 1071 627 1137 639
rect 1167 915 1229 927
rect 1167 639 1183 915
rect 1217 639 1229 915
rect 1167 627 1229 639
rect -1229 397 -1167 409
rect -1229 121 -1217 397
rect -1183 121 -1167 397
rect -1229 109 -1167 121
rect -1137 397 -1071 409
rect -1137 121 -1121 397
rect -1087 121 -1071 397
rect -1137 109 -1071 121
rect -1041 397 -975 409
rect -1041 121 -1025 397
rect -991 121 -975 397
rect -1041 109 -975 121
rect -945 397 -879 409
rect -945 121 -929 397
rect -895 121 -879 397
rect -945 109 -879 121
rect -849 397 -783 409
rect -849 121 -833 397
rect -799 121 -783 397
rect -849 109 -783 121
rect -753 397 -687 409
rect -753 121 -737 397
rect -703 121 -687 397
rect -753 109 -687 121
rect -657 397 -591 409
rect -657 121 -641 397
rect -607 121 -591 397
rect -657 109 -591 121
rect -561 397 -495 409
rect -561 121 -545 397
rect -511 121 -495 397
rect -561 109 -495 121
rect -465 397 -399 409
rect -465 121 -449 397
rect -415 121 -399 397
rect -465 109 -399 121
rect -369 397 -303 409
rect -369 121 -353 397
rect -319 121 -303 397
rect -369 109 -303 121
rect -273 397 -207 409
rect -273 121 -257 397
rect -223 121 -207 397
rect -273 109 -207 121
rect -177 397 -111 409
rect -177 121 -161 397
rect -127 121 -111 397
rect -177 109 -111 121
rect -81 397 -15 409
rect -81 121 -65 397
rect -31 121 -15 397
rect -81 109 -15 121
rect 15 397 81 409
rect 15 121 31 397
rect 65 121 81 397
rect 15 109 81 121
rect 111 397 177 409
rect 111 121 127 397
rect 161 121 177 397
rect 111 109 177 121
rect 207 397 273 409
rect 207 121 223 397
rect 257 121 273 397
rect 207 109 273 121
rect 303 397 369 409
rect 303 121 319 397
rect 353 121 369 397
rect 303 109 369 121
rect 399 397 465 409
rect 399 121 415 397
rect 449 121 465 397
rect 399 109 465 121
rect 495 397 561 409
rect 495 121 511 397
rect 545 121 561 397
rect 495 109 561 121
rect 591 397 657 409
rect 591 121 607 397
rect 641 121 657 397
rect 591 109 657 121
rect 687 397 753 409
rect 687 121 703 397
rect 737 121 753 397
rect 687 109 753 121
rect 783 397 849 409
rect 783 121 799 397
rect 833 121 849 397
rect 783 109 849 121
rect 879 397 945 409
rect 879 121 895 397
rect 929 121 945 397
rect 879 109 945 121
rect 975 397 1041 409
rect 975 121 991 397
rect 1025 121 1041 397
rect 975 109 1041 121
rect 1071 397 1137 409
rect 1071 121 1087 397
rect 1121 121 1137 397
rect 1071 109 1137 121
rect 1167 397 1229 409
rect 1167 121 1183 397
rect 1217 121 1229 397
rect 1167 109 1229 121
rect -1229 -121 -1167 -109
rect -1229 -397 -1217 -121
rect -1183 -397 -1167 -121
rect -1229 -409 -1167 -397
rect -1137 -121 -1071 -109
rect -1137 -397 -1121 -121
rect -1087 -397 -1071 -121
rect -1137 -409 -1071 -397
rect -1041 -121 -975 -109
rect -1041 -397 -1025 -121
rect -991 -397 -975 -121
rect -1041 -409 -975 -397
rect -945 -121 -879 -109
rect -945 -397 -929 -121
rect -895 -397 -879 -121
rect -945 -409 -879 -397
rect -849 -121 -783 -109
rect -849 -397 -833 -121
rect -799 -397 -783 -121
rect -849 -409 -783 -397
rect -753 -121 -687 -109
rect -753 -397 -737 -121
rect -703 -397 -687 -121
rect -753 -409 -687 -397
rect -657 -121 -591 -109
rect -657 -397 -641 -121
rect -607 -397 -591 -121
rect -657 -409 -591 -397
rect -561 -121 -495 -109
rect -561 -397 -545 -121
rect -511 -397 -495 -121
rect -561 -409 -495 -397
rect -465 -121 -399 -109
rect -465 -397 -449 -121
rect -415 -397 -399 -121
rect -465 -409 -399 -397
rect -369 -121 -303 -109
rect -369 -397 -353 -121
rect -319 -397 -303 -121
rect -369 -409 -303 -397
rect -273 -121 -207 -109
rect -273 -397 -257 -121
rect -223 -397 -207 -121
rect -273 -409 -207 -397
rect -177 -121 -111 -109
rect -177 -397 -161 -121
rect -127 -397 -111 -121
rect -177 -409 -111 -397
rect -81 -121 -15 -109
rect -81 -397 -65 -121
rect -31 -397 -15 -121
rect -81 -409 -15 -397
rect 15 -121 81 -109
rect 15 -397 31 -121
rect 65 -397 81 -121
rect 15 -409 81 -397
rect 111 -121 177 -109
rect 111 -397 127 -121
rect 161 -397 177 -121
rect 111 -409 177 -397
rect 207 -121 273 -109
rect 207 -397 223 -121
rect 257 -397 273 -121
rect 207 -409 273 -397
rect 303 -121 369 -109
rect 303 -397 319 -121
rect 353 -397 369 -121
rect 303 -409 369 -397
rect 399 -121 465 -109
rect 399 -397 415 -121
rect 449 -397 465 -121
rect 399 -409 465 -397
rect 495 -121 561 -109
rect 495 -397 511 -121
rect 545 -397 561 -121
rect 495 -409 561 -397
rect 591 -121 657 -109
rect 591 -397 607 -121
rect 641 -397 657 -121
rect 591 -409 657 -397
rect 687 -121 753 -109
rect 687 -397 703 -121
rect 737 -397 753 -121
rect 687 -409 753 -397
rect 783 -121 849 -109
rect 783 -397 799 -121
rect 833 -397 849 -121
rect 783 -409 849 -397
rect 879 -121 945 -109
rect 879 -397 895 -121
rect 929 -397 945 -121
rect 879 -409 945 -397
rect 975 -121 1041 -109
rect 975 -397 991 -121
rect 1025 -397 1041 -121
rect 975 -409 1041 -397
rect 1071 -121 1137 -109
rect 1071 -397 1087 -121
rect 1121 -397 1137 -121
rect 1071 -409 1137 -397
rect 1167 -121 1229 -109
rect 1167 -397 1183 -121
rect 1217 -397 1229 -121
rect 1167 -409 1229 -397
rect -1229 -639 -1167 -627
rect -1229 -915 -1217 -639
rect -1183 -915 -1167 -639
rect -1229 -927 -1167 -915
rect -1137 -639 -1071 -627
rect -1137 -915 -1121 -639
rect -1087 -915 -1071 -639
rect -1137 -927 -1071 -915
rect -1041 -639 -975 -627
rect -1041 -915 -1025 -639
rect -991 -915 -975 -639
rect -1041 -927 -975 -915
rect -945 -639 -879 -627
rect -945 -915 -929 -639
rect -895 -915 -879 -639
rect -945 -927 -879 -915
rect -849 -639 -783 -627
rect -849 -915 -833 -639
rect -799 -915 -783 -639
rect -849 -927 -783 -915
rect -753 -639 -687 -627
rect -753 -915 -737 -639
rect -703 -915 -687 -639
rect -753 -927 -687 -915
rect -657 -639 -591 -627
rect -657 -915 -641 -639
rect -607 -915 -591 -639
rect -657 -927 -591 -915
rect -561 -639 -495 -627
rect -561 -915 -545 -639
rect -511 -915 -495 -639
rect -561 -927 -495 -915
rect -465 -639 -399 -627
rect -465 -915 -449 -639
rect -415 -915 -399 -639
rect -465 -927 -399 -915
rect -369 -639 -303 -627
rect -369 -915 -353 -639
rect -319 -915 -303 -639
rect -369 -927 -303 -915
rect -273 -639 -207 -627
rect -273 -915 -257 -639
rect -223 -915 -207 -639
rect -273 -927 -207 -915
rect -177 -639 -111 -627
rect -177 -915 -161 -639
rect -127 -915 -111 -639
rect -177 -927 -111 -915
rect -81 -639 -15 -627
rect -81 -915 -65 -639
rect -31 -915 -15 -639
rect -81 -927 -15 -915
rect 15 -639 81 -627
rect 15 -915 31 -639
rect 65 -915 81 -639
rect 15 -927 81 -915
rect 111 -639 177 -627
rect 111 -915 127 -639
rect 161 -915 177 -639
rect 111 -927 177 -915
rect 207 -639 273 -627
rect 207 -915 223 -639
rect 257 -915 273 -639
rect 207 -927 273 -915
rect 303 -639 369 -627
rect 303 -915 319 -639
rect 353 -915 369 -639
rect 303 -927 369 -915
rect 399 -639 465 -627
rect 399 -915 415 -639
rect 449 -915 465 -639
rect 399 -927 465 -915
rect 495 -639 561 -627
rect 495 -915 511 -639
rect 545 -915 561 -639
rect 495 -927 561 -915
rect 591 -639 657 -627
rect 591 -915 607 -639
rect 641 -915 657 -639
rect 591 -927 657 -915
rect 687 -639 753 -627
rect 687 -915 703 -639
rect 737 -915 753 -639
rect 687 -927 753 -915
rect 783 -639 849 -627
rect 783 -915 799 -639
rect 833 -915 849 -639
rect 783 -927 849 -915
rect 879 -639 945 -627
rect 879 -915 895 -639
rect 929 -915 945 -639
rect 879 -927 945 -915
rect 975 -639 1041 -627
rect 975 -915 991 -639
rect 1025 -915 1041 -639
rect 975 -927 1041 -915
rect 1071 -639 1137 -627
rect 1071 -915 1087 -639
rect 1121 -915 1137 -639
rect 1071 -927 1137 -915
rect 1167 -639 1229 -627
rect 1167 -915 1183 -639
rect 1217 -915 1229 -639
rect 1167 -927 1229 -915
<< ndiffc >>
rect -1217 639 -1183 915
rect -1121 639 -1087 915
rect -1025 639 -991 915
rect -929 639 -895 915
rect -833 639 -799 915
rect -737 639 -703 915
rect -641 639 -607 915
rect -545 639 -511 915
rect -449 639 -415 915
rect -353 639 -319 915
rect -257 639 -223 915
rect -161 639 -127 915
rect -65 639 -31 915
rect 31 639 65 915
rect 127 639 161 915
rect 223 639 257 915
rect 319 639 353 915
rect 415 639 449 915
rect 511 639 545 915
rect 607 639 641 915
rect 703 639 737 915
rect 799 639 833 915
rect 895 639 929 915
rect 991 639 1025 915
rect 1087 639 1121 915
rect 1183 639 1217 915
rect -1217 121 -1183 397
rect -1121 121 -1087 397
rect -1025 121 -991 397
rect -929 121 -895 397
rect -833 121 -799 397
rect -737 121 -703 397
rect -641 121 -607 397
rect -545 121 -511 397
rect -449 121 -415 397
rect -353 121 -319 397
rect -257 121 -223 397
rect -161 121 -127 397
rect -65 121 -31 397
rect 31 121 65 397
rect 127 121 161 397
rect 223 121 257 397
rect 319 121 353 397
rect 415 121 449 397
rect 511 121 545 397
rect 607 121 641 397
rect 703 121 737 397
rect 799 121 833 397
rect 895 121 929 397
rect 991 121 1025 397
rect 1087 121 1121 397
rect 1183 121 1217 397
rect -1217 -397 -1183 -121
rect -1121 -397 -1087 -121
rect -1025 -397 -991 -121
rect -929 -397 -895 -121
rect -833 -397 -799 -121
rect -737 -397 -703 -121
rect -641 -397 -607 -121
rect -545 -397 -511 -121
rect -449 -397 -415 -121
rect -353 -397 -319 -121
rect -257 -397 -223 -121
rect -161 -397 -127 -121
rect -65 -397 -31 -121
rect 31 -397 65 -121
rect 127 -397 161 -121
rect 223 -397 257 -121
rect 319 -397 353 -121
rect 415 -397 449 -121
rect 511 -397 545 -121
rect 607 -397 641 -121
rect 703 -397 737 -121
rect 799 -397 833 -121
rect 895 -397 929 -121
rect 991 -397 1025 -121
rect 1087 -397 1121 -121
rect 1183 -397 1217 -121
rect -1217 -915 -1183 -639
rect -1121 -915 -1087 -639
rect -1025 -915 -991 -639
rect -929 -915 -895 -639
rect -833 -915 -799 -639
rect -737 -915 -703 -639
rect -641 -915 -607 -639
rect -545 -915 -511 -639
rect -449 -915 -415 -639
rect -353 -915 -319 -639
rect -257 -915 -223 -639
rect -161 -915 -127 -639
rect -65 -915 -31 -639
rect 31 -915 65 -639
rect 127 -915 161 -639
rect 223 -915 257 -639
rect 319 -915 353 -639
rect 415 -915 449 -639
rect 511 -915 545 -639
rect 607 -915 641 -639
rect 703 -915 737 -639
rect 799 -915 833 -639
rect 895 -915 929 -639
rect 991 -915 1025 -639
rect 1087 -915 1121 -639
rect 1183 -915 1217 -639
<< psubdiff >>
rect -1331 1067 -1235 1101
rect 1235 1067 1331 1101
rect -1331 1005 -1297 1067
rect 1297 1005 1331 1067
rect -1331 -1067 -1297 -1005
rect 1297 -1067 1331 -1005
rect -1331 -1101 -1235 -1067
rect 1235 -1101 1331 -1067
<< psubdiffcont >>
rect -1235 1067 1235 1101
rect -1331 -1005 -1297 1005
rect 1297 -1005 1331 1005
rect -1235 -1101 1235 -1067
<< poly >>
rect -1185 999 -1119 1015
rect -1185 965 -1169 999
rect -1135 965 -1119 999
rect -1185 949 -1119 965
rect -993 999 -927 1015
rect -993 965 -977 999
rect -943 965 -927 999
rect -1167 927 -1137 949
rect -1071 927 -1041 953
rect -993 949 -927 965
rect -801 999 -735 1015
rect -801 965 -785 999
rect -751 965 -735 999
rect -975 927 -945 949
rect -879 927 -849 953
rect -801 949 -735 965
rect -609 999 -543 1015
rect -609 965 -593 999
rect -559 965 -543 999
rect -783 927 -753 949
rect -687 927 -657 953
rect -609 949 -543 965
rect -417 999 -351 1015
rect -417 965 -401 999
rect -367 965 -351 999
rect -591 927 -561 949
rect -495 927 -465 953
rect -417 949 -351 965
rect -225 999 -159 1015
rect -225 965 -209 999
rect -175 965 -159 999
rect -399 927 -369 949
rect -303 927 -273 953
rect -225 949 -159 965
rect -33 999 33 1015
rect -33 965 -17 999
rect 17 965 33 999
rect -207 927 -177 949
rect -111 927 -81 953
rect -33 949 33 965
rect 159 999 225 1015
rect 159 965 175 999
rect 209 965 225 999
rect -15 927 15 949
rect 81 927 111 953
rect 159 949 225 965
rect 351 999 417 1015
rect 351 965 367 999
rect 401 965 417 999
rect 177 927 207 949
rect 273 927 303 953
rect 351 949 417 965
rect 543 999 609 1015
rect 543 965 559 999
rect 593 965 609 999
rect 369 927 399 949
rect 465 927 495 953
rect 543 949 609 965
rect 735 999 801 1015
rect 735 965 751 999
rect 785 965 801 999
rect 561 927 591 949
rect 657 927 687 953
rect 735 949 801 965
rect 927 999 993 1015
rect 927 965 943 999
rect 977 965 993 999
rect 753 927 783 949
rect 849 927 879 953
rect 927 949 993 965
rect 1119 999 1185 1015
rect 1119 965 1135 999
rect 1169 965 1185 999
rect 945 927 975 949
rect 1041 927 1071 953
rect 1119 949 1185 965
rect 1137 927 1167 949
rect -1167 601 -1137 627
rect -1071 605 -1041 627
rect -1089 589 -1023 605
rect -975 601 -945 627
rect -879 605 -849 627
rect -1089 555 -1073 589
rect -1039 555 -1023 589
rect -1089 539 -1023 555
rect -897 589 -831 605
rect -783 601 -753 627
rect -687 605 -657 627
rect -897 555 -881 589
rect -847 555 -831 589
rect -897 539 -831 555
rect -705 589 -639 605
rect -591 601 -561 627
rect -495 605 -465 627
rect -705 555 -689 589
rect -655 555 -639 589
rect -705 539 -639 555
rect -513 589 -447 605
rect -399 601 -369 627
rect -303 605 -273 627
rect -513 555 -497 589
rect -463 555 -447 589
rect -513 539 -447 555
rect -321 589 -255 605
rect -207 601 -177 627
rect -111 605 -81 627
rect -321 555 -305 589
rect -271 555 -255 589
rect -321 539 -255 555
rect -129 589 -63 605
rect -15 601 15 627
rect 81 605 111 627
rect -129 555 -113 589
rect -79 555 -63 589
rect -129 539 -63 555
rect 63 589 129 605
rect 177 601 207 627
rect 273 605 303 627
rect 63 555 79 589
rect 113 555 129 589
rect 63 539 129 555
rect 255 589 321 605
rect 369 601 399 627
rect 465 605 495 627
rect 255 555 271 589
rect 305 555 321 589
rect 255 539 321 555
rect 447 589 513 605
rect 561 601 591 627
rect 657 605 687 627
rect 447 555 463 589
rect 497 555 513 589
rect 447 539 513 555
rect 639 589 705 605
rect 753 601 783 627
rect 849 605 879 627
rect 639 555 655 589
rect 689 555 705 589
rect 639 539 705 555
rect 831 589 897 605
rect 945 601 975 627
rect 1041 605 1071 627
rect 831 555 847 589
rect 881 555 897 589
rect 831 539 897 555
rect 1023 589 1089 605
rect 1137 601 1167 627
rect 1023 555 1039 589
rect 1073 555 1089 589
rect 1023 539 1089 555
rect -1089 481 -1023 497
rect -1089 447 -1073 481
rect -1039 447 -1023 481
rect -1167 409 -1137 435
rect -1089 431 -1023 447
rect -897 481 -831 497
rect -897 447 -881 481
rect -847 447 -831 481
rect -1071 409 -1041 431
rect -975 409 -945 435
rect -897 431 -831 447
rect -705 481 -639 497
rect -705 447 -689 481
rect -655 447 -639 481
rect -879 409 -849 431
rect -783 409 -753 435
rect -705 431 -639 447
rect -513 481 -447 497
rect -513 447 -497 481
rect -463 447 -447 481
rect -687 409 -657 431
rect -591 409 -561 435
rect -513 431 -447 447
rect -321 481 -255 497
rect -321 447 -305 481
rect -271 447 -255 481
rect -495 409 -465 431
rect -399 409 -369 435
rect -321 431 -255 447
rect -129 481 -63 497
rect -129 447 -113 481
rect -79 447 -63 481
rect -303 409 -273 431
rect -207 409 -177 435
rect -129 431 -63 447
rect 63 481 129 497
rect 63 447 79 481
rect 113 447 129 481
rect -111 409 -81 431
rect -15 409 15 435
rect 63 431 129 447
rect 255 481 321 497
rect 255 447 271 481
rect 305 447 321 481
rect 81 409 111 431
rect 177 409 207 435
rect 255 431 321 447
rect 447 481 513 497
rect 447 447 463 481
rect 497 447 513 481
rect 273 409 303 431
rect 369 409 399 435
rect 447 431 513 447
rect 639 481 705 497
rect 639 447 655 481
rect 689 447 705 481
rect 465 409 495 431
rect 561 409 591 435
rect 639 431 705 447
rect 831 481 897 497
rect 831 447 847 481
rect 881 447 897 481
rect 657 409 687 431
rect 753 409 783 435
rect 831 431 897 447
rect 1023 481 1089 497
rect 1023 447 1039 481
rect 1073 447 1089 481
rect 849 409 879 431
rect 945 409 975 435
rect 1023 431 1089 447
rect 1041 409 1071 431
rect 1137 409 1167 435
rect -1167 87 -1137 109
rect -1185 71 -1119 87
rect -1071 83 -1041 109
rect -975 87 -945 109
rect -1185 37 -1169 71
rect -1135 37 -1119 71
rect -1185 21 -1119 37
rect -993 71 -927 87
rect -879 83 -849 109
rect -783 87 -753 109
rect -993 37 -977 71
rect -943 37 -927 71
rect -993 21 -927 37
rect -801 71 -735 87
rect -687 83 -657 109
rect -591 87 -561 109
rect -801 37 -785 71
rect -751 37 -735 71
rect -801 21 -735 37
rect -609 71 -543 87
rect -495 83 -465 109
rect -399 87 -369 109
rect -609 37 -593 71
rect -559 37 -543 71
rect -609 21 -543 37
rect -417 71 -351 87
rect -303 83 -273 109
rect -207 87 -177 109
rect -417 37 -401 71
rect -367 37 -351 71
rect -417 21 -351 37
rect -225 71 -159 87
rect -111 83 -81 109
rect -15 87 15 109
rect -225 37 -209 71
rect -175 37 -159 71
rect -225 21 -159 37
rect -33 71 33 87
rect 81 83 111 109
rect 177 87 207 109
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 159 71 225 87
rect 273 83 303 109
rect 369 87 399 109
rect 159 37 175 71
rect 209 37 225 71
rect 159 21 225 37
rect 351 71 417 87
rect 465 83 495 109
rect 561 87 591 109
rect 351 37 367 71
rect 401 37 417 71
rect 351 21 417 37
rect 543 71 609 87
rect 657 83 687 109
rect 753 87 783 109
rect 543 37 559 71
rect 593 37 609 71
rect 543 21 609 37
rect 735 71 801 87
rect 849 83 879 109
rect 945 87 975 109
rect 735 37 751 71
rect 785 37 801 71
rect 735 21 801 37
rect 927 71 993 87
rect 1041 83 1071 109
rect 1137 87 1167 109
rect 927 37 943 71
rect 977 37 993 71
rect 927 21 993 37
rect 1119 71 1185 87
rect 1119 37 1135 71
rect 1169 37 1185 71
rect 1119 21 1185 37
rect -1185 -37 -1119 -21
rect -1185 -71 -1169 -37
rect -1135 -71 -1119 -37
rect -1185 -87 -1119 -71
rect -993 -37 -927 -21
rect -993 -71 -977 -37
rect -943 -71 -927 -37
rect -1167 -109 -1137 -87
rect -1071 -109 -1041 -83
rect -993 -87 -927 -71
rect -801 -37 -735 -21
rect -801 -71 -785 -37
rect -751 -71 -735 -37
rect -975 -109 -945 -87
rect -879 -109 -849 -83
rect -801 -87 -735 -71
rect -609 -37 -543 -21
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -783 -109 -753 -87
rect -687 -109 -657 -83
rect -609 -87 -543 -71
rect -417 -37 -351 -21
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -591 -109 -561 -87
rect -495 -109 -465 -83
rect -417 -87 -351 -71
rect -225 -37 -159 -21
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -399 -109 -369 -87
rect -303 -109 -273 -83
rect -225 -87 -159 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -207 -109 -177 -87
rect -111 -109 -81 -83
rect -33 -87 33 -71
rect 159 -37 225 -21
rect 159 -71 175 -37
rect 209 -71 225 -37
rect -15 -109 15 -87
rect 81 -109 111 -83
rect 159 -87 225 -71
rect 351 -37 417 -21
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 177 -109 207 -87
rect 273 -109 303 -83
rect 351 -87 417 -71
rect 543 -37 609 -21
rect 543 -71 559 -37
rect 593 -71 609 -37
rect 369 -109 399 -87
rect 465 -109 495 -83
rect 543 -87 609 -71
rect 735 -37 801 -21
rect 735 -71 751 -37
rect 785 -71 801 -37
rect 561 -109 591 -87
rect 657 -109 687 -83
rect 735 -87 801 -71
rect 927 -37 993 -21
rect 927 -71 943 -37
rect 977 -71 993 -37
rect 753 -109 783 -87
rect 849 -109 879 -83
rect 927 -87 993 -71
rect 1119 -37 1185 -21
rect 1119 -71 1135 -37
rect 1169 -71 1185 -37
rect 945 -109 975 -87
rect 1041 -109 1071 -83
rect 1119 -87 1185 -71
rect 1137 -109 1167 -87
rect -1167 -435 -1137 -409
rect -1071 -431 -1041 -409
rect -1089 -447 -1023 -431
rect -975 -435 -945 -409
rect -879 -431 -849 -409
rect -1089 -481 -1073 -447
rect -1039 -481 -1023 -447
rect -1089 -497 -1023 -481
rect -897 -447 -831 -431
rect -783 -435 -753 -409
rect -687 -431 -657 -409
rect -897 -481 -881 -447
rect -847 -481 -831 -447
rect -897 -497 -831 -481
rect -705 -447 -639 -431
rect -591 -435 -561 -409
rect -495 -431 -465 -409
rect -705 -481 -689 -447
rect -655 -481 -639 -447
rect -705 -497 -639 -481
rect -513 -447 -447 -431
rect -399 -435 -369 -409
rect -303 -431 -273 -409
rect -513 -481 -497 -447
rect -463 -481 -447 -447
rect -513 -497 -447 -481
rect -321 -447 -255 -431
rect -207 -435 -177 -409
rect -111 -431 -81 -409
rect -321 -481 -305 -447
rect -271 -481 -255 -447
rect -321 -497 -255 -481
rect -129 -447 -63 -431
rect -15 -435 15 -409
rect 81 -431 111 -409
rect -129 -481 -113 -447
rect -79 -481 -63 -447
rect -129 -497 -63 -481
rect 63 -447 129 -431
rect 177 -435 207 -409
rect 273 -431 303 -409
rect 63 -481 79 -447
rect 113 -481 129 -447
rect 63 -497 129 -481
rect 255 -447 321 -431
rect 369 -435 399 -409
rect 465 -431 495 -409
rect 255 -481 271 -447
rect 305 -481 321 -447
rect 255 -497 321 -481
rect 447 -447 513 -431
rect 561 -435 591 -409
rect 657 -431 687 -409
rect 447 -481 463 -447
rect 497 -481 513 -447
rect 447 -497 513 -481
rect 639 -447 705 -431
rect 753 -435 783 -409
rect 849 -431 879 -409
rect 639 -481 655 -447
rect 689 -481 705 -447
rect 639 -497 705 -481
rect 831 -447 897 -431
rect 945 -435 975 -409
rect 1041 -431 1071 -409
rect 831 -481 847 -447
rect 881 -481 897 -447
rect 831 -497 897 -481
rect 1023 -447 1089 -431
rect 1137 -435 1167 -409
rect 1023 -481 1039 -447
rect 1073 -481 1089 -447
rect 1023 -497 1089 -481
rect -1089 -555 -1023 -539
rect -1089 -589 -1073 -555
rect -1039 -589 -1023 -555
rect -1167 -627 -1137 -601
rect -1089 -605 -1023 -589
rect -897 -555 -831 -539
rect -897 -589 -881 -555
rect -847 -589 -831 -555
rect -1071 -627 -1041 -605
rect -975 -627 -945 -601
rect -897 -605 -831 -589
rect -705 -555 -639 -539
rect -705 -589 -689 -555
rect -655 -589 -639 -555
rect -879 -627 -849 -605
rect -783 -627 -753 -601
rect -705 -605 -639 -589
rect -513 -555 -447 -539
rect -513 -589 -497 -555
rect -463 -589 -447 -555
rect -687 -627 -657 -605
rect -591 -627 -561 -601
rect -513 -605 -447 -589
rect -321 -555 -255 -539
rect -321 -589 -305 -555
rect -271 -589 -255 -555
rect -495 -627 -465 -605
rect -399 -627 -369 -601
rect -321 -605 -255 -589
rect -129 -555 -63 -539
rect -129 -589 -113 -555
rect -79 -589 -63 -555
rect -303 -627 -273 -605
rect -207 -627 -177 -601
rect -129 -605 -63 -589
rect 63 -555 129 -539
rect 63 -589 79 -555
rect 113 -589 129 -555
rect -111 -627 -81 -605
rect -15 -627 15 -601
rect 63 -605 129 -589
rect 255 -555 321 -539
rect 255 -589 271 -555
rect 305 -589 321 -555
rect 81 -627 111 -605
rect 177 -627 207 -601
rect 255 -605 321 -589
rect 447 -555 513 -539
rect 447 -589 463 -555
rect 497 -589 513 -555
rect 273 -627 303 -605
rect 369 -627 399 -601
rect 447 -605 513 -589
rect 639 -555 705 -539
rect 639 -589 655 -555
rect 689 -589 705 -555
rect 465 -627 495 -605
rect 561 -627 591 -601
rect 639 -605 705 -589
rect 831 -555 897 -539
rect 831 -589 847 -555
rect 881 -589 897 -555
rect 657 -627 687 -605
rect 753 -627 783 -601
rect 831 -605 897 -589
rect 1023 -555 1089 -539
rect 1023 -589 1039 -555
rect 1073 -589 1089 -555
rect 849 -627 879 -605
rect 945 -627 975 -601
rect 1023 -605 1089 -589
rect 1041 -627 1071 -605
rect 1137 -627 1167 -601
rect -1167 -949 -1137 -927
rect -1185 -965 -1119 -949
rect -1071 -953 -1041 -927
rect -975 -949 -945 -927
rect -1185 -999 -1169 -965
rect -1135 -999 -1119 -965
rect -1185 -1015 -1119 -999
rect -993 -965 -927 -949
rect -879 -953 -849 -927
rect -783 -949 -753 -927
rect -993 -999 -977 -965
rect -943 -999 -927 -965
rect -993 -1015 -927 -999
rect -801 -965 -735 -949
rect -687 -953 -657 -927
rect -591 -949 -561 -927
rect -801 -999 -785 -965
rect -751 -999 -735 -965
rect -801 -1015 -735 -999
rect -609 -965 -543 -949
rect -495 -953 -465 -927
rect -399 -949 -369 -927
rect -609 -999 -593 -965
rect -559 -999 -543 -965
rect -609 -1015 -543 -999
rect -417 -965 -351 -949
rect -303 -953 -273 -927
rect -207 -949 -177 -927
rect -417 -999 -401 -965
rect -367 -999 -351 -965
rect -417 -1015 -351 -999
rect -225 -965 -159 -949
rect -111 -953 -81 -927
rect -15 -949 15 -927
rect -225 -999 -209 -965
rect -175 -999 -159 -965
rect -225 -1015 -159 -999
rect -33 -965 33 -949
rect 81 -953 111 -927
rect 177 -949 207 -927
rect -33 -999 -17 -965
rect 17 -999 33 -965
rect -33 -1015 33 -999
rect 159 -965 225 -949
rect 273 -953 303 -927
rect 369 -949 399 -927
rect 159 -999 175 -965
rect 209 -999 225 -965
rect 159 -1015 225 -999
rect 351 -965 417 -949
rect 465 -953 495 -927
rect 561 -949 591 -927
rect 351 -999 367 -965
rect 401 -999 417 -965
rect 351 -1015 417 -999
rect 543 -965 609 -949
rect 657 -953 687 -927
rect 753 -949 783 -927
rect 543 -999 559 -965
rect 593 -999 609 -965
rect 543 -1015 609 -999
rect 735 -965 801 -949
rect 849 -953 879 -927
rect 945 -949 975 -927
rect 735 -999 751 -965
rect 785 -999 801 -965
rect 735 -1015 801 -999
rect 927 -965 993 -949
rect 1041 -953 1071 -927
rect 1137 -949 1167 -927
rect 927 -999 943 -965
rect 977 -999 993 -965
rect 927 -1015 993 -999
rect 1119 -965 1185 -949
rect 1119 -999 1135 -965
rect 1169 -999 1185 -965
rect 1119 -1015 1185 -999
<< polycont >>
rect -1169 965 -1135 999
rect -977 965 -943 999
rect -785 965 -751 999
rect -593 965 -559 999
rect -401 965 -367 999
rect -209 965 -175 999
rect -17 965 17 999
rect 175 965 209 999
rect 367 965 401 999
rect 559 965 593 999
rect 751 965 785 999
rect 943 965 977 999
rect 1135 965 1169 999
rect -1073 555 -1039 589
rect -881 555 -847 589
rect -689 555 -655 589
rect -497 555 -463 589
rect -305 555 -271 589
rect -113 555 -79 589
rect 79 555 113 589
rect 271 555 305 589
rect 463 555 497 589
rect 655 555 689 589
rect 847 555 881 589
rect 1039 555 1073 589
rect -1073 447 -1039 481
rect -881 447 -847 481
rect -689 447 -655 481
rect -497 447 -463 481
rect -305 447 -271 481
rect -113 447 -79 481
rect 79 447 113 481
rect 271 447 305 481
rect 463 447 497 481
rect 655 447 689 481
rect 847 447 881 481
rect 1039 447 1073 481
rect -1169 37 -1135 71
rect -977 37 -943 71
rect -785 37 -751 71
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect 751 37 785 71
rect 943 37 977 71
rect 1135 37 1169 71
rect -1169 -71 -1135 -37
rect -977 -71 -943 -37
rect -785 -71 -751 -37
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect 751 -71 785 -37
rect 943 -71 977 -37
rect 1135 -71 1169 -37
rect -1073 -481 -1039 -447
rect -881 -481 -847 -447
rect -689 -481 -655 -447
rect -497 -481 -463 -447
rect -305 -481 -271 -447
rect -113 -481 -79 -447
rect 79 -481 113 -447
rect 271 -481 305 -447
rect 463 -481 497 -447
rect 655 -481 689 -447
rect 847 -481 881 -447
rect 1039 -481 1073 -447
rect -1073 -589 -1039 -555
rect -881 -589 -847 -555
rect -689 -589 -655 -555
rect -497 -589 -463 -555
rect -305 -589 -271 -555
rect -113 -589 -79 -555
rect 79 -589 113 -555
rect 271 -589 305 -555
rect 463 -589 497 -555
rect 655 -589 689 -555
rect 847 -589 881 -555
rect 1039 -589 1073 -555
rect -1169 -999 -1135 -965
rect -977 -999 -943 -965
rect -785 -999 -751 -965
rect -593 -999 -559 -965
rect -401 -999 -367 -965
rect -209 -999 -175 -965
rect -17 -999 17 -965
rect 175 -999 209 -965
rect 367 -999 401 -965
rect 559 -999 593 -965
rect 751 -999 785 -965
rect 943 -999 977 -965
rect 1135 -999 1169 -965
<< locali >>
rect -1331 1067 -1235 1101
rect 1235 1067 1331 1101
rect -1331 1005 -1297 1067
rect 1297 1005 1331 1067
rect -1185 965 -1169 999
rect -1135 965 -1119 999
rect -993 965 -977 999
rect -943 965 -927 999
rect -801 965 -785 999
rect -751 965 -735 999
rect -609 965 -593 999
rect -559 965 -543 999
rect -417 965 -401 999
rect -367 965 -351 999
rect -225 965 -209 999
rect -175 965 -159 999
rect -33 965 -17 999
rect 17 965 33 999
rect 159 965 175 999
rect 209 965 225 999
rect 351 965 367 999
rect 401 965 417 999
rect 543 965 559 999
rect 593 965 609 999
rect 735 965 751 999
rect 785 965 801 999
rect 927 965 943 999
rect 977 965 993 999
rect 1119 965 1135 999
rect 1169 965 1185 999
rect -1217 915 -1183 931
rect -1217 623 -1183 639
rect -1121 915 -1087 931
rect -1121 623 -1087 639
rect -1025 915 -991 931
rect -1025 623 -991 639
rect -929 915 -895 931
rect -929 623 -895 639
rect -833 915 -799 931
rect -833 623 -799 639
rect -737 915 -703 931
rect -737 623 -703 639
rect -641 915 -607 931
rect -641 623 -607 639
rect -545 915 -511 931
rect -545 623 -511 639
rect -449 915 -415 931
rect -449 623 -415 639
rect -353 915 -319 931
rect -353 623 -319 639
rect -257 915 -223 931
rect -257 623 -223 639
rect -161 915 -127 931
rect -161 623 -127 639
rect -65 915 -31 931
rect -65 623 -31 639
rect 31 915 65 931
rect 31 623 65 639
rect 127 915 161 931
rect 127 623 161 639
rect 223 915 257 931
rect 223 623 257 639
rect 319 915 353 931
rect 319 623 353 639
rect 415 915 449 931
rect 415 623 449 639
rect 511 915 545 931
rect 511 623 545 639
rect 607 915 641 931
rect 607 623 641 639
rect 703 915 737 931
rect 703 623 737 639
rect 799 915 833 931
rect 799 623 833 639
rect 895 915 929 931
rect 895 623 929 639
rect 991 915 1025 931
rect 991 623 1025 639
rect 1087 915 1121 931
rect 1087 623 1121 639
rect 1183 915 1217 931
rect 1183 623 1217 639
rect -1089 555 -1073 589
rect -1039 555 -1023 589
rect -897 555 -881 589
rect -847 555 -831 589
rect -705 555 -689 589
rect -655 555 -639 589
rect -513 555 -497 589
rect -463 555 -447 589
rect -321 555 -305 589
rect -271 555 -255 589
rect -129 555 -113 589
rect -79 555 -63 589
rect 63 555 79 589
rect 113 555 129 589
rect 255 555 271 589
rect 305 555 321 589
rect 447 555 463 589
rect 497 555 513 589
rect 639 555 655 589
rect 689 555 705 589
rect 831 555 847 589
rect 881 555 897 589
rect 1023 555 1039 589
rect 1073 555 1089 589
rect -1089 447 -1073 481
rect -1039 447 -1023 481
rect -897 447 -881 481
rect -847 447 -831 481
rect -705 447 -689 481
rect -655 447 -639 481
rect -513 447 -497 481
rect -463 447 -447 481
rect -321 447 -305 481
rect -271 447 -255 481
rect -129 447 -113 481
rect -79 447 -63 481
rect 63 447 79 481
rect 113 447 129 481
rect 255 447 271 481
rect 305 447 321 481
rect 447 447 463 481
rect 497 447 513 481
rect 639 447 655 481
rect 689 447 705 481
rect 831 447 847 481
rect 881 447 897 481
rect 1023 447 1039 481
rect 1073 447 1089 481
rect -1217 397 -1183 413
rect -1217 105 -1183 121
rect -1121 397 -1087 413
rect -1121 105 -1087 121
rect -1025 397 -991 413
rect -1025 105 -991 121
rect -929 397 -895 413
rect -929 105 -895 121
rect -833 397 -799 413
rect -833 105 -799 121
rect -737 397 -703 413
rect -737 105 -703 121
rect -641 397 -607 413
rect -641 105 -607 121
rect -545 397 -511 413
rect -545 105 -511 121
rect -449 397 -415 413
rect -449 105 -415 121
rect -353 397 -319 413
rect -353 105 -319 121
rect -257 397 -223 413
rect -257 105 -223 121
rect -161 397 -127 413
rect -161 105 -127 121
rect -65 397 -31 413
rect -65 105 -31 121
rect 31 397 65 413
rect 31 105 65 121
rect 127 397 161 413
rect 127 105 161 121
rect 223 397 257 413
rect 223 105 257 121
rect 319 397 353 413
rect 319 105 353 121
rect 415 397 449 413
rect 415 105 449 121
rect 511 397 545 413
rect 511 105 545 121
rect 607 397 641 413
rect 607 105 641 121
rect 703 397 737 413
rect 703 105 737 121
rect 799 397 833 413
rect 799 105 833 121
rect 895 397 929 413
rect 895 105 929 121
rect 991 397 1025 413
rect 991 105 1025 121
rect 1087 397 1121 413
rect 1087 105 1121 121
rect 1183 397 1217 413
rect 1183 105 1217 121
rect -1185 37 -1169 71
rect -1135 37 -1119 71
rect -993 37 -977 71
rect -943 37 -927 71
rect -801 37 -785 71
rect -751 37 -735 71
rect -609 37 -593 71
rect -559 37 -543 71
rect -417 37 -401 71
rect -367 37 -351 71
rect -225 37 -209 71
rect -175 37 -159 71
rect -33 37 -17 71
rect 17 37 33 71
rect 159 37 175 71
rect 209 37 225 71
rect 351 37 367 71
rect 401 37 417 71
rect 543 37 559 71
rect 593 37 609 71
rect 735 37 751 71
rect 785 37 801 71
rect 927 37 943 71
rect 977 37 993 71
rect 1119 37 1135 71
rect 1169 37 1185 71
rect -1185 -71 -1169 -37
rect -1135 -71 -1119 -37
rect -993 -71 -977 -37
rect -943 -71 -927 -37
rect -801 -71 -785 -37
rect -751 -71 -735 -37
rect -609 -71 -593 -37
rect -559 -71 -543 -37
rect -417 -71 -401 -37
rect -367 -71 -351 -37
rect -225 -71 -209 -37
rect -175 -71 -159 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 159 -71 175 -37
rect 209 -71 225 -37
rect 351 -71 367 -37
rect 401 -71 417 -37
rect 543 -71 559 -37
rect 593 -71 609 -37
rect 735 -71 751 -37
rect 785 -71 801 -37
rect 927 -71 943 -37
rect 977 -71 993 -37
rect 1119 -71 1135 -37
rect 1169 -71 1185 -37
rect -1217 -121 -1183 -105
rect -1217 -413 -1183 -397
rect -1121 -121 -1087 -105
rect -1121 -413 -1087 -397
rect -1025 -121 -991 -105
rect -1025 -413 -991 -397
rect -929 -121 -895 -105
rect -929 -413 -895 -397
rect -833 -121 -799 -105
rect -833 -413 -799 -397
rect -737 -121 -703 -105
rect -737 -413 -703 -397
rect -641 -121 -607 -105
rect -641 -413 -607 -397
rect -545 -121 -511 -105
rect -545 -413 -511 -397
rect -449 -121 -415 -105
rect -449 -413 -415 -397
rect -353 -121 -319 -105
rect -353 -413 -319 -397
rect -257 -121 -223 -105
rect -257 -413 -223 -397
rect -161 -121 -127 -105
rect -161 -413 -127 -397
rect -65 -121 -31 -105
rect -65 -413 -31 -397
rect 31 -121 65 -105
rect 31 -413 65 -397
rect 127 -121 161 -105
rect 127 -413 161 -397
rect 223 -121 257 -105
rect 223 -413 257 -397
rect 319 -121 353 -105
rect 319 -413 353 -397
rect 415 -121 449 -105
rect 415 -413 449 -397
rect 511 -121 545 -105
rect 511 -413 545 -397
rect 607 -121 641 -105
rect 607 -413 641 -397
rect 703 -121 737 -105
rect 703 -413 737 -397
rect 799 -121 833 -105
rect 799 -413 833 -397
rect 895 -121 929 -105
rect 895 -413 929 -397
rect 991 -121 1025 -105
rect 991 -413 1025 -397
rect 1087 -121 1121 -105
rect 1087 -413 1121 -397
rect 1183 -121 1217 -105
rect 1183 -413 1217 -397
rect -1089 -481 -1073 -447
rect -1039 -481 -1023 -447
rect -897 -481 -881 -447
rect -847 -481 -831 -447
rect -705 -481 -689 -447
rect -655 -481 -639 -447
rect -513 -481 -497 -447
rect -463 -481 -447 -447
rect -321 -481 -305 -447
rect -271 -481 -255 -447
rect -129 -481 -113 -447
rect -79 -481 -63 -447
rect 63 -481 79 -447
rect 113 -481 129 -447
rect 255 -481 271 -447
rect 305 -481 321 -447
rect 447 -481 463 -447
rect 497 -481 513 -447
rect 639 -481 655 -447
rect 689 -481 705 -447
rect 831 -481 847 -447
rect 881 -481 897 -447
rect 1023 -481 1039 -447
rect 1073 -481 1089 -447
rect -1089 -589 -1073 -555
rect -1039 -589 -1023 -555
rect -897 -589 -881 -555
rect -847 -589 -831 -555
rect -705 -589 -689 -555
rect -655 -589 -639 -555
rect -513 -589 -497 -555
rect -463 -589 -447 -555
rect -321 -589 -305 -555
rect -271 -589 -255 -555
rect -129 -589 -113 -555
rect -79 -589 -63 -555
rect 63 -589 79 -555
rect 113 -589 129 -555
rect 255 -589 271 -555
rect 305 -589 321 -555
rect 447 -589 463 -555
rect 497 -589 513 -555
rect 639 -589 655 -555
rect 689 -589 705 -555
rect 831 -589 847 -555
rect 881 -589 897 -555
rect 1023 -589 1039 -555
rect 1073 -589 1089 -555
rect -1217 -639 -1183 -623
rect -1217 -931 -1183 -915
rect -1121 -639 -1087 -623
rect -1121 -931 -1087 -915
rect -1025 -639 -991 -623
rect -1025 -931 -991 -915
rect -929 -639 -895 -623
rect -929 -931 -895 -915
rect -833 -639 -799 -623
rect -833 -931 -799 -915
rect -737 -639 -703 -623
rect -737 -931 -703 -915
rect -641 -639 -607 -623
rect -641 -931 -607 -915
rect -545 -639 -511 -623
rect -545 -931 -511 -915
rect -449 -639 -415 -623
rect -449 -931 -415 -915
rect -353 -639 -319 -623
rect -353 -931 -319 -915
rect -257 -639 -223 -623
rect -257 -931 -223 -915
rect -161 -639 -127 -623
rect -161 -931 -127 -915
rect -65 -639 -31 -623
rect -65 -931 -31 -915
rect 31 -639 65 -623
rect 31 -931 65 -915
rect 127 -639 161 -623
rect 127 -931 161 -915
rect 223 -639 257 -623
rect 223 -931 257 -915
rect 319 -639 353 -623
rect 319 -931 353 -915
rect 415 -639 449 -623
rect 415 -931 449 -915
rect 511 -639 545 -623
rect 511 -931 545 -915
rect 607 -639 641 -623
rect 607 -931 641 -915
rect 703 -639 737 -623
rect 703 -931 737 -915
rect 799 -639 833 -623
rect 799 -931 833 -915
rect 895 -639 929 -623
rect 895 -931 929 -915
rect 991 -639 1025 -623
rect 991 -931 1025 -915
rect 1087 -639 1121 -623
rect 1087 -931 1121 -915
rect 1183 -639 1217 -623
rect 1183 -931 1217 -915
rect -1185 -999 -1169 -965
rect -1135 -999 -1119 -965
rect -993 -999 -977 -965
rect -943 -999 -927 -965
rect -801 -999 -785 -965
rect -751 -999 -735 -965
rect -609 -999 -593 -965
rect -559 -999 -543 -965
rect -417 -999 -401 -965
rect -367 -999 -351 -965
rect -225 -999 -209 -965
rect -175 -999 -159 -965
rect -33 -999 -17 -965
rect 17 -999 33 -965
rect 159 -999 175 -965
rect 209 -999 225 -965
rect 351 -999 367 -965
rect 401 -999 417 -965
rect 543 -999 559 -965
rect 593 -999 609 -965
rect 735 -999 751 -965
rect 785 -999 801 -965
rect 927 -999 943 -965
rect 977 -999 993 -965
rect 1119 -999 1135 -965
rect 1169 -999 1185 -965
rect -1331 -1067 -1297 -1005
rect 1297 -1067 1331 -1005
rect -1331 -1101 -1235 -1067
rect 1235 -1101 1331 -1067
<< viali >>
rect -1169 965 -1135 999
rect -977 965 -943 999
rect -785 965 -751 999
rect -593 965 -559 999
rect -401 965 -367 999
rect -209 965 -175 999
rect -17 965 17 999
rect 175 965 209 999
rect 367 965 401 999
rect 559 965 593 999
rect 751 965 785 999
rect 943 965 977 999
rect 1135 965 1169 999
rect -1217 639 -1183 915
rect -1121 639 -1087 915
rect -1025 639 -991 915
rect -929 639 -895 915
rect -833 639 -799 915
rect -737 639 -703 915
rect -641 639 -607 915
rect -545 639 -511 915
rect -449 639 -415 915
rect -353 639 -319 915
rect -257 639 -223 915
rect -161 639 -127 915
rect -65 639 -31 915
rect 31 639 65 915
rect 127 639 161 915
rect 223 639 257 915
rect 319 639 353 915
rect 415 639 449 915
rect 511 639 545 915
rect 607 639 641 915
rect 703 639 737 915
rect 799 639 833 915
rect 895 639 929 915
rect 991 639 1025 915
rect 1087 639 1121 915
rect 1183 639 1217 915
rect -1073 555 -1039 589
rect -881 555 -847 589
rect -689 555 -655 589
rect -497 555 -463 589
rect -305 555 -271 589
rect -113 555 -79 589
rect 79 555 113 589
rect 271 555 305 589
rect 463 555 497 589
rect 655 555 689 589
rect 847 555 881 589
rect 1039 555 1073 589
rect -1073 447 -1039 481
rect -881 447 -847 481
rect -689 447 -655 481
rect -497 447 -463 481
rect -305 447 -271 481
rect -113 447 -79 481
rect 79 447 113 481
rect 271 447 305 481
rect 463 447 497 481
rect 655 447 689 481
rect 847 447 881 481
rect 1039 447 1073 481
rect -1217 121 -1183 397
rect -1121 121 -1087 397
rect -1025 121 -991 397
rect -929 121 -895 397
rect -833 121 -799 397
rect -737 121 -703 397
rect -641 121 -607 397
rect -545 121 -511 397
rect -449 121 -415 397
rect -353 121 -319 397
rect -257 121 -223 397
rect -161 121 -127 397
rect -65 121 -31 397
rect 31 121 65 397
rect 127 121 161 397
rect 223 121 257 397
rect 319 121 353 397
rect 415 121 449 397
rect 511 121 545 397
rect 607 121 641 397
rect 703 121 737 397
rect 799 121 833 397
rect 895 121 929 397
rect 991 121 1025 397
rect 1087 121 1121 397
rect 1183 121 1217 397
rect -1169 37 -1135 71
rect -977 37 -943 71
rect -785 37 -751 71
rect -593 37 -559 71
rect -401 37 -367 71
rect -209 37 -175 71
rect -17 37 17 71
rect 175 37 209 71
rect 367 37 401 71
rect 559 37 593 71
rect 751 37 785 71
rect 943 37 977 71
rect 1135 37 1169 71
rect -1169 -71 -1135 -37
rect -977 -71 -943 -37
rect -785 -71 -751 -37
rect -593 -71 -559 -37
rect -401 -71 -367 -37
rect -209 -71 -175 -37
rect -17 -71 17 -37
rect 175 -71 209 -37
rect 367 -71 401 -37
rect 559 -71 593 -37
rect 751 -71 785 -37
rect 943 -71 977 -37
rect 1135 -71 1169 -37
rect -1217 -397 -1183 -121
rect -1121 -397 -1087 -121
rect -1025 -397 -991 -121
rect -929 -397 -895 -121
rect -833 -397 -799 -121
rect -737 -397 -703 -121
rect -641 -397 -607 -121
rect -545 -397 -511 -121
rect -449 -397 -415 -121
rect -353 -397 -319 -121
rect -257 -397 -223 -121
rect -161 -397 -127 -121
rect -65 -397 -31 -121
rect 31 -397 65 -121
rect 127 -397 161 -121
rect 223 -397 257 -121
rect 319 -397 353 -121
rect 415 -397 449 -121
rect 511 -397 545 -121
rect 607 -397 641 -121
rect 703 -397 737 -121
rect 799 -397 833 -121
rect 895 -397 929 -121
rect 991 -397 1025 -121
rect 1087 -397 1121 -121
rect 1183 -397 1217 -121
rect -1073 -481 -1039 -447
rect -881 -481 -847 -447
rect -689 -481 -655 -447
rect -497 -481 -463 -447
rect -305 -481 -271 -447
rect -113 -481 -79 -447
rect 79 -481 113 -447
rect 271 -481 305 -447
rect 463 -481 497 -447
rect 655 -481 689 -447
rect 847 -481 881 -447
rect 1039 -481 1073 -447
rect -1073 -589 -1039 -555
rect -881 -589 -847 -555
rect -689 -589 -655 -555
rect -497 -589 -463 -555
rect -305 -589 -271 -555
rect -113 -589 -79 -555
rect 79 -589 113 -555
rect 271 -589 305 -555
rect 463 -589 497 -555
rect 655 -589 689 -555
rect 847 -589 881 -555
rect 1039 -589 1073 -555
rect -1217 -915 -1183 -639
rect -1121 -915 -1087 -639
rect -1025 -915 -991 -639
rect -929 -915 -895 -639
rect -833 -915 -799 -639
rect -737 -915 -703 -639
rect -641 -915 -607 -639
rect -545 -915 -511 -639
rect -449 -915 -415 -639
rect -353 -915 -319 -639
rect -257 -915 -223 -639
rect -161 -915 -127 -639
rect -65 -915 -31 -639
rect 31 -915 65 -639
rect 127 -915 161 -639
rect 223 -915 257 -639
rect 319 -915 353 -639
rect 415 -915 449 -639
rect 511 -915 545 -639
rect 607 -915 641 -639
rect 703 -915 737 -639
rect 799 -915 833 -639
rect 895 -915 929 -639
rect 991 -915 1025 -639
rect 1087 -915 1121 -639
rect 1183 -915 1217 -639
rect -1169 -999 -1135 -965
rect -977 -999 -943 -965
rect -785 -999 -751 -965
rect -593 -999 -559 -965
rect -401 -999 -367 -965
rect -209 -999 -175 -965
rect -17 -999 17 -965
rect 175 -999 209 -965
rect 367 -999 401 -965
rect 559 -999 593 -965
rect 751 -999 785 -965
rect 943 -999 977 -965
rect 1135 -999 1169 -965
<< metal1 >>
rect -1181 999 -1123 1005
rect -1181 965 -1169 999
rect -1135 965 -1123 999
rect -1181 959 -1123 965
rect -989 999 -931 1005
rect -989 965 -977 999
rect -943 965 -931 999
rect -989 959 -931 965
rect -797 999 -739 1005
rect -797 965 -785 999
rect -751 965 -739 999
rect -797 959 -739 965
rect -605 999 -547 1005
rect -605 965 -593 999
rect -559 965 -547 999
rect -605 959 -547 965
rect -413 999 -355 1005
rect -413 965 -401 999
rect -367 965 -355 999
rect -413 959 -355 965
rect -221 999 -163 1005
rect -221 965 -209 999
rect -175 965 -163 999
rect -221 959 -163 965
rect -29 999 29 1005
rect -29 965 -17 999
rect 17 965 29 999
rect -29 959 29 965
rect 163 999 221 1005
rect 163 965 175 999
rect 209 965 221 999
rect 163 959 221 965
rect 355 999 413 1005
rect 355 965 367 999
rect 401 965 413 999
rect 355 959 413 965
rect 547 999 605 1005
rect 547 965 559 999
rect 593 965 605 999
rect 547 959 605 965
rect 739 999 797 1005
rect 739 965 751 999
rect 785 965 797 999
rect 739 959 797 965
rect 931 999 989 1005
rect 931 965 943 999
rect 977 965 989 999
rect 931 959 989 965
rect 1123 999 1181 1005
rect 1123 965 1135 999
rect 1169 965 1181 999
rect 1123 959 1181 965
rect -1223 915 -1177 927
rect -1223 639 -1217 915
rect -1183 639 -1177 915
rect -1223 627 -1177 639
rect -1127 915 -1081 927
rect -1127 639 -1121 915
rect -1087 639 -1081 915
rect -1127 627 -1081 639
rect -1031 915 -985 927
rect -1031 639 -1025 915
rect -991 639 -985 915
rect -1031 627 -985 639
rect -935 915 -889 927
rect -935 639 -929 915
rect -895 639 -889 915
rect -935 627 -889 639
rect -839 915 -793 927
rect -839 639 -833 915
rect -799 639 -793 915
rect -839 627 -793 639
rect -743 915 -697 927
rect -743 639 -737 915
rect -703 639 -697 915
rect -743 627 -697 639
rect -647 915 -601 927
rect -647 639 -641 915
rect -607 639 -601 915
rect -647 627 -601 639
rect -551 915 -505 927
rect -551 639 -545 915
rect -511 639 -505 915
rect -551 627 -505 639
rect -455 915 -409 927
rect -455 639 -449 915
rect -415 639 -409 915
rect -455 627 -409 639
rect -359 915 -313 927
rect -359 639 -353 915
rect -319 639 -313 915
rect -359 627 -313 639
rect -263 915 -217 927
rect -263 639 -257 915
rect -223 639 -217 915
rect -263 627 -217 639
rect -167 915 -121 927
rect -167 639 -161 915
rect -127 639 -121 915
rect -167 627 -121 639
rect -71 915 -25 927
rect -71 639 -65 915
rect -31 639 -25 915
rect -71 627 -25 639
rect 25 915 71 927
rect 25 639 31 915
rect 65 639 71 915
rect 25 627 71 639
rect 121 915 167 927
rect 121 639 127 915
rect 161 639 167 915
rect 121 627 167 639
rect 217 915 263 927
rect 217 639 223 915
rect 257 639 263 915
rect 217 627 263 639
rect 313 915 359 927
rect 313 639 319 915
rect 353 639 359 915
rect 313 627 359 639
rect 409 915 455 927
rect 409 639 415 915
rect 449 639 455 915
rect 409 627 455 639
rect 505 915 551 927
rect 505 639 511 915
rect 545 639 551 915
rect 505 627 551 639
rect 601 915 647 927
rect 601 639 607 915
rect 641 639 647 915
rect 601 627 647 639
rect 697 915 743 927
rect 697 639 703 915
rect 737 639 743 915
rect 697 627 743 639
rect 793 915 839 927
rect 793 639 799 915
rect 833 639 839 915
rect 793 627 839 639
rect 889 915 935 927
rect 889 639 895 915
rect 929 639 935 915
rect 889 627 935 639
rect 985 915 1031 927
rect 985 639 991 915
rect 1025 639 1031 915
rect 985 627 1031 639
rect 1081 915 1127 927
rect 1081 639 1087 915
rect 1121 639 1127 915
rect 1081 627 1127 639
rect 1177 915 1223 927
rect 1177 639 1183 915
rect 1217 639 1223 915
rect 1177 627 1223 639
rect -1085 589 -1027 595
rect -1085 555 -1073 589
rect -1039 555 -1027 589
rect -1085 549 -1027 555
rect -893 589 -835 595
rect -893 555 -881 589
rect -847 555 -835 589
rect -893 549 -835 555
rect -701 589 -643 595
rect -701 555 -689 589
rect -655 555 -643 589
rect -701 549 -643 555
rect -509 589 -451 595
rect -509 555 -497 589
rect -463 555 -451 589
rect -509 549 -451 555
rect -317 589 -259 595
rect -317 555 -305 589
rect -271 555 -259 589
rect -317 549 -259 555
rect -125 589 -67 595
rect -125 555 -113 589
rect -79 555 -67 589
rect -125 549 -67 555
rect 67 589 125 595
rect 67 555 79 589
rect 113 555 125 589
rect 67 549 125 555
rect 259 589 317 595
rect 259 555 271 589
rect 305 555 317 589
rect 259 549 317 555
rect 451 589 509 595
rect 451 555 463 589
rect 497 555 509 589
rect 451 549 509 555
rect 643 589 701 595
rect 643 555 655 589
rect 689 555 701 589
rect 643 549 701 555
rect 835 589 893 595
rect 835 555 847 589
rect 881 555 893 589
rect 835 549 893 555
rect 1027 589 1085 595
rect 1027 555 1039 589
rect 1073 555 1085 589
rect 1027 549 1085 555
rect -1085 481 -1027 487
rect -1085 447 -1073 481
rect -1039 447 -1027 481
rect -1085 441 -1027 447
rect -893 481 -835 487
rect -893 447 -881 481
rect -847 447 -835 481
rect -893 441 -835 447
rect -701 481 -643 487
rect -701 447 -689 481
rect -655 447 -643 481
rect -701 441 -643 447
rect -509 481 -451 487
rect -509 447 -497 481
rect -463 447 -451 481
rect -509 441 -451 447
rect -317 481 -259 487
rect -317 447 -305 481
rect -271 447 -259 481
rect -317 441 -259 447
rect -125 481 -67 487
rect -125 447 -113 481
rect -79 447 -67 481
rect -125 441 -67 447
rect 67 481 125 487
rect 67 447 79 481
rect 113 447 125 481
rect 67 441 125 447
rect 259 481 317 487
rect 259 447 271 481
rect 305 447 317 481
rect 259 441 317 447
rect 451 481 509 487
rect 451 447 463 481
rect 497 447 509 481
rect 451 441 509 447
rect 643 481 701 487
rect 643 447 655 481
rect 689 447 701 481
rect 643 441 701 447
rect 835 481 893 487
rect 835 447 847 481
rect 881 447 893 481
rect 835 441 893 447
rect 1027 481 1085 487
rect 1027 447 1039 481
rect 1073 447 1085 481
rect 1027 441 1085 447
rect -1223 397 -1177 409
rect -1223 121 -1217 397
rect -1183 121 -1177 397
rect -1223 109 -1177 121
rect -1127 397 -1081 409
rect -1127 121 -1121 397
rect -1087 121 -1081 397
rect -1127 109 -1081 121
rect -1031 397 -985 409
rect -1031 121 -1025 397
rect -991 121 -985 397
rect -1031 109 -985 121
rect -935 397 -889 409
rect -935 121 -929 397
rect -895 121 -889 397
rect -935 109 -889 121
rect -839 397 -793 409
rect -839 121 -833 397
rect -799 121 -793 397
rect -839 109 -793 121
rect -743 397 -697 409
rect -743 121 -737 397
rect -703 121 -697 397
rect -743 109 -697 121
rect -647 397 -601 409
rect -647 121 -641 397
rect -607 121 -601 397
rect -647 109 -601 121
rect -551 397 -505 409
rect -551 121 -545 397
rect -511 121 -505 397
rect -551 109 -505 121
rect -455 397 -409 409
rect -455 121 -449 397
rect -415 121 -409 397
rect -455 109 -409 121
rect -359 397 -313 409
rect -359 121 -353 397
rect -319 121 -313 397
rect -359 109 -313 121
rect -263 397 -217 409
rect -263 121 -257 397
rect -223 121 -217 397
rect -263 109 -217 121
rect -167 397 -121 409
rect -167 121 -161 397
rect -127 121 -121 397
rect -167 109 -121 121
rect -71 397 -25 409
rect -71 121 -65 397
rect -31 121 -25 397
rect -71 109 -25 121
rect 25 397 71 409
rect 25 121 31 397
rect 65 121 71 397
rect 25 109 71 121
rect 121 397 167 409
rect 121 121 127 397
rect 161 121 167 397
rect 121 109 167 121
rect 217 397 263 409
rect 217 121 223 397
rect 257 121 263 397
rect 217 109 263 121
rect 313 397 359 409
rect 313 121 319 397
rect 353 121 359 397
rect 313 109 359 121
rect 409 397 455 409
rect 409 121 415 397
rect 449 121 455 397
rect 409 109 455 121
rect 505 397 551 409
rect 505 121 511 397
rect 545 121 551 397
rect 505 109 551 121
rect 601 397 647 409
rect 601 121 607 397
rect 641 121 647 397
rect 601 109 647 121
rect 697 397 743 409
rect 697 121 703 397
rect 737 121 743 397
rect 697 109 743 121
rect 793 397 839 409
rect 793 121 799 397
rect 833 121 839 397
rect 793 109 839 121
rect 889 397 935 409
rect 889 121 895 397
rect 929 121 935 397
rect 889 109 935 121
rect 985 397 1031 409
rect 985 121 991 397
rect 1025 121 1031 397
rect 985 109 1031 121
rect 1081 397 1127 409
rect 1081 121 1087 397
rect 1121 121 1127 397
rect 1081 109 1127 121
rect 1177 397 1223 409
rect 1177 121 1183 397
rect 1217 121 1223 397
rect 1177 109 1223 121
rect -1181 71 -1123 77
rect -1181 37 -1169 71
rect -1135 37 -1123 71
rect -1181 31 -1123 37
rect -989 71 -931 77
rect -989 37 -977 71
rect -943 37 -931 71
rect -989 31 -931 37
rect -797 71 -739 77
rect -797 37 -785 71
rect -751 37 -739 71
rect -797 31 -739 37
rect -605 71 -547 77
rect -605 37 -593 71
rect -559 37 -547 71
rect -605 31 -547 37
rect -413 71 -355 77
rect -413 37 -401 71
rect -367 37 -355 71
rect -413 31 -355 37
rect -221 71 -163 77
rect -221 37 -209 71
rect -175 37 -163 71
rect -221 31 -163 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 163 71 221 77
rect 163 37 175 71
rect 209 37 221 71
rect 163 31 221 37
rect 355 71 413 77
rect 355 37 367 71
rect 401 37 413 71
rect 355 31 413 37
rect 547 71 605 77
rect 547 37 559 71
rect 593 37 605 71
rect 547 31 605 37
rect 739 71 797 77
rect 739 37 751 71
rect 785 37 797 71
rect 739 31 797 37
rect 931 71 989 77
rect 931 37 943 71
rect 977 37 989 71
rect 931 31 989 37
rect 1123 71 1181 77
rect 1123 37 1135 71
rect 1169 37 1181 71
rect 1123 31 1181 37
rect -1181 -37 -1123 -31
rect -1181 -71 -1169 -37
rect -1135 -71 -1123 -37
rect -1181 -77 -1123 -71
rect -989 -37 -931 -31
rect -989 -71 -977 -37
rect -943 -71 -931 -37
rect -989 -77 -931 -71
rect -797 -37 -739 -31
rect -797 -71 -785 -37
rect -751 -71 -739 -37
rect -797 -77 -739 -71
rect -605 -37 -547 -31
rect -605 -71 -593 -37
rect -559 -71 -547 -37
rect -605 -77 -547 -71
rect -413 -37 -355 -31
rect -413 -71 -401 -37
rect -367 -71 -355 -37
rect -413 -77 -355 -71
rect -221 -37 -163 -31
rect -221 -71 -209 -37
rect -175 -71 -163 -37
rect -221 -77 -163 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 163 -37 221 -31
rect 163 -71 175 -37
rect 209 -71 221 -37
rect 163 -77 221 -71
rect 355 -37 413 -31
rect 355 -71 367 -37
rect 401 -71 413 -37
rect 355 -77 413 -71
rect 547 -37 605 -31
rect 547 -71 559 -37
rect 593 -71 605 -37
rect 547 -77 605 -71
rect 739 -37 797 -31
rect 739 -71 751 -37
rect 785 -71 797 -37
rect 739 -77 797 -71
rect 931 -37 989 -31
rect 931 -71 943 -37
rect 977 -71 989 -37
rect 931 -77 989 -71
rect 1123 -37 1181 -31
rect 1123 -71 1135 -37
rect 1169 -71 1181 -37
rect 1123 -77 1181 -71
rect -1223 -121 -1177 -109
rect -1223 -397 -1217 -121
rect -1183 -397 -1177 -121
rect -1223 -409 -1177 -397
rect -1127 -121 -1081 -109
rect -1127 -397 -1121 -121
rect -1087 -397 -1081 -121
rect -1127 -409 -1081 -397
rect -1031 -121 -985 -109
rect -1031 -397 -1025 -121
rect -991 -397 -985 -121
rect -1031 -409 -985 -397
rect -935 -121 -889 -109
rect -935 -397 -929 -121
rect -895 -397 -889 -121
rect -935 -409 -889 -397
rect -839 -121 -793 -109
rect -839 -397 -833 -121
rect -799 -397 -793 -121
rect -839 -409 -793 -397
rect -743 -121 -697 -109
rect -743 -397 -737 -121
rect -703 -397 -697 -121
rect -743 -409 -697 -397
rect -647 -121 -601 -109
rect -647 -397 -641 -121
rect -607 -397 -601 -121
rect -647 -409 -601 -397
rect -551 -121 -505 -109
rect -551 -397 -545 -121
rect -511 -397 -505 -121
rect -551 -409 -505 -397
rect -455 -121 -409 -109
rect -455 -397 -449 -121
rect -415 -397 -409 -121
rect -455 -409 -409 -397
rect -359 -121 -313 -109
rect -359 -397 -353 -121
rect -319 -397 -313 -121
rect -359 -409 -313 -397
rect -263 -121 -217 -109
rect -263 -397 -257 -121
rect -223 -397 -217 -121
rect -263 -409 -217 -397
rect -167 -121 -121 -109
rect -167 -397 -161 -121
rect -127 -397 -121 -121
rect -167 -409 -121 -397
rect -71 -121 -25 -109
rect -71 -397 -65 -121
rect -31 -397 -25 -121
rect -71 -409 -25 -397
rect 25 -121 71 -109
rect 25 -397 31 -121
rect 65 -397 71 -121
rect 25 -409 71 -397
rect 121 -121 167 -109
rect 121 -397 127 -121
rect 161 -397 167 -121
rect 121 -409 167 -397
rect 217 -121 263 -109
rect 217 -397 223 -121
rect 257 -397 263 -121
rect 217 -409 263 -397
rect 313 -121 359 -109
rect 313 -397 319 -121
rect 353 -397 359 -121
rect 313 -409 359 -397
rect 409 -121 455 -109
rect 409 -397 415 -121
rect 449 -397 455 -121
rect 409 -409 455 -397
rect 505 -121 551 -109
rect 505 -397 511 -121
rect 545 -397 551 -121
rect 505 -409 551 -397
rect 601 -121 647 -109
rect 601 -397 607 -121
rect 641 -397 647 -121
rect 601 -409 647 -397
rect 697 -121 743 -109
rect 697 -397 703 -121
rect 737 -397 743 -121
rect 697 -409 743 -397
rect 793 -121 839 -109
rect 793 -397 799 -121
rect 833 -397 839 -121
rect 793 -409 839 -397
rect 889 -121 935 -109
rect 889 -397 895 -121
rect 929 -397 935 -121
rect 889 -409 935 -397
rect 985 -121 1031 -109
rect 985 -397 991 -121
rect 1025 -397 1031 -121
rect 985 -409 1031 -397
rect 1081 -121 1127 -109
rect 1081 -397 1087 -121
rect 1121 -397 1127 -121
rect 1081 -409 1127 -397
rect 1177 -121 1223 -109
rect 1177 -397 1183 -121
rect 1217 -397 1223 -121
rect 1177 -409 1223 -397
rect -1085 -447 -1027 -441
rect -1085 -481 -1073 -447
rect -1039 -481 -1027 -447
rect -1085 -487 -1027 -481
rect -893 -447 -835 -441
rect -893 -481 -881 -447
rect -847 -481 -835 -447
rect -893 -487 -835 -481
rect -701 -447 -643 -441
rect -701 -481 -689 -447
rect -655 -481 -643 -447
rect -701 -487 -643 -481
rect -509 -447 -451 -441
rect -509 -481 -497 -447
rect -463 -481 -451 -447
rect -509 -487 -451 -481
rect -317 -447 -259 -441
rect -317 -481 -305 -447
rect -271 -481 -259 -447
rect -317 -487 -259 -481
rect -125 -447 -67 -441
rect -125 -481 -113 -447
rect -79 -481 -67 -447
rect -125 -487 -67 -481
rect 67 -447 125 -441
rect 67 -481 79 -447
rect 113 -481 125 -447
rect 67 -487 125 -481
rect 259 -447 317 -441
rect 259 -481 271 -447
rect 305 -481 317 -447
rect 259 -487 317 -481
rect 451 -447 509 -441
rect 451 -481 463 -447
rect 497 -481 509 -447
rect 451 -487 509 -481
rect 643 -447 701 -441
rect 643 -481 655 -447
rect 689 -481 701 -447
rect 643 -487 701 -481
rect 835 -447 893 -441
rect 835 -481 847 -447
rect 881 -481 893 -447
rect 835 -487 893 -481
rect 1027 -447 1085 -441
rect 1027 -481 1039 -447
rect 1073 -481 1085 -447
rect 1027 -487 1085 -481
rect -1085 -555 -1027 -549
rect -1085 -589 -1073 -555
rect -1039 -589 -1027 -555
rect -1085 -595 -1027 -589
rect -893 -555 -835 -549
rect -893 -589 -881 -555
rect -847 -589 -835 -555
rect -893 -595 -835 -589
rect -701 -555 -643 -549
rect -701 -589 -689 -555
rect -655 -589 -643 -555
rect -701 -595 -643 -589
rect -509 -555 -451 -549
rect -509 -589 -497 -555
rect -463 -589 -451 -555
rect -509 -595 -451 -589
rect -317 -555 -259 -549
rect -317 -589 -305 -555
rect -271 -589 -259 -555
rect -317 -595 -259 -589
rect -125 -555 -67 -549
rect -125 -589 -113 -555
rect -79 -589 -67 -555
rect -125 -595 -67 -589
rect 67 -555 125 -549
rect 67 -589 79 -555
rect 113 -589 125 -555
rect 67 -595 125 -589
rect 259 -555 317 -549
rect 259 -589 271 -555
rect 305 -589 317 -555
rect 259 -595 317 -589
rect 451 -555 509 -549
rect 451 -589 463 -555
rect 497 -589 509 -555
rect 451 -595 509 -589
rect 643 -555 701 -549
rect 643 -589 655 -555
rect 689 -589 701 -555
rect 643 -595 701 -589
rect 835 -555 893 -549
rect 835 -589 847 -555
rect 881 -589 893 -555
rect 835 -595 893 -589
rect 1027 -555 1085 -549
rect 1027 -589 1039 -555
rect 1073 -589 1085 -555
rect 1027 -595 1085 -589
rect -1223 -639 -1177 -627
rect -1223 -915 -1217 -639
rect -1183 -915 -1177 -639
rect -1223 -927 -1177 -915
rect -1127 -639 -1081 -627
rect -1127 -915 -1121 -639
rect -1087 -915 -1081 -639
rect -1127 -927 -1081 -915
rect -1031 -639 -985 -627
rect -1031 -915 -1025 -639
rect -991 -915 -985 -639
rect -1031 -927 -985 -915
rect -935 -639 -889 -627
rect -935 -915 -929 -639
rect -895 -915 -889 -639
rect -935 -927 -889 -915
rect -839 -639 -793 -627
rect -839 -915 -833 -639
rect -799 -915 -793 -639
rect -839 -927 -793 -915
rect -743 -639 -697 -627
rect -743 -915 -737 -639
rect -703 -915 -697 -639
rect -743 -927 -697 -915
rect -647 -639 -601 -627
rect -647 -915 -641 -639
rect -607 -915 -601 -639
rect -647 -927 -601 -915
rect -551 -639 -505 -627
rect -551 -915 -545 -639
rect -511 -915 -505 -639
rect -551 -927 -505 -915
rect -455 -639 -409 -627
rect -455 -915 -449 -639
rect -415 -915 -409 -639
rect -455 -927 -409 -915
rect -359 -639 -313 -627
rect -359 -915 -353 -639
rect -319 -915 -313 -639
rect -359 -927 -313 -915
rect -263 -639 -217 -627
rect -263 -915 -257 -639
rect -223 -915 -217 -639
rect -263 -927 -217 -915
rect -167 -639 -121 -627
rect -167 -915 -161 -639
rect -127 -915 -121 -639
rect -167 -927 -121 -915
rect -71 -639 -25 -627
rect -71 -915 -65 -639
rect -31 -915 -25 -639
rect -71 -927 -25 -915
rect 25 -639 71 -627
rect 25 -915 31 -639
rect 65 -915 71 -639
rect 25 -927 71 -915
rect 121 -639 167 -627
rect 121 -915 127 -639
rect 161 -915 167 -639
rect 121 -927 167 -915
rect 217 -639 263 -627
rect 217 -915 223 -639
rect 257 -915 263 -639
rect 217 -927 263 -915
rect 313 -639 359 -627
rect 313 -915 319 -639
rect 353 -915 359 -639
rect 313 -927 359 -915
rect 409 -639 455 -627
rect 409 -915 415 -639
rect 449 -915 455 -639
rect 409 -927 455 -915
rect 505 -639 551 -627
rect 505 -915 511 -639
rect 545 -915 551 -639
rect 505 -927 551 -915
rect 601 -639 647 -627
rect 601 -915 607 -639
rect 641 -915 647 -639
rect 601 -927 647 -915
rect 697 -639 743 -627
rect 697 -915 703 -639
rect 737 -915 743 -639
rect 697 -927 743 -915
rect 793 -639 839 -627
rect 793 -915 799 -639
rect 833 -915 839 -639
rect 793 -927 839 -915
rect 889 -639 935 -627
rect 889 -915 895 -639
rect 929 -915 935 -639
rect 889 -927 935 -915
rect 985 -639 1031 -627
rect 985 -915 991 -639
rect 1025 -915 1031 -639
rect 985 -927 1031 -915
rect 1081 -639 1127 -627
rect 1081 -915 1087 -639
rect 1121 -915 1127 -639
rect 1081 -927 1127 -915
rect 1177 -639 1223 -627
rect 1177 -915 1183 -639
rect 1217 -915 1223 -639
rect 1177 -927 1223 -915
rect -1181 -965 -1123 -959
rect -1181 -999 -1169 -965
rect -1135 -999 -1123 -965
rect -1181 -1005 -1123 -999
rect -989 -965 -931 -959
rect -989 -999 -977 -965
rect -943 -999 -931 -965
rect -989 -1005 -931 -999
rect -797 -965 -739 -959
rect -797 -999 -785 -965
rect -751 -999 -739 -965
rect -797 -1005 -739 -999
rect -605 -965 -547 -959
rect -605 -999 -593 -965
rect -559 -999 -547 -965
rect -605 -1005 -547 -999
rect -413 -965 -355 -959
rect -413 -999 -401 -965
rect -367 -999 -355 -965
rect -413 -1005 -355 -999
rect -221 -965 -163 -959
rect -221 -999 -209 -965
rect -175 -999 -163 -965
rect -221 -1005 -163 -999
rect -29 -965 29 -959
rect -29 -999 -17 -965
rect 17 -999 29 -965
rect -29 -1005 29 -999
rect 163 -965 221 -959
rect 163 -999 175 -965
rect 209 -999 221 -965
rect 163 -1005 221 -999
rect 355 -965 413 -959
rect 355 -999 367 -965
rect 401 -999 413 -965
rect 355 -1005 413 -999
rect 547 -965 605 -959
rect 547 -999 559 -965
rect 593 -999 605 -965
rect 547 -1005 605 -999
rect 739 -965 797 -959
rect 739 -999 751 -965
rect 785 -999 797 -965
rect 739 -1005 797 -999
rect 931 -965 989 -959
rect 931 -999 943 -965
rect 977 -999 989 -965
rect 931 -1005 989 -999
rect 1123 -965 1181 -959
rect 1123 -999 1135 -965
rect 1169 -999 1181 -965
rect 1123 -1005 1181 -999
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1314 -1084 1314 1084
string parameters w 1.5 l 0.15 m 4 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
