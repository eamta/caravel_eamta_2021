magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 9043 4969 9078 4986
rect 12787 4969 12822 4986
rect 9007 4952 9078 4969
rect 12751 4952 12822 4969
rect 8674 4916 8709 4933
rect 8638 4899 8709 4916
rect 8305 4863 8340 4880
rect 8269 4846 8340 4863
rect 7936 4810 7971 4827
rect 7900 4793 7971 4810
rect 7567 4757 7602 4774
rect 7531 4740 7602 4757
rect 7198 4687 7233 4721
rect 6829 4634 6864 4668
rect 6460 4598 6495 4615
rect 6424 4581 6495 4598
rect 6055 4545 6091 4548
rect 607 4476 625 4528
rect 635 4476 653 4528
rect 4351 4476 4369 4528
rect 4379 4476 4397 4528
rect 5686 4522 6091 4545
rect 6125 4528 6399 4562
rect 6125 4522 6371 4528
rect 5291 4492 5686 4518
rect 5784 4509 6010 4522
rect 5722 4500 6072 4509
rect 6091 4500 6337 4522
rect 5722 4494 6337 4500
rect 5722 4490 6125 4494
rect 5319 4489 6125 4490
rect 6199 4489 6321 4494
rect 6345 4489 6371 4522
rect 5317 4488 6371 4489
rect 5722 4476 5737 4488
rect 6057 4476 6072 4488
rect 5722 4475 6072 4476
rect 5353 4446 5703 4456
rect 607 4440 625 4446
rect 635 4440 653 4446
rect 4351 4440 4369 4446
rect 4379 4440 4397 4446
rect 5353 4442 5388 4446
rect 1493 4402 1511 4440
rect 659 4356 668 4399
rect 506 4288 614 4345
rect 659 4322 805 4356
rect 556 4255 682 4288
rect 867 4282 1064 4356
rect 879 4278 996 4282
rect 576 4251 602 4255
rect 889 4252 996 4278
rect 1487 4256 1511 4402
rect 1521 4374 1539 4440
rect 1515 4284 1539 4374
rect 4403 4351 4412 4399
rect 4035 4348 4158 4350
rect 3924 4288 4158 4348
rect 4308 4306 4312 4331
rect 4403 4322 4461 4351
rect 4491 4322 4549 4351
rect 4711 4350 4745 4360
rect 4799 4350 4833 4384
rect 4984 4369 5107 4403
rect 5237 4402 5255 4440
rect 5231 4374 5255 4402
rect 5265 4374 5283 4440
rect 5334 4439 5467 4442
rect 5317 4404 5467 4439
rect 5669 4404 5680 4415
rect 5688 4404 5703 4446
rect 5317 4400 5603 4404
rect 5311 4394 5370 4400
rect 5387 4394 5603 4400
rect 5311 4374 5603 4394
rect 5669 4374 5703 4404
rect 5722 4404 5756 4475
rect 5822 4446 5972 4465
rect 6038 4446 6072 4475
rect 6091 4446 6125 4488
rect 6424 4466 6494 4581
rect 6606 4513 6664 4519
rect 6606 4479 6618 4513
rect 6606 4473 6664 4479
rect 6233 4454 6299 4460
rect 6249 4450 6283 4454
rect 5879 4441 6249 4446
rect 5840 4440 6249 4441
rect 5722 4374 5737 4404
rect 5231 4369 5387 4374
rect 4415 4318 4449 4322
rect 4503 4318 4537 4322
rect 4611 4316 4845 4350
rect 4850 4339 4902 4350
rect 4939 4341 4965 4350
rect 4984 4341 5018 4369
rect 4861 4327 4891 4339
rect 4939 4334 5018 4341
rect 4850 4316 4902 4327
rect 4939 4322 4965 4334
rect 4611 4306 4650 4316
rect 4711 4306 4745 4316
rect 4212 4297 4246 4306
rect 4300 4297 4358 4306
rect 4212 4288 4596 4297
rect 4611 4294 4745 4306
rect 4611 4288 4757 4294
rect 3924 4280 4103 4288
rect 4158 4286 4757 4288
rect 4158 4282 4845 4286
rect 610 4251 636 4252
rect 610 4233 645 4251
rect 810 4244 996 4252
rect 810 4241 862 4244
rect 691 4236 801 4240
rect 207 4166 226 4231
rect 574 4218 645 4233
rect 679 4229 813 4236
rect 821 4229 851 4241
rect 679 4218 862 4229
rect 241 4170 414 4197
rect 515 4186 567 4197
rect 526 4174 556 4186
rect 241 4102 268 4170
rect 315 4163 367 4170
rect 515 4163 567 4174
rect 341 4111 356 4153
rect 384 4152 444 4156
rect 384 4124 416 4128
rect 383 4102 398 4111
rect 402 4102 416 4124
rect 430 4102 444 4152
rect 557 4102 567 4163
rect 574 4102 644 4218
rect 889 4214 996 4244
rect 1159 4214 1250 4232
rect 1717 4216 1802 4250
rect 1908 4216 2127 4248
rect 3924 4244 3925 4280
rect 4024 4244 4058 4280
rect 4158 4278 4745 4282
rect 4799 4278 4833 4282
rect 4112 4252 4740 4278
rect 4112 4244 4165 4252
rect 3877 4233 4165 4244
rect 4173 4233 4193 4251
rect 4210 4233 4740 4252
rect 4757 4244 4823 4248
rect 3841 4227 4740 4233
rect 713 4184 779 4202
rect 821 4184 851 4208
rect 718 4168 851 4184
rect 779 4164 851 4168
rect 779 4156 784 4164
rect 779 4150 814 4156
rect 752 4136 814 4150
rect 752 4134 813 4136
rect 756 4130 801 4134
rect 205 4074 644 4102
rect 728 4082 745 4124
rect 756 4110 773 4130
rect 821 4110 851 4164
rect 926 4127 960 4145
rect 1143 4127 1250 4214
rect 1722 4180 1734 4182
rect 1314 4127 1329 4174
rect 1410 4146 1417 4158
rect 1348 4127 1429 4146
rect 926 4091 996 4127
rect 1143 4112 1429 4127
rect 1444 4135 1538 4146
rect 1572 4145 1624 4146
rect 1572 4135 1657 4145
rect 1976 4142 1988 4180
rect 3508 4174 3543 4191
rect 3472 4157 3543 4174
rect 3734 4176 4740 4227
rect 4861 4198 4865 4306
rect 4950 4232 4965 4318
rect 4984 4232 5018 4334
rect 5039 4318 5052 4369
rect 5231 4280 5255 4369
rect 5259 4284 5299 4369
rect 5266 4280 5299 4284
rect 5300 4285 5387 4369
rect 5393 4344 5495 4374
rect 5519 4354 5549 4374
rect 5561 4354 5737 4374
rect 5519 4344 5737 4354
rect 5393 4320 5737 4344
rect 5393 4310 5495 4320
rect 5507 4314 5737 4320
rect 5393 4306 5507 4310
rect 5519 4306 5737 4314
rect 5756 4326 5824 4374
rect 5840 4339 5859 4440
rect 5879 4438 6249 4440
rect 5879 4413 6251 4438
rect 5868 4410 6251 4413
rect 6281 4416 6299 4438
rect 5868 4379 6249 4410
rect 6281 4379 6331 4416
rect 5868 4378 6251 4379
rect 5868 4373 5887 4378
rect 5925 4373 5930 4378
rect 5868 4367 5926 4373
rect 5947 4364 5966 4378
rect 6013 4366 6081 4378
rect 5947 4352 5992 4364
rect 5947 4330 5993 4352
rect 5836 4326 5893 4328
rect 5756 4306 5893 4326
rect 5925 4314 5993 4330
rect 5399 4285 5467 4306
rect 5300 4284 5467 4285
rect 5473 4295 5519 4306
rect 5549 4304 5595 4306
rect 5055 4256 5255 4280
rect 5027 4232 5283 4252
rect 4903 4228 5283 4232
rect 4903 4214 5232 4228
rect 5300 4214 5387 4284
rect 5461 4273 5462 4284
rect 5473 4273 5535 4295
rect 5555 4286 5595 4304
rect 5669 4294 5756 4306
rect 5561 4273 5595 4286
rect 4883 4182 4885 4204
rect 4887 4182 5387 4214
rect 1444 4112 1451 4135
rect 1461 4128 1527 4135
rect 1583 4127 1657 4135
rect 2028 4134 2188 4144
rect 2028 4133 2069 4134
rect 1687 4127 1698 4133
rect 2039 4127 2069 4133
rect 2111 4133 2188 4134
rect 2250 4133 2302 4144
rect 2338 4143 2362 4144
rect 1583 4123 2029 4127
rect 1572 4112 2029 4123
rect 1143 4091 1382 4112
rect 943 4090 1086 4091
rect 1106 4090 1382 4091
rect 184 4062 644 4074
rect 724 4069 758 4080
rect 770 4069 800 4080
rect 812 4069 846 4080
rect 205 4046 644 4062
rect 722 4057 770 4069
rect 800 4065 858 4069
rect 809 4059 858 4065
rect 800 4057 858 4059
rect 724 4054 770 4057
rect 724 4046 767 4054
rect 812 4046 858 4057
rect 178 4039 913 4046
rect 178 4034 926 4039
rect 205 4021 926 4034
rect 943 4038 1382 4090
rect 1383 4038 1416 4112
rect 1466 4066 1580 4078
rect 1466 4056 1562 4066
rect 1490 4038 1562 4056
rect 1607 4059 2029 4112
rect 2039 4110 2101 4127
rect 2111 4120 2177 4133
rect 2261 4121 2291 4133
rect 2250 4112 2291 4121
rect 2351 4112 2362 4123
rect 2480 4121 2657 4142
rect 3139 4121 3174 4138
rect 2250 4110 2362 4112
rect 2039 4093 2046 4110
rect 2039 4059 2067 4093
rect 943 4021 1429 4038
rect 1434 4036 1578 4038
rect 1434 4032 1605 4036
rect 1607 4032 2067 4059
rect 2154 4040 2181 4058
rect 2261 4040 2262 4078
rect 2328 4067 2362 4110
rect 2734 4068 2945 4121
rect 3103 4104 3174 4121
rect 2333 4062 2362 4067
rect 2328 4040 2362 4048
rect 1434 4027 2067 4032
rect 205 4012 1429 4021
rect 1445 4017 1475 4027
rect 1483 4018 2067 4027
rect 1483 4017 2047 4018
rect 1445 4015 2047 4017
rect 205 3956 644 4012
rect 737 3966 767 4012
rect 812 4004 1429 4012
rect 1434 4004 2047 4015
rect 812 3988 1382 4004
rect 825 3974 858 3988
rect 171 3938 644 3956
rect 171 3922 192 3938
rect 205 3932 644 3938
rect 724 3938 767 3966
rect 724 3932 787 3938
rect 800 3932 858 3974
rect 869 3932 1382 3988
rect 205 3922 1382 3932
rect 1383 3983 1416 4004
rect 1490 3998 1517 4004
rect 1490 3994 1584 3998
rect 1383 3922 1429 3983
rect 1508 3978 1584 3994
rect 1590 3997 2047 4004
rect 2052 3997 2067 4018
rect 1508 3970 1588 3978
rect 1462 3967 1500 3970
rect 1462 3964 1496 3967
rect 1462 3963 1500 3964
rect 1508 3963 1530 3970
rect 1533 3964 1588 3970
rect 1450 3956 1509 3963
rect 1432 3922 1509 3956
rect 1517 3928 1530 3963
rect 1538 3963 1588 3964
rect 1590 3963 2067 3997
rect 2086 4033 2362 4040
rect 2365 4033 2691 4068
rect 2086 4032 2691 4033
rect 2734 4051 2805 4068
rect 2086 4023 2717 4032
rect 2734 4023 2804 4051
rect 2086 4006 2804 4023
rect 2086 3979 2120 4006
rect 2154 3992 2181 4006
rect 2261 3992 2262 4006
rect 2172 3983 2181 3992
rect 2128 3979 2282 3983
rect 2328 3979 2362 4006
rect 2365 3979 2804 4006
rect 1538 3948 2067 3963
rect 1550 3946 2067 3948
rect 2092 3946 2097 3979
rect 2109 3970 2804 3979
rect 2916 3983 2974 3989
rect 2109 3952 2805 3970
rect 2916 3963 2928 3983
rect 2916 3952 2930 3963
rect 2960 3952 2962 3963
rect 3103 3952 3173 4104
rect 3285 4036 3343 4042
rect 3285 4002 3297 4036
rect 3285 3996 3343 4002
rect 2109 3946 3173 3952
rect 1550 3945 3173 3946
rect 1550 3934 2067 3945
rect 2086 3934 2191 3945
rect 1550 3928 2191 3934
rect 2197 3938 2278 3945
rect 2294 3938 3173 3945
rect 1550 3922 1584 3928
rect 1590 3922 2120 3928
rect 2126 3922 2185 3928
rect 2197 3922 3173 3938
rect 181 3916 3173 3922
rect 181 3915 3174 3916
rect 144 3911 3174 3915
rect 144 3904 2295 3911
rect 144 3899 2294 3904
rect 144 3898 2302 3899
rect 144 3896 644 3898
rect 679 3896 2302 3898
rect 144 3895 2302 3896
rect 2328 3895 3174 3911
rect 144 3888 3174 3895
rect 144 3884 702 3888
rect 711 3885 782 3888
rect 711 3884 745 3885
rect 757 3884 782 3885
rect 799 3885 846 3888
rect 799 3884 833 3885
rect 144 3876 755 3884
rect 144 3846 644 3876
rect 652 3846 786 3876
rect 144 3840 653 3846
rect 664 3842 786 3846
rect 787 3872 845 3884
rect 852 3872 2120 3888
rect 787 3846 2120 3872
rect 787 3842 798 3846
rect 799 3842 2120 3846
rect 664 3840 2120 3842
rect 2126 3879 2197 3888
rect 2202 3879 2260 3888
rect 2126 3858 2260 3879
rect 2126 3857 2282 3858
rect 2288 3857 2322 3861
rect 2328 3857 3174 3888
rect 3241 3874 3299 3917
rect 3329 3874 3387 3917
rect 3472 3899 3542 4157
rect 3734 4125 4758 4176
rect 4805 4161 4834 4176
rect 4805 4125 4819 4161
rect 4841 4146 5387 4182
rect 5455 4200 5460 4273
rect 5461 4217 5601 4273
rect 5649 4228 5717 4294
rect 5722 4228 5771 4294
rect 5824 4228 5893 4306
rect 5924 4300 5993 4314
rect 5924 4289 5992 4300
rect 6038 4289 6081 4366
rect 6091 4289 6125 4378
rect 6135 4289 6159 4378
rect 6167 4300 6169 4366
rect 6171 4289 6175 4378
rect 6181 4375 6251 4378
rect 6281 4375 6339 4379
rect 6407 4375 6494 4466
rect 6181 4289 6494 4375
rect 5924 4288 6494 4289
rect 5924 4262 5958 4288
rect 5959 4284 5992 4288
rect 6038 4284 6081 4288
rect 5925 4250 5958 4262
rect 5669 4217 5703 4228
rect 5722 4217 5756 4228
rect 5824 4217 5871 4228
rect 5461 4216 5871 4217
rect 4841 4127 5401 4146
rect 5430 4127 5442 4146
rect 5455 4127 5496 4200
rect 5543 4127 5549 4216
rect 5592 4213 5601 4216
rect 5588 4127 5601 4213
rect 5669 4127 5703 4216
rect 5722 4127 5756 4216
rect 5824 4179 5828 4216
rect 5836 4186 5870 4208
rect 5905 4204 5952 4217
rect 5836 4179 5882 4186
rect 5824 4170 5882 4179
rect 5905 4170 5955 4204
rect 5824 4144 5955 4170
rect 6038 4144 6072 4284
rect 5772 4134 5970 4144
rect 5772 4133 5813 4134
rect 5783 4127 5813 4133
rect 5824 4127 5970 4134
rect 5994 4133 6072 4144
rect 4841 4125 5773 4127
rect 3734 4098 4763 4125
rect 4805 4098 5773 4125
rect 3654 4089 3712 4095
rect 3734 4091 4758 4098
rect 4805 4091 4819 4098
rect 4841 4091 5773 4098
rect 3654 4055 3666 4089
rect 3654 4049 3712 4055
rect 3734 4048 5773 4091
rect 5783 4110 5970 4127
rect 6005 4121 6035 4133
rect 5994 4112 6035 4121
rect 6038 4112 6072 4133
rect 6091 4112 6125 4288
rect 6135 4284 6159 4288
rect 6195 4280 6207 4288
rect 6199 4260 6203 4280
rect 6213 4246 6494 4288
rect 6606 4313 6664 4319
rect 6606 4279 6618 4313
rect 6606 4273 6664 4279
rect 6205 4211 6494 4246
rect 6205 4201 6495 4211
rect 6193 4177 6495 4201
rect 6795 4196 6810 4615
rect 6829 4264 6863 4634
rect 6975 4566 7033 4572
rect 6975 4532 6987 4566
rect 6975 4526 7033 4532
rect 6975 4366 7033 4372
rect 6975 4332 6987 4366
rect 6975 4326 7033 4332
rect 6829 4230 6864 4264
rect 7164 4249 7179 4668
rect 7198 4317 7232 4687
rect 7344 4619 7402 4625
rect 7344 4585 7356 4619
rect 7344 4579 7402 4585
rect 7344 4419 7402 4425
rect 7344 4385 7356 4419
rect 7344 4379 7402 4385
rect 7198 4283 7233 4317
rect 7531 4283 7601 4740
rect 7713 4672 7771 4678
rect 7713 4638 7725 4672
rect 7713 4632 7771 4638
rect 7900 4423 7970 4793
rect 8082 4725 8140 4731
rect 8082 4691 8094 4725
rect 8082 4685 8140 4691
rect 8082 4525 8140 4531
rect 8082 4491 8094 4525
rect 8082 4485 8140 4491
rect 7900 4389 7971 4423
rect 8269 4389 8339 4846
rect 8451 4778 8509 4784
rect 8451 4744 8463 4778
rect 8451 4738 8509 4744
rect 8638 4529 8708 4899
rect 8820 4831 8878 4837
rect 8820 4797 8832 4831
rect 8820 4791 8878 4797
rect 8820 4631 8878 4637
rect 8820 4597 8832 4631
rect 8820 4591 8878 4597
rect 8638 4495 8709 4529
rect 9007 4495 9077 4952
rect 12418 4916 12453 4933
rect 12382 4899 12453 4916
rect 9189 4884 9247 4890
rect 9189 4850 9201 4884
rect 12049 4863 12084 4880
rect 9189 4844 9247 4850
rect 12013 4846 12084 4863
rect 11680 4810 11715 4827
rect 9176 4545 9429 4799
rect 11644 4793 11715 4810
rect 11311 4757 11346 4774
rect 11275 4740 11346 4757
rect 10942 4687 10977 4721
rect 10573 4634 10608 4668
rect 10204 4598 10239 4615
rect 10168 4581 10239 4598
rect 9189 4542 9201 4545
rect 9189 4536 9247 4542
rect 8451 4470 8509 4476
rect 8451 4436 8463 4470
rect 8638 4459 8691 4495
rect 9007 4459 9060 4495
rect 9430 4492 9683 4545
rect 9835 4528 9870 4562
rect 9466 4475 9501 4492
rect 9043 4440 9132 4457
rect 9139 4456 9297 4474
rect 9139 4440 9351 4456
rect 9432 4440 9447 4456
rect 9097 4439 9447 4440
rect 8451 4430 8509 4436
rect 9007 4422 9447 4439
rect 7713 4364 7771 4370
rect 7713 4330 7725 4364
rect 7900 4353 7953 4389
rect 8269 4353 8322 4389
rect 8728 4387 8763 4403
rect 9007 4387 9131 4422
rect 8728 4386 9131 4387
rect 9221 4386 9323 4388
rect 8323 4351 8691 4386
rect 8305 4334 8691 4351
rect 8728 4369 9114 4386
rect 8694 4334 8709 4350
rect 8323 4333 8709 4334
rect 8728 4333 8762 4369
rect 9007 4360 9114 4369
rect 8852 4333 8954 4335
rect 7713 4324 7771 4330
rect 8269 4297 8709 4333
rect 8770 4299 8796 4333
rect 8839 4299 8967 4333
rect 8024 4288 8709 4297
rect 7531 4251 7584 4283
rect 7954 4263 8709 4288
rect 7663 4251 7821 4262
rect 7900 4251 8709 4263
rect 7531 4247 7621 4251
rect 7567 4233 7621 4247
rect 7655 4233 8709 4251
rect 7531 4227 8709 4233
rect 6193 4139 6477 4177
rect 7252 4175 7287 4191
rect 7478 4182 8709 4227
rect 8728 4182 8762 4299
rect 8874 4289 8886 4299
rect 8870 4267 8920 4289
rect 9007 4283 9131 4360
rect 9139 4352 9165 4386
rect 9217 4352 9327 4386
rect 9243 4342 9255 4352
rect 9239 4320 9289 4342
rect 9379 4327 9393 4386
rect 9239 4314 9301 4320
rect 9239 4304 9293 4314
rect 8870 4261 8932 4267
rect 8870 4251 8924 4261
rect 8808 4237 8866 4251
rect 8808 4233 8878 4237
rect 8808 4231 8866 4233
rect 8808 4229 8832 4231
rect 8888 4229 8918 4251
rect 8808 4217 8904 4229
rect 8830 4197 8900 4217
rect 8830 4182 8882 4197
rect 8930 4187 8944 4197
rect 8924 4185 8944 4187
rect 8924 4182 8948 4185
rect 8956 4182 8964 4233
rect 8965 4182 8976 4229
rect 8990 4182 9131 4283
rect 9177 4290 9235 4295
rect 9177 4286 9247 4290
rect 9177 4284 9235 4286
rect 9177 4273 9201 4284
rect 9235 4273 9245 4284
rect 9257 4273 9287 4304
rect 9177 4261 9282 4273
rect 9199 4250 9269 4261
rect 9199 4234 9251 4250
rect 9199 4219 9245 4234
rect 9299 4231 9313 4241
rect 9157 4203 9165 4207
rect 9177 4203 9191 4207
rect 9203 4203 9245 4219
rect 9293 4229 9313 4231
rect 7478 4175 9131 4182
rect 7252 4174 9131 4175
rect 6205 4127 6477 4139
rect 5994 4110 6125 4112
rect 5783 4093 5790 4110
rect 5783 4048 5811 4093
rect 3734 4040 5811 4048
rect 5824 4063 5828 4110
rect 5836 4098 5870 4110
rect 5924 4098 5943 4110
rect 5836 4063 5845 4098
rect 5924 4076 5970 4089
rect 6038 4078 6125 4110
rect 5824 4048 5845 4063
rect 5864 4048 5870 4076
rect 5874 4048 5876 4076
rect 5924 4058 5982 4076
rect 5824 4040 5882 4048
rect 5902 4042 5904 4048
rect 5898 4040 5904 4042
rect 5912 4040 5982 4058
rect 6038 4048 6072 4078
rect 6077 4068 6125 4078
rect 6193 4121 6477 4127
rect 6883 4122 6918 4138
rect 7216 4122 9131 4174
rect 6883 4121 9131 4122
rect 6193 4068 6239 4121
rect 6281 4068 6327 4121
rect 6407 4068 6441 4121
rect 6478 4069 6731 4121
rect 6847 4104 9131 4121
rect 6793 4069 6917 4104
rect 7198 4093 9131 4104
rect 9145 4093 9197 4203
rect 9205 4191 9245 4203
rect 9265 4203 9279 4207
rect 9265 4202 9285 4203
rect 9257 4191 9285 4202
rect 9205 4105 9285 4191
rect 9205 4093 9225 4105
rect 9245 4093 9285 4105
rect 9293 4105 9317 4229
rect 9293 4093 9313 4105
rect 9325 4093 9333 4277
rect 9334 4093 9345 4273
rect 7198 4084 9291 4093
rect 9325 4084 9340 4093
rect 6478 4068 6917 4069
rect 7007 4068 7109 4070
rect 6077 4062 6477 4068
rect 6091 4048 6477 4062
rect 6038 4040 6477 4048
rect 3734 4023 6477 4040
rect 6478 4042 6900 4068
rect 6478 4023 6917 4042
rect 6925 4034 6951 4068
rect 6994 4034 7122 4068
rect 7029 4024 7041 4034
rect 3734 4008 6917 4023
rect 3731 4006 6917 4008
rect 3731 3997 5790 4006
rect 5796 3997 5811 4006
rect 3731 3979 5811 3997
rect 5824 3983 5882 4006
rect 5902 4002 5904 4006
rect 5912 3992 5970 4006
rect 5916 3983 5970 3992
rect 6038 3987 6917 4006
rect 5984 3983 6917 3987
rect 7025 4002 7075 4024
rect 7164 4018 7179 4068
rect 7025 3996 7087 4002
rect 7025 3986 7079 3996
rect 5824 3979 6917 3983
rect 3731 3972 6917 3979
rect 3731 3954 5811 3972
rect 5824 3966 6917 3972
rect 3731 3946 5823 3954
rect 5836 3946 5841 3966
rect 5853 3953 6917 3966
rect 5846 3946 6917 3953
rect 6963 3972 7021 3986
rect 6963 3968 7033 3972
rect 6963 3966 7021 3968
rect 6963 3964 6987 3966
rect 7043 3964 7073 3986
rect 6963 3952 7059 3964
rect 3731 3945 6917 3946
rect 3731 3938 5823 3945
rect 5830 3938 6018 3945
rect 6038 3938 6917 3945
rect 3731 3932 6917 3938
rect 3731 3930 6106 3932
rect 3734 3929 6106 3930
rect 3734 3909 5173 3929
rect 5176 3909 5280 3929
rect 5294 3928 6106 3929
rect 6109 3928 6917 3932
rect 5294 3916 6917 3928
rect 6985 3932 7055 3952
rect 6985 3916 7037 3932
rect 7085 3922 7099 3932
rect 7079 3920 7099 3922
rect 7079 3917 7103 3920
rect 7111 3917 7119 3968
rect 7120 3917 7131 3964
rect 5294 3911 6918 3916
rect 5294 3909 6018 3911
rect 6022 3909 6026 3911
rect 6038 3909 6918 3911
rect 3734 3901 6918 3909
rect 6985 3904 7031 3916
rect 6985 3901 7065 3904
rect 3472 3897 3579 3899
rect 3253 3870 3287 3874
rect 3341 3870 3375 3874
rect 2126 3846 3174 3857
rect 2126 3845 2291 3846
rect 2126 3843 2248 3845
rect 2126 3840 2197 3843
rect 144 3748 644 3840
rect 664 3837 2197 3840
rect 2200 3837 2248 3843
rect 2254 3840 2291 3845
rect 664 3830 2248 3837
rect 2276 3834 2291 3840
rect 2294 3834 2322 3846
rect 2276 3830 2322 3834
rect 664 3827 2197 3830
rect 664 3812 2185 3827
rect 659 3800 2185 3812
rect 2191 3809 2197 3827
rect 2192 3800 2197 3809
rect 2200 3800 2248 3830
rect 2254 3812 2322 3830
rect 2276 3800 2322 3812
rect 659 3799 2322 3800
rect 2328 3799 3174 3846
rect 659 3781 3174 3799
rect 659 3778 2120 3781
rect 659 3774 2067 3778
rect 2086 3774 2120 3778
rect 2126 3777 3174 3781
rect 2140 3774 2143 3777
rect 2146 3774 3174 3777
rect 659 3753 3174 3774
rect 650 3748 3174 3753
rect 144 3738 3174 3748
rect 144 3734 2195 3738
rect 2200 3734 3174 3738
rect 3193 3836 3409 3863
rect 3455 3846 3579 3897
rect 3734 3883 6106 3901
rect 6109 3883 6918 3901
rect 6989 3898 7065 3901
rect 6943 3894 6952 3898
rect 6963 3894 6977 3898
rect 6989 3894 7031 3898
rect 7037 3894 7065 3898
rect 3734 3879 6918 3883
rect 3734 3875 6046 3879
rect 3734 3857 6026 3875
rect 6038 3861 6052 3875
rect 6032 3857 6052 3861
rect 6072 3863 6918 3879
rect 6931 3863 6983 3894
rect 6991 3882 7031 3894
rect 7051 3893 7071 3894
rect 7043 3882 7071 3893
rect 6991 3874 7071 3882
rect 7077 3874 7131 3917
rect 6997 3870 7073 3874
rect 7085 3870 7119 3874
rect 7031 3863 7073 3870
rect 7145 3863 7179 4018
rect 7198 4059 9340 4084
rect 7198 3968 9131 4059
rect 9145 4038 9191 4059
rect 9208 4049 9340 4059
rect 9203 4038 9340 4049
rect 9145 4035 9340 4038
rect 9145 4023 9305 4035
rect 9157 4019 9191 4023
rect 9136 3995 9194 3997
rect 9203 3992 9233 4023
rect 9239 4012 9305 4023
rect 9239 3996 9293 4012
rect 9132 3985 9219 3991
rect 9132 3978 9182 3985
rect 9198 3982 9219 3985
rect 9198 3978 9247 3982
rect 9132 3968 9185 3978
rect 9198 3976 9219 3978
rect 7198 3957 9193 3968
rect 7198 3944 9150 3957
rect 9180 3944 9193 3957
rect 9201 3944 9220 3976
rect 9306 3944 9340 4035
rect 9359 4040 9393 4327
rect 9413 4040 9447 4422
rect 9466 4040 9500 4475
rect 9612 4407 9670 4413
rect 9612 4373 9624 4407
rect 9612 4367 9670 4373
rect 9359 4006 9394 4040
rect 9413 4006 9427 4040
rect 9455 4006 9714 4040
rect 9801 4021 9816 4509
rect 7198 3929 9351 3944
rect 7198 3910 9077 3929
rect 9097 3928 9351 3929
rect 9359 3928 9393 4006
rect 9413 3944 9447 4006
rect 9097 3926 9393 3928
rect 9097 3923 9185 3926
rect 9097 3910 9131 3923
rect 9150 3910 9180 3923
rect 9193 3910 9393 3926
rect 9432 3910 9447 3944
rect 7198 3895 9060 3910
rect 9063 3895 9077 3910
rect 7198 3874 9077 3895
rect 9092 3874 9131 3910
rect 9186 3908 9232 3910
rect 9192 3874 9226 3908
rect 7198 3863 9078 3874
rect 6072 3859 9078 3863
rect 6072 3857 8655 3859
rect 3734 3846 8655 3857
rect 3193 3829 3228 3836
rect 3270 3829 3358 3836
rect 3455 3830 8655 3846
rect 3455 3829 8720 3830
rect 3193 3734 3227 3829
rect 3285 3819 3297 3829
rect 3472 3827 6918 3829
rect 3472 3823 5929 3827
rect 3285 3796 3347 3819
rect 3293 3786 3347 3796
rect 3351 3767 3385 3768
rect 3339 3761 3397 3767
rect 3339 3734 3351 3761
rect 3472 3756 4403 3823
rect 4408 3817 5930 3823
rect 5931 3817 6918 3827
rect 4408 3781 6918 3817
rect 6931 3804 6972 3829
rect 7003 3816 7125 3829
rect 7019 3810 7125 3816
rect 7145 3810 7179 3829
rect 7198 3810 8720 3829
rect 7019 3804 8720 3810
rect 4408 3780 5864 3781
rect 5868 3780 6918 3781
rect 4408 3778 6918 3780
rect 4408 3756 5811 3778
rect 3472 3749 5811 3756
rect 3472 3743 4448 3749
rect 3455 3740 4448 3743
rect 4449 3740 5811 3749
rect 3455 3734 5811 3740
rect 144 3706 3174 3734
rect 144 3688 622 3706
rect 650 3702 698 3706
rect 711 3704 2067 3706
rect 644 3690 698 3702
rect 638 3688 698 3690
rect 144 3661 570 3688
rect 602 3684 698 3688
rect 602 3662 684 3684
rect 704 3674 705 3704
rect 711 3700 798 3704
rect 726 3696 798 3700
rect 732 3690 733 3696
rect 738 3690 798 3696
rect 726 3688 798 3690
rect 799 3688 2067 3704
rect 726 3684 786 3688
rect 726 3674 784 3684
rect 798 3674 833 3688
rect 840 3684 2067 3688
rect 852 3674 2067 3684
rect 726 3663 2067 3674
rect 726 3662 772 3663
rect 778 3662 2067 3663
rect 596 3661 2067 3662
rect 144 3655 2067 3661
rect 144 3654 564 3655
rect 144 3651 569 3654
rect 144 3643 570 3651
rect 596 3643 2067 3655
rect 144 3633 2067 3643
rect 2081 3702 2120 3706
rect 2081 3674 2121 3702
rect 2127 3688 3174 3706
rect 3175 3706 5811 3734
rect 5817 3767 6918 3778
rect 6937 3782 6971 3804
rect 7025 3795 8748 3804
rect 7025 3788 7179 3795
rect 7187 3788 8748 3795
rect 7025 3786 8748 3788
rect 6937 3767 6972 3782
rect 6975 3767 7033 3772
rect 5817 3766 5878 3767
rect 5880 3766 6926 3767
rect 5817 3730 5864 3766
rect 5878 3761 6926 3766
rect 6937 3766 7033 3767
rect 5878 3734 6930 3761
rect 6937 3734 6995 3766
rect 7004 3734 7037 3766
rect 7038 3734 7072 3786
rect 7091 3776 8748 3786
rect 7091 3768 7125 3776
rect 7091 3767 7129 3768
rect 7083 3761 7141 3767
rect 7145 3761 7179 3776
rect 7079 3742 7179 3761
rect 7079 3734 7125 3742
rect 7145 3734 7179 3742
rect 7198 3753 8748 3776
rect 7198 3740 8061 3753
rect 8106 3740 8147 3753
rect 8199 3740 8748 3753
rect 7198 3734 8159 3740
rect 5817 3726 5870 3730
rect 5878 3726 8159 3734
rect 5817 3725 5882 3726
rect 5817 3706 5870 3725
rect 3175 3702 5870 3706
rect 5890 3722 8159 3726
rect 5890 3702 8174 3722
rect 3175 3700 5876 3702
rect 2127 3686 2215 3688
rect 2234 3686 3174 3688
rect 2127 3677 3174 3686
rect 2127 3674 2195 3677
rect 2200 3674 2280 3677
rect 2288 3674 2322 3677
rect 2328 3674 3174 3677
rect 2081 3633 2120 3674
rect 2127 3673 3174 3674
rect 2127 3652 2215 3673
rect 2234 3652 3174 3673
rect 2127 3633 3174 3652
rect 144 3586 3174 3633
rect 144 3582 684 3586
rect 144 3578 696 3582
rect 144 3569 698 3578
rect 707 3569 848 3586
rect 144 3550 644 3569
rect 167 3530 201 3550
rect 167 3502 188 3530
rect 190 3519 201 3530
rect 193 3502 201 3519
rect 227 3530 644 3550
rect 646 3532 698 3569
rect 713 3568 848 3569
rect 713 3556 726 3568
rect 738 3565 848 3568
rect 770 3560 848 3565
rect 738 3558 848 3560
rect 852 3564 1701 3586
rect 1717 3575 1731 3586
rect 1740 3581 2215 3586
rect 2222 3585 2294 3586
rect 1745 3578 2215 3581
rect 2240 3584 2294 3585
rect 2348 3584 3174 3586
rect 2240 3580 3174 3584
rect 2261 3578 3174 3580
rect 1745 3575 2184 3578
rect 2190 3575 2224 3578
rect 1717 3564 1732 3575
rect 1745 3569 2224 3575
rect 1745 3564 2240 3569
rect 738 3556 804 3558
rect 713 3552 804 3556
rect 738 3550 804 3552
rect 852 3550 1697 3564
rect 1717 3560 2240 3564
rect 2261 3566 2291 3578
rect 2261 3560 2282 3566
rect 2292 3560 2333 3566
rect 738 3548 818 3550
rect 227 3502 275 3530
rect 281 3521 309 3530
rect 311 3525 415 3530
rect 327 3521 364 3525
rect 369 3521 403 3525
rect 369 3505 406 3521
rect 483 3517 678 3530
rect 685 3528 698 3532
rect 717 3531 818 3548
rect 717 3528 802 3531
rect 804 3528 818 3531
rect 685 3524 818 3528
rect 852 3542 1122 3550
rect 1143 3546 1697 3550
rect 1698 3552 2240 3560
rect 2348 3558 3174 3578
rect 2348 3556 2382 3558
rect 1698 3550 2224 3552
rect 1698 3546 2184 3550
rect 1143 3544 2184 3546
rect 2190 3548 2224 3550
rect 2296 3550 2382 3556
rect 2296 3548 2342 3550
rect 2190 3544 2199 3548
rect 2296 3544 2308 3548
rect 2348 3544 2382 3550
rect 852 3525 996 3542
rect 1143 3530 2382 3544
rect 1023 3525 1042 3530
rect 704 3520 744 3522
rect 745 3520 814 3524
rect 704 3517 745 3520
rect 483 3506 745 3517
rect 752 3517 814 3520
rect 752 3516 818 3517
rect 756 3510 814 3516
rect 852 3514 1026 3525
rect 341 3502 435 3505
rect 483 3502 644 3506
rect 144 3464 644 3502
rect 678 3500 745 3506
rect 852 3501 998 3514
rect 1045 3501 1075 3530
rect 1143 3527 1698 3530
rect 1745 3528 2291 3530
rect 2292 3528 2382 3530
rect 2402 3554 2436 3558
rect 2455 3554 2500 3558
rect 2402 3530 2500 3554
rect 2402 3528 2436 3530
rect 1745 3527 2413 3528
rect 1143 3519 2413 3527
rect 1143 3516 2380 3519
rect 1143 3512 2358 3516
rect 2421 3512 2436 3528
rect 1143 3508 2436 3512
rect 1143 3501 2445 3508
rect 657 3490 664 3492
rect 678 3490 842 3500
rect 852 3494 2445 3501
rect 678 3488 846 3490
rect 698 3479 704 3488
rect 710 3482 846 3488
rect 710 3479 758 3482
rect 698 3469 758 3479
rect 764 3479 792 3482
rect 798 3479 846 3482
rect 764 3469 846 3479
rect 852 3469 2184 3494
rect 698 3467 2184 3469
rect 2230 3491 2251 3494
rect 2230 3484 2286 3491
rect 2230 3469 2298 3484
rect 2328 3482 2382 3494
rect 2395 3482 2445 3494
rect 2230 3467 2310 3469
rect 2328 3468 2445 3482
rect 2455 3480 2500 3530
rect 2519 3480 2553 3558
rect 2613 3555 2635 3558
rect 2613 3548 2769 3555
rect 2619 3530 2769 3548
rect 2770 3539 3174 3558
rect 2771 3538 3174 3539
rect 3193 3538 3227 3700
rect 3325 3693 3463 3700
rect 3307 3689 3463 3693
rect 3295 3681 3463 3689
rect 3472 3681 5876 3700
rect 3229 3677 5876 3681
rect 3229 3674 5811 3677
rect 5817 3674 5876 3677
rect 5884 3700 8174 3702
rect 5884 3689 6971 3700
rect 5884 3686 5972 3689
rect 5978 3686 6971 3689
rect 5884 3681 6971 3686
rect 7017 3688 8159 3700
rect 8213 3698 8748 3740
rect 8213 3690 8430 3698
rect 7017 3683 8078 3688
rect 8113 3684 8145 3686
rect 7017 3682 7207 3683
rect 7216 3682 8078 3683
rect 7017 3681 8078 3682
rect 5884 3674 8078 3681
rect 3229 3666 5870 3674
rect 3229 3647 3281 3666
rect 3295 3647 3441 3666
rect 3472 3652 5870 3666
rect 5890 3673 8078 3674
rect 5890 3664 5972 3673
rect 5978 3666 8078 3673
rect 8168 3668 8179 3679
rect 5978 3664 7012 3666
rect 7038 3664 8078 3666
rect 5890 3652 8078 3664
rect 8177 3652 8179 3668
rect 8216 3652 8430 3690
rect 3472 3650 8145 3652
rect 3229 3538 3263 3647
rect 3295 3572 3317 3647
rect 3472 3630 8137 3650
rect 3395 3613 3433 3617
rect 3337 3572 3341 3613
rect 3395 3595 3455 3613
rect 3295 3538 3341 3572
rect 3371 3572 3375 3579
rect 3383 3572 3455 3595
rect 3371 3545 3455 3572
rect 3472 3595 6918 3630
rect 6924 3595 6971 3630
rect 3472 3578 6971 3595
rect 3472 3575 5970 3578
rect 3472 3569 5980 3575
rect 5984 3569 6971 3578
rect 3472 3565 6971 3569
rect 3472 3556 6082 3565
rect 6091 3558 6971 3565
rect 6091 3556 6192 3558
rect 3472 3555 6192 3556
rect 6193 3555 6251 3558
rect 3472 3550 6251 3555
rect 3383 3538 3437 3545
rect 2771 3530 3226 3538
rect 2597 3527 2663 3530
rect 2455 3475 2553 3480
rect 2665 3497 2723 3503
rect 2665 3484 2677 3497
rect 2771 3485 3174 3530
rect 2770 3484 3174 3485
rect 2665 3482 2711 3484
rect 2770 3482 3156 3484
rect 3159 3482 3174 3484
rect 3193 3529 3226 3530
rect 3229 3529 3471 3538
rect 3472 3535 6029 3550
rect 3472 3530 5970 3535
rect 5984 3530 6029 3535
rect 3472 3529 4808 3530
rect 3193 3501 4808 3529
rect 4811 3501 4814 3530
rect 4817 3501 4820 3530
rect 4841 3528 6029 3530
rect 6036 3543 6251 3550
rect 6036 3531 6126 3543
rect 6036 3528 6082 3531
rect 6086 3530 6126 3531
rect 6146 3530 6251 3543
rect 6084 3528 6244 3530
rect 4841 3527 6244 3528
rect 4841 3517 6146 3527
rect 4841 3501 6125 3517
rect 3193 3499 6125 3501
rect 6126 3509 6146 3517
rect 6156 3513 6244 3527
rect 6263 3529 6971 3558
rect 6973 3529 7007 3630
rect 7038 3626 8137 3630
rect 8164 3626 8430 3652
rect 7038 3618 8430 3626
rect 7038 3611 8078 3618
rect 7038 3592 8097 3611
rect 7038 3558 8121 3592
rect 8145 3561 8179 3618
rect 8186 3617 8430 3618
rect 8186 3586 8233 3617
rect 8199 3561 8233 3586
rect 8234 3570 8252 3602
rect 7038 3540 8109 3558
rect 8124 3548 8314 3561
rect 8124 3540 8333 3548
rect 8360 3540 8394 3617
rect 8585 3546 8748 3698
rect 8767 3736 8825 3742
rect 8767 3702 8779 3736
rect 8767 3696 8825 3702
rect 8956 3600 8971 3859
rect 8990 3633 9024 3859
rect 9043 3840 9078 3859
rect 9092 3840 9238 3874
rect 9136 3683 9194 3689
rect 9136 3649 9148 3683
rect 9136 3643 9194 3649
rect 9306 3643 9340 3910
rect 9325 3633 9340 3643
rect 9359 3633 9393 3910
rect 9466 3817 9500 4006
rect 9674 3987 9714 4006
rect 9790 3987 9816 4021
rect 9835 3987 9869 4528
rect 9981 4460 10039 4466
rect 9981 4426 9993 4460
rect 9981 4420 10039 4426
rect 10168 4211 10238 4581
rect 10350 4513 10408 4519
rect 10350 4479 10362 4513
rect 10350 4473 10408 4479
rect 10350 4313 10408 4319
rect 10350 4279 10362 4313
rect 10350 4273 10408 4279
rect 10168 4177 10239 4211
rect 10539 4196 10554 4615
rect 10573 4264 10607 4634
rect 10719 4566 10777 4572
rect 10719 4532 10731 4566
rect 10719 4526 10777 4532
rect 10719 4366 10777 4372
rect 10719 4332 10731 4366
rect 10719 4326 10777 4332
rect 10573 4230 10608 4264
rect 10908 4249 10923 4668
rect 10942 4317 10976 4687
rect 11088 4619 11146 4625
rect 11088 4585 11100 4619
rect 11088 4579 11146 4585
rect 11088 4419 11146 4425
rect 11088 4385 11100 4419
rect 11088 4379 11146 4385
rect 10942 4283 10977 4317
rect 11275 4283 11345 4740
rect 11457 4672 11515 4678
rect 11457 4638 11469 4672
rect 11457 4632 11515 4638
rect 11644 4423 11714 4793
rect 11826 4725 11884 4731
rect 11826 4691 11838 4725
rect 11826 4685 11884 4691
rect 11826 4525 11884 4531
rect 11826 4491 11838 4525
rect 11826 4485 11884 4491
rect 11644 4389 11715 4423
rect 12013 4389 12083 4846
rect 12195 4778 12253 4784
rect 12195 4744 12207 4778
rect 12195 4738 12253 4744
rect 12382 4529 12452 4899
rect 12564 4831 12622 4837
rect 12564 4797 12576 4831
rect 12564 4791 12622 4797
rect 12564 4631 12622 4637
rect 12564 4597 12576 4631
rect 12564 4591 12622 4597
rect 12382 4495 12453 4529
rect 12751 4495 12821 4952
rect 12933 4884 12991 4890
rect 12933 4850 12945 4884
rect 12933 4844 12991 4850
rect 12933 4576 12991 4582
rect 12933 4542 12945 4576
rect 12933 4536 12991 4542
rect 12195 4470 12253 4476
rect 12195 4436 12207 4470
rect 12382 4459 12435 4495
rect 12751 4459 12804 4495
rect 12195 4430 12253 4436
rect 11457 4364 11515 4370
rect 11457 4330 11469 4364
rect 11644 4353 11697 4389
rect 12013 4353 12066 4389
rect 11457 4324 11515 4330
rect 11275 4247 11328 4283
rect 10168 4141 10221 4177
rect 9937 4021 9977 4041
rect 10043 4021 10083 4041
rect 9937 4019 9983 4021
rect 9949 4015 9983 4019
rect 10037 4019 10083 4021
rect 10037 4015 10071 4019
rect 9568 3978 9580 3985
rect 9568 3972 9598 3978
rect 9568 3966 9601 3972
rect 9675 3966 9714 3987
rect 9728 3966 9768 3987
rect 9824 3981 10078 3987
rect 9824 3970 10065 3981
rect 9580 3962 9601 3966
rect 9694 3957 9709 3966
rect 9505 3938 9563 3944
rect 9566 3938 9567 3954
rect 9501 3904 9538 3938
rect 9551 3928 9567 3938
rect 9505 3898 9563 3904
rect 9608 3895 9609 3935
rect 9612 3919 9670 3925
rect 9612 3904 9624 3919
rect 9641 3904 9674 3919
rect 9612 3895 9674 3904
rect 9608 3885 9674 3895
rect 9612 3879 9670 3885
rect 9574 3857 9595 3861
rect 9574 3854 9607 3857
rect 9574 3851 9601 3854
rect 9528 3845 9595 3851
rect 9528 3817 9561 3845
rect 9675 3817 9709 3957
rect 9728 3953 9763 3966
rect 9824 3953 10078 3970
rect 9466 3783 9720 3817
rect 9461 3677 9519 3706
rect 9549 3677 9607 3706
rect 9473 3673 9507 3677
rect 9561 3673 9595 3677
rect 9519 3652 9585 3664
rect 9675 3652 9709 3783
rect 9423 3639 9709 3652
rect 9423 3633 9458 3639
rect 8990 3618 9458 3633
rect 9479 3630 9709 3639
rect 9501 3629 9709 3630
rect 9490 3618 9709 3629
rect 8990 3597 9457 3618
rect 9505 3602 9517 3618
rect 9523 3602 9567 3608
rect 8990 3560 9005 3597
rect 9018 3560 9457 3597
rect 9501 3580 9567 3602
rect 9675 3590 9709 3618
rect 8990 3547 9457 3560
rect 9675 3560 9686 3571
rect 9694 3560 9709 3590
rect 7038 3530 8430 3540
rect 7038 3529 8334 3530
rect 6263 3527 8334 3529
rect 8360 3527 8394 3530
rect 8419 3527 8430 3530
rect 8585 3530 8971 3546
rect 8585 3527 8748 3530
rect 6263 3524 8494 3527
rect 6263 3514 8119 3524
rect 8145 3514 8494 3524
rect 6156 3509 6251 3513
rect 6126 3499 6251 3509
rect 3193 3497 6251 3499
rect 6263 3503 8494 3514
rect 3193 3494 6180 3497
rect 3193 3482 5970 3494
rect 5984 3491 6029 3494
rect 6038 3491 6082 3494
rect 6091 3491 6126 3494
rect 2665 3475 2723 3482
rect 2770 3475 5970 3482
rect 2455 3468 5970 3475
rect 2328 3467 5970 3468
rect 5974 3484 6030 3491
rect 6038 3484 6164 3491
rect 5974 3475 6164 3484
rect 6190 3475 6256 3497
rect 6263 3482 6649 3503
rect 6669 3482 6703 3503
rect 6710 3491 8494 3503
rect 8585 3512 8656 3527
rect 8936 3512 8971 3530
rect 6710 3490 8568 3491
rect 6714 3488 8568 3490
rect 8585 3488 8655 3512
rect 6714 3484 8655 3488
rect 6722 3482 8655 3484
rect 6263 3475 8655 3482
rect 8937 3493 8971 3512
rect 9018 3528 9457 3547
rect 9569 3550 9627 3556
rect 9569 3530 9581 3550
rect 9675 3530 9709 3560
rect 9565 3528 9583 3530
rect 9613 3528 9631 3530
rect 9675 3528 9686 3530
rect 9018 3519 9686 3528
rect 9018 3516 9653 3519
rect 9018 3508 9631 3516
rect 9018 3507 9663 3508
rect 9018 3500 9693 3507
rect 9694 3500 9709 3530
rect 9018 3494 9709 3500
rect 9728 3652 9762 3953
rect 9782 3817 9816 3953
rect 9835 3870 9869 3953
rect 9981 3938 9993 3953
rect 10010 3938 10043 3953
rect 10044 3952 10078 3953
rect 9981 3932 10039 3938
rect 10044 3904 10221 3952
rect 10061 3891 10221 3904
rect 9874 3885 9932 3891
rect 9870 3870 9907 3885
rect 10044 3870 10221 3891
rect 10412 3882 10447 3916
rect 9835 3836 10221 3870
rect 10413 3863 10447 3882
rect 9776 3804 9816 3817
rect 9842 3804 9876 3808
rect 9801 3802 9816 3804
rect 9805 3783 9816 3802
rect 9830 3802 9876 3804
rect 9930 3802 9964 3808
rect 9830 3783 9870 3802
rect 10044 3800 10221 3836
rect 10243 3814 10301 3820
rect 9842 3749 9850 3783
rect 9018 3493 9457 3494
rect 8937 3488 8948 3493
rect 8956 3488 8971 3493
rect 5974 3467 8655 3475
rect 698 3466 792 3467
rect 798 3466 8655 3467
rect 676 3464 767 3466
rect 144 3462 664 3464
rect 144 3460 644 3462
rect 698 3460 792 3464
rect 798 3460 8142 3466
rect 144 3458 8142 3460
rect 144 3446 2787 3458
rect 2788 3454 8142 3458
rect 8145 3454 8655 3466
rect 2788 3446 8655 3454
rect 8745 3446 8847 3478
rect 8937 3458 8971 3488
rect 8937 3450 8948 3458
rect 8956 3450 8971 3458
rect 8937 3446 8971 3450
rect 8990 3446 9457 3493
rect 9533 3469 9583 3494
rect 9525 3458 9583 3469
rect 9613 3469 9663 3494
rect 9728 3475 9773 3652
rect 9830 3624 9888 3653
rect 9918 3624 9976 3653
rect 10044 3635 10131 3800
rect 10243 3780 10255 3814
rect 10243 3774 10301 3780
rect 9842 3620 9876 3624
rect 9930 3620 9964 3624
rect 9888 3599 9954 3611
rect 10044 3599 10178 3635
rect 9792 3586 10178 3599
rect 9792 3571 9827 3586
rect 9848 3577 10178 3586
rect 9870 3576 10178 3577
rect 9859 3571 10178 3576
rect 9792 3565 10178 3571
rect 9792 3475 9826 3565
rect 9874 3543 9886 3565
rect 9892 3543 10042 3555
rect 9874 3537 10042 3543
rect 9892 3530 10042 3537
rect 9870 3527 9936 3530
rect 9938 3497 9996 3503
rect 9938 3484 9950 3497
rect 9938 3482 9984 3484
rect 10044 3482 10178 3565
rect 10199 3562 10257 3575
rect 10287 3562 10345 3575
rect 10413 3560 10424 3571
rect 10432 3560 10447 3863
rect 10413 3530 10447 3560
rect 10243 3524 10301 3530
rect 10243 3490 10255 3524
rect 10413 3519 10424 3530
rect 10243 3484 10301 3490
rect 10413 3488 10424 3499
rect 10413 3482 10427 3488
rect 10432 3482 10447 3530
rect 10466 3829 10501 3863
rect 10781 3829 10816 3863
rect 10466 3529 10500 3829
rect 10782 3810 10816 3829
rect 10612 3761 10670 3767
rect 10612 3727 10624 3761
rect 10612 3721 10670 3727
rect 10598 3681 10736 3711
rect 10502 3647 10554 3681
rect 10568 3647 10714 3681
rect 10782 3647 10790 3715
rect 10801 3681 10816 3810
rect 10835 3776 10870 3810
rect 11150 3776 11185 3810
rect 10835 3682 10869 3776
rect 11151 3757 11185 3776
rect 11537 3757 11590 3758
rect 10981 3708 11039 3714
rect 10981 3684 10993 3708
rect 10981 3682 10995 3684
rect 11025 3682 11027 3684
rect 11170 3682 11185 3757
rect 11204 3723 11239 3757
rect 11519 3723 11590 3757
rect 11204 3682 11238 3723
rect 11520 3722 11590 3723
rect 11537 3688 11608 3722
rect 10835 3681 11257 3682
rect 10817 3647 11257 3681
rect 10502 3529 10536 3647
rect 10568 3561 10590 3647
rect 10668 3613 10706 3617
rect 10610 3561 10614 3613
rect 10668 3595 10728 3613
rect 10568 3529 10626 3561
rect 10644 3545 10648 3579
rect 10656 3545 10728 3595
rect 10784 3561 10816 3647
rect 10656 3529 10714 3545
rect 10782 3529 10816 3561
rect 10818 3603 11257 3647
rect 11350 3655 11408 3661
rect 11350 3621 11362 3655
rect 11350 3615 11408 3621
rect 11537 3611 11607 3688
rect 11719 3620 11777 3626
rect 11336 3603 11474 3605
rect 11520 3603 11528 3609
rect 11537 3603 11626 3611
rect 10818 3529 11626 3603
rect 11719 3586 11731 3620
rect 11719 3580 11777 3586
rect 11705 3540 11843 3561
rect 11705 3539 11774 3540
rect 10466 3482 11626 3529
rect 9938 3475 9996 3482
rect 10044 3475 11626 3482
rect 11675 3514 11863 3539
rect 11889 3514 11923 3626
rect 11675 3480 11923 3514
rect 9613 3458 9671 3469
rect 9525 3446 9571 3458
rect 9625 3446 9671 3458
rect 9728 3458 11626 3475
rect 9728 3447 9773 3458
rect 9739 3446 9773 3447
rect 9792 3454 10000 3458
rect 9792 3446 10024 3454
rect 10061 3446 11626 3458
rect 144 3444 11626 3446
rect 144 3418 11643 3444
rect 11650 3418 11671 3480
rect 144 3412 11671 3418
rect 144 3406 6196 3412
rect 144 3399 2184 3406
rect 144 3394 1382 3399
rect 1383 3394 1429 3399
rect 1445 3398 1517 3399
rect 1445 3394 1583 3398
rect 144 3386 1436 3394
rect 144 3368 644 3386
rect 664 3373 1436 3386
rect 1444 3373 1494 3394
rect 144 3358 658 3368
rect 664 3367 1494 3373
rect 1517 3367 1583 3394
rect 1590 3383 2184 3399
rect 2252 3383 2320 3406
rect 1590 3379 2320 3383
rect 2328 3397 5970 3406
rect 2328 3389 2787 3397
rect 2788 3389 5970 3397
rect 2328 3382 5970 3389
rect 5995 3387 6082 3406
rect 6091 3397 6196 3406
rect 6208 3397 6297 3412
rect 6317 3406 9671 3412
rect 9694 3406 9709 3412
rect 6317 3400 9457 3406
rect 6317 3397 8852 3400
rect 6091 3394 8852 3397
rect 6084 3387 8852 3394
rect 5984 3382 8852 3387
rect 2328 3379 8852 3382
rect 1590 3372 8852 3379
rect 8919 3394 8930 3400
rect 8937 3394 8971 3400
rect 8919 3390 8971 3394
rect 8990 3390 9457 3400
rect 9525 3394 9540 3406
rect 9641 3394 9671 3406
rect 664 3364 1496 3367
rect 1517 3364 1584 3367
rect 144 3340 644 3358
rect 144 3332 658 3340
rect 664 3332 1382 3364
rect 144 3309 1382 3332
rect 1383 3309 1429 3364
rect 1436 3358 1496 3364
rect 1524 3363 1584 3364
rect 1590 3364 8886 3372
rect 1590 3363 5928 3364
rect 1525 3361 5928 3363
rect 1536 3358 5928 3361
rect 1436 3336 1511 3358
rect 1432 3330 1511 3336
rect 1517 3345 5928 3358
rect 1517 3330 2191 3345
rect 2197 3338 2312 3345
rect 1432 3309 1496 3330
rect 1536 3322 1584 3330
rect 1590 3322 2191 3330
rect 1536 3311 2191 3322
rect 2208 3311 2312 3338
rect 1536 3309 2312 3311
rect 144 3304 2312 3309
rect 2328 3329 5928 3345
rect 144 3298 2310 3304
rect 144 3296 658 3298
rect 144 3278 644 3296
rect 664 3295 2310 3298
rect 664 3284 710 3295
rect 711 3289 2310 3295
rect 2328 3289 5126 3329
rect 711 3285 732 3289
rect 745 3285 826 3289
rect 833 3285 2260 3289
rect 2264 3285 2298 3289
rect 711 3284 745 3285
rect 752 3284 833 3285
rect 840 3284 2260 3285
rect 664 3282 2260 3284
rect 650 3278 2260 3282
rect 144 3258 2260 3278
rect 2274 3267 2308 3271
rect 2310 3270 5126 3289
rect 5180 3319 5928 3329
rect 5931 3358 8886 3364
rect 5931 3354 5972 3358
rect 5984 3354 8886 3358
rect 5931 3353 8886 3354
rect 5931 3319 6082 3353
rect 6091 3330 6180 3353
rect 6091 3320 6130 3330
rect 5180 3289 6082 3319
rect 6084 3319 6130 3320
rect 6132 3319 6180 3330
rect 6084 3301 6180 3319
rect 6185 3338 6299 3353
rect 6185 3330 6297 3338
rect 6300 3330 8886 3353
rect 6185 3322 8886 3330
rect 6185 3301 6244 3322
rect 6084 3296 6244 3301
rect 6250 3296 8886 3322
rect 6084 3289 8886 3296
rect 5180 3285 6086 3289
rect 5180 3277 6029 3285
rect 5192 3271 6029 3277
rect 6038 3279 6086 3285
rect 6091 3279 8886 3289
rect 6038 3272 8886 3279
rect 8919 3358 9457 3390
rect 9459 3372 9521 3394
rect 9525 3385 9583 3394
rect 9525 3372 9584 3385
rect 9459 3364 9585 3372
rect 9613 3364 9671 3394
rect 9477 3358 9585 3364
rect 8919 3338 8971 3358
rect 8990 3338 9457 3358
rect 9525 3344 9585 3358
rect 8919 3330 9457 3338
rect 9505 3332 9585 3344
rect 8919 3273 8971 3330
rect 6038 3271 8179 3272
rect 5192 3270 8179 3271
rect 2310 3267 5145 3270
rect 144 3150 644 3258
rect 650 3246 704 3258
rect 705 3252 786 3258
rect 787 3257 2260 3258
rect 2262 3261 2320 3267
rect 2262 3257 2322 3261
rect 2328 3257 5145 3267
rect 787 3252 2258 3257
rect 2263 3255 5145 3257
rect 2268 3254 5145 3255
rect 705 3246 2258 3252
rect 650 3245 2258 3246
rect 650 3227 2248 3245
rect 650 3208 2185 3227
rect 650 3202 786 3208
rect 787 3202 798 3208
rect 799 3202 2185 3208
rect 650 3192 2185 3202
rect 650 3178 786 3192
rect 792 3178 793 3192
rect 799 3181 2185 3192
rect 2186 3200 2248 3227
rect 2274 3223 5145 3254
rect 2274 3210 4442 3223
rect 4450 3210 5145 3223
rect 2186 3196 2268 3200
rect 2274 3196 5145 3210
rect 2186 3181 5145 3196
rect 799 3178 5145 3181
rect 650 3176 5145 3178
rect 650 3150 4442 3176
rect 4450 3173 5145 3176
rect 4455 3156 5145 3173
rect 5150 3156 5184 3270
rect 5192 3268 8142 3270
rect 8145 3268 8179 3270
rect 5192 3258 8179 3268
rect 5192 3256 8142 3258
rect 8145 3256 8179 3258
rect 5192 3255 8179 3256
rect 5188 3215 8179 3255
rect 5188 3205 6244 3215
rect 6246 3210 8179 3215
rect 8181 3270 8886 3272
rect 8181 3210 8889 3270
rect 8898 3266 8971 3273
rect 6246 3205 8889 3210
rect 5188 3202 8889 3205
rect 5188 3192 6113 3202
rect 6118 3192 6252 3202
rect 5188 3189 6252 3192
rect 5188 3156 6256 3189
rect 4455 3155 6256 3156
rect 6263 3176 8889 3202
rect 6263 3170 8176 3176
rect 8181 3170 8889 3176
rect 6263 3156 8889 3170
rect 8894 3239 8971 3266
rect 8894 3156 8901 3239
rect 8919 3210 8971 3239
rect 8990 3222 9457 3330
rect 9501 3320 9585 3332
rect 9641 3320 9671 3364
rect 9501 3304 9671 3320
rect 9505 3298 9582 3304
rect 8986 3221 9457 3222
rect 8978 3210 9457 3221
rect 8919 3156 9457 3210
rect 4455 3153 6252 3155
rect 6263 3153 9457 3156
rect 4455 3150 9457 3153
rect 144 3140 9457 3150
rect 9459 3294 9493 3298
rect 9459 3273 9505 3294
rect 9525 3289 9582 3298
rect 9583 3289 9671 3304
rect 9459 3270 9499 3273
rect 9459 3245 9493 3270
rect 9504 3257 9505 3273
rect 9523 3285 9571 3289
rect 9583 3288 9609 3289
rect 9523 3276 9551 3285
rect 9583 3276 9593 3288
rect 9625 3285 9659 3289
rect 9523 3258 9595 3276
rect 9675 3270 9709 3406
rect 9739 3387 9773 3412
rect 9792 3387 9826 3412
rect 9906 3387 9940 3404
rect 9994 3387 10028 3404
rect 10061 3387 11671 3412
rect 9647 3266 9709 3270
rect 9547 3257 9595 3258
rect 9459 3140 9507 3245
rect 9547 3242 9607 3257
rect 9635 3251 9709 3266
rect 9549 3140 9551 3242
rect 9565 3192 9607 3242
rect 9609 3208 9631 3242
rect 9613 3202 9627 3208
rect 9592 3177 9607 3192
rect 9635 3174 9665 3251
rect 9561 3140 9595 3174
rect 9635 3140 9661 3174
rect 9675 3140 9709 3251
rect 9728 3378 11671 3387
rect 9728 3353 10040 3378
rect 10061 3370 11671 3378
rect 10043 3353 11671 3370
rect 11675 3411 11725 3480
rect 11775 3472 11821 3480
rect 11762 3454 11763 3459
rect 11775 3454 11835 3472
rect 11675 3361 11733 3411
rect 11751 3404 11755 3438
rect 11762 3412 11835 3454
rect 11763 3395 11821 3412
rect 11829 3404 11843 3412
rect 11827 3395 11843 3404
rect 11763 3378 11845 3395
rect 11763 3372 11841 3378
rect 11763 3361 11821 3372
rect 11675 3359 11757 3361
rect 11763 3359 11845 3361
rect 11687 3357 11721 3359
rect 11723 3357 11757 3359
rect 11769 3357 11809 3359
rect 11811 3357 11845 3359
rect 11687 3355 11769 3357
rect 11775 3355 11857 3357
rect 9728 3249 9773 3353
rect 9792 3254 9826 3353
rect 9906 3319 9953 3332
rect 9846 3316 9900 3319
rect 9906 3316 9954 3319
rect 9846 3296 9954 3316
rect 9979 3314 9994 3348
rect 10010 3330 10040 3353
rect 9894 3291 9954 3296
rect 9874 3285 9954 3291
rect 9836 3266 9857 3270
rect 9836 3254 9863 3266
rect 9792 3249 9863 3254
rect 9870 3265 9954 3285
rect 9997 3283 10040 3330
rect 10044 3283 11671 3353
rect 11711 3346 11769 3355
rect 11799 3347 11857 3355
rect 11799 3346 11851 3347
rect 11697 3344 11851 3346
rect 11697 3331 11845 3344
rect 11697 3312 11799 3331
rect 9994 3280 11671 3283
rect 9870 3251 9956 3265
rect 9874 3249 9891 3251
rect 9899 3249 9945 3251
rect 9952 3249 9956 3251
rect 9994 3249 10040 3280
rect 10044 3249 11671 3280
rect 9728 3236 11671 3249
rect 9728 3227 9982 3236
rect 10021 3227 11671 3236
rect 9728 3215 11671 3227
rect 9728 3153 9773 3215
rect 9792 3208 9857 3215
rect 9792 3181 9876 3208
rect 9899 3204 10042 3215
rect 9877 3181 9882 3204
rect 9792 3153 9882 3181
rect 9905 3163 9910 3204
rect 9911 3202 10042 3204
rect 9911 3195 9987 3202
rect 9911 3189 9996 3195
rect 9911 3181 10000 3189
rect 9911 3163 9998 3181
rect 9899 3155 9998 3163
rect 9899 3153 9987 3155
rect 9728 3147 9882 3153
rect 9884 3147 9998 3153
rect 9728 3140 9998 3147
rect 144 3123 9998 3140
rect 10021 3139 10042 3202
rect 10044 3210 11671 3215
rect 11711 3278 11799 3312
rect 11805 3319 11845 3331
rect 11855 3331 11873 3335
rect 11855 3319 11885 3331
rect 11711 3210 11791 3278
rect 11805 3210 11885 3319
rect 11889 3210 11923 3480
rect 10044 3176 11885 3210
rect 11891 3176 11923 3210
rect 11925 3418 11977 3480
rect 11925 3415 11987 3418
rect 12347 3415 12382 3433
rect 144 3112 2067 3123
rect 2072 3112 2132 3123
rect 2144 3114 5495 3123
rect 144 3110 2132 3112
rect 144 3106 2120 3110
rect 144 3102 610 3106
rect 650 3102 698 3106
rect 144 3100 616 3102
rect 144 3088 622 3100
rect 644 3090 704 3102
rect 711 3100 732 3106
rect 738 3090 798 3106
rect 638 3088 704 3090
rect 726 3088 798 3090
rect 799 3098 820 3106
rect 828 3102 2120 3106
rect 2134 3103 5495 3114
rect 5526 3103 5560 3123
rect 5562 3106 9235 3123
rect 5562 3103 5706 3106
rect 5717 3103 5811 3106
rect 5816 3103 5864 3106
rect 2134 3102 5864 3103
rect 828 3098 2067 3102
rect 799 3088 2067 3098
rect 144 3074 570 3088
rect 576 3084 610 3088
rect 638 3084 698 3088
rect 726 3084 786 3088
rect 799 3086 833 3088
rect 638 3074 684 3084
rect 726 3074 784 3084
rect 798 3074 833 3086
rect 840 3084 2067 3088
rect 852 3077 2070 3084
rect 2072 3077 2132 3102
rect 852 3074 2132 3077
rect 2134 3087 2268 3102
rect 2274 3096 5864 3102
rect 5869 3099 5880 3106
rect 5888 3103 9235 3106
rect 9306 3103 9340 3123
rect 9359 3122 9405 3123
rect 9423 3122 9998 3123
rect 9359 3114 9998 3122
rect 9359 3103 9394 3114
rect 9417 3106 9998 3114
rect 9417 3103 9629 3106
rect 5888 3099 9629 3103
rect 5869 3098 9629 3099
rect 5869 3096 6243 3098
rect 2274 3088 6243 3096
rect 2274 3087 4403 3088
rect 2134 3084 4403 3087
rect 4408 3084 4442 3088
rect 144 3062 625 3074
rect 635 3062 684 3074
rect 698 3062 2120 3074
rect 144 3060 2120 3062
rect 144 3043 570 3060
rect 596 3043 2120 3060
rect 2134 3062 2180 3084
rect 2183 3083 4398 3084
rect 2183 3077 2274 3083
rect 2276 3077 2278 3083
rect 2280 3077 4398 3083
rect 2183 3074 2278 3077
rect 2288 3074 2322 3077
rect 2328 3074 4398 3077
rect 2183 3062 4398 3074
rect 4466 3062 5876 3088
rect 5891 3087 6243 3088
rect 6263 3089 9629 3098
rect 6263 3088 9623 3089
rect 9635 3088 9998 3106
rect 6263 3087 8142 3088
rect 5891 3086 8142 3087
rect 5903 3082 6078 3086
rect 5931 3077 6078 3082
rect 5931 3074 5978 3077
rect 5984 3074 6025 3077
rect 5931 3073 6025 3074
rect 6032 3073 6067 3077
rect 5931 3062 5965 3073
rect 5976 3062 6067 3073
rect 6079 3062 8142 3086
rect 2134 3058 5876 3062
rect 2134 3052 5874 3058
rect 5880 3053 8142 3062
rect 5880 3052 6243 3053
rect 2134 3050 6243 3052
rect 2134 3043 4398 3050
rect 4433 3046 6243 3050
rect 144 3030 4398 3043
rect 144 2994 4399 3030
rect 4428 3028 6243 3046
rect 6287 3034 8142 3053
rect 6299 3030 8142 3034
rect 4428 3020 6052 3028
rect 6086 3024 6243 3028
rect 6098 3020 6243 3024
rect 4428 3018 6082 3020
rect 4428 3005 5914 3018
rect 4417 2994 5914 3005
rect 144 2986 4398 2994
rect 144 2981 684 2986
rect 144 2970 678 2981
rect 698 2978 2186 2986
rect 2220 2978 4398 2986
rect 4428 2980 4433 2994
rect 707 2975 2184 2978
rect 2236 2976 2240 2978
rect 707 2974 2186 2975
rect 707 2970 848 2974
rect 852 2970 2186 2974
rect 144 2950 696 2970
rect 698 2969 2186 2970
rect 2220 2970 2236 2975
rect 2278 2970 2282 2976
rect 2346 2974 4398 2978
rect 4442 2974 5914 2994
rect 2346 2970 4405 2974
rect 4455 2971 4650 2974
rect 4418 2970 4650 2971
rect 4656 2970 5914 2974
rect 2220 2969 4398 2970
rect 698 2968 782 2969
rect 784 2968 4398 2969
rect 698 2958 4398 2968
rect 698 2950 804 2958
rect 848 2952 2500 2958
rect 848 2950 2186 2952
rect 2190 2950 2500 2952
rect 167 2940 201 2950
rect 214 2940 644 2950
rect 646 2940 696 2950
rect 167 2930 696 2940
rect 167 2818 188 2930
rect 190 2919 201 2930
rect 193 2829 201 2919
rect 190 2818 201 2829
rect 167 2785 201 2818
rect 214 2920 696 2930
rect 726 2931 818 2950
rect 848 2946 2184 2950
rect 2190 2948 2224 2950
rect 852 2940 2184 2946
rect 726 2922 802 2931
rect 804 2924 818 2931
rect 828 2938 2184 2940
rect 2294 2938 2342 2950
rect 2348 2938 2382 2950
rect 2388 2940 2436 2950
rect 2441 2940 2500 2950
rect 2505 2940 2553 2958
rect 2583 2954 2587 2958
rect 2599 2954 4398 2958
rect 2388 2938 2438 2940
rect 828 2930 2438 2938
rect 2441 2930 2553 2940
rect 2556 2950 4398 2954
rect 4418 2967 4600 2970
rect 4418 2958 4599 2967
rect 4418 2953 4590 2958
rect 4400 2950 4590 2953
rect 4592 2950 4599 2958
rect 4602 2950 5914 2970
rect 2556 2938 5914 2950
rect 5931 3012 5965 3018
rect 5984 3014 6082 3018
rect 5984 3012 6090 3014
rect 5931 2990 5967 3012
rect 5984 3006 6082 3012
rect 6108 3011 6113 3020
rect 5972 2999 6082 3006
rect 6102 2999 6113 3011
rect 6132 3012 6243 3020
rect 6132 3009 6294 3012
rect 6300 3009 8142 3030
rect 6132 3004 8142 3009
rect 8145 3028 8179 3088
rect 8181 3046 9618 3088
rect 9635 3086 9672 3088
rect 9647 3082 9652 3086
rect 8181 3028 9611 3046
rect 8145 3026 9611 3028
rect 8145 3004 9618 3026
rect 6132 2999 9618 3004
rect 5972 2996 9618 2999
rect 5976 2994 9618 2996
rect 5976 2990 8142 2994
rect 5931 2970 5965 2990
rect 5982 2986 8142 2990
rect 5984 2970 6029 2986
rect 5931 2960 6029 2970
rect 6048 2977 8142 2986
rect 8145 2977 8179 2994
rect 8186 2986 9618 2994
rect 9675 2990 9719 3088
rect 9728 3036 9772 3088
rect 9792 3087 9826 3088
rect 9842 3087 9882 3088
rect 9899 3087 9998 3088
rect 10044 3122 11671 3176
rect 11733 3146 11751 3164
rect 11769 3156 11797 3176
rect 11767 3146 11797 3156
rect 11733 3130 11797 3146
rect 11801 3130 11873 3176
rect 11751 3122 11873 3130
rect 10044 3090 11885 3122
rect 10044 3087 11626 3090
rect 9792 3086 11626 3087
rect 9792 3078 9826 3086
rect 9781 3058 9826 3078
rect 9830 3064 11626 3086
rect 9830 3058 10960 3064
rect 9792 3053 10960 3058
rect 9842 3036 9898 3053
rect 9728 3020 9792 3036
rect 9852 3029 9898 3036
rect 9830 3024 9898 3029
rect 8198 2977 9618 2986
rect 6048 2972 6122 2977
rect 6126 2974 9618 2977
rect 6126 2972 8142 2974
rect 6048 2965 8142 2972
rect 6048 2960 6082 2965
rect 5931 2952 6088 2960
rect 5931 2939 5965 2952
rect 5984 2939 6029 2952
rect 6038 2948 6088 2952
rect 6048 2939 6088 2948
rect 6126 2955 6243 2965
rect 6249 2955 6283 2965
rect 6126 2943 6283 2955
rect 5931 2938 6029 2939
rect 6030 2938 6088 2939
rect 6132 2938 6283 2943
rect 2556 2930 6283 2938
rect 852 2929 2382 2930
rect 214 2917 678 2920
rect 704 2917 802 2922
rect 214 2916 818 2917
rect 852 2916 2380 2929
rect 214 2910 756 2916
rect 214 2908 744 2910
rect 752 2908 786 2910
rect 214 2906 786 2908
rect 214 2870 644 2906
rect 678 2898 786 2906
rect 852 2898 2376 2916
rect 2407 2910 2436 2930
rect 2398 2907 2436 2910
rect 2382 2898 2436 2907
rect 678 2890 756 2898
rect 852 2894 2436 2898
rect 852 2890 2184 2894
rect 2284 2890 2286 2891
rect 2348 2890 2382 2894
rect 678 2888 758 2890
rect 706 2879 758 2888
rect 798 2879 2184 2890
rect 2264 2883 2298 2890
rect 2250 2879 2298 2883
rect 2338 2879 2386 2890
rect 698 2870 758 2879
rect 786 2870 2184 2879
rect 214 2867 2184 2870
rect 2238 2869 2298 2879
rect 2326 2869 2386 2879
rect 2441 2885 2500 2930
rect 2505 2885 2553 2930
rect 2597 2927 2663 2930
rect 2614 2896 2648 2919
rect 2625 2894 2648 2896
rect 2614 2885 2648 2894
rect 2663 2885 2711 2907
rect 2748 2898 6243 2930
rect 2723 2885 2727 2897
rect 2757 2894 6243 2898
rect 2757 2890 5914 2894
rect 2757 2885 5915 2890
rect 2441 2869 5915 2885
rect 5942 2885 6243 2894
rect 6249 2885 6283 2930
rect 6300 2949 8142 2965
rect 8145 2971 8179 2974
rect 8198 2971 9618 2974
rect 8145 2953 9618 2971
rect 9685 2961 9719 2990
rect 9726 3014 9806 3020
rect 9726 2986 9772 3014
rect 9776 2986 9834 3014
rect 8144 2950 9618 2953
rect 8145 2949 9618 2950
rect 6300 2941 9618 2949
rect 6300 2911 8511 2941
rect 8567 2928 9618 2941
rect 9664 2939 9719 2961
rect 9728 2939 9772 2986
rect 9799 2984 9834 2986
rect 9799 2970 9829 2984
rect 9840 2977 9898 3024
rect 9900 3036 9987 3053
rect 9900 3024 9934 3036
rect 9940 3024 9987 3036
rect 9900 2977 9987 3024
rect 9799 2967 9816 2970
rect 9840 2967 9987 2977
rect 10044 3040 10960 3053
rect 10999 3058 11043 3064
rect 11059 3058 11085 3064
rect 10999 3046 11025 3058
rect 11057 3046 11105 3058
rect 11041 3040 11105 3046
rect 10044 3036 10967 3040
rect 11037 3036 11105 3040
rect 10044 2971 10987 3036
rect 11019 3030 11105 3036
rect 11026 3021 11083 3030
rect 11041 2980 11083 3021
rect 11091 2996 11105 3030
rect 9787 2962 9987 2967
rect 9799 2943 9816 2962
rect 9840 2943 9987 2962
rect 9786 2939 9816 2943
rect 9818 2939 9820 2943
rect 9840 2940 9898 2943
rect 9900 2940 9987 2943
rect 8567 2917 9660 2928
rect 9664 2927 9772 2939
rect 9784 2927 9832 2939
rect 6300 2909 8510 2911
rect 6300 2885 8511 2909
rect 5942 2880 8511 2885
rect 2238 2867 2310 2869
rect 2327 2867 2398 2869
rect 214 2858 2398 2867
rect 214 2856 1698 2858
rect 1703 2856 2398 2858
rect 2441 2858 5927 2869
rect 2441 2856 2500 2858
rect 2505 2856 2727 2858
rect 2748 2856 5927 2858
rect 5942 2860 8101 2880
rect 8110 2860 8142 2880
rect 5942 2856 8142 2860
rect 8144 2856 8511 2880
rect 8567 2905 9618 2917
rect 9619 2905 9649 2917
rect 8567 2894 9660 2905
rect 8567 2884 9618 2894
rect 214 2850 8511 2856
rect 214 2836 8512 2850
rect 8523 2836 8545 2864
rect 214 2831 8545 2836
rect 214 2830 8523 2831
rect 214 2821 8512 2830
rect 214 2812 8511 2821
rect 214 2786 886 2812
rect 890 2788 904 2812
rect 912 2804 1698 2812
rect 1731 2807 2436 2812
rect 1703 2806 2436 2807
rect 1703 2804 2184 2806
rect 912 2799 2184 2804
rect 912 2786 1436 2799
rect 214 2785 644 2786
rect 167 2782 644 2785
rect 167 2762 188 2782
rect 214 2768 644 2782
rect 216 2762 644 2768
rect 167 2751 199 2762
rect 205 2751 644 2762
rect 216 2678 644 2751
rect 650 2784 1436 2786
rect 650 2744 886 2784
rect 912 2773 1436 2784
rect 1444 2773 1494 2799
rect 1650 2780 2184 2799
rect 2204 2804 2219 2806
rect 2238 2804 2436 2806
rect 2446 2804 2500 2812
rect 2505 2804 2553 2812
rect 2204 2782 2438 2804
rect 2452 2797 2553 2804
rect 2568 2797 2602 2812
rect 2607 2797 2614 2812
rect 2619 2797 2667 2812
rect 2707 2804 2741 2812
rect 2748 2804 2767 2812
rect 2707 2797 2767 2804
rect 2774 2804 6131 2812
rect 6132 2804 6296 2812
rect 2774 2797 6296 2804
rect 6300 2797 6307 2812
rect 6311 2797 8511 2812
rect 1536 2776 1570 2777
rect 1650 2774 1698 2780
rect 1703 2774 2184 2780
rect 912 2772 1494 2773
rect 1524 2772 1582 2773
rect 1596 2772 1604 2774
rect 912 2768 1610 2772
rect 1634 2768 2184 2774
rect 912 2764 2184 2768
rect 912 2758 1698 2764
rect 912 2750 1610 2758
rect 912 2749 1412 2750
rect 912 2748 1382 2749
rect 904 2744 1382 2748
rect 650 2738 1382 2744
rect 1400 2738 1406 2749
rect 1420 2740 1610 2750
rect 1650 2740 1698 2758
rect 1420 2738 1698 2740
rect 650 2729 1416 2738
rect 650 2695 874 2729
rect 650 2678 710 2695
rect 712 2689 874 2695
rect 724 2685 732 2689
rect 738 2685 874 2689
rect 720 2680 874 2685
rect 720 2678 838 2680
rect 840 2678 874 2680
rect 216 2670 874 2678
rect 886 2690 1416 2729
rect 1436 2730 1698 2738
rect 1436 2694 1610 2730
rect 1650 2710 1698 2730
rect 1703 2710 2184 2764
rect 2196 2768 2438 2782
rect 2441 2789 8511 2797
rect 8567 2818 9685 2884
rect 8567 2804 9249 2818
rect 9316 2816 9685 2818
rect 9686 2875 9772 2927
rect 9786 2924 9832 2927
rect 9840 2937 9987 2940
rect 10033 2937 10987 2971
rect 11068 2965 11083 2980
rect 9840 2927 9898 2937
rect 9786 2913 9829 2924
rect 9786 2884 9832 2913
rect 9840 2912 9886 2927
rect 9900 2912 9987 2937
rect 9840 2909 9987 2912
rect 9840 2896 9898 2909
rect 9900 2896 9987 2909
rect 9840 2884 9987 2896
rect 9786 2875 9987 2884
rect 10044 2928 10987 2937
rect 11037 2928 11071 2962
rect 11151 2928 11185 3064
rect 10044 2920 11185 2928
rect 10044 2875 10051 2920
rect 9686 2841 9987 2875
rect 10010 2864 10051 2875
rect 10021 2852 10051 2864
rect 10054 2911 11185 2920
rect 10054 2909 10714 2911
rect 10054 2884 10708 2909
rect 10054 2855 10730 2884
rect 10782 2855 10816 2911
rect 10835 2855 10869 2911
rect 10899 2909 10903 2911
rect 10915 2909 11185 2911
rect 10899 2894 11185 2909
rect 10915 2856 10995 2894
rect 11025 2886 11083 2894
rect 11007 2856 11083 2886
rect 10915 2855 10937 2856
rect 11007 2855 11037 2856
rect 10054 2852 10749 2855
rect 10010 2850 10749 2852
rect 10010 2841 10764 2850
rect 9686 2820 9772 2841
rect 9786 2820 9829 2841
rect 9686 2816 9829 2820
rect 9832 2838 9886 2841
rect 9900 2838 9934 2841
rect 9832 2816 9934 2838
rect 8567 2789 9299 2804
rect 2441 2769 8494 2789
rect 8531 2780 9299 2789
rect 8531 2776 9196 2780
rect 9215 2776 9249 2780
rect 2441 2768 8516 2769
rect 2196 2764 8516 2768
rect 8531 2764 9271 2776
rect 2196 2758 9271 2764
rect 2196 2748 2436 2758
rect 2204 2744 2436 2748
rect 2441 2755 9271 2758
rect 2441 2753 8561 2755
rect 2441 2744 2556 2753
rect 2204 2740 2556 2744
rect 2568 2740 2667 2753
rect 2668 2740 2673 2753
rect 2694 2744 6296 2753
rect 2690 2740 6296 2744
rect 6300 2740 8561 2753
rect 2204 2738 2562 2740
rect 2204 2727 2436 2738
rect 2441 2733 2562 2738
rect 2568 2733 2602 2740
rect 2607 2733 2614 2740
rect 2441 2727 2614 2733
rect 2204 2726 2614 2727
rect 2619 2726 2667 2740
rect 2673 2738 8561 2740
rect 2673 2730 6131 2738
rect 1650 2708 2184 2710
rect 1650 2704 2206 2708
rect 2214 2704 2436 2726
rect 1650 2699 2436 2704
rect 1650 2698 2240 2699
rect 2250 2698 2436 2699
rect 1650 2695 2436 2698
rect 1650 2694 2250 2695
rect 886 2676 1426 2690
rect 1436 2676 2250 2694
rect 2252 2689 2436 2695
rect 2264 2688 2336 2689
rect 2264 2685 2320 2688
rect 2352 2685 2386 2689
rect 886 2672 2250 2676
rect 216 2668 872 2670
rect 886 2668 1588 2672
rect 216 2658 886 2668
rect 912 2664 1588 2668
rect 1589 2666 1614 2672
rect 1650 2667 2250 2672
rect 2296 2679 2320 2685
rect 2388 2680 2436 2689
rect 2296 2676 2356 2679
rect 2360 2676 2436 2680
rect 2441 2676 2500 2726
rect 2505 2704 2556 2726
rect 2568 2722 2602 2726
rect 2502 2696 2568 2704
rect 2583 2702 2598 2711
rect 2582 2700 2598 2702
rect 2607 2705 2667 2726
rect 2690 2727 6131 2730
rect 6132 2735 8561 2738
rect 6132 2730 8480 2735
rect 6132 2727 6296 2730
rect 2690 2726 6296 2727
rect 2690 2722 6131 2726
rect 2690 2717 5927 2722
rect 5931 2717 6128 2722
rect 6132 2719 6296 2726
rect 2607 2698 2671 2705
rect 2590 2696 2671 2698
rect 2690 2699 6128 2717
rect 6131 2714 6296 2719
rect 6300 2719 8480 2730
rect 6300 2714 8141 2719
rect 6131 2704 8141 2714
rect 8142 2704 8480 2719
rect 8550 2734 8561 2735
rect 8567 2752 9271 2755
rect 8567 2734 9208 2752
rect 8550 2731 9208 2734
rect 9215 2748 9271 2752
rect 9281 2748 9315 2752
rect 8550 2717 9196 2731
rect 2296 2671 2500 2676
rect 2274 2667 2500 2671
rect 1589 2664 1628 2666
rect 912 2661 1628 2664
rect 912 2660 1602 2661
rect 216 2554 644 2658
rect 650 2656 684 2658
rect 690 2656 698 2658
rect 650 2584 698 2656
rect 720 2652 786 2658
rect 788 2656 860 2658
rect 788 2652 874 2656
rect 725 2642 874 2652
rect 738 2615 874 2642
rect 738 2608 886 2615
rect 738 2584 786 2608
rect 792 2602 814 2608
rect 820 2602 886 2608
rect 826 2584 886 2602
rect 650 2580 886 2584
rect 912 2586 1382 2660
rect 1392 2593 1528 2660
rect 1536 2654 1602 2660
rect 1604 2654 1628 2661
rect 1536 2620 1628 2654
rect 1534 2595 1628 2620
rect 1534 2593 1562 2595
rect 1392 2589 1474 2593
rect 1392 2586 1452 2589
rect 912 2580 1452 2586
rect 650 2556 1452 2580
rect 1462 2580 1474 2589
rect 1480 2592 1534 2593
rect 1536 2592 1562 2593
rect 1480 2583 1528 2592
rect 1534 2589 1562 2592
rect 1534 2583 1544 2589
rect 1480 2580 1544 2583
rect 1550 2580 1562 2589
rect 1568 2580 1628 2595
rect 1462 2579 1628 2580
rect 650 2554 1386 2556
rect 216 2548 1386 2554
rect 216 2544 1383 2548
rect 1392 2544 1452 2556
rect 1458 2570 1560 2579
rect 1568 2570 1628 2579
rect 1650 2658 2220 2667
rect 2230 2664 2250 2667
rect 2261 2666 2500 2667
rect 2505 2695 2553 2696
rect 2590 2695 2673 2696
rect 2505 2670 2673 2695
rect 2690 2695 6116 2699
rect 6131 2696 8480 2704
rect 2690 2685 6082 2695
rect 6128 2692 6131 2696
rect 6125 2691 6131 2692
rect 6132 2693 8480 2696
rect 6132 2691 8499 2693
rect 6125 2685 6130 2691
rect 6131 2685 8499 2691
rect 2690 2680 6106 2685
rect 6125 2680 8499 2685
rect 8516 2687 9196 2717
rect 8516 2683 8565 2687
rect 8567 2683 9196 2687
rect 2505 2668 2568 2670
rect 2505 2666 2553 2668
rect 2585 2666 2678 2670
rect 2261 2664 2436 2666
rect 2230 2661 2436 2664
rect 1650 2656 2232 2658
rect 1650 2578 2234 2656
rect 2261 2642 2436 2661
rect 2240 2592 2250 2620
rect 2262 2608 2436 2642
rect 2262 2601 2358 2608
rect 2360 2601 2436 2608
rect 2262 2578 2436 2601
rect 1650 2570 2436 2578
rect 1458 2550 2436 2570
rect 2441 2664 2553 2666
rect 2441 2661 2570 2664
rect 2582 2661 2678 2666
rect 2441 2645 2596 2661
rect 2597 2651 2678 2661
rect 2690 2658 8499 2680
rect 8550 2682 9196 2683
rect 9215 2715 9242 2748
rect 9244 2715 9315 2748
rect 9215 2682 9315 2715
rect 8550 2666 9190 2682
rect 2690 2654 4428 2658
rect 2624 2646 2678 2651
rect 2701 2646 2706 2654
rect 2721 2648 4428 2654
rect 2719 2646 4428 2648
rect 2624 2645 4428 2646
rect 2441 2608 2602 2645
rect 2618 2636 4428 2645
rect 2618 2626 2701 2636
rect 2723 2633 4428 2636
rect 2721 2632 4428 2633
rect 2618 2623 2725 2626
rect 2734 2623 4428 2632
rect 2618 2620 4428 2623
rect 4436 2649 8141 2658
rect 8145 2649 8499 2658
rect 4436 2643 8499 2649
rect 8519 2663 9190 2666
rect 9215 2663 9230 2682
rect 9244 2663 9315 2682
rect 9316 2738 9645 2816
rect 9685 2805 9832 2816
rect 9665 2759 9832 2805
rect 9665 2746 9733 2759
rect 9738 2750 9787 2759
rect 9807 2755 9820 2759
rect 9738 2746 9814 2750
rect 9665 2738 9814 2746
rect 9316 2727 9618 2738
rect 9685 2727 9814 2738
rect 9835 2738 9934 2816
rect 9835 2731 9887 2738
rect 9840 2727 9887 2731
rect 9316 2726 9887 2727
rect 9316 2663 9618 2726
rect 8519 2648 9230 2663
rect 9247 2658 9618 2663
rect 8519 2646 9190 2648
rect 8519 2643 8845 2646
rect 4436 2632 8845 2643
rect 8906 2639 9190 2646
rect 4436 2622 8839 2632
rect 4436 2620 8838 2622
rect 2618 2617 8518 2620
rect 8519 2619 8838 2620
rect 8519 2617 8849 2619
rect 2618 2609 8849 2617
rect 2441 2604 2603 2608
rect 2618 2605 8480 2609
rect 2441 2592 2609 2604
rect 2618 2602 8482 2605
rect 8550 2603 8849 2609
rect 2618 2592 2725 2602
rect 2734 2592 8482 2602
rect 8549 2601 8849 2603
rect 2441 2550 2603 2592
rect 1458 2546 2603 2550
rect 1476 2545 2603 2546
rect 1480 2544 2603 2545
rect 2624 2583 8482 2592
rect 8537 2583 8851 2601
rect 2624 2576 8851 2583
rect 2624 2574 6166 2576
rect 2624 2570 2727 2574
rect 2624 2556 2734 2570
rect 2757 2556 6166 2574
rect 2624 2555 6166 2556
rect 2624 2544 2703 2555
rect 2727 2550 6166 2555
rect 6167 2570 8141 2576
rect 8156 2570 8851 2576
rect 8906 2570 8907 2639
rect 8919 2630 9190 2639
rect 9247 2630 9271 2658
rect 6167 2566 8907 2570
rect 8918 2593 9190 2630
rect 8918 2570 9052 2593
rect 9055 2592 9074 2593
rect 9108 2573 9154 2593
rect 9253 2592 9271 2630
rect 9281 2592 9299 2658
rect 9327 2632 9618 2658
rect 9333 2628 9618 2632
rect 9333 2610 9601 2628
rect 9607 2617 9618 2628
rect 9685 2722 9787 2726
rect 9685 2718 9772 2722
rect 9685 2712 9788 2718
rect 9799 2712 9829 2726
rect 9685 2628 9719 2712
rect 9726 2700 9829 2712
rect 9840 2722 9852 2726
rect 9840 2706 9844 2722
rect 9866 2702 9886 2726
rect 9726 2688 9806 2700
rect 9726 2687 9772 2688
rect 9776 2687 9806 2688
rect 9726 2678 9806 2687
rect 9730 2672 9788 2678
rect 9685 2617 9696 2628
rect 9704 2610 9719 2628
rect 9738 2662 9772 2672
rect 9738 2644 9753 2662
rect 9761 2651 9772 2662
rect 9856 2649 9875 2693
rect 9900 2683 9934 2738
rect 9940 2812 9987 2841
rect 10054 2823 10764 2841
rect 10782 2831 11041 2855
rect 10054 2821 10782 2823
rect 10787 2821 11041 2831
rect 10054 2812 10725 2821
rect 9940 2769 10725 2812
rect 10782 2793 10826 2821
rect 10835 2802 10869 2821
rect 10981 2818 11041 2821
rect 10977 2802 11041 2818
rect 11151 2802 11185 2894
rect 11204 3011 11626 3064
rect 11637 3088 11885 3090
rect 11891 3088 11923 3122
rect 11204 2841 11618 3011
rect 11204 2805 11607 2841
rect 11204 2802 11238 2805
rect 11306 2803 11364 2805
rect 11376 2803 11452 2805
rect 11520 2804 11607 2805
rect 11637 2822 11671 3088
rect 11751 3080 11797 3088
rect 11751 3054 11785 3080
rect 11833 3062 11885 3088
rect 11697 3028 11785 3054
rect 11839 3028 11885 3062
rect 11889 3028 11923 3088
rect 11925 3077 12023 3415
rect 12311 3400 12382 3415
rect 12311 3283 12381 3400
rect 12493 3332 12551 3338
rect 12493 3298 12505 3332
rect 12493 3292 12551 3298
rect 12124 3277 12182 3283
rect 12124 3243 12136 3277
rect 12124 3237 12182 3243
rect 12294 3209 12381 3283
rect 13797 3215 13832 3249
rect 12068 3193 12126 3207
rect 12068 3173 12092 3193
rect 12180 3173 12214 3207
rect 12080 3139 12226 3173
rect 12294 3156 12392 3209
rect 13798 3196 13832 3215
rect 12080 3115 12094 3139
rect 11925 3028 12040 3077
rect 12136 3043 12198 3077
rect 12164 3037 12198 3043
rect 12294 3037 12733 3156
rect 13113 3103 13148 3121
rect 13077 3088 13148 3103
rect 11693 2994 11885 3028
rect 11739 2986 11799 2994
rect 11739 2971 11796 2986
rect 11855 2971 11885 2994
rect 11737 2967 11785 2971
rect 11797 2970 11823 2971
rect 11737 2958 11763 2967
rect 11797 2958 11805 2970
rect 11855 2967 11873 2971
rect 11687 2939 11705 2943
rect 11737 2940 11809 2958
rect 11761 2939 11809 2940
rect 11675 2822 11725 2939
rect 11761 2924 11821 2939
rect 11779 2874 11821 2924
rect 11829 2890 11843 2924
rect 11806 2859 11821 2874
rect 11775 2822 11809 2856
rect 11889 2822 11923 3026
rect 11942 2905 12040 3028
rect 12120 2975 12154 3003
rect 12294 2975 12308 3037
rect 12108 2941 12254 2975
rect 12120 2905 12154 2941
rect 11953 2840 12040 2905
rect 12152 2871 12210 2877
rect 12152 2842 12164 2871
rect 12311 2852 12733 3037
rect 12744 3033 12779 3067
rect 12152 2840 12186 2842
rect 11953 2837 12186 2840
rect 11953 2831 12210 2837
rect 11953 2822 12184 2831
rect 11637 2804 11661 2822
rect 11675 2804 11923 2822
rect 11970 2804 12184 2822
rect 11376 2802 11406 2803
rect 10835 2793 11054 2802
rect 10737 2769 10759 2793
rect 10782 2787 11075 2793
rect 10782 2777 10933 2787
rect 10941 2777 10971 2787
rect 10977 2777 11075 2787
rect 11151 2778 11410 2802
rect 10782 2770 10971 2777
rect 10973 2770 11075 2777
rect 10782 2769 11075 2770
rect 9940 2752 10759 2769
rect 10802 2768 11075 2769
rect 11094 2768 11151 2770
rect 11156 2768 11410 2778
rect 10802 2759 10879 2768
rect 10883 2759 10933 2768
rect 10802 2753 10933 2759
rect 9940 2744 10141 2752
rect 10155 2748 10267 2752
rect 10151 2744 10267 2748
rect 9940 2732 9987 2744
rect 10029 2736 10267 2744
rect 10029 2732 10255 2736
rect 9940 2702 10021 2732
rect 9896 2665 9934 2683
rect 9953 2666 10021 2702
rect 10054 2718 10255 2732
rect 10054 2713 10197 2718
rect 10054 2706 10201 2713
rect 10209 2706 10255 2718
rect 10265 2706 10267 2736
rect 10054 2702 10101 2706
rect 10054 2693 10097 2702
rect 10107 2693 10143 2706
rect 10054 2682 10143 2693
rect 10151 2697 10175 2706
rect 10183 2697 10185 2706
rect 10054 2675 10145 2682
rect 10151 2675 10185 2697
rect 10054 2666 10185 2675
rect 9884 2659 9942 2665
rect 9953 2659 9987 2666
rect 10054 2659 10175 2666
rect 10187 2659 10191 2706
rect 10197 2659 10267 2706
rect 10269 2726 10356 2752
rect 10269 2708 10355 2726
rect 10269 2666 10303 2708
rect 10309 2677 10355 2708
rect 10423 2694 10759 2752
rect 10803 2735 10933 2753
rect 10792 2716 10949 2735
rect 11007 2716 11041 2768
rect 11060 2716 11094 2768
rect 11170 2734 11195 2768
rect 10792 2706 11089 2716
rect 10792 2703 11094 2706
rect 10423 2682 10725 2694
rect 10771 2687 11094 2703
rect 10771 2682 10826 2687
rect 10835 2682 11094 2687
rect 10423 2681 10708 2682
rect 10771 2681 10839 2682
rect 10845 2681 10879 2682
rect 10309 2666 10356 2677
rect 10269 2659 10356 2666
rect 9884 2649 9934 2659
rect 9939 2654 10197 2659
rect 9939 2649 9987 2654
rect 10021 2650 10161 2654
rect 10209 2653 10356 2659
rect 9772 2644 9992 2649
rect 9738 2615 9992 2644
rect 10021 2644 10249 2650
rect 10265 2644 10356 2653
rect 10021 2636 10356 2644
rect 10021 2628 10303 2636
rect 10035 2625 10303 2628
rect 10054 2620 10141 2625
rect 10054 2619 10157 2620
rect 9738 2610 9772 2615
rect 9856 2610 9875 2615
rect 9900 2610 9968 2615
rect 9333 2598 9623 2610
rect 9680 2609 9968 2610
rect 10071 2609 10141 2619
rect 9680 2598 9900 2609
rect 9333 2593 9900 2598
rect 9333 2586 9530 2593
rect 9564 2592 9900 2593
rect 9905 2592 9934 2609
rect 9939 2592 9987 2609
rect 9564 2591 9987 2592
rect 9564 2586 9934 2591
rect 9333 2578 9934 2586
rect 9939 2578 9987 2591
rect 10054 2586 10065 2597
rect 10071 2592 10097 2609
rect 10107 2596 10141 2609
rect 10255 2606 10303 2625
rect 10322 2606 10356 2636
rect 10423 2606 10724 2681
rect 10771 2669 10879 2681
rect 10249 2596 10303 2606
rect 10308 2598 10356 2606
rect 10404 2603 10724 2606
rect 10793 2603 10879 2669
rect 10881 2681 10931 2682
rect 10881 2661 10939 2681
rect 10887 2659 10939 2661
rect 10991 2666 11003 2682
rect 11007 2666 11053 2682
rect 10991 2660 11049 2666
rect 10891 2657 10939 2659
rect 10404 2598 10725 2603
rect 10308 2596 10725 2598
rect 10107 2592 10725 2596
rect 10071 2591 10725 2592
rect 10073 2586 10088 2591
rect 10054 2578 10088 2586
rect 9333 2576 9992 2578
rect 9333 2573 9444 2576
rect 9530 2573 9896 2576
rect 9108 2570 9190 2573
rect 8918 2566 9190 2570
rect 6167 2556 9190 2566
rect 6167 2550 8516 2556
rect 2727 2545 8516 2550
rect 2727 2544 8128 2545
rect 8129 2544 8516 2545
rect 8537 2544 9190 2556
rect 9333 2557 9896 2573
rect 9930 2557 9992 2576
rect 10049 2557 10097 2578
rect 10107 2572 10725 2591
rect 10107 2562 10418 2572
rect 10423 2566 10725 2572
rect 10107 2557 10207 2562
rect 10255 2557 10387 2562
rect 9333 2556 10387 2557
rect 9333 2544 9992 2556
rect 10049 2544 10387 2556
rect 216 2523 10387 2544
rect 216 2443 230 2523
rect 286 2520 9973 2523
rect 9987 2520 10387 2523
rect 300 2510 10387 2520
rect 10440 2544 10725 2566
rect 10792 2587 10839 2603
rect 10845 2587 10879 2603
rect 10893 2628 10939 2657
rect 10959 2628 10961 2632
rect 10973 2628 10993 2632
rect 10893 2598 10913 2628
rect 10921 2603 10933 2628
rect 10925 2598 10933 2603
rect 10947 2598 10993 2628
rect 10893 2591 10939 2598
rect 10893 2587 10913 2591
rect 10925 2587 10927 2591
rect 10792 2578 10879 2587
rect 10792 2553 10883 2578
rect 10792 2544 10826 2553
rect 10833 2544 10879 2553
rect 10883 2544 10913 2553
rect 10440 2519 10913 2544
rect 10922 2538 10943 2544
rect 10947 2538 10997 2598
rect 10440 2510 10919 2519
rect 10925 2510 10935 2538
rect 10959 2534 10969 2538
rect 10973 2534 10993 2538
rect 440 2470 458 2504
rect 462 2500 522 2510
rect 542 2509 890 2510
rect 926 2509 1383 2510
rect 542 2506 1383 2509
rect 542 2500 610 2506
rect 652 2500 698 2506
rect 462 2498 491 2500
rect 542 2498 608 2500
rect 652 2498 696 2500
rect 476 2488 534 2498
rect 542 2488 622 2498
rect 652 2496 710 2498
rect 740 2496 798 2506
rect 828 2496 886 2506
rect 926 2500 1383 2506
rect 650 2494 710 2496
rect 738 2494 798 2496
rect 826 2494 886 2496
rect 652 2488 710 2494
rect 740 2488 798 2494
rect 828 2488 886 2494
rect 929 2498 1383 2500
rect 1392 2498 1452 2510
rect 1472 2508 1616 2510
rect 929 2496 1452 2498
rect 454 2468 458 2470
rect 564 2468 614 2488
rect 652 2468 702 2488
rect 364 2462 608 2468
rect 652 2462 696 2468
rect 740 2462 790 2488
rect 828 2486 878 2488
rect 798 2462 878 2486
rect 929 2462 1382 2496
rect 1392 2492 1452 2496
rect 1394 2486 1452 2492
rect 1482 2502 1616 2508
rect 1482 2496 1552 2502
rect 1562 2498 1616 2502
rect 1562 2496 1590 2498
rect 1482 2486 1540 2496
rect 1568 2495 1622 2496
rect 1625 2495 1628 2510
rect 1646 2506 1751 2510
rect 1568 2492 1628 2495
rect 1570 2486 1628 2492
rect 364 2450 1382 2462
rect 364 2448 692 2450
rect 696 2448 790 2450
rect 828 2448 878 2450
rect 364 2443 564 2448
rect 596 2443 652 2448
rect 216 2439 652 2443
rect 696 2439 740 2448
rect 890 2444 1382 2450
rect 1392 2482 1416 2486
rect 1582 2482 1590 2486
rect 1392 2444 1406 2482
rect 1528 2458 1646 2468
rect 1650 2458 1751 2506
rect 1646 2444 1751 2458
rect 746 2439 850 2440
rect 890 2439 1406 2444
rect 216 2437 663 2439
rect 685 2437 850 2439
rect 879 2437 1406 2439
rect 216 2428 1406 2437
rect 1427 2440 1645 2444
rect 1427 2434 1588 2440
rect 1590 2434 1645 2440
rect 1427 2433 1645 2434
rect 216 2370 630 2428
rect 912 2427 1406 2428
rect 912 2426 934 2427
rect 935 2426 1406 2427
rect 1430 2426 1634 2433
rect 1646 2426 1660 2444
rect 1668 2443 1751 2444
rect 1768 2483 1929 2510
rect 1948 2504 1962 2510
rect 2019 2504 2120 2510
rect 2150 2506 2603 2510
rect 1948 2494 1984 2504
rect 1768 2443 1828 2483
rect 1845 2476 1938 2483
rect 1845 2459 1850 2476
rect 1856 2449 1938 2476
rect 1856 2443 1918 2449
rect 1962 2443 1984 2494
rect 1990 2478 2012 2504
rect 2019 2484 2067 2504
rect 2019 2478 2070 2484
rect 1990 2472 2070 2478
rect 1990 2453 2012 2472
rect 2019 2468 2070 2472
rect 2072 2468 2120 2504
rect 2174 2487 2234 2506
rect 2262 2487 2334 2506
rect 2348 2496 2436 2506
rect 2360 2492 2436 2496
rect 2186 2483 2246 2487
rect 2274 2483 2334 2487
rect 2362 2486 2436 2492
rect 2188 2477 2246 2483
rect 2276 2477 2334 2483
rect 2374 2482 2436 2486
rect 2200 2474 2234 2477
rect 2288 2474 2322 2477
rect 2200 2473 2322 2474
rect 2019 2454 2130 2468
rect 2232 2464 2298 2473
rect 2388 2468 2436 2482
rect 2441 2504 2603 2506
rect 2624 2508 2691 2510
rect 2624 2504 2637 2508
rect 2441 2498 2609 2504
rect 2441 2497 2553 2498
rect 2555 2497 2609 2498
rect 2618 2497 2637 2504
rect 2638 2498 2691 2508
rect 2643 2497 2691 2498
rect 2757 2508 8141 2510
rect 2757 2506 6243 2508
rect 2757 2497 5863 2506
rect 2441 2494 5863 2497
rect 5874 2494 6243 2506
rect 2441 2488 6243 2494
rect 2441 2486 4433 2488
rect 2441 2482 2496 2486
rect 2441 2468 2489 2482
rect 2232 2462 2312 2464
rect 2378 2462 2489 2468
rect 2505 2468 4433 2486
rect 2505 2463 4398 2468
rect 4452 2464 5874 2488
rect 5891 2486 5919 2488
rect 5931 2487 5970 2488
rect 5979 2487 6018 2488
rect 5931 2486 6018 2487
rect 5903 2482 5908 2486
rect 2019 2453 2070 2454
rect 1990 2444 2070 2453
rect 1990 2443 2012 2444
rect 2019 2443 2070 2444
rect 2072 2443 2120 2454
rect 2136 2443 2489 2462
rect 2508 2458 4398 2463
rect 2519 2453 4398 2458
rect 2555 2446 2603 2453
rect 2643 2450 2691 2453
rect 2643 2446 2697 2450
rect 2569 2443 2603 2446
rect 2657 2443 2697 2446
rect 1668 2439 2489 2443
rect 2555 2441 2603 2443
rect 1668 2437 2185 2439
rect 2203 2437 2489 2439
rect 1668 2434 2489 2437
rect 2543 2434 2603 2441
rect 2643 2441 2697 2443
rect 1668 2428 2496 2434
rect 2555 2430 2615 2434
rect 2643 2430 2703 2441
rect 1668 2426 2170 2428
rect 2214 2426 2216 2428
rect 696 2412 768 2418
rect 912 2417 2170 2426
rect 912 2412 946 2417
rect 1328 2412 2170 2417
rect 2230 2418 2278 2428
rect 2230 2412 2332 2418
rect 2388 2412 2436 2428
rect 2438 2424 2496 2428
rect 2557 2424 2615 2430
rect 2657 2426 2703 2430
rect 2645 2424 2703 2426
rect 2757 2426 4398 2453
rect 4404 2438 4428 2464
rect 4452 2438 5857 2464
rect 4404 2436 5857 2438
rect 4404 2426 5860 2436
rect 5863 2426 5874 2464
rect 652 2402 768 2412
rect 652 2396 834 2402
rect 696 2394 834 2396
rect 848 2398 890 2412
rect 912 2398 1210 2412
rect 848 2396 1210 2398
rect 1254 2400 2170 2412
rect 1254 2396 1452 2400
rect 1562 2396 1590 2400
rect 1634 2396 2170 2400
rect 2174 2396 2332 2412
rect 2376 2396 2436 2412
rect 696 2388 782 2394
rect 710 2378 782 2388
rect 214 2340 630 2370
rect 726 2360 738 2370
rect 768 2368 782 2378
rect 784 2368 832 2394
rect 848 2374 1056 2396
rect 1312 2394 1378 2396
rect 912 2370 934 2374
rect 935 2370 946 2374
rect 1392 2370 1406 2396
rect 1438 2376 1452 2396
rect 1590 2370 1604 2396
rect 1646 2370 1660 2396
rect 770 2360 782 2368
rect 174 2298 188 2340
rect 214 2306 696 2340
rect 726 2336 788 2360
rect 798 2358 832 2368
rect 848 2346 1084 2370
rect 1284 2366 1406 2370
rect 1668 2356 2170 2396
rect 2204 2390 2332 2396
rect 2204 2370 2220 2390
rect 2228 2382 2332 2390
rect 2228 2380 2294 2382
rect 2332 2380 2336 2382
rect 2204 2362 2318 2370
rect 738 2334 788 2336
rect 740 2330 788 2334
rect 740 2318 756 2330
rect 760 2326 788 2330
rect 912 2337 946 2346
rect 1028 2340 1084 2346
rect 1334 2340 2170 2356
rect 1334 2337 1338 2340
rect 706 2310 756 2318
rect 214 2270 630 2306
rect 706 2298 782 2310
rect 912 2298 1351 2337
rect 1518 2333 1562 2340
rect 1590 2333 1634 2340
rect 1668 2338 2170 2340
rect 2388 2338 2436 2396
rect 1507 2322 1573 2333
rect 1579 2322 1645 2333
rect 1668 2329 2399 2338
rect 1668 2327 2387 2329
rect 1668 2322 2376 2327
rect 1357 2298 1368 2309
rect 1590 2298 1604 2322
rect 1650 2317 2376 2322
rect 1650 2310 2406 2317
rect 2407 2310 2436 2338
rect 1650 2304 2436 2310
rect 1650 2298 2170 2304
rect 2182 2298 2436 2304
rect 638 2270 694 2298
rect 706 2279 756 2298
rect 798 2279 832 2290
rect 698 2270 756 2279
rect 786 2270 844 2279
rect 214 2256 844 2270
rect 912 2268 1368 2298
rect 1650 2294 2436 2298
rect 2441 2412 2489 2424
rect 2569 2421 2603 2424
rect 2645 2422 2695 2424
rect 2645 2421 2725 2422
rect 2559 2420 2725 2421
rect 2559 2412 2584 2420
rect 2441 2409 2505 2412
rect 2556 2409 2584 2412
rect 2601 2412 2725 2420
rect 2601 2409 2734 2412
rect 2757 2409 5874 2426
rect 2441 2396 5874 2409
rect 912 2260 1351 2268
rect 1357 2260 1368 2268
rect 912 2256 1368 2260
rect 1458 2256 1560 2288
rect 1590 2256 1604 2268
rect 1650 2262 2170 2294
rect 2246 2279 2296 2294
rect 1650 2256 1684 2262
rect 1694 2258 2170 2262
rect 1703 2256 2170 2258
rect 2238 2268 2296 2279
rect 2326 2279 2376 2294
rect 2441 2285 2489 2396
rect 2505 2394 5874 2396
rect 2505 2392 4345 2394
rect 4350 2392 4398 2394
rect 2505 2375 4398 2392
rect 4452 2387 4526 2394
rect 4528 2387 4650 2394
rect 4442 2386 4650 2387
rect 4452 2381 4650 2386
rect 4464 2377 4650 2381
rect 2505 2285 2539 2375
rect 2559 2370 2647 2375
rect 2757 2374 4398 2375
rect 4428 2374 4650 2377
rect 2757 2370 4405 2374
rect 4466 2371 4650 2374
rect 2599 2365 2647 2370
rect 2738 2365 4405 2370
rect 2599 2364 4405 2365
rect 2542 2358 4405 2364
rect 2542 2350 4345 2358
rect 4350 2353 4405 2358
rect 4418 2367 4650 2371
rect 4418 2358 4578 2367
rect 4418 2353 4590 2358
rect 4350 2350 4590 2353
rect 4599 2350 4650 2367
rect 4655 2382 5874 2394
rect 5931 2424 5965 2486
rect 5984 2483 6018 2486
rect 6037 2487 6086 2488
rect 6098 2487 6243 2488
rect 6249 2498 8141 2508
rect 8156 2498 8497 2510
rect 6249 2488 8497 2498
rect 6249 2487 8141 2488
rect 6037 2486 8141 2487
rect 5984 2482 6025 2483
rect 5984 2474 6018 2482
rect 6037 2474 6072 2486
rect 5984 2458 6072 2474
rect 6079 2459 8141 2486
rect 6086 2458 8141 2459
rect 5984 2440 6042 2458
rect 6048 2453 8141 2458
rect 6098 2441 6243 2453
rect 5974 2430 6042 2440
rect 6086 2436 6243 2441
rect 5974 2424 6034 2430
rect 6086 2426 6101 2436
rect 6125 2426 6243 2436
rect 6287 2434 8141 2453
rect 6086 2424 6243 2426
rect 5931 2420 6034 2424
rect 5931 2419 6048 2420
rect 5931 2400 6032 2419
rect 5931 2392 5965 2400
rect 5968 2396 6032 2400
rect 5931 2390 5967 2392
rect 5972 2390 6032 2396
rect 4655 2350 5898 2382
rect 2542 2340 2755 2350
rect 2542 2322 2556 2340
rect 2583 2337 2663 2340
rect 2597 2327 2663 2337
rect 2584 2308 2598 2322
rect 2600 2306 2614 2319
rect 2634 2306 2648 2319
rect 2600 2285 2648 2306
rect 2663 2294 2686 2307
rect 2734 2298 2755 2340
rect 2757 2349 4405 2350
rect 4418 2349 5898 2350
rect 5931 2353 5965 2390
rect 5982 2387 6032 2390
rect 5982 2386 6048 2387
rect 5984 2367 6018 2386
rect 6055 2377 6090 2392
rect 6094 2377 6113 2424
rect 5931 2349 5974 2353
rect 5984 2349 6022 2367
rect 6043 2362 6113 2377
rect 6122 2412 6243 2424
rect 6297 2426 8141 2434
rect 8145 2426 8497 2488
rect 8550 2503 9623 2510
rect 9648 2504 9846 2510
rect 9880 2509 9920 2510
rect 8550 2469 9195 2503
rect 9333 2488 9623 2503
rect 9650 2498 9846 2504
rect 9869 2498 9920 2509
rect 9650 2496 9719 2498
rect 9650 2490 9734 2496
rect 9738 2490 9772 2498
rect 9661 2488 9772 2490
rect 9333 2477 9604 2488
rect 6122 2396 6254 2412
rect 6297 2399 8497 2426
rect 8525 2467 9195 2469
rect 9201 2469 9604 2477
rect 9201 2467 9249 2469
rect 8525 2437 9254 2467
rect 9272 2437 9604 2469
rect 9676 2468 9772 2488
rect 9672 2464 9772 2468
rect 9852 2470 9880 2498
rect 9886 2470 9920 2498
rect 9852 2466 9920 2470
rect 9846 2464 9920 2466
rect 9672 2456 9796 2464
rect 9672 2450 9734 2456
rect 9672 2440 9719 2450
rect 8525 2433 9604 2437
rect 8525 2423 9195 2433
rect 9201 2423 9235 2433
rect 6055 2353 6072 2362
rect 6028 2352 6072 2353
rect 6028 2349 6052 2352
rect 6055 2349 6072 2352
rect 2757 2341 5898 2349
rect 2757 2333 4790 2341
rect 2757 2324 4593 2333
rect 4599 2332 4790 2333
rect 4821 2332 4881 2341
rect 4599 2324 4881 2332
rect 4921 2331 4981 2341
rect 2757 2322 4881 2324
rect 2757 2315 4790 2322
rect 4821 2321 4881 2322
rect 4935 2321 4981 2331
rect 4821 2319 4879 2321
rect 2757 2294 4664 2315
rect 4666 2294 4790 2315
rect 4813 2308 4834 2319
rect 4835 2315 4949 2319
rect 4966 2317 4981 2321
rect 5024 2338 5898 2341
rect 5928 2339 6074 2349
rect 5928 2338 6022 2339
rect 6028 2338 6088 2339
rect 6122 2338 6243 2396
rect 5024 2320 6243 2338
rect 4835 2312 4961 2315
rect 4969 2312 4975 2317
rect 4835 2309 4981 2312
rect 2663 2285 2697 2294
rect 2757 2285 4357 2294
rect 2326 2268 2384 2279
rect 2238 2256 2292 2268
rect 2332 2256 2384 2268
rect 2441 2276 4357 2285
rect 4364 2290 4664 2294
rect 4364 2284 4398 2290
rect 4366 2276 4398 2284
rect 2441 2268 4398 2276
rect 2441 2256 2486 2268
rect 2505 2257 2713 2268
rect 2505 2256 2709 2257
rect 2734 2256 4398 2268
rect 214 2248 866 2256
rect 879 2252 4398 2256
rect 879 2248 4384 2252
rect 4388 2248 4398 2252
rect 4400 2282 4448 2290
rect 4482 2282 4664 2290
rect 4680 2290 4790 2294
rect 4680 2284 4767 2290
rect 4400 2280 4664 2282
rect 4683 2280 4767 2284
rect 4800 2281 4834 2308
rect 4847 2305 4909 2309
rect 4879 2297 4909 2305
rect 4935 2308 4961 2309
rect 4935 2305 4969 2308
rect 5024 2305 5874 2320
rect 5875 2305 5905 2320
rect 4901 2287 4902 2297
rect 4935 2290 4951 2305
rect 5024 2304 5912 2305
rect 5928 2304 6243 2320
rect 5024 2294 5916 2304
rect 5928 2294 6022 2304
rect 4865 2281 4874 2287
rect 4901 2281 4923 2287
rect 4400 2264 4767 2280
rect 4772 2268 4795 2280
rect 4800 2268 4823 2281
rect 4861 2274 4927 2281
rect 4930 2277 4951 2290
rect 4969 2281 4996 2290
rect 5024 2284 5874 2294
rect 5928 2284 5933 2293
rect 4861 2271 4996 2274
rect 4400 2252 4801 2264
rect 4400 2250 4767 2252
rect 4400 2248 4672 2250
rect 214 2238 872 2248
rect 879 2245 4550 2248
rect 214 2233 886 2238
rect 890 2233 4550 2245
rect 4558 2235 4672 2248
rect 4678 2246 4767 2250
rect 214 2232 4550 2233
rect 4564 2232 4672 2235
rect 214 2228 4672 2232
rect 4683 2236 4767 2246
rect 4779 2236 4801 2252
rect 4877 2247 4925 2271
rect 4891 2237 4925 2247
rect 4946 2240 4963 2271
rect 4683 2234 4801 2236
rect 4683 2231 4823 2234
rect 4955 2231 4996 2234
rect 4683 2230 4795 2231
rect 4683 2228 4767 2230
rect 214 2222 4767 2228
rect 214 2168 644 2222
rect 216 2084 644 2168
rect 650 2199 874 2222
rect 875 2199 1428 2222
rect 1590 2218 1604 2222
rect 1650 2218 1684 2222
rect 650 2184 1428 2199
rect 650 2154 886 2184
rect 912 2160 1428 2184
rect 1494 2182 1530 2188
rect 1582 2182 1684 2218
rect 1448 2173 1530 2182
rect 1536 2173 1684 2182
rect 1436 2168 1684 2173
rect 1436 2160 1511 2168
rect 1524 2160 1684 2168
rect 912 2159 1398 2160
rect 912 2154 1368 2159
rect 650 2148 1368 2154
rect 1428 2150 1684 2160
rect 1398 2148 1400 2149
rect 1429 2148 1684 2150
rect 650 2139 1402 2148
rect 650 2099 874 2139
rect 650 2084 698 2099
rect 710 2095 732 2099
rect 738 2086 786 2099
rect 798 2095 820 2099
rect 826 2090 874 2099
rect 216 2078 698 2084
rect 720 2078 786 2086
rect 788 2078 874 2090
rect 216 2070 874 2078
rect 886 2138 1402 2139
rect 886 2116 1400 2138
rect 1436 2132 1684 2148
rect 886 2098 1402 2116
rect 1436 2104 1604 2132
rect 1646 2120 1684 2132
rect 1703 2220 2422 2222
rect 2432 2220 2500 2222
rect 2505 2220 2668 2222
rect 1703 2216 2426 2220
rect 1703 2214 2205 2216
rect 1703 2204 2236 2214
rect 2238 2204 2426 2216
rect 2432 2214 2486 2220
rect 2500 2216 2668 2220
rect 2500 2214 2602 2216
rect 1703 2174 2438 2204
rect 2452 2197 2548 2214
rect 2554 2197 2602 2214
rect 2607 2197 2614 2216
rect 2619 2214 2636 2216
rect 2734 2214 2757 2222
rect 2619 2197 2653 2214
rect 2707 2197 2757 2214
rect 2774 2216 4767 2222
rect 4772 2216 4795 2230
rect 2774 2214 4795 2216
rect 2774 2203 4767 2214
rect 2774 2197 4758 2203
rect 2441 2188 4758 2197
rect 4800 2189 4823 2231
rect 4875 2221 4929 2231
rect 4930 2224 4996 2231
rect 5024 2228 5909 2284
rect 5918 2248 5933 2284
rect 5940 2288 6022 2294
rect 6028 2294 6088 2304
rect 6127 2298 6243 2304
rect 6142 2296 6243 2298
rect 6127 2294 6243 2296
rect 6297 2394 8510 2399
rect 6297 2371 8141 2394
rect 8145 2371 8179 2394
rect 8196 2387 8510 2394
rect 8196 2385 8497 2387
rect 8498 2385 8510 2387
rect 8196 2371 8510 2385
rect 8525 2396 9235 2423
rect 8525 2379 9195 2396
rect 6297 2324 8088 2371
rect 8094 2367 8129 2371
rect 8094 2324 8128 2367
rect 8145 2353 8510 2371
rect 8144 2349 8510 2353
rect 8531 2351 8532 2379
rect 8565 2375 9195 2379
rect 8547 2365 9195 2375
rect 8544 2351 9195 2365
rect 6297 2321 8128 2324
rect 6297 2311 7361 2321
rect 5940 2275 6018 2288
rect 6028 2285 6286 2294
rect 6297 2285 6975 2311
rect 6028 2280 6975 2285
rect 6976 2280 7003 2311
rect 7038 2294 7072 2311
rect 7091 2299 7149 2311
rect 7081 2294 7149 2299
rect 7155 2294 7361 2311
rect 7038 2290 7193 2294
rect 7199 2290 7232 2294
rect 7038 2289 7187 2290
rect 7205 2289 7232 2290
rect 7038 2281 7194 2289
rect 6028 2275 6964 2280
rect 5940 2266 6964 2275
rect 6984 2272 6991 2276
rect 7004 2272 7018 2276
rect 6972 2266 7018 2272
rect 5940 2265 7018 2266
rect 7038 2272 7081 2281
rect 7091 2272 7194 2281
rect 7038 2265 7194 2272
rect 7205 2268 7235 2289
rect 7205 2265 7228 2268
rect 7239 2265 7273 2294
rect 7283 2265 7339 2294
rect 5940 2262 6964 2265
rect 6972 2262 7339 2265
rect 5940 2256 7339 2262
rect 5940 2255 7283 2256
rect 7292 2255 7326 2256
rect 5940 2248 7326 2255
rect 4902 2196 4929 2221
rect 5024 2210 5719 2228
rect 5773 2220 5909 2228
rect 5742 2216 5909 2220
rect 5912 2241 7326 2248
rect 5912 2226 6286 2241
rect 6297 2230 6307 2241
rect 6309 2230 7326 2241
rect 6297 2226 7326 2230
rect 7360 2228 7361 2294
rect 7372 2294 8128 2321
rect 7372 2238 7394 2294
rect 7400 2292 8128 2294
rect 8132 2341 8510 2349
rect 7400 2290 8123 2292
rect 7400 2278 8101 2290
rect 8132 2286 8497 2341
rect 8565 2319 9195 2351
rect 7400 2266 7452 2278
rect 7460 2274 8101 2278
rect 7407 2234 7441 2266
rect 7460 2258 8094 2274
rect 8128 2258 8497 2286
rect 7460 2251 8077 2258
rect 7460 2246 8065 2251
rect 7450 2234 8065 2246
rect 7407 2228 8065 2234
rect 5912 2220 6102 2226
rect 6122 2220 6244 2226
rect 5912 2216 6244 2220
rect 5024 2206 5505 2210
rect 4983 2200 5505 2206
rect 5573 2203 5719 2210
rect 4983 2196 5452 2200
rect 5024 2189 5452 2196
rect 4787 2188 4945 2189
rect 2441 2178 4558 2188
rect 4564 2178 4596 2188
rect 1703 2168 2426 2174
rect 1703 2148 2432 2168
rect 1703 2120 2170 2148
rect 2190 2146 2432 2148
rect 2441 2163 4596 2178
rect 4602 2186 4945 2188
rect 4602 2164 4758 2186
rect 4787 2180 4945 2186
rect 4763 2179 4945 2180
rect 4763 2172 4973 2179
rect 5018 2178 5452 2189
rect 4763 2164 4987 2172
rect 4602 2163 4987 2164
rect 2441 2148 2548 2163
rect 2554 2148 2640 2163
rect 2190 2136 2438 2146
rect 2202 2132 2438 2136
rect 2204 2130 2384 2132
rect 2386 2130 2438 2132
rect 2204 2127 2438 2130
rect 2441 2142 2640 2148
rect 2650 2142 2653 2163
rect 2654 2142 2659 2163
rect 2707 2158 4987 2163
rect 2688 2154 4987 2158
rect 2676 2150 4987 2154
rect 5024 2150 5452 2178
rect 2441 2140 2666 2142
rect 2441 2138 2602 2140
rect 2441 2130 2539 2138
rect 2540 2133 2573 2138
rect 2585 2133 2602 2138
rect 2607 2133 2614 2140
rect 2540 2132 2614 2133
rect 2540 2130 2556 2132
rect 2561 2130 2614 2132
rect 2441 2127 2614 2130
rect 2204 2126 2614 2127
rect 2619 2129 2666 2140
rect 2676 2135 5452 2150
rect 2619 2126 2667 2129
rect 1646 2108 2170 2120
rect 2214 2114 2384 2126
rect 2214 2110 2230 2114
rect 1434 2102 1604 2104
rect 1650 2104 2170 2108
rect 2172 2104 2206 2108
rect 2214 2104 2232 2110
rect 1650 2102 2232 2104
rect 1434 2098 2232 2102
rect 2238 2099 2295 2114
rect 2296 2099 2384 2114
rect 2388 2122 2426 2126
rect 886 2090 1412 2098
rect 886 2076 1426 2090
rect 1434 2078 2218 2098
rect 2250 2095 2284 2099
rect 2296 2098 2322 2099
rect 1434 2076 2232 2078
rect 886 2072 1614 2076
rect 216 2059 872 2070
rect 886 2061 1368 2072
rect 1380 2061 1614 2072
rect 886 2060 1614 2061
rect 886 2059 1368 2060
rect 216 2058 1368 2059
rect 216 1954 630 2058
rect 638 2032 684 2058
rect 720 2054 786 2058
rect 720 2052 784 2054
rect 788 2052 860 2058
rect 726 2032 860 2052
rect 638 2000 664 2032
rect 738 2018 838 2032
rect 738 2012 800 2018
rect 738 2002 784 2012
rect 820 2002 838 2018
rect 778 2000 838 2002
rect 857 2000 872 2015
rect 638 1960 696 2000
rect 726 1984 872 2000
rect 726 1960 784 1984
rect 814 1980 872 1984
rect 912 1980 1368 2058
rect 1380 1980 1438 2060
rect 1442 2005 1520 2060
rect 1524 2034 1526 2060
rect 1530 2034 1614 2060
rect 1442 2002 1460 2005
rect 1448 1989 1460 2002
rect 1480 2002 1520 2005
rect 1526 2005 1614 2034
rect 1480 1996 1514 2002
rect 1526 1996 1556 2005
rect 1568 1996 1614 2005
rect 1468 1993 1514 1996
rect 1524 1993 1526 1996
rect 814 1960 1438 1980
rect 650 1954 664 1960
rect 857 1956 1438 1960
rect 1468 1980 1526 1993
rect 1536 1989 1548 1996
rect 1556 1980 1614 1996
rect 1650 2042 2232 2076
rect 2240 2064 2250 2092
rect 2296 2086 2306 2098
rect 2338 2095 2372 2099
rect 2260 2067 2308 2086
rect 2388 2080 2422 2122
rect 2360 2076 2422 2080
rect 2441 2078 2486 2126
rect 2260 2052 2320 2067
rect 1650 2032 1684 2042
rect 1694 2032 2232 2042
rect 1650 2028 2232 2032
rect 2262 2038 2320 2052
rect 2322 2038 2344 2052
rect 2348 2038 2422 2076
rect 1650 1996 2170 2028
rect 2172 1996 2220 2028
rect 2240 2002 2250 2030
rect 2262 2028 2422 2038
rect 2436 2028 2486 2078
rect 2262 1996 2264 2028
rect 2268 2002 2344 2028
rect 2348 2002 2378 2028
rect 2305 1996 2378 2002
rect 2388 1996 2422 2028
rect 2441 1996 2486 2028
rect 2505 2064 2539 2126
rect 2540 2102 2556 2126
rect 2568 2122 2667 2126
rect 2583 2106 2598 2111
rect 2602 2106 2667 2122
rect 2676 2110 4736 2135
rect 4770 2126 4804 2130
rect 4758 2110 4816 2126
rect 4895 2125 4929 2135
rect 4883 2120 4929 2125
rect 2583 2102 2602 2106
rect 2582 2101 2602 2102
rect 2607 2101 2667 2106
rect 2582 2100 2598 2101
rect 2602 2095 2667 2101
rect 2549 2064 2570 2080
rect 2505 2002 2570 2064
rect 2583 2075 2667 2095
rect 2673 2093 4736 2110
rect 2673 2076 4755 2093
rect 2583 2061 2669 2075
rect 2676 2072 4755 2076
rect 2676 2066 4620 2072
rect 2676 2064 2753 2066
rect 2585 2018 2602 2055
rect 2582 2002 2589 2013
rect 2590 2002 2602 2018
rect 2612 2046 2664 2061
rect 2665 2046 2669 2061
rect 2688 2060 2753 2064
rect 2690 2055 2753 2060
rect 2757 2058 4620 2066
rect 2757 2055 4384 2058
rect 2690 2054 4384 2055
rect 2719 2046 2753 2054
rect 2757 2046 4384 2054
rect 2612 2033 2701 2046
rect 2723 2042 4384 2046
rect 2734 2036 4384 2042
rect 2734 2033 2755 2036
rect 2612 2030 2755 2033
rect 2757 2030 4384 2036
rect 2612 2026 4384 2030
rect 2612 2014 2677 2026
rect 2683 2020 4384 2026
rect 4402 2020 4403 2058
rect 4424 2038 4620 2058
rect 4638 2069 4755 2072
rect 4770 2087 4821 2110
rect 4837 2087 4843 2093
rect 4876 2087 4929 2120
rect 4770 2069 4815 2087
rect 4818 2069 4821 2087
rect 4638 2050 4821 2069
rect 4833 2053 4843 2087
rect 4849 2072 4929 2087
rect 4934 2120 4941 2135
rect 4983 2124 5452 2135
rect 5457 2180 5505 2200
rect 5585 2199 5619 2203
rect 5661 2186 5711 2203
rect 5733 2186 5901 2216
rect 5457 2148 5527 2180
rect 5528 2148 5555 2180
rect 5661 2176 5901 2186
rect 5661 2175 5728 2176
rect 5599 2165 5728 2175
rect 5457 2136 5559 2148
rect 5565 2136 5571 2152
rect 5599 2141 5605 2165
rect 5613 2158 5728 2165
rect 5733 2161 5901 2176
rect 5738 2158 5901 2161
rect 4976 2120 5446 2124
rect 5457 2120 5571 2136
rect 4934 2102 4940 2120
rect 4965 2108 4971 2119
rect 4976 2106 5452 2120
rect 4849 2069 4922 2072
rect 4934 2069 4941 2102
rect 4973 2082 5452 2106
rect 5457 2082 5505 2120
rect 4973 2073 5505 2082
rect 5512 2073 5571 2120
rect 5613 2138 5901 2158
rect 5909 2214 6244 2216
rect 5909 2207 6190 2214
rect 5909 2204 6110 2207
rect 6122 2204 6190 2207
rect 5909 2201 6190 2204
rect 5909 2141 5918 2201
rect 5928 2181 6190 2201
rect 5921 2159 6190 2181
rect 5921 2155 6079 2159
rect 5921 2141 6074 2155
rect 5909 2138 6074 2141
rect 5613 2131 5772 2138
rect 5613 2115 5671 2131
rect 5687 2115 5772 2131
rect 5625 2103 5629 2115
rect 5656 2100 5671 2115
rect 5704 2073 5772 2115
rect 5773 2127 5894 2138
rect 5909 2127 5933 2138
rect 5934 2136 6074 2138
rect 6085 2148 6190 2159
rect 6085 2138 6131 2148
rect 5934 2127 6070 2136
rect 6085 2132 6125 2138
rect 6142 2137 6190 2148
rect 6195 2148 6244 2214
rect 6264 2206 6267 2226
rect 6286 2221 7326 2226
rect 6286 2179 7018 2221
rect 7038 2179 7140 2221
rect 7239 2218 7326 2221
rect 7233 2212 7326 2218
rect 7407 2212 7450 2228
rect 7460 2222 8065 2228
rect 8069 2222 8077 2251
rect 8094 2232 8128 2258
rect 8132 2239 8497 2258
rect 8567 2252 9195 2319
rect 8578 2247 8689 2252
rect 8578 2241 8667 2247
rect 8578 2239 8612 2241
rect 8631 2239 8665 2241
rect 8132 2237 8501 2239
rect 8132 2232 8480 2237
rect 8519 2233 8705 2239
rect 8733 2233 8739 2239
rect 8742 2233 9195 2252
rect 8094 2224 8480 2232
rect 8094 2222 8131 2224
rect 8132 2222 8480 2224
rect 7460 2212 8480 2222
rect 7233 2201 7359 2212
rect 7398 2205 8480 2212
rect 8497 2205 9195 2233
rect 7398 2202 7556 2205
rect 7562 2203 7708 2205
rect 7571 2202 7652 2203
rect 7661 2202 7695 2203
rect 7160 2191 7163 2201
rect 7160 2179 7177 2191
rect 7233 2187 7348 2201
rect 7398 2199 7570 2202
rect 7571 2199 7695 2202
rect 7398 2187 7695 2199
rect 7233 2184 7695 2187
rect 7239 2179 7695 2184
rect 6286 2178 7695 2179
rect 6195 2137 6243 2148
rect 6264 2144 6267 2172
rect 6286 2168 7407 2178
rect 7412 2168 7695 2178
rect 6286 2166 7350 2168
rect 6285 2152 7350 2166
rect 6264 2143 6271 2144
rect 6142 2136 6243 2137
rect 6085 2127 6131 2132
rect 6142 2127 6190 2136
rect 5773 2126 6190 2127
rect 5773 2080 5894 2126
rect 5934 2122 5955 2126
rect 5980 2122 6022 2126
rect 6034 2122 6043 2126
rect 5968 2118 6032 2122
rect 5968 2112 6044 2118
rect 5968 2098 6048 2112
rect 6055 2110 6090 2126
rect 6097 2122 6131 2126
rect 6055 2100 6085 2110
rect 6097 2108 6102 2122
rect 5968 2088 6032 2098
rect 6034 2088 6048 2098
rect 5998 2082 6032 2088
rect 5773 2073 5872 2080
rect 4973 2072 5872 2073
rect 4849 2060 4941 2069
rect 4976 2069 5872 2072
rect 4976 2068 5874 2069
rect 4849 2053 4934 2060
rect 4837 2050 4843 2053
rect 4638 2047 4843 2050
rect 4424 2026 4615 2038
rect 4638 2032 4839 2047
rect 4638 2026 4736 2032
rect 4424 2022 4515 2026
rect 4518 2022 4736 2026
rect 4424 2020 4504 2022
rect 4518 2020 4598 2022
rect 4602 2020 4736 2022
rect 4739 2020 4839 2032
rect 4876 2030 4934 2053
rect 4964 2045 4971 2060
rect 4976 2058 5728 2068
rect 5738 2058 5756 2068
rect 5784 2058 5874 2068
rect 4976 2046 5874 2058
rect 4976 2045 5077 2046
rect 4964 2042 5077 2045
rect 4964 2030 4986 2042
rect 4888 2026 4922 2030
rect 2683 2014 4602 2020
rect 2618 2012 4602 2014
rect 2618 2005 2689 2012
rect 2618 2002 2709 2005
rect 2734 2002 2755 2012
rect 2757 2008 4602 2012
rect 4638 2008 4736 2020
rect 4799 2019 4839 2020
rect 5007 2019 5077 2042
rect 5162 2042 5357 2046
rect 4775 2016 4839 2017
rect 2757 2002 2764 2008
rect 2774 2002 4736 2008
rect 4781 2015 4839 2016
rect 4893 2015 4927 2019
rect 1650 1994 2232 1996
rect 1650 1980 1684 1994
rect 1468 1978 1684 1980
rect 1703 1984 2232 1994
rect 2262 1984 2422 1996
rect 1703 1978 2422 1984
rect 1468 1956 2422 1978
rect 2436 1956 2494 1996
rect 857 1954 1426 1956
rect 1476 1954 1560 1956
rect 1568 1954 2170 1956
rect 2172 1954 2422 1956
rect 2441 1954 2486 1956
rect 2505 1954 2589 2002
rect 2624 1992 4770 2002
rect 4781 1994 4851 2015
rect 4887 2002 4939 2015
rect 4893 2000 4939 2002
rect 4893 1996 4927 2000
rect 4934 1996 4939 2000
rect 4781 1992 4808 1994
rect 4809 1992 4851 1994
rect 2624 1984 4736 1992
rect 2624 1980 2713 1984
rect 2757 1983 4736 1984
rect 4781 1986 4816 1992
rect 4837 1986 4851 1992
rect 4781 1983 4851 1986
rect 4881 1983 4939 1996
rect 5007 1983 5105 2019
rect 2757 1980 5105 1983
rect 5162 1996 5172 2042
rect 5174 2032 5357 2042
rect 5185 2020 5357 2032
rect 5185 2002 5214 2020
rect 5223 2016 5257 2020
rect 5262 2011 5302 2020
rect 5262 2002 5308 2011
rect 5311 2002 5330 2020
rect 5342 2016 5345 2020
rect 5185 1996 5256 2002
rect 5262 1996 5311 2002
rect 5162 1992 5311 1996
rect 5376 1997 5379 2046
rect 5162 1980 5220 1992
rect 2624 1965 2734 1980
rect 2624 1954 2689 1965
rect 2713 1956 2734 1965
rect 2757 1976 5220 1980
rect 2757 1966 4510 1976
rect 4540 1966 5220 1976
rect 5250 1980 5308 1992
rect 5376 1988 5387 1997
rect 5390 1992 5410 2046
rect 5412 2039 5874 2046
rect 5958 2044 5980 2082
rect 5986 2078 6032 2082
rect 5986 2072 6008 2078
rect 5412 2030 5464 2039
rect 5471 2030 5558 2039
rect 5421 2026 5458 2030
rect 5471 2029 5511 2030
rect 5567 2029 5874 2039
rect 5687 2028 5874 2029
rect 5421 2003 5446 2026
rect 5435 1993 5446 2003
rect 5710 2002 5728 2028
rect 5738 2002 5756 2028
rect 5790 2008 5857 2028
rect 5863 2020 5874 2028
rect 6142 2038 6190 2126
rect 6142 2027 6153 2038
rect 5863 2017 6080 2020
rect 5922 2010 6080 2017
rect 5922 2008 6094 2010
rect 6161 2008 6190 2038
rect 5790 1993 6190 2008
rect 5399 1988 5410 1992
rect 5376 1980 5410 1988
rect 5826 1986 6190 1993
rect 5840 1980 6190 1986
rect 6195 2132 6243 2136
rect 6256 2136 6271 2143
rect 6285 2142 6472 2152
rect 6485 2144 6654 2152
rect 6666 2145 7350 2152
rect 6666 2144 7194 2145
rect 6485 2142 7194 2144
rect 6256 2132 6277 2136
rect 6285 2132 6479 2142
rect 6485 2136 6500 2142
rect 6508 2136 7194 2142
rect 6195 2066 6277 2132
rect 6297 2118 6479 2132
rect 6511 2135 7194 2136
rect 6511 2129 7018 2135
rect 6297 2116 6472 2118
rect 6195 2059 6243 2066
rect 6270 2059 6271 2066
rect 6298 2059 6299 2116
rect 6311 2113 6472 2116
rect 6511 2113 6648 2129
rect 6311 2106 6478 2113
rect 6319 2103 6353 2106
rect 6355 2103 6365 2106
rect 6319 2102 6365 2103
rect 6319 2100 6353 2102
rect 6355 2100 6365 2102
rect 6387 2100 6478 2106
rect 6319 2066 6478 2100
rect 6337 2059 6437 2066
rect 6441 2065 6478 2066
rect 6508 2081 6648 2113
rect 6654 2099 7018 2129
rect 7071 2119 7206 2135
rect 7071 2116 7125 2119
rect 7147 2116 7155 2119
rect 7159 2116 7206 2119
rect 7249 2126 7350 2145
rect 7360 2126 7406 2168
rect 7407 2126 7441 2168
rect 7460 2132 7494 2168
rect 7503 2160 7524 2168
rect 7608 2165 7695 2168
rect 7602 2159 7695 2165
rect 7776 2198 8497 2205
rect 7776 2188 8480 2198
rect 7776 2159 8077 2188
rect 8132 2170 8480 2188
rect 8597 2179 8612 2205
rect 8631 2179 8665 2205
rect 8756 2199 9195 2205
rect 9201 2363 9235 2396
rect 9307 2395 9604 2433
rect 9685 2436 9719 2440
rect 9738 2436 9796 2456
rect 9846 2454 9880 2464
rect 9886 2454 9920 2464
rect 9846 2441 9920 2454
rect 9685 2431 9796 2436
rect 9840 2436 9920 2441
rect 9651 2409 9678 2413
rect 9685 2409 9800 2431
rect 9316 2385 9604 2395
rect 9632 2397 9800 2409
rect 9632 2396 9719 2397
rect 9316 2370 9598 2385
rect 9282 2363 9309 2367
rect 9201 2315 9229 2363
rect 9201 2199 9235 2315
rect 9263 2273 9309 2363
rect 9316 2307 9604 2370
rect 9281 2269 9309 2273
rect 9315 2251 9604 2307
rect 9303 2213 9604 2251
rect 8756 2179 9235 2199
rect 8497 2176 9235 2179
rect 8497 2171 9195 2176
rect 9201 2171 9235 2176
rect 8132 2169 8142 2170
rect 7460 2126 7503 2132
rect 7602 2131 7699 2159
rect 7767 2149 8075 2159
rect 7608 2126 7668 2131
rect 7767 2127 8071 2149
rect 7249 2117 7546 2126
rect 7568 2117 7668 2126
rect 7249 2116 7668 2117
rect 6654 2081 6726 2099
rect 6508 2076 6726 2081
rect 6508 2066 6559 2076
rect 6564 2066 6612 2076
rect 6639 2066 6726 2076
rect 6766 2094 6848 2099
rect 6880 2094 7018 2099
rect 7061 2115 7668 2116
rect 7719 2125 8071 2127
rect 7719 2115 7776 2125
rect 7781 2118 8071 2125
rect 7781 2115 8074 2118
rect 7061 2110 7652 2115
rect 7061 2099 7406 2110
rect 7061 2095 7071 2099
rect 7091 2097 7406 2099
rect 7422 2106 7652 2110
rect 7793 2108 8074 2115
rect 6766 2091 6826 2094
rect 6880 2091 6981 2094
rect 6766 2083 6829 2091
rect 6859 2083 6981 2091
rect 7013 2088 7018 2094
rect 7047 2091 7052 2095
rect 7091 2092 7350 2097
rect 7422 2093 7666 2106
rect 7411 2092 7666 2093
rect 7059 2091 7085 2092
rect 6766 2082 6981 2083
rect 6766 2075 6826 2082
rect 6508 2065 6654 2066
rect 6441 2064 6654 2065
rect 6441 2060 6559 2064
rect 6453 2059 6559 2060
rect 6195 2054 6559 2059
rect 6195 2038 6243 2054
rect 6195 2025 6244 2038
rect 6277 2028 6307 2054
rect 6337 2036 6425 2054
rect 6441 2048 6559 2054
rect 6441 2038 6508 2048
rect 6511 2038 6559 2048
rect 6564 2038 6612 2064
rect 6666 2063 6738 2066
rect 6768 2063 6826 2075
rect 6326 2025 6428 2036
rect 6441 2026 6500 2038
rect 6511 2036 6612 2038
rect 6664 2056 6826 2063
rect 6880 2056 7003 2082
rect 6664 2053 7003 2056
rect 6664 2050 6724 2053
rect 6664 2049 6726 2050
rect 6664 2040 6724 2049
rect 6768 2046 7003 2053
rect 7035 2069 7085 2091
rect 7091 2082 7441 2092
rect 7123 2081 7148 2082
rect 7093 2069 7095 2080
rect 7124 2079 7148 2081
rect 7035 2051 7095 2069
rect 6664 2036 6770 2040
rect 6511 2029 6559 2036
rect 6195 1980 6243 2025
rect 6327 2019 6417 2025
rect 6525 2019 6559 2029
rect 6327 2009 6365 2019
rect 6395 2009 6417 2019
rect 6327 2002 6353 2009
rect 6327 1991 6441 2002
rect 6511 1996 6522 2007
rect 6530 1996 6559 2019
rect 5250 1966 5446 1980
rect 2757 1956 5446 1966
rect 2713 1954 2755 1956
rect 2757 1955 4736 1956
rect 2757 1954 4586 1955
rect 4598 1954 4736 1955
rect 4762 1954 4973 1956
rect 5007 1954 5446 1956
rect 5790 1967 6243 1980
rect 6291 1967 6353 1988
rect 6387 1967 6463 1988
rect 6511 1980 6559 1996
rect 6564 2006 6612 2036
rect 6722 2016 6770 2036
rect 6706 2015 6772 2016
rect 6722 2006 6770 2015
rect 6775 2012 6796 2046
rect 6880 2006 7003 2046
rect 7047 2039 7095 2051
rect 6564 1996 6633 2006
rect 6663 2002 7003 2006
rect 7035 2003 7095 2039
rect 7135 2069 7169 2079
rect 7176 2069 7195 2081
rect 7135 2057 7195 2069
rect 7135 2013 7183 2057
rect 6663 1996 6981 2002
rect 7035 2001 7093 2003
rect 7137 2001 7148 2013
rect 7149 2008 7183 2013
rect 7149 2003 7195 2008
rect 6564 1980 6981 1996
rect 7033 1994 7148 2001
rect 7155 1997 7195 2003
rect 7149 1994 7195 1997
rect 7049 1991 7195 1994
rect 7061 1988 7095 1991
rect 7149 1988 7175 1991
rect 7061 1987 7125 1988
rect 7149 1987 7183 1988
rect 6511 1976 6981 1980
rect 6511 1972 6880 1976
rect 6894 1972 6981 1976
rect 6511 1967 6633 1972
rect 5790 1956 6633 1967
rect 5790 1954 6229 1956
rect 6291 1954 6463 1956
rect 6511 1954 6633 1956
rect 6663 1954 6844 1972
rect 6880 1970 6981 1972
rect 216 1949 6810 1954
rect 216 1944 4778 1949
rect 4793 1944 4839 1949
rect 4842 1944 4851 1949
rect 4893 1944 6810 1949
rect 6818 1944 6844 1954
rect 6864 1954 6981 1970
rect 7091 1963 7173 1987
rect 7075 1954 7173 1963
rect 7249 1954 7297 2082
rect 7302 1954 7350 2082
rect 7444 2076 7524 2092
rect 7458 2066 7524 2076
rect 7460 2063 7520 2066
rect 7531 2063 7548 2092
rect 7618 2063 7666 2092
rect 7430 2053 7714 2063
rect 7430 2042 7719 2053
rect 7424 2039 7719 2042
rect 7793 2039 8088 2108
rect 8145 2072 8179 2170
rect 8226 2162 8480 2170
rect 8559 2170 8717 2171
rect 8739 2170 9235 2171
rect 8226 2122 8440 2162
rect 8559 2148 9235 2170
rect 8559 2145 9195 2148
rect 8597 2135 8612 2145
rect 8631 2135 8665 2145
rect 8756 2144 9195 2145
rect 8188 2099 8440 2122
rect 8631 2107 8646 2135
rect 8742 2133 9195 2144
rect 9201 2133 9235 2148
rect 9316 2186 9604 2213
rect 9610 2201 9611 2339
rect 9632 2229 9678 2396
rect 9685 2371 9719 2396
rect 9720 2380 9800 2397
rect 9730 2377 9800 2380
rect 9726 2371 9800 2377
rect 9685 2353 9800 2371
rect 9650 2225 9678 2229
rect 9684 2337 9800 2353
rect 9840 2426 9880 2436
rect 9886 2426 9920 2436
rect 9939 2441 9973 2510
rect 10054 2498 10088 2510
rect 10107 2504 10141 2510
rect 10225 2504 10342 2510
rect 10440 2504 10708 2510
rect 10107 2498 10361 2504
rect 10054 2480 10361 2498
rect 10366 2503 10708 2504
rect 10366 2493 10725 2503
rect 10377 2481 10407 2493
rect 10418 2481 10725 2493
rect 10053 2476 10361 2480
rect 10054 2470 10187 2476
rect 10203 2470 10361 2476
rect 10366 2470 10725 2481
rect 10054 2441 10141 2470
rect 10253 2468 10289 2470
rect 10308 2468 10342 2470
rect 10249 2460 10289 2468
rect 10297 2460 10342 2468
rect 10249 2454 10342 2460
rect 10249 2444 10289 2454
rect 9939 2426 9986 2441
rect 9840 2396 9920 2426
rect 9928 2396 9986 2426
rect 9684 2203 9804 2337
rect 9684 2198 9772 2203
rect 9672 2186 9772 2198
rect 9316 2181 9639 2186
rect 9654 2182 9818 2186
rect 9672 2181 9818 2182
rect 9316 2169 9818 2181
rect 9316 2159 9772 2169
rect 9316 2152 9598 2159
rect 9612 2156 9772 2159
rect 9612 2152 9812 2156
rect 9316 2133 9604 2152
rect 9685 2148 9796 2152
rect 9685 2142 9734 2148
rect 8742 2131 9239 2133
rect 8742 2116 9208 2131
rect 9243 2128 9604 2133
rect 9672 2132 9719 2142
rect 9685 2128 9719 2132
rect 9738 2128 9796 2148
rect 9243 2127 9599 2128
rect 8665 2115 9208 2116
rect 8665 2111 9178 2115
rect 8742 2107 9178 2111
rect 8631 2099 9178 2107
rect 9181 2099 9201 2115
rect 9235 2114 9599 2127
rect 9235 2099 9604 2114
rect 8188 2088 8246 2099
rect 8182 2078 8246 2088
rect 8346 2089 8404 2099
rect 8631 2092 9182 2099
rect 8346 2082 8440 2089
rect 8631 2082 9181 2092
rect 7424 2038 8088 2039
rect 7407 2029 8088 2038
rect 8146 2035 8179 2072
rect 8196 2069 8246 2078
rect 8355 2075 8440 2082
rect 8196 2068 8262 2069
rect 8346 2053 8440 2075
rect 8742 2076 9181 2082
rect 9201 2076 9235 2099
rect 9333 2082 9604 2099
rect 9685 2088 9796 2128
rect 9840 2124 9880 2396
rect 9886 2124 9920 2396
rect 9840 2118 9920 2124
rect 9840 2106 9880 2118
rect 9852 2090 9880 2102
rect 9333 2078 9599 2082
rect 9685 2080 9772 2088
rect 9832 2080 9880 2090
rect 9886 2080 9920 2118
rect 9316 2076 9587 2078
rect 8742 2053 9587 2076
rect 9647 2074 9812 2080
rect 9832 2074 9920 2080
rect 8146 2034 8188 2035
rect 8242 2034 8276 2035
rect 8146 2031 8179 2034
rect 7407 2027 7462 2029
rect 7492 2028 7516 2029
rect 7407 2023 7464 2027
rect 7493 2026 7516 2028
rect 7416 2016 7452 2023
rect 7462 2016 7464 2023
rect 7416 2008 7464 2016
rect 6864 1944 6982 1954
rect 6997 1944 7376 1954
rect 7379 1948 7400 1954
rect 7404 1950 7464 2008
rect 7498 2016 7538 2026
rect 7550 2016 7564 2028
rect 7498 2004 7564 2016
rect 7404 1948 7462 1950
rect 7470 1948 7488 2002
rect 7498 1960 7552 2004
rect 7498 1948 7516 1960
rect 7518 1950 7552 1960
rect 216 1938 7376 1944
rect 216 1933 6794 1938
rect 286 1920 6794 1933
rect 6796 1922 7376 1938
rect 7382 1922 7392 1948
rect 7393 1938 7400 1948
rect 7416 1944 7532 1948
rect 7418 1938 7544 1944
rect 7430 1934 7494 1938
rect 7518 1934 7544 1938
rect 7462 1926 7494 1934
rect 6796 1920 7400 1922
rect 7470 1920 7488 1926
rect 300 1916 4598 1920
rect 300 1911 2320 1916
rect 2326 1911 4598 1916
rect 300 1910 4598 1911
rect 462 1908 477 1910
rect 857 1908 872 1910
rect 462 1898 520 1908
rect 470 1878 520 1898
rect 550 1878 608 1908
rect 246 1868 320 1878
rect 350 1858 608 1878
rect 638 1858 696 1908
rect 726 1878 784 1908
rect 814 1898 872 1908
rect 926 1900 1368 1910
rect 814 1878 864 1898
rect 929 1878 1368 1900
rect 1380 1898 1422 1910
rect 1476 1898 1526 1910
rect 1380 1896 1438 1898
rect 1468 1896 1590 1898
rect 1392 1892 1402 1896
rect 726 1868 890 1878
rect 726 1858 784 1868
rect 814 1858 864 1868
rect 350 1852 550 1858
rect 920 1848 1368 1878
rect 929 1844 1368 1848
rect 1650 1844 1684 1910
rect 929 1836 1386 1844
rect 1427 1836 1479 1844
rect 1515 1839 1631 1844
rect 1579 1836 1631 1839
rect 1668 1836 1684 1844
rect 1703 1836 1737 1910
rect 1768 1836 1771 1910
rect 1827 1909 1856 1910
rect 1863 1909 1902 1910
rect 1827 1893 1902 1909
rect 1918 1893 1948 1910
rect 1845 1859 1948 1893
rect 2019 1878 2053 1910
rect 2072 1878 2106 1910
rect 2174 1887 2175 1910
rect 2262 1902 2264 1910
rect 2262 1899 2274 1902
rect 2262 1887 2279 1899
rect 2348 1896 2374 1910
rect 1990 1876 2130 1878
rect 2006 1872 2130 1876
rect 1845 1843 1911 1859
rect 1918 1843 1948 1859
rect 2019 1864 2130 1872
rect 2019 1844 2056 1864
rect 1887 1836 1902 1843
rect 929 1827 1737 1836
rect 1334 1810 1737 1827
rect 156 1764 158 1796
rect 184 1792 186 1796
rect 156 1698 174 1764
rect 184 1716 202 1792
rect 216 1778 320 1806
rect 350 1796 424 1806
rect 490 1780 608 1806
rect 638 1796 768 1806
rect 834 1796 890 1806
rect 920 1796 1170 1806
rect 1240 1796 1366 1804
rect 1668 1796 1737 1810
rect 1756 1796 1814 1836
rect 1844 1796 1902 1836
rect 696 1788 768 1796
rect 1668 1781 1683 1796
rect 1703 1791 1737 1796
rect 1768 1791 1771 1796
rect 1887 1791 1902 1796
rect 2019 1828 2053 1844
rect 2072 1828 2106 1864
rect 2019 1796 2106 1828
rect 2019 1791 2053 1796
rect 1703 1786 2030 1791
rect 2038 1786 2053 1791
rect 1703 1785 2053 1786
rect 1703 1776 1902 1785
rect 1907 1780 2053 1785
rect 1918 1776 2053 1780
rect 440 1760 474 1769
rect 814 1768 818 1769
rect 1703 1757 2053 1776
rect 2072 1786 2106 1796
rect 2388 1796 2422 1910
rect 2214 1790 2280 1792
rect 978 1722 1028 1756
rect 1620 1722 1668 1748
rect 1680 1722 1714 1756
rect 1768 1722 1802 1756
rect 1856 1722 1890 1756
rect 1902 1722 2056 1748
rect 2072 1723 2087 1786
rect 2095 1785 2106 1786
rect 2388 1785 2399 1796
rect 2168 1738 2326 1756
rect 2407 1748 2422 1796
rect 2441 1892 2482 1910
rect 2505 1908 2589 1910
rect 2624 1908 2677 1910
rect 2505 1897 2539 1908
rect 2555 1897 2589 1908
rect 2643 1897 2677 1908
rect 2757 1908 4598 1910
rect 4604 1908 4636 1920
rect 2757 1898 4636 1908
rect 2757 1897 4384 1898
rect 2505 1896 4384 1897
rect 2441 1848 2475 1892
rect 2505 1878 2529 1896
rect 2494 1868 2529 1878
rect 2543 1874 4384 1896
rect 4452 1888 4510 1898
rect 2543 1868 3744 1874
rect 3759 1868 3772 1874
rect 3802 1868 4384 1874
rect 4386 1868 4510 1888
rect 4540 1868 4598 1898
rect 2505 1863 3852 1868
rect 2555 1851 2601 1863
rect 2441 1836 2456 1848
rect 2471 1847 2475 1848
rect 2464 1836 2475 1847
rect 2441 1748 2475 1836
rect 2543 1846 2601 1851
rect 2677 1846 2689 1851
rect 2543 1836 2558 1846
rect 2582 1836 2601 1846
rect 2674 1836 2689 1846
rect 2543 1834 2601 1836
rect 2631 1834 2689 1836
rect 2757 1848 3852 1863
rect 2757 1840 3818 1848
rect 2583 1756 2584 1794
rect 2631 1786 2681 1834
rect 2757 1806 3796 1840
rect 3804 1806 3818 1840
rect 3864 1806 3898 1868
rect 3917 1836 4339 1868
rect 4350 1836 4384 1868
rect 4452 1864 4498 1868
rect 4410 1838 4498 1864
rect 4552 1838 4598 1868
rect 4602 1838 4636 1898
rect 4638 1914 6612 1920
rect 6617 1914 6643 1920
rect 6772 1914 6783 1920
rect 6796 1915 7175 1920
rect 6796 1914 7199 1915
rect 4638 1910 7199 1914
rect 7249 1910 7253 1920
rect 7263 1913 7297 1920
rect 4638 1908 4736 1910
rect 4742 1908 4753 1910
rect 4638 1838 4753 1908
rect 4410 1836 4598 1838
rect 4655 1836 4753 1838
rect 4833 1881 4911 1887
rect 4833 1876 4927 1881
rect 4833 1853 4911 1876
rect 4833 1846 4861 1853
rect 4877 1847 4911 1853
rect 5007 1847 5446 1910
rect 5790 1898 5861 1910
rect 5790 1877 5860 1898
rect 4833 1837 4879 1846
rect 3917 1806 4753 1836
rect 4829 1809 4879 1837
rect 2757 1804 4753 1806
rect 2757 1796 4446 1804
rect 2757 1790 3820 1796
rect 2757 1772 3774 1790
rect 3781 1775 3796 1790
rect 3864 1782 3898 1796
rect 2599 1756 2633 1760
rect 2583 1753 2649 1756
rect 2583 1748 2584 1753
rect 2119 1727 2373 1738
rect 2072 1722 2086 1723
rect 2130 1722 2326 1727
rect 2332 1722 2362 1727
rect 2407 1722 2424 1748
rect 2441 1722 2512 1748
rect 2542 1740 2584 1748
rect 2650 1740 2734 1748
rect 2542 1722 2734 1740
rect 2757 1740 3784 1772
rect 3834 1748 3898 1782
rect 3917 1748 4331 1796
rect 4350 1748 4384 1796
rect 4428 1784 4446 1796
rect 4396 1749 4446 1784
rect 4452 1796 4512 1804
rect 4540 1796 4753 1804
rect 4452 1781 4509 1796
rect 4552 1793 4598 1796
rect 4568 1781 4598 1793
rect 4464 1780 4536 1781
rect 4464 1777 4526 1780
rect 4568 1777 4586 1781
rect 4476 1768 4526 1777
rect 4388 1748 4446 1749
rect 2757 1730 3160 1740
rect 2757 1722 2764 1730
rect 2774 1722 3160 1730
rect 298 1711 361 1722
rect 597 1716 737 1722
rect 597 1711 608 1716
rect 696 1711 737 1716
rect 773 1711 825 1722
rect 879 1711 931 1722
rect 951 1711 1028 1722
rect 1199 1721 1335 1722
rect 298 1694 350 1711
rect 520 1699 550 1702
rect 520 1694 561 1699
rect 298 1692 561 1694
rect 608 1692 638 1702
rect 696 1699 726 1711
rect 784 1699 814 1711
rect 890 1699 920 1711
rect 962 1699 1028 1711
rect 1155 1711 1335 1721
rect 1507 1711 1559 1722
rect 1579 1711 1631 1722
rect 1155 1708 1283 1711
rect 1155 1701 1286 1708
rect 685 1692 737 1699
rect 773 1692 825 1699
rect 298 1688 864 1692
rect 879 1688 931 1699
rect 951 1690 1028 1699
rect 1152 1699 1286 1701
rect 1294 1699 1324 1711
rect 1518 1699 1548 1711
rect 1590 1699 1620 1711
rect 951 1688 1018 1690
rect 1152 1688 1335 1699
rect 1507 1688 1559 1699
rect 1579 1689 1631 1699
rect 1646 1689 1902 1722
rect 1903 1689 2031 1722
rect 2045 1711 3160 1722
rect 2056 1706 3160 1711
rect 2056 1704 2422 1706
rect 2056 1699 2086 1704
rect 2248 1699 2278 1704
rect 2332 1699 2362 1704
rect 2424 1700 3160 1706
rect 2424 1699 3050 1700
rect 2045 1689 2097 1699
rect 2237 1694 2289 1699
rect 2321 1694 2373 1699
rect 2413 1694 3050 1699
rect 2122 1689 3050 1694
rect 1579 1688 3050 1689
rect 3126 1694 3160 1700
rect 470 1648 520 1688
rect 462 1642 520 1648
rect 550 1642 608 1688
rect 638 1642 696 1688
rect 726 1642 784 1688
rect 814 1648 864 1688
rect 1887 1686 1902 1688
rect 2122 1686 2668 1688
rect 1616 1685 2668 1686
rect 2757 1685 2764 1688
rect 1616 1681 2764 1685
rect 2774 1681 2844 1688
rect 814 1642 872 1648
rect 920 1642 984 1660
rect 1186 1654 1252 1674
rect 1616 1668 2844 1681
rect 1202 1650 1236 1654
rect 462 1640 477 1642
rect 440 1582 458 1640
rect 462 1627 486 1640
rect 468 1610 486 1627
rect 650 1610 684 1636
rect 857 1627 872 1642
rect 1186 1640 1252 1650
rect 1616 1648 2122 1668
rect 1444 1646 1518 1648
rect 1412 1640 1612 1644
rect 1616 1640 2144 1648
rect 2168 1640 2202 1654
rect 2236 1640 2290 1654
rect 2324 1640 2378 1654
rect 2405 1644 2844 1668
rect 3126 1651 3140 1694
rect 3145 1651 3160 1694
rect 3126 1648 3160 1651
rect 3179 1738 3646 1740
rect 3650 1738 3708 1740
rect 3744 1738 3784 1740
rect 3864 1738 3898 1748
rect 3902 1738 4446 1748
rect 3179 1722 3629 1738
rect 3650 1734 4446 1738
rect 4474 1756 4526 1768
rect 4474 1734 4542 1756
rect 4602 1748 4636 1796
rect 4655 1776 4753 1796
rect 4821 1796 4879 1809
rect 4909 1809 4959 1846
rect 5007 1836 5018 1847
rect 5024 1836 5446 1847
rect 4909 1796 4967 1809
rect 4821 1785 4867 1796
rect 4952 1785 4967 1796
rect 5007 1796 5446 1836
rect 5007 1785 5021 1796
rect 4821 1776 4967 1785
rect 5024 1776 5446 1796
rect 4655 1764 4816 1776
rect 4821 1764 5446 1776
rect 4655 1751 5446 1764
rect 4655 1748 4753 1751
rect 3650 1722 4438 1734
rect 4488 1722 4556 1734
rect 4558 1722 4753 1748
rect 4821 1734 4872 1751
rect 3179 1721 3632 1722
rect 3179 1648 3213 1721
rect 3229 1704 3632 1721
rect 3650 1711 4636 1722
rect 4655 1717 4778 1722
rect 4821 1719 4879 1734
rect 4921 1731 4955 1751
rect 5024 1722 5446 1751
rect 5457 1876 5860 1877
rect 5457 1847 5492 1876
rect 5457 1843 5784 1847
rect 5457 1722 5491 1843
rect 5773 1836 5784 1843
rect 5790 1836 5860 1876
rect 5557 1796 5707 1833
rect 5773 1796 5860 1836
rect 5773 1785 5784 1796
rect 5790 1781 5860 1796
rect 5615 1760 5617 1769
rect 5647 1760 5649 1769
rect 5615 1756 5649 1760
rect 5599 1741 5665 1756
rect 5773 1748 5860 1781
rect 6142 1836 6153 1847
rect 6161 1836 6176 1910
rect 5537 1722 5727 1725
rect 5773 1722 5928 1748
rect 5940 1722 5974 1756
rect 6028 1722 6062 1756
rect 6142 1748 6176 1836
rect 6195 1748 6229 1910
rect 6309 1876 6343 1880
rect 6397 1876 6431 1880
rect 6297 1836 6312 1851
rect 6428 1836 6443 1851
rect 6297 1796 6355 1836
rect 6385 1796 6443 1836
rect 6297 1781 6312 1796
rect 6428 1781 6443 1796
rect 6074 1743 6297 1748
rect 6309 1743 6343 1756
rect 6397 1743 6431 1756
rect 6511 1748 6545 1910
rect 6564 1870 6599 1910
rect 6612 1904 6818 1910
rect 6612 1886 6832 1904
rect 6633 1881 6832 1886
rect 6834 1881 6864 1910
rect 6622 1870 6875 1881
rect 6880 1870 6981 1910
rect 6564 1762 6598 1870
rect 6706 1854 6724 1870
rect 6674 1823 6724 1854
rect 6666 1806 6724 1823
rect 6754 1854 6772 1870
rect 6880 1869 6968 1870
rect 7268 1869 7297 1913
rect 6880 1861 6981 1869
rect 7249 1861 7297 1869
rect 6754 1823 6804 1854
rect 6754 1806 6812 1823
rect 6666 1781 6712 1806
rect 6678 1762 6712 1781
rect 6766 1791 6812 1806
rect 6880 1817 7297 1861
rect 7302 1868 7350 1920
rect 7484 1910 7506 1916
rect 7444 1906 7510 1910
rect 7444 1904 7520 1906
rect 7531 1904 7548 1934
rect 7444 1900 7510 1904
rect 7444 1876 7458 1900
rect 7460 1876 7508 1900
rect 7474 1868 7508 1876
rect 7618 1870 7666 2029
rect 7302 1862 7351 1868
rect 7410 1864 7618 1868
rect 7632 1864 7666 1870
rect 7671 1921 7719 2029
rect 7793 2020 8088 2029
rect 8145 2020 8179 2031
rect 8230 2021 8259 2031
rect 8244 2020 8259 2021
rect 8346 2020 8458 2053
rect 7793 1993 8458 2020
rect 8505 2048 9587 2053
rect 8505 2043 8663 2048
rect 8742 2046 9587 2048
rect 9604 2065 9920 2074
rect 9939 2381 9986 2396
rect 10041 2426 10141 2441
rect 10172 2426 10187 2441
rect 10041 2396 10187 2426
rect 10255 2413 10289 2444
rect 10041 2381 10141 2396
rect 10172 2381 10187 2396
rect 10209 2396 10289 2413
rect 10297 2426 10342 2454
rect 10423 2451 10712 2470
rect 10811 2451 10826 2510
rect 10845 2451 10879 2510
rect 11007 2506 11041 2660
rect 11060 2632 11094 2682
rect 11168 2663 11195 2734
rect 11204 2749 11238 2768
rect 11350 2765 11410 2768
rect 11346 2749 11410 2765
rect 11520 2785 11608 2804
rect 11675 2803 12184 2804
rect 11617 2788 12184 2803
rect 11617 2785 11843 2788
rect 11520 2771 11843 2785
rect 11520 2770 11837 2771
rect 11889 2770 12184 2788
rect 11204 2740 11423 2749
rect 11204 2734 11444 2740
rect 11204 2717 11302 2734
rect 11342 2717 11444 2734
rect 11520 2728 11832 2770
rect 11889 2740 11923 2770
rect 11520 2725 11825 2728
rect 11204 2715 11444 2717
rect 11463 2715 11520 2717
rect 11525 2715 11825 2725
rect 11204 2706 11248 2715
rect 11204 2700 11264 2706
rect 11202 2666 11268 2700
rect 11204 2663 11264 2666
rect 11376 2663 11410 2715
rect 11429 2663 11463 2715
rect 11537 2708 11825 2715
rect 11168 2653 11458 2663
rect 11168 2650 11463 2653
rect 11047 2616 11094 2632
rect 11140 2632 11463 2650
rect 11140 2629 11195 2632
rect 11204 2629 11463 2632
rect 11140 2628 11208 2629
rect 11214 2628 11248 2629
rect 11262 2628 11282 2629
rect 11140 2616 11248 2628
rect 11047 2538 11093 2616
rect 11162 2550 11248 2616
rect 11250 2604 11308 2628
rect 11360 2613 11372 2629
rect 11376 2613 11422 2629
rect 11360 2607 11418 2613
rect 11162 2538 11208 2550
rect 11047 2534 11094 2538
rect 11180 2534 11208 2538
rect 11214 2534 11248 2550
rect 11262 2575 11308 2604
rect 11328 2575 11330 2579
rect 11342 2575 11362 2579
rect 11262 2534 11282 2575
rect 11290 2550 11302 2575
rect 11294 2538 11302 2550
rect 11316 2538 11362 2575
rect 11294 2534 11296 2538
rect 11060 2516 11094 2534
rect 10991 2500 11049 2506
rect 10991 2485 11003 2500
rect 11007 2485 11053 2500
rect 10987 2466 11053 2485
rect 10991 2460 11049 2466
rect 11007 2451 11041 2460
rect 10423 2434 10708 2451
rect 10297 2413 10347 2426
rect 10297 2396 10355 2413
rect 9939 2106 9973 2381
rect 10054 2162 10141 2381
rect 10053 2128 10141 2162
rect 10054 2116 10088 2128
rect 10073 2107 10088 2116
rect 9939 2097 9954 2106
rect 9939 2065 9968 2097
rect 10059 2075 10088 2107
rect 10107 2103 10141 2128
rect 10209 2116 10241 2396
rect 10107 2075 10165 2103
rect 10059 2069 10165 2075
rect 9604 2059 9968 2065
rect 9604 2054 9880 2059
rect 9884 2054 9920 2059
rect 9604 2046 9920 2054
rect 8505 2041 8677 2043
rect 8505 1993 8725 2041
rect 8742 2023 8826 2046
rect 8964 2023 9604 2046
rect 8742 2020 9604 2023
rect 9685 2020 9719 2046
rect 9738 2020 9772 2046
rect 9832 2020 9866 2046
rect 9880 2025 9920 2046
rect 9939 2025 9968 2059
rect 10073 2052 10097 2069
rect 10107 2052 10165 2069
rect 10255 2052 10289 2396
rect 10308 2381 10355 2396
rect 10410 2381 10422 2423
rect 10423 2381 10694 2434
rect 10879 2417 11041 2451
rect 11060 2450 11087 2516
rect 11168 2506 11248 2534
rect 11322 2512 11334 2538
rect 11322 2510 11330 2512
rect 11168 2500 11264 2506
rect 11328 2500 11330 2510
rect 11060 2417 11094 2450
rect 11168 2432 11195 2500
rect 11202 2466 11248 2500
rect 11252 2466 11282 2500
rect 11342 2481 11362 2538
rect 11206 2460 11264 2466
rect 11060 2398 11075 2417
rect 11180 2398 11195 2432
rect 11214 2398 11248 2460
rect 11376 2453 11410 2607
rect 11429 2579 11463 2629
rect 11537 2597 11832 2708
rect 11889 2679 11933 2740
rect 11970 2708 12184 2770
rect 12341 2752 12356 2852
rect 12267 2735 12356 2752
rect 12375 2735 12409 2852
rect 12521 2818 12579 2824
rect 12521 2784 12533 2818
rect 12521 2778 12579 2784
rect 12375 2734 12390 2735
rect 12710 2734 12725 2852
rect 12744 2734 12778 3033
rect 12890 2965 12948 2971
rect 12890 2931 12902 2965
rect 12890 2925 12948 2931
rect 12890 2765 12948 2771
rect 12890 2736 12902 2765
rect 12890 2734 12924 2736
rect 11944 2702 12184 2708
rect 11940 2699 12184 2702
rect 12285 2731 12924 2734
rect 12285 2725 12948 2731
rect 11940 2679 11971 2699
rect 11988 2679 11990 2690
rect 11889 2672 12184 2679
rect 11898 2643 12184 2672
rect 11878 2609 12184 2643
rect 12285 2646 12922 2725
rect 13077 2646 13147 3088
rect 13259 3020 13317 3026
rect 13259 2986 13271 3020
rect 13259 2980 13317 2986
rect 13259 2712 13317 2718
rect 13259 2678 13271 2712
rect 13259 2672 13317 2678
rect 12285 2612 12570 2646
rect 12656 2630 12671 2634
rect 11416 2563 11463 2579
rect 11509 2563 11832 2597
rect 11416 2485 11462 2563
rect 11531 2485 11832 2563
rect 11416 2481 11463 2485
rect 11547 2481 11832 2485
rect 11429 2463 11463 2481
rect 11360 2447 11418 2453
rect 11360 2432 11372 2447
rect 11376 2432 11422 2447
rect 11356 2413 11422 2432
rect 11360 2407 11418 2413
rect 11376 2398 11410 2407
rect 10879 2383 11075 2398
rect 10308 2053 10342 2381
rect 10423 2291 10490 2381
rect 11248 2364 11410 2398
rect 11429 2397 11456 2463
rect 11537 2453 11832 2481
rect 11900 2557 12201 2609
rect 12285 2575 12563 2612
rect 12644 2591 12671 2630
rect 12708 2602 12922 2646
rect 13005 2629 13147 2646
rect 13077 2628 13130 2629
rect 12682 2596 12922 2602
rect 11900 2491 12194 2557
rect 12275 2546 12563 2575
rect 12637 2573 12671 2591
rect 12678 2593 12922 2596
rect 13023 2593 13130 2628
rect 12678 2573 12709 2593
rect 13023 2592 13176 2593
rect 13209 2592 13367 2610
rect 13448 2592 13463 3122
rect 13482 2592 13516 3176
rect 13628 3147 13686 3153
rect 13628 3113 13640 3147
rect 13628 3107 13686 3113
rect 13628 2659 13686 2665
rect 13628 2630 13640 2659
rect 13628 2626 13662 2630
rect 13624 2625 13662 2626
rect 13628 2619 13686 2625
rect 12726 2573 12728 2584
rect 13023 2576 13367 2592
rect 13370 2576 13401 2592
rect 13516 2591 13624 2592
rect 12275 2515 12570 2546
rect 12637 2537 12922 2573
rect 12275 2491 12569 2515
rect 12616 2503 12922 2537
rect 13023 2558 13313 2576
rect 13516 2558 13590 2591
rect 13023 2506 13308 2558
rect 13516 2530 13590 2557
rect 13394 2524 13409 2528
rect 11900 2469 12201 2491
rect 11537 2441 11831 2453
rect 11900 2441 12200 2469
rect 12247 2457 12569 2491
rect 11537 2410 11832 2441
rect 11916 2428 12200 2441
rect 11429 2364 11463 2397
rect 11537 2379 11825 2410
rect 11429 2345 11444 2364
rect 11248 2330 11444 2345
rect 11547 2344 11825 2379
rect 11906 2379 12200 2428
rect 12269 2379 12569 2457
rect 11906 2357 12201 2379
rect 12285 2375 12569 2379
rect 10624 2301 10658 2319
rect 11547 2311 11832 2344
rect 11906 2326 12194 2357
rect 10624 2291 10694 2301
rect 10423 2265 10694 2291
rect 11547 2275 11815 2311
rect 11916 2291 12194 2326
rect 12275 2335 12569 2375
rect 12638 2451 12939 2503
rect 13023 2469 13301 2506
rect 12638 2385 12932 2451
rect 13013 2440 13301 2469
rect 13382 2463 13409 2524
rect 13482 2524 13504 2528
rect 13516 2524 13658 2530
rect 13482 2523 13516 2524
rect 13578 2523 13658 2524
rect 13817 2523 13832 3196
rect 13851 3162 13886 3196
rect 13851 2523 13885 3162
rect 13997 3094 14055 3100
rect 13997 3060 14009 3094
rect 13997 3054 14055 3060
rect 14167 2891 14201 2909
rect 14167 2855 14237 2891
rect 14184 2821 14255 2855
rect 14535 2821 14570 2855
rect 13997 2606 14055 2612
rect 13997 2572 14009 2606
rect 13997 2566 14055 2572
rect 13420 2490 13478 2496
rect 13013 2409 13308 2440
rect 13380 2431 13409 2463
rect 13416 2456 13447 2490
rect 13469 2489 13482 2490
rect 13851 2489 13866 2523
rect 13420 2450 13478 2456
rect 13815 2434 13914 2487
rect 14184 2470 14254 2821
rect 14536 2802 14570 2821
rect 14366 2753 14424 2759
rect 14366 2719 14378 2753
rect 14366 2713 14424 2719
rect 14366 2553 14424 2559
rect 14366 2519 14378 2553
rect 14366 2513 14424 2519
rect 14184 2434 14237 2470
rect 13013 2385 13307 2409
rect 13354 2397 13409 2431
rect 14555 2417 14570 2802
rect 14589 2768 14624 2802
rect 14589 2417 14623 2768
rect 12638 2363 12939 2385
rect 12638 2335 12938 2363
rect 12985 2351 13307 2385
rect 12275 2304 12570 2335
rect 12654 2322 12938 2335
rect 11916 2268 12201 2291
rect 12275 2273 12563 2304
rect 10423 2255 10712 2265
rect 10992 2256 11027 2265
rect 11730 2258 12201 2268
rect 10423 2221 10694 2255
rect 10791 2231 11027 2256
rect 10791 2221 10826 2231
rect 10423 2109 10711 2221
rect 10792 2169 10826 2221
rect 10993 2212 11027 2231
rect 11916 2222 12184 2258
rect 12285 2238 12563 2273
rect 12644 2273 12938 2322
rect 13007 2273 13307 2351
rect 12644 2251 12939 2273
rect 13023 2269 13307 2273
rect 11012 2202 11027 2212
rect 11046 2202 11081 2212
rect 11361 2203 11396 2212
rect 11784 2204 11819 2213
rect 10845 2197 11099 2202
rect 10845 2169 10919 2197
rect 10792 2168 10919 2169
rect 10941 2168 11099 2197
rect 11160 2178 11396 2203
rect 11617 2195 11819 2204
rect 11160 2168 11195 2178
rect 10792 2163 10881 2168
rect 10819 2145 10835 2163
rect 10422 2075 10711 2109
rect 10423 2063 10711 2075
rect 10440 2054 10711 2063
rect 10308 2052 10323 2053
rect 10428 2052 10711 2054
rect 9884 2020 9954 2025
rect 8742 2019 9954 2020
rect 8742 2012 9920 2019
rect 8742 2010 9604 2012
rect 9665 2011 9824 2012
rect 9832 2011 9920 2012
rect 9665 2010 9920 2011
rect 8742 2003 9646 2010
rect 9666 2003 9920 2010
rect 8742 1999 9920 2003
rect 9939 2009 9954 2019
rect 9939 1999 9973 2009
rect 10018 1999 10711 2052
rect 10792 2129 10835 2145
rect 10845 2134 10885 2163
rect 10845 2129 10879 2134
rect 10792 2123 10881 2129
rect 10792 2113 10826 2123
rect 10845 2113 10879 2123
rect 10792 2047 10879 2113
rect 10993 2106 11027 2168
rect 11046 2106 11080 2168
rect 11161 2116 11195 2168
rect 11362 2159 11396 2178
rect 11547 2170 11819 2195
rect 11381 2149 11396 2159
rect 11415 2149 11450 2159
rect 11214 2144 11468 2149
rect 11214 2116 11288 2144
rect 11161 2115 11288 2116
rect 11310 2115 11468 2144
rect 11547 2118 11818 2170
rect 11916 2169 12170 2222
rect 12285 2205 12570 2238
rect 12644 2220 12932 2251
rect 12285 2169 12553 2205
rect 12654 2185 12932 2220
rect 13013 2229 13307 2269
rect 13376 2241 13443 2397
rect 14589 2383 14604 2417
rect 15291 2275 15344 2785
rect 13375 2240 13409 2241
rect 13375 2229 13416 2240
rect 13482 2229 13522 2240
rect 13013 2198 13308 2229
rect 13375 2216 13409 2229
rect 15660 2222 15713 2679
rect 11904 2118 11933 2150
rect 11161 2110 11250 2115
rect 10991 2100 11080 2106
rect 10791 2013 10879 2047
rect 10893 2028 10925 2079
rect 10991 2066 11027 2100
rect 11046 2066 11080 2100
rect 11188 2092 11204 2110
rect 10991 2060 11080 2066
rect 8742 1998 10711 1999
rect 8742 1993 10718 1998
rect 7793 1986 8457 1993
rect 7793 1976 8202 1986
rect 7793 1974 8088 1976
rect 8154 1974 8202 1976
rect 8242 1974 8302 1986
rect 8356 1974 8457 1986
rect 7793 1973 8457 1974
rect 7785 1970 8457 1973
rect 8674 1970 8725 1987
rect 7785 1959 8725 1970
rect 7785 1953 8709 1959
rect 8742 1957 9077 1993
rect 7785 1942 8708 1953
rect 7785 1940 8089 1942
rect 8136 1940 8708 1942
rect 7785 1921 7833 1940
rect 7873 1935 7921 1940
rect 7873 1921 7933 1935
rect 7987 1921 8088 1940
rect 7671 1887 7720 1921
rect 7773 1917 8088 1921
rect 8154 1919 8202 1940
rect 8242 1919 8302 1940
rect 8356 1934 8708 1940
rect 8154 1917 8302 1919
rect 8305 1917 8708 1934
rect 7773 1900 8708 1917
rect 7773 1895 8339 1900
rect 7787 1891 8339 1895
rect 7779 1887 8339 1891
rect 7671 1864 7719 1887
rect 7791 1885 7933 1887
rect 7799 1881 7833 1885
rect 7887 1881 7921 1885
rect 7987 1881 8339 1887
rect 7936 1864 8339 1881
rect 7410 1862 8339 1864
rect 7302 1853 8339 1862
rect 7302 1847 7971 1853
rect 7302 1834 7970 1847
rect 7302 1817 7350 1834
rect 6880 1815 6950 1817
rect 6766 1776 6800 1791
rect 6880 1783 7283 1815
rect 6880 1781 6968 1783
rect 7144 1781 7249 1783
rect 6766 1762 6812 1776
rect 6880 1762 6967 1781
rect 7268 1775 7283 1783
rect 7302 1776 7337 1817
rect 7475 1808 7488 1834
rect 7503 1808 7516 1834
rect 7531 1808 7970 1834
rect 7350 1800 7970 1808
rect 7398 1776 7970 1800
rect 7302 1775 7970 1776
rect 6564 1748 6967 1762
rect 6443 1743 6967 1748
rect 7198 1747 7249 1775
rect 6074 1728 6967 1743
rect 6074 1722 6666 1728
rect 6678 1722 6712 1728
rect 6766 1722 6967 1728
rect 7057 1722 7159 1747
rect 7232 1741 7249 1747
rect 7283 1741 7970 1775
rect 7987 1755 8339 1853
rect 7215 1722 7232 1741
rect 7249 1722 7283 1741
rect 7302 1722 7336 1741
rect 7480 1732 7510 1741
rect 7514 1726 7970 1741
rect 7475 1722 7488 1726
rect 4896 1719 5860 1722
rect 4655 1715 4753 1717
rect 4833 1715 4867 1719
rect 3650 1704 4558 1711
rect 3229 1688 3648 1704
rect 3650 1688 3656 1704
rect 3240 1672 3274 1676
rect 3321 1672 3396 1688
rect 3416 1672 3450 1676
rect 2405 1640 3036 1644
rect 3068 1640 3213 1648
rect 468 1582 508 1610
rect 474 1576 508 1582
rect 562 1582 618 1610
rect 644 1582 684 1610
rect 562 1576 625 1582
rect 181 1565 408 1576
rect 181 1553 205 1565
rect 216 1553 408 1565
rect 440 1562 625 1576
rect 181 1542 408 1553
rect 462 1542 625 1562
rect 274 1517 308 1542
rect 262 1502 308 1517
rect 174 1472 216 1492
rect 262 1472 320 1502
rect 262 1466 308 1472
rect 350 1469 356 1502
rect 362 1469 396 1542
rect 474 1494 508 1542
rect 350 1466 396 1469
rect 262 1458 277 1466
rect 350 1458 371 1466
rect 262 1454 320 1458
rect 326 1454 408 1458
rect 270 1452 320 1454
rect 350 1452 400 1454
rect 188 1404 238 1420
rect 268 1404 318 1420
rect 180 1399 238 1404
rect 305 1400 326 1404
rect 399 1400 414 1404
rect 440 1402 458 1494
rect 468 1458 508 1494
rect 462 1424 508 1458
rect 462 1406 514 1424
rect 550 1410 556 1425
rect 562 1424 596 1542
rect 607 1530 625 1542
rect 635 1576 684 1582
rect 738 1576 772 1610
rect 826 1576 860 1610
rect 934 1606 984 1638
rect 1186 1624 1232 1640
rect 1616 1628 2122 1640
rect 2405 1632 2844 1640
rect 3126 1632 3160 1640
rect 2405 1630 3039 1632
rect 1152 1612 1178 1616
rect 1232 1612 1266 1616
rect 1440 1612 1612 1616
rect 1152 1610 1190 1612
rect 926 1588 984 1606
rect 926 1576 972 1588
rect 1026 1576 1060 1610
rect 1144 1609 1190 1610
rect 1220 1609 1267 1612
rect 1632 1610 1938 1628
rect 2028 1612 2116 1620
rect 2196 1619 2202 1626
rect 2190 1610 2205 1619
rect 2236 1612 2242 1626
rect 2284 1612 2290 1626
rect 2324 1612 2330 1626
rect 2372 1612 2378 1626
rect 2405 1615 3042 1630
rect 2412 1612 2418 1615
rect 2460 1612 2466 1615
rect 2500 1612 2506 1615
rect 2548 1612 2554 1615
rect 2588 1612 2594 1615
rect 2724 1612 2776 1615
rect 2810 1612 3042 1615
rect 3065 1620 3160 1632
rect 3065 1612 3162 1620
rect 1144 1596 1184 1609
rect 1226 1596 1266 1609
rect 1144 1576 1178 1596
rect 1232 1576 1266 1596
rect 1474 1594 1646 1610
rect 1318 1588 1646 1594
rect 1318 1582 1596 1588
rect 1318 1576 1674 1582
rect 1680 1576 1714 1610
rect 1720 1590 1762 1610
rect 1768 1600 1814 1610
rect 2028 1600 2082 1610
rect 1768 1596 2082 1600
rect 2190 1604 2236 1610
rect 2290 1604 2324 1610
rect 2378 1604 2412 1610
rect 1720 1576 1762 1582
rect 1768 1576 2150 1596
rect 2190 1576 2248 1604
rect 2278 1576 2336 1604
rect 2366 1576 2424 1604
rect 2466 1576 2500 1610
rect 2554 1576 2611 1610
rect 2724 1582 2776 1606
rect 2810 1604 3160 1612
rect 2810 1598 3162 1604
rect 2810 1582 2864 1598
rect 2898 1582 2932 1598
rect 2776 1578 2810 1582
rect 2864 1578 2898 1582
rect 635 1542 872 1576
rect 904 1552 1072 1576
rect 900 1542 1098 1552
rect 1110 1546 1278 1576
rect 1283 1572 1386 1576
rect 1387 1572 1439 1576
rect 1474 1572 1814 1576
rect 1283 1565 1814 1572
rect 1294 1560 1814 1565
rect 1294 1553 1574 1560
rect 1590 1553 1620 1560
rect 1283 1548 1574 1553
rect 1283 1546 1335 1548
rect 1106 1542 1335 1546
rect 1340 1542 1574 1548
rect 1579 1542 1631 1553
rect 1646 1546 1814 1560
rect 1960 1574 2116 1576
rect 2133 1574 2611 1576
rect 1960 1546 2128 1574
rect 2133 1565 2174 1574
rect 2144 1553 2174 1565
rect 1642 1542 1840 1546
rect 1982 1542 2128 1546
rect 2133 1544 2185 1553
rect 2190 1548 2611 1574
rect 2190 1544 2600 1548
rect 2133 1542 2600 1544
rect 635 1530 684 1542
rect 738 1530 772 1542
rect 826 1530 872 1542
rect 638 1500 696 1530
rect 726 1500 784 1530
rect 814 1500 872 1530
rect 607 1494 625 1500
rect 635 1494 684 1500
rect 644 1466 684 1494
rect 704 1466 705 1470
rect 726 1466 772 1500
rect 821 1494 872 1500
rect 792 1466 793 1494
rect 820 1485 872 1494
rect 926 1530 972 1542
rect 1026 1530 1072 1542
rect 926 1516 984 1530
rect 1014 1516 1072 1530
rect 1132 1534 1278 1542
rect 1132 1530 1253 1534
rect 1263 1530 1278 1534
rect 1132 1522 1278 1530
rect 1340 1530 1386 1542
rect 1440 1530 1474 1542
rect 1528 1530 1574 1542
rect 1253 1520 1262 1522
rect 926 1510 1118 1516
rect 1132 1510 1162 1520
rect 926 1508 1162 1510
rect 1238 1508 1278 1520
rect 926 1500 1178 1508
rect 926 1490 972 1500
rect 978 1494 1020 1500
rect 1026 1496 1178 1500
rect 1026 1494 1147 1496
rect 1026 1490 1072 1494
rect 650 1454 684 1466
rect 696 1454 717 1466
rect 650 1442 717 1454
rect 732 1454 772 1466
rect 784 1454 805 1466
rect 732 1442 805 1454
rect 820 1454 860 1485
rect 562 1410 602 1424
rect 650 1410 711 1442
rect 732 1410 799 1442
rect 820 1410 866 1454
rect 875 1426 925 1474
rect 926 1464 955 1490
rect 1057 1488 1072 1490
rect 978 1480 1020 1488
rect 1057 1485 1090 1488
rect 1066 1480 1090 1485
rect 1132 1482 1147 1494
rect 1173 1494 1178 1496
rect 1173 1492 1184 1494
rect 978 1466 1090 1480
rect 1130 1480 1147 1482
rect 1130 1466 1155 1480
rect 926 1454 972 1464
rect 926 1436 984 1454
rect 1013 1436 1072 1466
rect 1132 1445 1155 1466
rect 1169 1446 1184 1492
rect 1232 1476 1278 1508
rect 1340 1500 1398 1530
rect 1428 1500 1486 1530
rect 1516 1500 1574 1530
rect 1668 1534 1714 1542
rect 1668 1530 1683 1534
rect 1726 1530 1756 1542
rect 1768 1534 1814 1542
rect 1799 1530 1814 1534
rect 1668 1522 1814 1530
rect 1982 1530 2028 1542
rect 2082 1530 2128 1542
rect 2190 1536 2600 1542
rect 1676 1520 1726 1522
rect 1207 1466 1278 1476
rect 1294 1470 1324 1500
rect 1340 1470 1395 1500
rect 1440 1482 1474 1500
rect 1528 1494 1574 1500
rect 1493 1482 1511 1494
rect 1521 1485 1574 1494
rect 1668 1500 1726 1520
rect 1756 1520 1806 1522
rect 1756 1508 1814 1520
rect 1982 1508 2040 1530
rect 1756 1500 2040 1508
rect 2070 1500 2128 1530
rect 2174 1506 2190 1510
rect 2198 1506 2248 1536
rect 2174 1500 2248 1506
rect 2278 1500 2336 1536
rect 2374 1506 2424 1536
rect 2366 1500 2424 1506
rect 2454 1500 2512 1536
rect 2542 1506 2592 1536
rect 2542 1500 2600 1506
rect 1521 1482 1562 1485
rect 1455 1481 1518 1482
rect 1521 1481 1539 1482
rect 1548 1481 1574 1482
rect 1455 1470 1574 1481
rect 1294 1466 1329 1470
rect 1352 1466 1363 1470
rect 1201 1465 1278 1466
rect 1196 1454 1278 1465
rect 1158 1445 1184 1446
rect 934 1426 1005 1436
rect 1014 1430 1064 1436
rect 1132 1433 1184 1445
rect 1201 1442 1278 1454
rect 1283 1451 1339 1466
rect 1493 1454 1511 1470
rect 1521 1466 1539 1470
rect 1521 1454 1548 1466
rect 1201 1440 1241 1442
rect 1201 1436 1245 1440
rect 1253 1436 1278 1442
rect 1132 1430 1190 1433
rect 1201 1430 1278 1436
rect 1289 1432 1329 1451
rect 1555 1442 1596 1454
rect 1486 1436 1509 1438
rect 1014 1426 1089 1430
rect 873 1424 925 1426
rect 955 1424 1013 1426
rect 873 1410 920 1424
rect 961 1410 1013 1424
rect 1026 1410 1035 1426
rect 1055 1411 1089 1426
rect 1144 1418 1147 1430
rect 1152 1426 1178 1430
rect 1195 1426 1266 1430
rect 1195 1418 1274 1426
rect 1186 1414 1274 1418
rect 1055 1410 1101 1411
rect 462 1402 486 1406
rect 508 1403 514 1406
rect 180 1366 189 1399
rect 201 1389 238 1399
rect 216 1370 238 1389
rect 268 1370 326 1400
rect 180 1362 196 1366
rect 180 1358 208 1362
rect 280 1358 314 1370
rect 320 1358 326 1370
rect 356 1358 414 1400
rect 462 1400 477 1402
rect 520 1400 1101 1410
rect 1158 1402 1274 1414
rect 1289 1408 1324 1432
rect 1567 1430 1590 1442
rect 1668 1432 1814 1500
rect 1982 1482 2028 1500
rect 2082 1485 2128 1500
rect 2190 1498 2236 1500
rect 2290 1498 2324 1500
rect 2366 1498 2412 1500
rect 2466 1498 2500 1500
rect 2554 1498 2600 1500
rect 2190 1485 2205 1498
rect 2366 1495 2379 1498
rect 2585 1495 2600 1498
rect 2688 1495 2722 1566
rect 2724 1554 2728 1578
rect 2770 1573 2822 1578
rect 2852 1573 2910 1578
rect 2770 1554 2816 1573
rect 2858 1554 2904 1573
rect 2942 1564 3008 1596
rect 3145 1570 3162 1598
rect 3179 1579 3213 1640
rect 3228 1663 3286 1672
rect 3316 1663 3462 1672
rect 3228 1648 3274 1663
rect 3316 1657 3409 1663
rect 3321 1648 3409 1657
rect 3228 1618 3286 1648
rect 3316 1647 3409 1648
rect 3416 1650 3450 1663
rect 3316 1618 3374 1647
rect 3228 1603 3274 1618
rect 3416 1613 3421 1650
rect 3228 1579 3237 1603
rect 3240 1579 3274 1603
rect 3495 1591 3529 1688
rect 3495 1587 3516 1591
rect 3495 1579 3529 1587
rect 3179 1568 3462 1579
rect 3179 1566 3222 1568
rect 3228 1566 3462 1568
rect 2776 1498 2810 1554
rect 2864 1498 2898 1554
rect 3179 1551 3462 1566
rect 3516 1575 3529 1579
rect 3548 1575 3582 1688
rect 3662 1666 3708 1704
rect 3744 1681 3774 1704
rect 3738 1678 3784 1681
rect 3738 1666 3789 1678
rect 3662 1662 3682 1666
rect 3731 1662 3774 1666
rect 3666 1644 3780 1662
rect 3666 1640 3744 1644
rect 3694 1612 3752 1634
rect 3694 1594 3706 1612
rect 3731 1597 3752 1612
rect 3708 1594 3752 1597
rect 3694 1588 3752 1594
rect 3516 1551 3582 1575
rect 3179 1550 3582 1551
rect 3744 1550 3750 1578
rect 3759 1560 3780 1644
rect 3864 1588 3898 1704
rect 3179 1545 3802 1550
rect 2756 1495 2822 1498
rect 2082 1482 2116 1485
rect 1982 1468 2128 1482
rect 2190 1468 2205 1483
rect 2028 1440 2081 1452
rect 2190 1446 2248 1468
rect 2278 1446 2336 1468
rect 2337 1446 2600 1495
rect 2676 1464 2822 1495
rect 2852 1464 2910 1498
rect 3240 1497 3274 1545
rect 3328 1497 3362 1545
rect 3416 1497 3450 1545
rect 3528 1497 3802 1545
rect 3805 1539 3857 1550
rect 3816 1503 3846 1539
rect 2776 1460 2810 1464
rect 2864 1460 2898 1464
rect 2190 1442 2249 1446
rect 2278 1442 2600 1446
rect 2190 1438 2600 1442
rect 1632 1431 1726 1432
rect 1756 1431 1814 1432
rect 1632 1430 1814 1431
rect 1511 1428 1515 1430
rect 1561 1428 1603 1430
rect 1632 1428 1729 1430
rect 1756 1428 1814 1430
rect 1844 1428 1934 1438
rect 1981 1436 2070 1438
rect 1509 1426 1635 1428
rect 1487 1424 1635 1426
rect 1646 1424 1649 1428
rect 1655 1424 1743 1428
rect 1487 1422 1743 1424
rect 1756 1422 1806 1428
rect 1487 1416 1806 1422
rect 1487 1414 1814 1416
rect 1487 1413 1563 1414
rect 1487 1411 1511 1413
rect 1515 1411 1548 1413
rect 1326 1408 1341 1411
rect 462 1398 1101 1400
rect 462 1394 1055 1398
rect 1086 1396 1101 1398
rect 180 1354 414 1358
rect 468 1354 614 1394
rect 638 1376 805 1394
rect 638 1372 705 1376
rect 638 1354 688 1372
rect 747 1354 797 1376
rect 814 1354 864 1394
rect 867 1392 1055 1394
rect 867 1382 1072 1392
rect 1098 1382 1101 1396
rect 1186 1392 1274 1402
rect 1195 1388 1274 1392
rect 867 1354 1101 1382
rect 1186 1376 1274 1388
rect 1283 1376 1341 1408
rect 1487 1402 1548 1411
rect 1597 1408 1814 1414
rect 1597 1402 1723 1408
rect 1726 1402 1814 1408
rect 1509 1396 1548 1402
rect 1561 1398 1743 1402
rect 1186 1368 1253 1376
rect 1203 1366 1253 1368
rect 1283 1366 1333 1376
rect 1509 1366 1567 1396
rect 1597 1394 1743 1398
rect 1597 1382 1723 1394
rect 1726 1382 1743 1394
rect 1756 1382 1814 1402
rect 1844 1382 1894 1416
rect 1902 1382 1934 1428
rect 2028 1422 2081 1430
rect 2115 1422 2116 1430
rect 2190 1427 2689 1438
rect 2724 1436 2776 1460
rect 2810 1444 2864 1460
rect 2898 1444 2932 1460
rect 2942 1446 3008 1478
rect 3179 1476 3462 1497
rect 3179 1474 3222 1476
rect 3228 1474 3462 1476
rect 3145 1444 3162 1472
rect 2810 1438 3162 1444
rect 3179 1463 3462 1474
rect 3516 1492 3802 1497
rect 3805 1492 3857 1503
rect 3516 1467 3582 1492
rect 3516 1463 3529 1467
rect 3548 1466 3582 1467
rect 2810 1430 3160 1438
rect 2190 1420 2405 1427
rect 2424 1425 2425 1427
rect 2407 1420 2425 1425
rect 2190 1416 2425 1420
rect 2460 1425 2466 1427
rect 2490 1425 2512 1427
rect 2460 1417 2512 1425
rect 2542 1420 2689 1427
rect 2724 1427 2776 1430
rect 2810 1427 3042 1430
rect 2724 1426 3042 1427
rect 2774 1421 2852 1426
rect 2548 1417 2668 1420
rect 2437 1416 2668 1417
rect 2000 1402 2069 1414
rect 2086 1402 2122 1414
rect 2203 1402 2437 1416
rect 2462 1402 2512 1416
rect 2542 1402 2592 1416
rect 2774 1410 2863 1421
rect 2908 1412 3042 1426
rect 3096 1422 3162 1430
rect 3110 1421 3140 1422
rect 3099 1410 3140 1421
rect 2774 1402 2844 1410
rect 3126 1402 3140 1410
rect 3145 1402 3160 1422
rect 3179 1402 3213 1463
rect 2000 1394 2081 1402
rect 2086 1394 2144 1402
rect 1950 1382 1984 1388
rect 2000 1382 2069 1394
rect 2086 1382 2122 1394
rect 2168 1388 2202 1402
rect 2203 1400 2622 1402
rect 2203 1391 2466 1400
rect 2500 1391 2554 1400
rect 2588 1391 2622 1400
rect 2724 1398 3036 1402
rect 2774 1391 2844 1398
rect 3068 1394 3213 1402
rect 2203 1388 2844 1391
rect 1597 1374 2149 1382
rect 2203 1374 2437 1388
rect 1597 1370 2261 1374
rect 1203 1354 1324 1366
rect 1509 1358 1555 1366
rect 1597 1358 1643 1370
rect 1509 1354 1643 1358
rect 1655 1366 2261 1370
rect 2291 1366 2349 1374
rect 2379 1366 2437 1374
rect 1655 1354 2218 1366
rect 2248 1354 2261 1366
rect 2332 1354 2349 1366
rect 2407 1354 2437 1366
rect 2441 1378 2844 1388
rect 2441 1376 2952 1378
rect 2441 1366 3036 1376
rect 2441 1357 2764 1366
rect 2441 1354 2553 1357
rect 2650 1354 2734 1357
rect 2757 1354 2764 1357
rect 2774 1354 3036 1366
rect 180 1336 1117 1354
rect 154 1294 174 1328
rect 180 1320 1034 1336
rect 1043 1332 1093 1336
rect 180 1290 414 1320
rect 468 1309 614 1320
rect 480 1305 514 1309
rect 576 1305 602 1309
rect 821 1308 851 1320
rect 890 1308 893 1320
rect 925 1310 955 1320
rect 962 1318 1012 1320
rect 1021 1318 1028 1320
rect 962 1310 997 1318
rect 1098 1308 1117 1336
rect 1152 1350 1367 1354
rect 1509 1353 2185 1354
rect 1152 1341 1363 1350
rect 1152 1320 1158 1341
rect 1160 1338 1363 1341
rect 1509 1338 2149 1353
rect 2203 1342 3050 1354
rect 3126 1348 3140 1394
rect 3145 1348 3160 1394
rect 3126 1342 3160 1348
rect 2248 1338 2291 1342
rect 2332 1338 2379 1342
rect 1160 1334 1286 1338
rect 1176 1331 1283 1334
rect 1294 1331 1324 1338
rect 1518 1331 1548 1338
rect 1567 1331 1620 1338
rect 1646 1336 2422 1338
rect 2424 1336 3160 1342
rect 1646 1334 3160 1336
rect 1646 1331 2422 1334
rect 2424 1331 3160 1334
rect 1176 1330 1631 1331
rect 1242 1321 1631 1330
rect 1646 1321 3160 1331
rect 1199 1320 3160 1321
rect 1294 1310 1324 1320
rect 750 1306 852 1308
rect 180 1287 238 1290
rect 268 1287 326 1290
rect 356 1287 414 1290
rect 490 1287 526 1304
rect 556 1287 608 1304
rect 610 1287 960 1306
rect 180 1278 960 1287
rect 1341 1280 1366 1320
rect 1396 1290 1461 1308
rect 1491 1290 1518 1308
rect 180 1263 638 1278
rect 679 1272 862 1278
rect 879 1272 931 1278
rect 949 1272 960 1278
rect 180 1251 189 1263
rect 192 1260 638 1263
rect 192 1256 196 1260
rect 180 1236 195 1251
rect 207 1247 638 1260
rect 745 1256 768 1272
rect 207 1236 644 1247
rect 713 1238 768 1256
rect 784 1242 801 1272
rect 784 1240 818 1242
rect 180 1224 644 1236
rect 188 1214 644 1224
rect 718 1222 779 1238
rect 890 1236 893 1272
rect 926 1236 960 1272
rect 1253 1256 1283 1280
rect 1518 1266 1533 1290
rect 1210 1246 1333 1256
rect 1541 1248 1548 1290
rect 1671 1285 1714 1320
rect 1717 1285 1902 1320
rect 1905 1286 1939 1320
rect 1993 1286 2027 1320
rect 2069 1315 2127 1320
rect 2130 1315 2291 1320
rect 2332 1315 2379 1320
rect 2069 1304 2302 1315
rect 2321 1304 2390 1315
rect 1905 1285 1951 1286
rect 1981 1285 2039 1286
rect 1671 1271 2053 1285
rect 2069 1271 2106 1304
rect 2115 1294 2195 1304
rect 2115 1292 2261 1294
rect 2115 1271 2195 1292
rect 1671 1270 2195 1271
rect 1671 1263 2053 1270
rect 1668 1251 2053 1263
rect 2069 1258 2087 1270
rect 2069 1256 2106 1258
rect 1210 1238 1363 1246
rect 1210 1236 1282 1238
rect 216 1156 644 1214
rect 920 1215 1056 1236
rect 1203 1224 1253 1236
rect 1283 1232 1363 1238
rect 1583 1236 1590 1248
rect 1668 1244 1737 1251
rect 1668 1236 1701 1244
rect 1703 1236 1737 1244
rect 1768 1236 1805 1251
rect 1856 1244 2053 1251
rect 1859 1236 2053 1244
rect 1668 1232 1737 1236
rect 1283 1224 1737 1232
rect 1195 1215 1253 1224
rect 1267 1222 1737 1224
rect 1283 1215 1737 1222
rect 920 1206 1737 1215
rect 1756 1206 1814 1236
rect 1844 1217 1953 1236
rect 1827 1206 1953 1217
rect 2019 1206 2053 1236
rect 752 1204 768 1206
rect 752 1188 813 1204
rect 752 1184 802 1188
rect 821 1184 851 1206
rect 205 1144 644 1156
rect 646 1144 696 1184
rect 205 1142 696 1144
rect 136 1134 696 1142
rect 726 1182 768 1184
rect 784 1182 802 1184
rect 814 1182 864 1184
rect 726 1170 864 1182
rect 726 1144 776 1170
rect 814 1144 864 1170
rect 890 1164 893 1206
rect 926 1200 1429 1206
rect 1430 1200 1620 1206
rect 1668 1200 1684 1206
rect 926 1181 1698 1200
rect 1703 1181 1737 1206
rect 1768 1181 1805 1206
rect 1827 1199 1856 1206
rect 1859 1199 1902 1206
rect 1827 1183 1902 1199
rect 1918 1183 1948 1206
rect 1845 1181 1948 1183
rect 1951 1181 1981 1206
rect 1990 1198 2053 1206
rect 2072 1198 2106 1256
rect 2214 1236 2219 1252
rect 2332 1250 2333 1304
rect 2388 1252 2390 1304
rect 2407 1252 2422 1320
rect 2111 1202 2140 1224
rect 2214 1202 2280 1232
rect 2388 1208 2422 1252
rect 2441 1216 2475 1320
rect 2541 1305 2542 1320
rect 2757 1312 2764 1320
rect 2774 1312 3160 1320
rect 2583 1289 2584 1305
rect 2757 1302 3160 1312
rect 3179 1321 3213 1394
rect 3228 1439 3237 1463
rect 3240 1439 3274 1463
rect 3228 1424 3274 1439
rect 3495 1455 3529 1463
rect 3536 1455 3582 1466
rect 3744 1464 3750 1492
rect 3495 1451 3516 1455
rect 3303 1424 3328 1429
rect 3371 1424 3409 1433
rect 3228 1370 3286 1424
rect 3303 1420 3409 1424
rect 3299 1408 3409 1420
rect 3416 1408 3421 1429
rect 3299 1382 3462 1408
rect 3316 1370 3462 1382
rect 3240 1366 3274 1370
rect 3321 1361 3387 1370
rect 3416 1366 3450 1370
rect 3321 1354 3358 1361
rect 3495 1354 3529 1451
rect 3548 1354 3582 1455
rect 3694 1448 3752 1454
rect 3694 1430 3706 1448
rect 3731 1430 3752 1448
rect 3694 1408 3752 1430
rect 3759 1402 3780 1482
rect 3883 1454 3898 1588
rect 3666 1380 3780 1402
rect 3662 1376 3682 1380
rect 3744 1376 3774 1380
rect 3229 1338 3648 1354
rect 3650 1338 3656 1354
rect 3662 1338 3708 1376
rect 3738 1364 3789 1376
rect 3738 1361 3784 1364
rect 3744 1338 3784 1361
rect 3864 1338 3898 1454
rect 3917 1699 4558 1704
rect 4568 1699 4636 1711
rect 3917 1694 4636 1699
rect 4666 1694 4753 1715
rect 4879 1697 5860 1719
rect 3917 1688 4753 1694
rect 4896 1690 5860 1697
rect 5906 1690 6074 1722
rect 6108 1690 7400 1722
rect 7470 1716 7488 1722
rect 7462 1713 7492 1716
rect 7503 1713 7970 1726
rect 7416 1694 7440 1698
rect 7462 1694 7970 1713
rect 7984 1711 8339 1755
rect 4896 1688 7400 1690
rect 3917 1685 4331 1688
rect 3917 1672 4303 1685
rect 4316 1672 4331 1685
rect 3917 1656 4331 1672
rect 4350 1656 4384 1688
rect 4388 1672 4438 1688
rect 4492 1684 4558 1688
rect 4519 1672 4534 1684
rect 4388 1656 4446 1672
rect 4476 1656 4534 1672
rect 4602 1656 4636 1688
rect 3917 1632 4636 1656
rect 4666 1632 4753 1688
rect 4870 1654 4927 1681
rect 5024 1662 5446 1688
rect 4882 1650 4911 1654
rect 4861 1647 4927 1650
rect 3917 1631 4753 1632
rect 4934 1631 4964 1646
rect 3917 1615 4636 1631
rect 3917 1603 3951 1615
rect 4019 1613 4077 1615
rect 4107 1613 4165 1615
rect 4031 1609 4065 1613
rect 4119 1609 4153 1613
rect 3917 1602 4187 1603
rect 4190 1602 4202 1615
rect 3917 1598 4202 1602
rect 3917 1574 4206 1598
rect 4218 1574 4230 1615
rect 4250 1600 4636 1615
rect 4672 1606 4753 1631
rect 4250 1596 4303 1600
rect 4233 1574 4303 1596
rect 4316 1598 4636 1600
rect 4316 1588 4436 1598
rect 4440 1588 4446 1598
rect 4316 1574 4446 1588
rect 4478 1581 4522 1598
rect 4528 1596 4636 1598
rect 4478 1574 4525 1581
rect 4528 1574 4638 1596
rect 3917 1569 4340 1574
rect 4388 1569 4534 1574
rect 3917 1473 3951 1569
rect 4014 1544 4144 1569
rect 4018 1541 4147 1544
rect 4184 1541 4202 1569
rect 4212 1541 4230 1569
rect 4233 1564 4340 1569
rect 4394 1564 4400 1569
rect 4233 1562 4320 1564
rect 4428 1562 4440 1569
rect 4233 1541 4340 1562
rect 4018 1535 4064 1541
rect 4025 1529 4064 1535
rect 4025 1507 4052 1529
rect 4059 1525 4064 1529
rect 4094 1539 4140 1541
rect 4094 1525 4144 1539
rect 4106 1517 4144 1525
rect 4018 1483 4052 1507
rect 4059 1501 4064 1517
rect 4094 1507 4144 1517
rect 4075 1501 4144 1507
rect 4059 1483 4144 1501
rect 4184 1507 4340 1541
rect 4006 1473 4152 1483
rect 4184 1473 4202 1507
rect 4212 1473 4230 1507
rect 4233 1473 4340 1507
rect 4394 1560 4440 1562
rect 4394 1554 4468 1560
rect 4470 1554 4516 1569
rect 4570 1564 4638 1574
rect 4394 1531 4516 1554
rect 4394 1511 4440 1531
rect 4444 1511 4516 1531
rect 4394 1488 4516 1511
rect 4394 1482 4468 1488
rect 4394 1473 4440 1482
rect 4470 1478 4516 1488
rect 4602 1478 4638 1564
rect 4670 1579 4753 1606
rect 4770 1579 4787 1610
rect 4888 1579 4922 1616
rect 5001 1612 5010 1616
rect 5001 1600 5022 1612
rect 4976 1579 5022 1600
rect 5035 1579 5069 1662
rect 4670 1551 4838 1579
rect 4854 1551 5022 1579
rect 5030 1572 5069 1579
rect 5088 1572 5122 1662
rect 5188 1646 5338 1662
rect 5198 1640 5328 1646
rect 5198 1634 5248 1640
rect 5278 1634 5328 1640
rect 5198 1626 5328 1634
rect 5234 1612 5292 1626
rect 5234 1610 5246 1612
rect 5230 1594 5296 1610
rect 5334 1600 5338 1646
rect 5404 1628 5438 1662
rect 5390 1600 5438 1628
rect 5457 1616 5491 1688
rect 5559 1676 5574 1688
rect 5690 1676 5705 1688
rect 5457 1603 5492 1616
rect 5512 1603 5525 1616
rect 5537 1603 5546 1616
rect 5559 1613 5617 1676
rect 5647 1613 5705 1676
rect 5773 1656 5860 1688
rect 5928 1676 5943 1688
rect 6059 1676 6074 1688
rect 5928 1656 5986 1676
rect 6016 1656 6074 1676
rect 6142 1656 6176 1688
rect 5773 1646 6176 1656
rect 5773 1642 5861 1646
rect 5928 1642 6176 1646
rect 5571 1609 5605 1613
rect 5659 1609 5693 1613
rect 5710 1603 5728 1640
rect 5457 1600 5728 1603
rect 5234 1588 5292 1594
rect 5196 1572 5218 1576
rect 5272 1572 5306 1584
rect 5038 1556 5069 1572
rect 5027 1551 5069 1556
rect 4670 1545 5069 1551
rect 5084 1550 5123 1572
rect 5196 1560 5224 1572
rect 5260 1563 5312 1572
rect 5266 1560 5312 1563
rect 5327 1560 5340 1600
rect 5404 1599 5728 1600
rect 5738 1599 5756 1640
rect 5773 1622 6176 1642
rect 5773 1604 5974 1622
rect 6028 1604 6074 1622
rect 6142 1616 6176 1622
rect 6195 1676 6230 1688
rect 6297 1676 6967 1688
rect 7075 1679 7141 1688
rect 6195 1675 6967 1676
rect 6195 1616 6229 1675
rect 6297 1654 6355 1675
rect 6385 1665 6967 1675
rect 7075 1665 7093 1668
rect 7145 1665 7179 1688
rect 7198 1665 7232 1688
rect 7249 1665 7283 1688
rect 6385 1663 7175 1665
rect 7179 1663 7221 1665
rect 6385 1654 7221 1663
rect 7232 1654 7283 1665
rect 6297 1631 7187 1654
rect 7198 1631 7221 1654
rect 6306 1626 6975 1631
rect 6976 1626 7003 1631
rect 6306 1616 6967 1626
rect 6975 1620 6976 1626
rect 7035 1620 7093 1631
rect 7111 1626 7181 1631
rect 7198 1626 7232 1631
rect 5773 1601 5986 1604
rect 6016 1601 6074 1604
rect 5773 1599 6074 1601
rect 5404 1588 6074 1599
rect 5412 1564 5438 1588
rect 5457 1575 6074 1588
rect 5457 1569 5580 1575
rect 5588 1574 6074 1575
rect 6091 1604 6176 1616
rect 6187 1604 6967 1616
rect 6091 1582 6967 1604
rect 6971 1618 7093 1620
rect 6971 1604 7071 1618
rect 6971 1601 7075 1604
rect 6971 1586 7081 1601
rect 6091 1574 6125 1582
rect 6142 1574 6176 1582
rect 6195 1574 6229 1582
rect 6315 1580 6967 1582
rect 7035 1581 7081 1586
rect 7123 1581 7232 1626
rect 5588 1569 6233 1574
rect 5457 1564 5492 1569
rect 5512 1564 5525 1569
rect 5184 1550 5218 1560
rect 5272 1550 5306 1560
rect 5084 1546 5375 1550
rect 5412 1546 5492 1564
rect 5500 1546 5558 1564
rect 5686 1563 5986 1569
rect 6016 1563 6066 1569
rect 6072 1563 6233 1569
rect 5599 1546 5665 1559
rect 5686 1546 6233 1563
rect 4670 1516 4740 1545
rect 4758 1516 4816 1545
rect 4876 1522 4934 1545
rect 4964 1522 5022 1545
rect 5084 1529 6233 1546
rect 4888 1518 4922 1522
rect 4976 1518 5010 1522
rect 4685 1512 4716 1516
rect 4770 1512 4804 1516
rect 5084 1499 5860 1529
rect 5866 1520 6233 1529
rect 6283 1520 6286 1574
rect 6315 1573 6975 1580
rect 6297 1557 6309 1561
rect 6315 1557 6355 1573
rect 6385 1557 6975 1573
rect 6297 1528 6343 1557
rect 6397 1552 6975 1557
rect 6976 1554 7003 1580
rect 7031 1572 7106 1581
rect 7107 1572 7232 1581
rect 7031 1570 7232 1572
rect 7030 1563 7232 1570
rect 7249 1567 7283 1654
rect 7302 1612 7336 1688
rect 7404 1679 7462 1694
rect 7470 1679 7970 1694
rect 7404 1673 7452 1679
rect 7340 1639 7452 1673
rect 7470 1640 7488 1679
rect 7382 1633 7402 1639
rect 7404 1623 7406 1639
rect 7410 1629 7452 1639
rect 7410 1623 7456 1629
rect 7366 1612 7468 1623
rect 7498 1612 7970 1679
rect 7302 1605 7970 1612
rect 7302 1601 7337 1605
rect 7347 1603 7970 1605
rect 7987 1702 8339 1711
rect 8356 1702 8708 1900
rect 7987 1658 8708 1702
rect 7987 1656 8339 1658
rect 8356 1656 8708 1658
rect 7987 1645 8708 1656
rect 8725 1649 9077 1957
rect 7987 1624 8691 1645
rect 8742 1637 9077 1649
rect 7987 1622 8346 1624
rect 8356 1622 8691 1624
rect 7987 1614 8339 1622
rect 8346 1614 8691 1622
rect 7347 1601 7977 1603
rect 7030 1554 7181 1563
rect 6976 1552 7018 1554
rect 6397 1550 7018 1552
rect 7030 1550 7194 1554
rect 6397 1548 7030 1550
rect 7031 1548 7052 1550
rect 7060 1548 7194 1550
rect 6397 1528 7018 1548
rect 7019 1538 7194 1548
rect 7198 1538 7232 1563
rect 7019 1535 7232 1538
rect 5866 1506 5968 1520
rect 5984 1514 6233 1520
rect 6270 1514 6295 1520
rect 6297 1514 6366 1528
rect 6407 1516 7018 1528
rect 5984 1510 6366 1514
rect 5984 1506 6233 1510
rect 6249 1506 6366 1510
rect 5872 1499 5940 1506
rect 4719 1480 4838 1497
rect 4854 1484 5069 1497
rect 4470 1473 4522 1478
rect 3917 1462 4340 1473
rect 3917 1450 3952 1462
rect 3960 1450 4340 1462
rect 3917 1439 4340 1450
rect 4388 1461 4534 1473
rect 4388 1444 4550 1461
rect 4570 1444 4638 1478
rect 4683 1478 4838 1480
rect 4683 1474 4758 1478
rect 4683 1463 4769 1474
rect 4930 1463 5035 1484
rect 4683 1444 4753 1463
rect 5038 1457 5069 1484
rect 5084 1494 5940 1499
rect 5946 1494 6072 1506
rect 6088 1494 6125 1506
rect 6142 1494 6366 1506
rect 5084 1492 6072 1494
rect 5084 1482 5142 1492
rect 5172 1486 5230 1492
rect 5296 1491 6072 1492
rect 5272 1486 6072 1491
rect 5172 1484 6072 1486
rect 5172 1482 5860 1484
rect 5088 1478 5130 1482
rect 5184 1478 5218 1482
rect 5272 1478 5306 1482
rect 5088 1457 5122 1478
rect 5317 1457 5860 1482
rect 5934 1482 6072 1484
rect 5934 1473 6008 1482
rect 6022 1473 6072 1482
rect 5928 1467 6074 1473
rect 6091 1467 6190 1494
rect 5868 1461 5926 1467
rect 5928 1461 6190 1467
rect 3917 1427 3951 1439
rect 4031 1429 4065 1433
rect 4119 1429 4153 1433
rect 4019 1427 4077 1429
rect 4107 1427 4165 1429
rect 4184 1427 4202 1439
rect 4206 1427 4340 1439
rect 3917 1420 4340 1427
rect 4350 1420 4753 1444
rect 3917 1404 4753 1420
rect 4984 1429 5035 1457
rect 4984 1423 5027 1429
rect 5038 1423 5068 1457
rect 5080 1423 5860 1457
rect 5864 1454 5898 1461
rect 5902 1454 6190 1461
rect 5864 1428 6190 1454
rect 6195 1480 6366 1494
rect 6387 1497 7018 1516
rect 7030 1504 7065 1535
rect 7072 1529 7232 1535
rect 7238 1549 7283 1567
rect 7300 1578 7977 1601
rect 7987 1588 8346 1614
rect 8356 1589 8691 1614
rect 8708 1590 9077 1637
rect 9094 1991 10718 1993
rect 9094 1976 9866 1991
rect 9880 1986 10711 1991
rect 9094 1958 9565 1976
rect 9596 1968 9866 1976
rect 9618 1958 9866 1968
rect 9094 1940 9564 1958
rect 9738 1947 9764 1958
rect 9832 1957 9866 1958
rect 9916 1970 10711 1986
rect 9916 1963 10719 1970
rect 10792 1969 10826 2013
rect 10845 1997 10879 2013
rect 10947 2001 10979 2028
rect 10845 1969 10903 1997
rect 10792 1963 10903 1969
rect 9916 1957 10711 1963
rect 9094 1597 9429 1940
rect 9463 1674 9564 1940
rect 9636 1916 9664 1938
rect 9708 1916 9764 1947
rect 9772 1924 10711 1957
rect 9636 1900 9676 1916
rect 9706 1900 9764 1916
rect 9636 1873 9764 1900
rect 9618 1823 9764 1873
rect 9832 1923 10711 1924
rect 9832 1896 9866 1923
rect 9916 1919 10711 1923
rect 10811 1929 10835 1963
rect 10845 1929 10903 1963
rect 10811 1923 10881 1929
rect 9916 1903 10694 1919
rect 9638 1822 9664 1823
rect 9624 1810 9670 1819
rect 9624 1809 9678 1810
rect 9706 1809 9758 1819
rect 9624 1795 9690 1809
rect 9707 1807 9772 1809
rect 9630 1776 9690 1795
rect 9708 1795 9772 1807
rect 9708 1776 9766 1795
rect 9630 1742 9766 1776
rect 9630 1726 9690 1742
rect 9630 1674 9678 1726
rect 9718 1674 9766 1742
rect 9463 1640 9565 1674
rect 9618 1656 9778 1674
rect 9618 1641 9824 1656
rect 9612 1640 9824 1641
rect 9832 1640 9880 1896
rect 9916 1887 10711 1903
rect 10071 1880 10711 1887
rect 10071 1869 10694 1880
rect 10811 1869 10826 1923
rect 10071 1861 10711 1869
rect 10792 1861 10826 1869
rect 10845 1861 10879 1923
rect 10993 1906 11027 2060
rect 11046 1906 11080 2060
rect 11161 2076 11204 2092
rect 11214 2081 11254 2110
rect 11214 2076 11248 2081
rect 11161 2070 11250 2076
rect 11161 2060 11195 2070
rect 11214 2060 11248 2070
rect 11161 1994 11248 2060
rect 11362 2053 11396 2115
rect 11415 2053 11449 2115
rect 11547 2104 11813 2118
rect 11904 2112 11988 2118
rect 11530 2075 11813 2104
rect 11926 2085 11942 2112
rect 11899 2079 11942 2085
rect 11974 2079 11976 2090
rect 12100 2089 12134 2107
rect 12285 2098 12424 2169
rect 12654 2162 12939 2185
rect 13013 2167 13291 2198
rect 13375 2186 13500 2216
rect 12468 2152 12939 2162
rect 12654 2116 12922 2152
rect 13023 2133 13291 2167
rect 13356 2182 13514 2186
rect 13356 2152 13504 2182
rect 13375 2142 13409 2152
rect 13416 2148 13447 2152
rect 13420 2142 13478 2148
rect 12987 2132 13291 2133
rect 12654 2108 12908 2116
rect 12522 2098 12557 2107
rect 12100 2079 12170 2089
rect 11530 2057 11818 2075
rect 11360 2047 11449 2053
rect 11160 1960 11248 1994
rect 11262 1975 11294 2026
rect 11360 2013 11396 2047
rect 11415 2013 11449 2047
rect 11547 2039 11818 2057
rect 11360 2007 11449 2013
rect 10991 1900 11080 1906
rect 10991 1895 11027 1900
rect 10987 1866 11027 1895
rect 11046 1868 11080 1900
rect 11161 1916 11195 1960
rect 11214 1944 11248 1960
rect 11316 1948 11348 1975
rect 11214 1916 11272 1944
rect 11362 1922 11396 2007
rect 11161 1910 11272 1916
rect 11161 1902 11204 1910
rect 11214 1902 11272 1910
rect 11161 1876 11272 1902
rect 11316 1885 11396 1922
rect 11328 1881 11396 1885
rect 11161 1870 11250 1876
rect 11161 1868 11195 1870
rect 11214 1868 11248 1870
rect 11362 1868 11396 1881
rect 11046 1866 11084 1868
rect 10991 1862 11081 1866
rect 11142 1862 11396 1868
rect 10991 1861 11396 1862
rect 10071 1860 11396 1861
rect 10071 1844 11027 1860
rect 10071 1834 10493 1844
rect 10623 1827 11027 1844
rect 11046 1853 11396 1860
rect 11415 1921 11449 2007
rect 11530 1974 11818 2039
rect 11899 2053 12170 2079
rect 12285 2053 12557 2098
rect 11899 2043 12188 2053
rect 12249 2046 12557 2053
rect 12618 2099 12908 2108
rect 12987 2099 13308 2132
rect 13382 2122 13409 2142
rect 13416 2132 13482 2142
rect 12618 2063 12925 2099
rect 12618 2046 12776 2063
rect 11899 2009 12170 2043
rect 11899 2008 12188 2009
rect 11898 1993 12188 2008
rect 12249 1993 12556 2046
rect 12642 2006 12671 2044
rect 12855 2012 12925 2063
rect 11898 1974 12187 1993
rect 11530 1955 11831 1974
rect 11529 1940 11831 1955
rect 11880 1940 12187 1974
rect 12268 1951 12556 1993
rect 12664 1979 12671 2006
rect 11529 1921 11818 1940
rect 11415 1887 11462 1921
rect 11517 1907 11818 1921
rect 11511 1887 11818 1907
rect 11899 1897 12187 1940
rect 12285 1925 12556 1951
rect 11415 1853 11449 1887
rect 11046 1847 11449 1853
rect 11046 1834 11396 1847
rect 10623 1817 10826 1827
rect 10845 1817 10879 1827
rect 10845 1815 10860 1817
rect 10677 1798 10860 1815
rect 10440 1783 10860 1798
rect 10879 1798 11027 1815
rect 11046 1808 11080 1834
rect 11180 1813 11195 1834
rect 11161 1808 11195 1813
rect 11214 1808 11248 1834
rect 11356 1813 11396 1834
rect 11415 1813 11449 1847
rect 11360 1808 11449 1813
rect 11046 1807 11449 1808
rect 11530 1807 11818 1887
rect 11898 1863 12187 1897
rect 12263 1879 12556 1925
rect 12637 1973 12671 1979
rect 12680 1973 12714 2006
rect 12838 1973 12925 2012
rect 12637 1947 12925 1973
rect 13023 2080 13295 2099
rect 13380 2090 13409 2122
rect 13380 2084 13464 2090
rect 13402 2080 13418 2084
rect 13023 2057 13313 2080
rect 13402 2069 13479 2080
rect 13402 2057 13468 2069
rect 13023 2056 13562 2057
rect 13576 2056 13610 2090
rect 13023 2046 13610 2056
rect 13023 2002 13294 2046
rect 13406 2044 13464 2046
rect 13023 1992 13295 2002
rect 13023 1963 13313 1992
rect 13005 1958 13313 1963
rect 13362 1968 13508 2002
rect 13362 1958 13409 1968
rect 13005 1947 13294 1958
rect 12637 1937 12926 1947
rect 12637 1913 12944 1937
rect 12268 1867 12556 1879
rect 11046 1800 11396 1807
rect 11046 1798 11081 1800
rect 11142 1799 11300 1800
rect 11322 1799 11396 1800
rect 10879 1793 11099 1798
rect 10440 1781 10712 1783
rect 10308 1728 10343 1762
rect 9939 1675 9974 1709
rect 9463 1639 9564 1640
rect 9570 1639 9880 1640
rect 9463 1622 9880 1639
rect 9905 1622 9920 1656
rect 9463 1605 9604 1622
rect 9094 1596 9463 1597
rect 8708 1589 9060 1590
rect 7987 1579 8339 1588
rect 8356 1583 8708 1589
rect 8742 1586 9060 1589
rect 9111 1586 9463 1596
rect 9477 1595 9604 1605
rect 8742 1583 9463 1586
rect 8356 1580 9463 1583
rect 7300 1573 7337 1578
rect 7394 1576 7446 1578
rect 7300 1550 7352 1573
rect 7410 1571 7446 1576
rect 7400 1566 7446 1571
rect 7448 1566 7506 1572
rect 7514 1569 7977 1578
rect 7994 1569 8339 1579
rect 7400 1550 7510 1566
rect 7514 1559 7970 1569
rect 7977 1559 8339 1569
rect 7514 1550 7977 1559
rect 7292 1549 7977 1550
rect 7238 1539 7977 1549
rect 7238 1533 7953 1539
rect 7072 1513 7118 1529
rect 7125 1513 7232 1529
rect 7072 1504 7232 1513
rect 7030 1497 7232 1504
rect 7249 1525 7953 1533
rect 7970 1525 7977 1539
rect 7994 1525 8339 1559
rect 7249 1517 7970 1525
rect 7977 1517 8339 1525
rect 7249 1516 7953 1517
rect 7249 1511 7352 1516
rect 7354 1511 7394 1516
rect 7400 1511 7446 1516
rect 7249 1507 7346 1511
rect 7354 1507 7398 1511
rect 7400 1507 7434 1511
rect 7448 1510 7506 1516
rect 6387 1485 7228 1497
rect 6195 1464 6256 1480
rect 6286 1469 6366 1480
rect 6385 1469 7228 1485
rect 6286 1464 7228 1469
rect 7249 1473 7340 1507
rect 7354 1489 7424 1507
rect 7348 1482 7424 1489
rect 7444 1504 7510 1510
rect 7514 1504 7953 1516
rect 7444 1498 7953 1504
rect 7444 1482 7510 1498
rect 7514 1483 7953 1498
rect 7970 1507 7977 1517
rect 7994 1507 8339 1517
rect 7970 1483 8339 1507
rect 7514 1482 7970 1483
rect 7348 1477 7970 1482
rect 7977 1477 8339 1483
rect 7348 1473 8339 1477
rect 7249 1467 8339 1473
rect 7249 1466 7283 1467
rect 7292 1466 7336 1467
rect 6195 1433 6244 1464
rect 6251 1433 6256 1464
rect 6297 1463 7228 1464
rect 7232 1463 7239 1465
rect 7249 1464 7336 1466
rect 7340 1464 7406 1467
rect 7416 1464 8339 1467
rect 7249 1463 8339 1464
rect 6297 1458 6977 1463
rect 6984 1458 7018 1463
rect 7030 1458 7106 1463
rect 6297 1435 7106 1458
rect 6297 1433 6366 1435
rect 6193 1428 6366 1433
rect 6385 1429 7106 1435
rect 7135 1429 7232 1463
rect 5864 1427 6125 1428
rect 4930 1404 4969 1418
rect 3917 1394 4965 1404
rect 3917 1387 4320 1394
rect 4331 1387 4350 1394
rect 4352 1387 4965 1394
rect 3917 1370 4965 1387
rect 3917 1352 4753 1370
rect 4896 1361 4927 1370
rect 4772 1352 4821 1360
rect 4902 1355 4923 1361
rect 4930 1352 4965 1370
rect 3917 1338 4787 1352
rect 3229 1321 3632 1338
rect 3179 1320 3632 1321
rect 3650 1330 4787 1338
rect 4874 1342 4901 1351
rect 4931 1342 4965 1352
rect 3179 1304 3629 1320
rect 3650 1318 4789 1330
rect 4833 1323 4867 1327
rect 4874 1323 4965 1342
rect 3650 1304 4753 1318
rect 4772 1308 4789 1318
rect 3179 1302 3646 1304
rect 3650 1302 3708 1304
rect 3744 1302 3774 1304
rect 2583 1286 2649 1289
rect 2583 1248 2584 1286
rect 2599 1282 2633 1286
rect 2757 1281 3774 1302
rect 3841 1291 4753 1304
rect 4821 1302 4873 1323
rect 4757 1291 4873 1302
rect 4874 1308 4967 1323
rect 4984 1308 5018 1423
rect 5035 1380 5069 1423
rect 5088 1389 5122 1423
rect 5266 1414 5296 1423
rect 5300 1420 5860 1423
rect 5868 1421 5926 1427
rect 5928 1420 5930 1427
rect 5934 1420 6125 1427
rect 6142 1420 6176 1428
rect 5300 1417 6176 1420
rect 6193 1419 6355 1428
rect 6385 1420 7232 1429
rect 6385 1419 6967 1420
rect 6193 1417 6344 1419
rect 5300 1416 6344 1417
rect 5088 1380 5136 1389
rect 5168 1380 5170 1398
rect 5300 1395 6114 1416
rect 5266 1386 6114 1395
rect 6142 1392 6176 1416
rect 6125 1386 6176 1392
rect 6193 1412 6244 1416
rect 6193 1391 6239 1412
rect 6281 1391 6286 1416
rect 6293 1391 6343 1416
rect 6397 1411 6967 1419
rect 6971 1411 7232 1420
rect 7239 1462 8339 1463
rect 8346 1569 9463 1580
rect 9480 1586 9604 1595
rect 9674 1616 9708 1620
rect 9674 1592 9756 1616
rect 9658 1588 9756 1592
rect 9674 1586 9796 1588
rect 8346 1555 9429 1569
rect 8346 1553 8709 1555
rect 8346 1489 8390 1553
rect 8638 1551 8709 1553
rect 8724 1551 9429 1555
rect 8638 1549 9429 1551
rect 8638 1533 8691 1549
rect 8427 1497 8691 1533
rect 8742 1543 9429 1549
rect 9480 1560 9587 1586
rect 9480 1552 9598 1560
rect 9612 1552 9638 1586
rect 9647 1575 9800 1586
rect 9650 1563 9800 1575
rect 9647 1552 9800 1563
rect 9832 1552 9880 1622
rect 8742 1535 9463 1543
rect 8742 1499 9440 1535
rect 8742 1497 9429 1499
rect 8427 1489 9429 1497
rect 8346 1463 9429 1489
rect 9480 1490 9604 1552
rect 9690 1548 9722 1552
rect 9728 1542 9760 1552
rect 9846 1542 9880 1552
rect 9672 1532 9762 1542
rect 9712 1524 9762 1532
rect 9712 1520 9778 1524
rect 9712 1504 9766 1520
rect 9730 1495 9760 1504
rect 9708 1490 9784 1495
rect 9852 1490 9880 1542
rect 9480 1483 9587 1490
rect 7239 1455 8322 1462
rect 7239 1411 7283 1455
rect 6397 1400 7221 1411
rect 6397 1391 6968 1400
rect 5266 1380 5882 1386
rect 4874 1291 4901 1308
rect 4931 1291 5018 1308
rect 5024 1364 5882 1380
rect 5912 1384 5933 1386
rect 5940 1384 5974 1386
rect 5912 1364 5974 1384
rect 5024 1352 5870 1364
rect 5918 1361 5974 1364
rect 5024 1338 5860 1352
rect 5924 1338 5974 1361
rect 6016 1338 6022 1386
rect 6038 1338 6125 1386
rect 5024 1327 6106 1338
rect 5024 1315 6074 1327
rect 6076 1315 6106 1327
rect 5024 1304 6106 1315
rect 6142 1304 6176 1386
rect 5024 1291 5860 1304
rect 3841 1290 4736 1291
rect 4746 1290 5860 1291
rect 3841 1281 5860 1290
rect 2631 1256 2649 1278
rect 2757 1256 5860 1281
rect 2441 1208 2505 1216
rect 2631 1208 2681 1256
rect 2362 1206 2422 1208
rect 2111 1198 2161 1202
rect 2214 1198 2219 1202
rect 1990 1195 2362 1198
rect 1990 1193 2314 1195
rect 1990 1188 2342 1193
rect 1990 1181 2069 1188
rect 2072 1181 2087 1188
rect 926 1178 2101 1181
rect 2108 1178 2342 1188
rect 926 1166 2342 1178
rect 2354 1177 2362 1195
rect 2351 1166 2362 1177
rect 926 1164 1382 1166
rect 726 1134 784 1144
rect 814 1134 872 1144
rect 136 1100 174 1134
rect 205 1126 644 1134
rect 650 1126 684 1134
rect 737 1126 767 1134
rect 770 1126 784 1134
rect 850 1126 890 1134
rect 904 1130 1382 1164
rect 926 1126 1382 1130
rect 205 1123 1382 1126
rect 205 1122 890 1123
rect 926 1122 1382 1123
rect 1383 1156 1417 1166
rect 1423 1156 1429 1166
rect 1607 1164 2362 1166
rect 1383 1146 1429 1156
rect 1458 1156 1514 1164
rect 1583 1156 1598 1162
rect 1458 1146 1526 1156
rect 1568 1146 1602 1156
rect 1607 1148 2053 1164
rect 2072 1148 2106 1164
rect 2186 1155 2220 1159
rect 2274 1155 2308 1160
rect 1607 1146 2029 1148
rect 1383 1122 1426 1146
rect 1429 1141 1438 1146
rect 1458 1130 2029 1146
rect 1468 1122 2029 1130
rect 2038 1147 2053 1148
rect 2038 1122 2067 1147
rect 2069 1140 2130 1148
rect 2174 1140 2232 1155
rect 2069 1139 2232 1140
rect 2069 1126 2220 1139
rect 2262 1126 2320 1155
rect 2328 1146 2362 1164
rect 2388 1146 2422 1206
rect 2436 1206 2505 1208
rect 2543 1206 2601 1208
rect 2631 1206 2689 1208
rect 2436 1194 2475 1206
rect 2441 1182 2475 1194
rect 2328 1138 2422 1146
rect 2436 1174 2475 1182
rect 2543 1196 2563 1206
rect 2582 1196 2601 1206
rect 2543 1179 2601 1196
rect 2643 1191 2689 1206
rect 2757 1206 5861 1256
rect 2643 1179 2677 1191
rect 2757 1179 5870 1206
rect 2505 1178 5870 1179
rect 5874 1178 5882 1304
rect 5912 1292 5986 1304
rect 6016 1293 6037 1304
rect 6038 1293 6074 1304
rect 6016 1292 6022 1293
rect 5937 1283 5970 1292
rect 5927 1246 5970 1283
rect 5972 1246 5992 1252
rect 5927 1236 6034 1246
rect 2436 1146 2486 1174
rect 2505 1168 5882 1178
rect 2505 1166 2529 1168
rect 2505 1146 2524 1166
rect 2533 1148 5882 1168
rect 5936 1177 5970 1236
rect 5974 1212 6034 1236
rect 5974 1202 6024 1212
rect 6038 1177 6072 1293
rect 5936 1168 6086 1177
rect 6091 1168 6125 1304
rect 5936 1164 6125 1168
rect 2533 1146 5870 1148
rect 2436 1138 2482 1146
rect 2505 1145 5870 1146
rect 2505 1138 2589 1145
rect 2613 1138 2677 1145
rect 2328 1132 2677 1138
rect 2328 1126 2374 1132
rect 2388 1126 2677 1132
rect 2069 1122 2339 1126
rect 2348 1124 2677 1126
rect 2689 1124 2734 1145
rect 2348 1122 2734 1124
rect 2757 1144 5870 1145
rect 5874 1144 5882 1148
rect 5958 1146 6125 1164
rect 5958 1144 6126 1146
rect 6132 1144 6176 1304
rect 2757 1134 6176 1144
rect 2757 1129 6086 1134
rect 2757 1122 5596 1129
rect 205 1113 5596 1122
rect 205 1111 5481 1113
rect 205 1109 2069 1111
rect 2072 1109 5481 1111
rect 5500 1109 5558 1113
rect 5562 1109 5596 1113
rect 5600 1118 5646 1129
rect 5669 1124 5703 1129
rect 5600 1109 5637 1118
rect 5669 1109 5717 1124
rect 5722 1109 5756 1129
rect 5763 1109 5797 1129
rect 5816 1126 6086 1129
rect 6091 1126 6176 1134
rect 6185 1388 6968 1391
rect 6971 1388 7221 1400
rect 6185 1382 7221 1388
rect 7232 1401 7239 1411
rect 7249 1401 7283 1411
rect 6185 1377 7206 1382
rect 7232 1377 7283 1401
rect 6185 1370 7030 1377
rect 7060 1370 7194 1377
rect 6185 1333 6975 1370
rect 6185 1213 6229 1333
rect 6281 1248 6286 1333
rect 6293 1323 6355 1333
rect 6377 1323 6975 1333
rect 6293 1321 6975 1323
rect 6976 1345 7003 1370
rect 7065 1363 7131 1370
rect 7145 1366 7194 1370
rect 7198 1371 7232 1377
rect 7239 1371 7283 1377
rect 7198 1370 7228 1371
rect 7232 1370 7283 1371
rect 7065 1345 7141 1363
rect 6976 1329 7141 1345
rect 6976 1321 7105 1329
rect 7145 1327 7179 1366
rect 7198 1343 7283 1370
rect 7198 1339 7233 1343
rect 7239 1339 7283 1343
rect 7292 1449 8322 1455
rect 7292 1445 7971 1449
rect 7977 1445 8322 1449
rect 7292 1444 8322 1445
rect 8346 1453 8691 1463
rect 8742 1458 9429 1463
rect 8742 1453 9182 1458
rect 8346 1444 9182 1453
rect 7292 1443 9182 1444
rect 7292 1430 7953 1443
rect 7292 1371 7336 1430
rect 7382 1404 7394 1430
rect 7404 1423 7406 1430
rect 7410 1427 7953 1430
rect 7977 1429 9182 1443
rect 7977 1427 8702 1429
rect 7410 1423 8702 1427
rect 7404 1414 8702 1423
rect 7404 1408 7462 1414
rect 7470 1408 8702 1414
rect 7372 1398 7394 1404
rect 7410 1398 7462 1408
rect 7492 1407 8702 1408
rect 7492 1398 8074 1407
rect 7372 1376 7462 1398
rect 7498 1394 8074 1398
rect 7494 1391 8074 1394
rect 7372 1371 7452 1376
rect 7483 1371 7492 1375
rect 7494 1374 8075 1391
rect 8094 1374 8128 1407
rect 8132 1374 8188 1407
rect 8190 1374 8199 1407
rect 8232 1389 8276 1407
rect 8280 1389 8288 1407
rect 8230 1376 8288 1389
rect 8305 1393 8702 1407
rect 8305 1388 8691 1393
rect 8230 1374 8320 1376
rect 8346 1374 8691 1388
rect 8742 1380 9182 1429
rect 9201 1387 9235 1458
rect 9265 1387 9271 1458
rect 9343 1451 9397 1458
rect 9463 1457 9587 1483
rect 9612 1486 9812 1490
rect 9612 1473 9784 1486
rect 9612 1457 9818 1473
rect 9463 1456 9818 1457
rect 9832 1456 9880 1490
rect 9281 1437 9339 1451
rect 9281 1433 9351 1437
rect 9281 1431 9339 1433
rect 9281 1429 9305 1431
rect 9361 1429 9391 1451
rect 9463 1446 9880 1456
rect 9281 1417 9377 1429
rect 9293 1391 9299 1417
rect 9303 1397 9373 1417
rect 8742 1377 9190 1380
rect 7494 1371 8074 1374
rect 7292 1357 8074 1371
rect 7292 1339 8075 1357
rect 8132 1354 8691 1374
rect 7198 1337 8075 1339
rect 7125 1323 7179 1327
rect 7113 1321 7179 1323
rect 7239 1321 7283 1337
rect 7292 1321 7336 1337
rect 7356 1321 7370 1337
rect 7372 1321 8075 1337
rect 6293 1320 8075 1321
rect 6293 1305 6343 1320
rect 6293 1295 6355 1305
rect 6377 1304 8075 1320
rect 6377 1302 7510 1304
rect 6377 1295 7528 1302
rect 6293 1292 7528 1295
rect 6293 1289 6355 1292
rect 6363 1289 7528 1292
rect 6293 1272 7528 1289
rect 7531 1272 8075 1304
rect 6293 1255 8075 1272
rect 6293 1248 6355 1255
rect 6363 1249 8075 1255
rect 6281 1218 6355 1248
rect 6385 1246 8075 1249
rect 6385 1239 7652 1246
rect 6391 1234 7652 1239
rect 6391 1221 7540 1234
rect 6185 1174 6239 1213
rect 6293 1179 6355 1218
rect 6397 1213 7540 1221
rect 6387 1208 7540 1213
rect 7548 1208 7562 1234
rect 7608 1208 7652 1234
rect 6376 1196 6385 1207
rect 6387 1195 7652 1208
rect 6387 1179 6465 1195
rect 6501 1179 7652 1195
rect 6249 1174 7652 1179
rect 6185 1172 7494 1174
rect 6185 1168 7506 1172
rect 7516 1168 7546 1174
rect 7608 1168 7652 1174
rect 7661 1221 8075 1246
rect 8094 1238 8128 1348
rect 8132 1340 8324 1354
rect 8346 1352 8691 1354
rect 8132 1293 8188 1340
rect 8190 1293 8199 1340
rect 8232 1308 8310 1340
rect 8232 1306 8288 1308
rect 8226 1293 8288 1306
rect 8142 1283 8200 1293
rect 8208 1283 8288 1293
rect 8142 1277 8288 1283
rect 8142 1261 8284 1277
rect 8296 1261 8310 1265
rect 8142 1251 8282 1261
rect 8154 1249 8279 1251
rect 8290 1249 8310 1261
rect 8312 1261 8330 1265
rect 8312 1249 8342 1261
rect 8154 1247 8182 1249
rect 8188 1247 8276 1249
rect 8172 1238 8182 1246
rect 8188 1238 8269 1247
rect 8290 1238 8342 1249
rect 7661 1168 8083 1221
rect 8088 1204 8342 1238
rect 8346 1206 8497 1352
rect 8567 1345 8617 1351
rect 8543 1327 8617 1345
rect 8543 1323 8601 1327
rect 8623 1323 8653 1345
rect 8543 1311 8639 1323
rect 8565 1307 8635 1311
rect 8555 1291 8635 1307
rect 8659 1305 8679 1307
rect 8659 1291 8683 1305
rect 8691 1291 8699 1327
rect 8700 1291 8711 1323
rect 8540 1280 8711 1291
rect 8551 1279 8711 1280
rect 8356 1204 8497 1206
rect 8088 1191 8128 1204
rect 8154 1196 8266 1204
rect 8150 1195 8266 1196
rect 8150 1191 8276 1195
rect 6185 1145 8083 1168
rect 6185 1134 6283 1145
rect 6293 1134 6339 1145
rect 6356 1143 6455 1145
rect 6185 1126 6339 1134
rect 5816 1119 6339 1126
rect 6353 1125 6455 1143
rect 6341 1119 6455 1125
rect 5816 1111 6455 1119
rect 6501 1142 8083 1145
rect 8094 1144 8128 1191
rect 8142 1170 8282 1191
rect 8142 1154 8200 1170
rect 8208 1164 8282 1170
rect 8142 1144 8194 1154
rect 8202 1144 8282 1164
rect 8290 1144 8342 1204
rect 8346 1155 8497 1204
rect 8511 1257 8711 1279
rect 8511 1189 8563 1257
rect 8571 1245 8651 1257
rect 8571 1233 8591 1245
rect 8577 1229 8591 1233
rect 8611 1233 8651 1245
rect 8659 1245 8683 1257
rect 8659 1233 8679 1245
rect 8611 1229 8653 1233
rect 8587 1227 8653 1229
rect 8655 1227 8657 1233
rect 8665 1229 8679 1233
rect 8691 1229 8699 1257
rect 8700 1233 8711 1257
rect 8583 1195 8657 1227
rect 8581 1189 8679 1195
rect 8511 1175 8679 1189
rect 8511 1163 8657 1175
rect 8346 1144 8480 1155
rect 8094 1142 8480 1144
rect 5816 1110 6475 1111
rect 5816 1109 5870 1110
rect 5874 1109 6475 1110
rect 6501 1110 8480 1142
rect 8483 1117 8497 1155
rect 8519 1157 8569 1163
rect 8577 1161 8655 1163
rect 8577 1159 8645 1161
rect 8577 1157 8643 1159
rect 8519 1155 8643 1157
rect 8519 1151 8591 1155
rect 8519 1117 8617 1151
rect 8637 1117 8671 1127
rect 6501 1109 8128 1110
rect 191 1102 8128 1109
rect 8142 1102 8194 1110
rect 8202 1102 8330 1110
rect 8331 1102 8342 1110
rect 8356 1103 8480 1110
rect 8356 1102 8497 1103
rect 191 1100 8497 1102
rect 178 1098 8497 1100
rect 178 1092 6475 1098
rect 178 1080 5965 1092
rect 191 1076 5965 1080
rect 191 1069 5428 1076
rect 5447 1069 5965 1076
rect 191 1066 5965 1069
rect 191 1050 696 1066
rect 178 1042 696 1050
rect 712 1042 772 1066
rect 178 1034 644 1042
rect 180 969 189 1004
rect 191 986 644 1034
rect 650 1012 684 1042
rect 720 1024 772 1042
rect 788 1060 5965 1066
rect 788 1058 2232 1060
rect 2261 1058 5965 1060
rect 788 1048 1438 1058
rect 1468 1053 2232 1058
rect 1448 1048 2232 1053
rect 788 1046 2232 1048
rect 2260 1056 5965 1058
rect 6006 1056 6008 1092
rect 6038 1090 6086 1092
rect 6018 1058 6086 1090
rect 6091 1058 6166 1092
rect 6018 1056 6166 1058
rect 6185 1086 6475 1092
rect 6478 1093 8497 1098
rect 8525 1093 8671 1117
rect 8725 1093 9190 1377
rect 9201 1376 9271 1387
rect 9303 1381 9355 1397
rect 9403 1387 9417 1397
rect 9397 1385 9417 1387
rect 9397 1381 9421 1385
rect 9429 1381 9437 1433
rect 9201 1347 9235 1376
rect 9303 1366 9349 1381
rect 9261 1359 9295 1363
rect 9307 1359 9349 1366
rect 9355 1363 9371 1367
rect 9355 1359 9383 1363
rect 9249 1347 9301 1359
rect 9309 1351 9349 1359
rect 9369 1351 9389 1359
rect 9309 1347 9329 1351
rect 9361 1347 9389 1351
rect 9397 1351 9437 1381
rect 9397 1347 9417 1351
rect 9429 1347 9437 1351
rect 9438 1347 9449 1429
rect 9201 1313 9216 1347
rect 9243 1339 9449 1347
rect 9463 1402 9604 1446
rect 9672 1434 9724 1446
rect 9772 1436 9786 1441
rect 9798 1436 9806 1446
rect 9672 1419 9718 1434
rect 9772 1431 9806 1436
rect 9630 1403 9638 1407
rect 9650 1403 9664 1407
rect 9676 1403 9718 1419
rect 9618 1402 9670 1403
rect 9678 1402 9718 1403
rect 9738 1403 9752 1407
rect 9738 1402 9758 1403
rect 9766 1402 9806 1431
rect 9807 1402 9818 1446
rect 9463 1368 9587 1402
rect 9612 1368 9818 1402
rect 9243 1335 9440 1339
rect 9243 1313 9443 1335
rect 9201 1199 9235 1313
rect 9249 1311 9301 1313
rect 9249 1283 9295 1311
rect 9321 1301 9395 1313
rect 9321 1283 9417 1301
rect 9249 1281 9417 1283
rect 9249 1279 9409 1281
rect 9249 1269 9395 1279
rect 9261 1265 9295 1269
rect 9337 1267 9389 1269
rect 9337 1265 9383 1267
rect 9337 1261 9379 1265
rect 9293 1245 9351 1251
rect 9289 1231 9355 1245
rect 9305 1201 9339 1231
rect 9293 1199 9351 1201
rect 9201 1183 9236 1199
rect 9278 1195 9366 1199
rect 9278 1188 9417 1195
rect 9289 1183 9417 1188
rect 9463 1183 9604 1368
rect 9618 1316 9670 1368
rect 9618 1300 9676 1316
rect 9678 1306 9758 1368
rect 9684 1300 9758 1306
rect 9618 1293 9758 1300
rect 9766 1305 9790 1368
rect 9766 1293 9786 1305
rect 9618 1277 9760 1293
rect 9762 1277 9764 1293
rect 9772 1289 9786 1293
rect 9798 1289 9806 1368
rect 9807 1293 9818 1368
rect 9618 1246 9764 1277
rect 9618 1235 9786 1246
rect 9618 1223 9764 1235
rect 9630 1219 9638 1223
rect 9712 1219 9762 1223
rect 9201 1173 9249 1183
rect 9289 1181 9604 1183
rect 9265 1173 9271 1176
rect 9297 1173 9604 1181
rect 9201 1165 9604 1173
rect 9265 1163 9301 1165
rect 9343 1163 9379 1165
rect 9261 1129 9295 1163
rect 9349 1129 9383 1163
rect 9463 1129 9604 1165
rect 9249 1095 9395 1129
rect 9401 1095 9417 1129
rect 6478 1086 9190 1093
rect 6185 1085 9190 1086
rect 6185 1075 8725 1085
rect 6185 1073 6339 1075
rect 6185 1069 6239 1073
rect 6185 1060 6230 1069
rect 788 1024 1382 1046
rect 650 986 690 1012
rect 711 1000 718 1012
rect 724 1000 1382 1024
rect 711 998 1382 1000
rect 711 990 860 998
rect 711 986 772 990
rect 778 986 860 990
rect 861 986 1382 998
rect 191 972 1382 986
rect 1383 1040 1428 1046
rect 1383 1006 1432 1040
rect 1438 1037 2170 1046
rect 1442 1033 2170 1037
rect 2172 1037 2220 1046
rect 2260 1043 6176 1056
rect 2236 1041 6176 1043
rect 6185 1041 6232 1060
rect 6249 1051 6339 1073
rect 6356 1069 6441 1075
rect 6233 1041 6238 1042
rect 6249 1041 6333 1051
rect 6334 1041 6339 1051
rect 2236 1040 6344 1041
rect 2260 1037 2320 1040
rect 2172 1033 2320 1037
rect 2328 1033 6339 1040
rect 1442 1028 6339 1033
rect 6362 1028 6367 1069
rect 6368 1058 6441 1069
rect 6368 1051 6453 1058
rect 6368 1043 6457 1051
rect 6368 1040 6455 1043
rect 6368 1037 6453 1040
rect 6368 1030 6441 1037
rect 6478 1030 6499 1075
rect 6368 1028 6499 1030
rect 1442 1022 6353 1028
rect 1442 1021 5914 1022
rect 5916 1021 5965 1022
rect 1442 1018 5965 1021
rect 1442 1017 1526 1018
rect 1383 994 1438 1006
rect 1442 996 1514 1017
rect 1448 994 1514 996
rect 1383 972 1514 994
rect 1536 1001 5965 1018
rect 5984 1017 6353 1022
rect 6356 1027 6499 1028
rect 6501 1068 8725 1075
rect 6501 1056 8128 1068
rect 8142 1059 8194 1068
rect 8202 1059 8282 1068
rect 8290 1059 8330 1068
rect 8142 1056 8330 1059
rect 8331 1056 8342 1068
rect 8356 1059 8725 1068
rect 8742 1076 9190 1085
rect 8356 1056 8480 1059
rect 6501 1049 8480 1056
rect 8549 1049 8583 1059
rect 8631 1057 8697 1059
rect 8637 1049 8697 1057
rect 8725 1049 8737 1059
rect 6501 1034 8725 1049
rect 6356 1024 6481 1027
rect 6356 1023 6402 1024
rect 6407 1023 6481 1024
rect 6356 1017 6481 1023
rect 6501 1022 8342 1034
rect 8356 1025 8725 1034
rect 8356 1022 8480 1025
rect 6501 1017 8128 1022
rect 5984 1009 8128 1017
rect 8142 1011 8253 1022
rect 8268 1011 8342 1022
rect 5984 1007 6449 1009
rect 5984 1001 6088 1007
rect 1536 999 6088 1001
rect 1536 976 2320 999
rect 2322 990 6088 999
rect 1528 975 2320 976
rect 2328 987 6086 990
rect 1528 974 2308 975
rect 2328 974 6076 987
rect 6091 986 6176 1007
rect 1528 972 2206 974
rect 191 969 1584 972
rect 144 966 1584 969
rect 1590 966 2206 972
rect 144 962 2206 966
rect 2214 971 2326 974
rect 2214 962 2294 971
rect 144 958 2294 962
rect 2296 965 2326 971
rect 2328 971 6072 974
rect 2328 965 6018 971
rect 2296 960 6018 965
rect 2296 958 6030 960
rect 144 954 6030 958
rect 144 952 6034 954
rect 144 948 644 952
rect 650 950 711 952
rect 712 950 6034 952
rect 650 948 690 950
rect 144 936 690 948
rect 711 947 5965 950
rect 710 943 5965 947
rect 698 936 2298 943
rect 144 926 684 936
rect 690 928 2298 936
rect 2304 938 5965 943
rect 5968 943 6034 950
rect 6038 943 6072 971
rect 6091 973 6126 986
rect 6132 973 6176 986
rect 6091 962 6176 973
rect 6185 1006 6449 1007
rect 6467 1006 8128 1009
rect 8154 1007 8162 1011
rect 8168 1007 8253 1011
rect 6185 983 8128 1006
rect 8168 1001 8248 1007
rect 8262 1001 8342 1011
rect 8168 998 8342 1001
rect 8164 988 8342 998
rect 6185 978 6232 983
rect 6233 978 6238 983
rect 6185 970 6238 978
rect 6180 966 6238 970
rect 6249 966 8128 983
rect 6091 947 6125 962
rect 6082 943 6125 947
rect 6132 945 6176 962
rect 6185 945 6230 966
rect 5968 938 6072 943
rect 6076 939 6128 943
rect 6130 939 6230 945
rect 6076 938 6230 939
rect 2304 931 5914 938
rect 5916 934 6072 938
rect 690 926 2322 928
rect 144 911 2322 926
rect 2328 911 5914 931
rect 144 881 5914 911
rect 144 835 2185 881
rect 2190 875 5914 881
rect 2190 874 4434 875
rect 4436 874 5914 875
rect 2190 871 5914 874
rect 5931 928 6072 934
rect 5931 920 6034 928
rect 6038 920 6072 928
rect 5931 888 6072 920
rect 5931 877 5965 888
rect 5931 874 5974 877
rect 5982 874 6072 888
rect 5931 873 6072 874
rect 5928 871 6072 873
rect 2190 868 6072 871
rect 6082 928 6230 938
rect 6082 924 6125 928
rect 6126 924 6230 928
rect 6249 924 6283 966
rect 6300 926 8128 966
rect 8154 954 8342 988
rect 6297 924 8128 926
rect 6082 895 8128 924
rect 8168 930 8342 954
rect 8168 920 8256 930
rect 8168 913 8248 920
rect 8168 911 8226 913
rect 8234 911 8248 913
rect 8168 901 8248 911
rect 8262 901 8342 930
rect 8346 901 8480 1022
rect 8505 989 8674 1025
rect 8742 1023 8849 1076
rect 8920 1036 9020 1076
rect 8920 1030 8964 1036
rect 8972 1030 8982 1036
rect 9000 1030 9020 1036
rect 9043 1030 9046 1076
rect 8581 955 8593 989
rect 8581 949 8639 955
rect 8168 897 8242 901
rect 8256 897 8330 901
rect 8168 895 8226 897
rect 8256 895 8314 897
rect 6082 890 8314 895
rect 6082 889 6122 890
rect 6126 889 6230 890
rect 6082 874 6128 889
rect 6132 874 6176 889
rect 6185 879 6230 889
rect 6249 879 6283 890
rect 6297 888 8314 890
rect 6297 879 8320 888
rect 6185 874 8320 879
rect 6082 871 8320 874
rect 6082 868 6128 871
rect 2190 862 6128 868
rect 6132 862 6176 871
rect 2190 858 6176 862
rect 6185 862 8320 871
rect 6185 861 8336 862
rect 6185 858 8128 861
rect 2190 845 8128 858
rect 2190 838 6232 845
rect 2190 837 6072 838
rect 2190 835 5914 837
rect 144 826 5914 835
rect 5928 826 5974 837
rect 5984 826 6062 837
rect 6082 826 6176 838
rect 144 820 6176 826
rect 6186 820 6232 838
rect 6249 820 6283 845
rect 6297 830 8128 845
rect 8132 837 8336 861
rect 8132 830 8324 837
rect 6297 829 8324 830
rect 8346 829 8380 901
rect 8382 829 8480 901
rect 8742 898 8838 1023
rect 8918 1020 8964 1030
rect 8918 996 8952 1020
rect 9000 1002 9066 1030
rect 9006 996 9066 1002
rect 8906 993 9066 996
rect 8874 981 9052 993
rect 8874 972 9032 981
rect 9071 976 9074 1076
rect 9094 1030 9190 1076
rect 9094 996 9106 1030
rect 8874 934 9034 972
rect 6297 828 8480 829
rect 6297 820 8173 828
rect 144 814 8173 820
rect 144 788 8100 814
rect 8128 812 8173 814
rect 8174 812 8178 828
rect 144 786 8083 788
rect 144 774 6140 786
rect 6142 774 6176 786
rect 6185 774 6232 786
rect 6249 774 8083 786
rect 8105 776 8128 812
rect 8132 811 8182 812
rect 8208 811 8212 828
rect 8220 822 8278 828
rect 8286 822 8300 828
rect 8220 820 8300 822
rect 8220 811 8292 820
rect 8346 811 8380 828
rect 8382 817 8480 828
rect 8768 853 8838 898
rect 8950 900 8962 934
rect 8950 894 9008 900
rect 9111 888 9190 1030
rect 9265 977 9271 1079
rect 9463 1074 9550 1129
rect 9570 1128 9604 1129
rect 9618 1195 9670 1219
rect 9706 1204 9764 1219
rect 9618 1192 9664 1195
rect 9708 1192 9764 1204
rect 9618 1176 9676 1192
rect 9706 1181 9764 1192
rect 9706 1176 9755 1181
rect 9618 1144 9755 1176
rect 9618 1128 9764 1144
rect 9832 1128 9866 1446
rect 9886 1144 9920 1622
rect 9570 1110 9866 1128
rect 9905 1110 9920 1144
rect 9939 1110 9973 1675
rect 10085 1607 10143 1613
rect 10085 1573 10097 1607
rect 10085 1567 10143 1573
rect 10085 1119 10143 1125
rect 9636 1108 9664 1110
rect 9630 1074 9664 1108
rect 9718 1108 9746 1110
rect 9718 1074 9752 1108
rect 9293 1045 9351 1051
rect 9293 1011 9305 1045
rect 9463 1040 9551 1074
rect 9618 1040 9764 1074
rect 9770 1051 9786 1074
rect 9293 1005 9351 1011
rect 9463 1005 9550 1040
rect 9480 909 9550 1005
rect 9662 992 9720 998
rect 9662 958 9674 992
rect 9832 983 9866 1110
rect 9939 1079 9954 1110
rect 10085 1085 10097 1119
rect 10085 1079 10143 1085
rect 9903 983 10156 1074
rect 10274 1002 10289 1709
rect 10308 1070 10342 1728
rect 10454 1660 10512 1666
rect 10454 1626 10466 1660
rect 10454 1620 10512 1626
rect 10641 1411 10711 1781
rect 10941 1764 11099 1793
rect 11142 1797 11396 1799
rect 11142 1774 11362 1797
rect 11157 1772 11248 1774
rect 11381 1772 11396 1797
rect 11157 1766 11250 1772
rect 11177 1764 11254 1766
rect 10823 1713 10881 1719
rect 10823 1679 10835 1713
rect 10823 1673 10881 1679
rect 10823 1513 10881 1519
rect 10823 1479 10835 1513
rect 10823 1473 10881 1479
rect 10641 1377 10712 1411
rect 11012 1396 11027 1764
rect 11046 1464 11080 1764
rect 11192 1745 11254 1764
rect 11362 1745 11396 1772
rect 11415 1755 11449 1807
rect 11415 1745 11450 1755
rect 11547 1747 11818 1807
rect 11192 1740 11468 1745
rect 11192 1732 11204 1740
rect 11214 1732 11468 1740
rect 11192 1726 11468 1732
rect 11214 1711 11468 1726
rect 11517 1711 11818 1747
rect 11180 1682 11194 1698
rect 11248 1694 11282 1698
rect 11236 1686 11294 1694
rect 11248 1677 11282 1686
rect 11192 1566 11250 1572
rect 11192 1532 11204 1566
rect 11192 1526 11250 1532
rect 11362 1526 11396 1711
rect 11046 1430 11081 1464
rect 11381 1449 11396 1526
rect 11415 1517 11449 1711
rect 11547 1702 11818 1711
rect 11899 1702 12187 1863
rect 12267 1835 12556 1867
rect 12234 1801 12556 1835
rect 12267 1775 12556 1801
rect 12636 1903 12944 1913
rect 12993 1903 13294 1947
rect 13375 1930 13409 1958
rect 12636 1791 12925 1903
rect 12268 1763 12556 1775
rect 12263 1717 12556 1763
rect 12603 1757 12925 1791
rect 13006 1763 13294 1903
rect 13341 1916 13409 1930
rect 13452 1916 13499 1947
rect 13341 1900 13420 1916
rect 13450 1900 13499 1916
rect 13341 1896 13499 1900
rect 13375 1873 13499 1896
rect 13362 1823 13508 1873
rect 13375 1819 13442 1823
rect 13368 1795 13442 1819
rect 12636 1729 12925 1757
rect 13005 1729 13294 1763
rect 12637 1717 12938 1729
rect 11547 1692 11819 1702
rect 11547 1658 11837 1692
rect 11886 1658 12187 1702
rect 11547 1622 11818 1658
rect 11561 1619 11619 1622
rect 11561 1585 11573 1619
rect 11561 1579 11619 1585
rect 11415 1483 11450 1517
rect 11748 1483 11818 1622
rect 11916 1649 12187 1658
rect 12285 1649 12556 1717
rect 12642 1698 12938 1717
rect 11916 1639 12188 1649
rect 11916 1605 12170 1639
rect 11916 1589 12188 1605
rect 12249 1596 12556 1649
rect 12654 1695 12938 1698
rect 12987 1695 13294 1729
rect 13375 1776 13442 1795
rect 13452 1795 13502 1819
rect 13452 1792 13499 1795
rect 13450 1776 13499 1792
rect 13375 1742 13499 1776
rect 13375 1708 13442 1742
rect 13450 1726 13490 1742
rect 12654 1601 12925 1695
rect 13006 1674 13294 1695
rect 13374 1674 13442 1708
rect 13462 1708 13490 1726
rect 13462 1674 13496 1708
rect 13006 1640 13307 1674
rect 13362 1651 13508 1674
rect 13514 1651 13530 1674
rect 13356 1640 13514 1651
rect 13006 1629 13294 1640
rect 13006 1620 13277 1629
rect 12654 1596 12908 1601
rect 12249 1589 12557 1596
rect 11916 1569 12170 1589
rect 11930 1564 11988 1569
rect 11930 1530 11942 1564
rect 12117 1553 12170 1569
rect 12285 1553 12539 1589
rect 12618 1585 12908 1596
rect 13006 1595 13289 1620
rect 11930 1524 11988 1530
rect 12285 1516 12424 1553
rect 12618 1543 12925 1585
rect 13023 1548 13289 1595
rect 13375 1598 13409 1640
rect 13375 1592 13464 1598
rect 13375 1558 13418 1592
rect 13375 1552 13464 1558
rect 13576 1552 13610 2046
rect 12618 1534 12926 1543
rect 12654 1498 12908 1534
rect 13023 1532 13277 1548
rect 13375 1542 13409 1552
rect 13023 1509 13294 1532
rect 13398 1531 13409 1542
rect 11748 1447 11801 1483
rect 13023 1473 13277 1509
rect 13023 1463 13076 1473
rect 10641 1341 10694 1377
rect 10454 1172 10512 1178
rect 10454 1138 10466 1172
rect 10491 1138 10512 1172
rect 10454 1132 10512 1138
rect 10519 1104 10540 1170
rect 10308 1036 10343 1070
rect 10505 1000 10694 1057
rect 9662 952 9720 958
rect 9767 936 9902 983
rect 9903 947 10325 983
rect 9111 873 9336 888
rect 9480 873 9533 909
rect 8768 851 8821 853
rect 8768 833 8838 851
rect 8950 833 8985 851
rect 8768 832 8985 833
rect 9024 832 9204 852
rect 8768 818 9204 832
rect 9265 818 9300 852
rect 9480 835 9590 873
rect 9705 820 9902 936
rect 8382 814 8444 817
rect 8382 811 8434 814
rect 144 765 8083 774
rect 144 760 5925 765
rect 144 716 630 760
rect 650 758 786 760
rect 787 758 5925 760
rect 650 754 798 758
rect 799 754 5925 758
rect 650 750 726 754
rect 738 750 798 754
rect 650 744 798 750
rect 638 742 798 744
rect 828 744 2192 754
rect 2200 744 5925 754
rect 828 742 2278 744
rect 638 738 786 742
rect 638 726 684 738
rect 692 726 784 738
rect 638 716 784 726
rect 814 716 828 740
rect 840 738 2278 742
rect 2279 742 5925 744
rect 2279 738 4384 742
rect 852 726 4384 738
rect 4388 738 5925 742
rect 5928 763 8083 765
rect 5928 744 6074 763
rect 6082 759 8083 763
rect 5928 738 6018 744
rect 6028 738 6074 744
rect 6086 757 8083 759
rect 6086 744 6232 757
rect 6086 738 6140 744
rect 6142 738 6176 744
rect 4388 726 6176 738
rect 852 716 6176 726
rect 144 707 6176 716
rect 6185 707 6232 744
rect 144 682 6232 707
rect 144 674 6076 682
rect 6086 678 6232 682
rect 6098 674 6176 678
rect 6185 674 6230 678
rect 6249 674 6283 757
rect 6297 717 8083 757
rect 6297 700 8125 717
rect 8132 700 8480 811
rect 8768 798 9058 818
rect 9266 799 9300 818
rect 8581 776 8596 797
rect 8768 794 8984 798
rect 8615 776 8984 794
rect 8525 775 8984 776
rect 8507 741 8984 775
rect 9285 756 9300 799
rect 8508 740 8984 741
rect 6297 692 8480 700
rect 6297 685 8083 692
rect 6297 674 8093 685
rect 144 646 8093 674
rect 8139 682 8480 692
rect 8525 682 8984 740
rect 8139 646 8984 682
rect 9064 646 9098 680
rect 9152 646 9186 680
rect 9266 646 9300 756
rect 9319 765 9354 799
rect 9319 646 9353 765
rect 11110 733 11145 767
rect 9465 697 9523 703
rect 9465 684 9477 697
rect 9465 682 9511 684
rect 9465 680 9523 682
rect 9461 663 9527 680
rect 9635 674 9669 703
rect 10021 674 10232 729
rect 11111 714 11145 733
rect 9465 657 9523 663
rect 9437 646 9551 654
rect 9635 646 9978 674
rect 144 623 9978 646
rect 144 614 644 623
rect 650 619 9978 623
rect 652 614 9978 619
rect 144 612 9978 614
rect 144 604 8099 612
rect 158 600 8099 604
rect 158 599 6975 600
rect 6990 599 7003 600
rect 158 584 7003 599
rect 7015 594 8099 600
rect 8139 594 9316 612
rect 9319 594 9353 612
rect 9395 600 9567 612
rect 7015 585 9353 594
rect 158 582 4384 584
rect 4395 583 7003 584
rect 7006 583 9353 585
rect 158 580 4394 582
rect 158 544 644 580
rect 649 576 710 580
rect 728 576 820 580
rect 649 570 820 576
rect 847 570 4394 580
rect 649 558 813 570
rect 847 558 2358 570
rect 650 554 798 558
rect 813 554 820 558
rect 852 554 2358 558
rect 2362 566 4394 570
rect 4395 578 9353 583
rect 4395 570 8119 578
rect 4395 566 5887 570
rect 2362 554 5887 566
rect 5891 568 8119 570
rect 8139 568 9353 578
rect 9433 574 9467 600
rect 9521 579 9555 600
rect 9491 574 9555 579
rect 9615 584 9621 600
rect 9635 584 9978 612
rect 650 544 813 554
rect 847 553 2351 554
rect 847 548 2353 553
rect 2362 548 5880 554
rect 5891 548 9353 568
rect 9491 566 9538 574
rect 826 544 2335 548
rect 158 542 786 544
rect 158 526 698 542
rect 726 537 786 542
rect 710 526 786 537
rect 792 537 813 544
rect 814 537 2335 544
rect 792 530 2335 537
rect 798 526 2335 530
rect 2342 544 5860 548
rect 5871 544 9353 548
rect 2342 542 5880 544
rect 5891 542 9353 544
rect 2342 534 9353 542
rect 2342 528 8077 534
rect 8086 528 8099 534
rect 8126 528 9353 534
rect 9423 532 9433 566
rect 9473 558 9541 566
rect 9441 538 9479 548
rect 9491 538 9541 558
rect 2342 526 9353 528
rect 158 510 9353 526
rect 158 500 5850 510
rect 5871 500 8132 510
rect 158 460 8132 500
rect 158 450 2220 460
rect 2228 450 2308 460
rect 158 448 2308 450
rect 2310 448 2319 460
rect 2328 449 5855 460
rect 5869 449 8132 460
rect 158 424 2320 448
rect 2328 439 8132 449
rect 2328 424 7927 439
rect 158 415 7927 424
rect 158 402 5855 415
rect 5869 409 7927 415
rect 7931 436 7989 439
rect 7998 436 8132 439
rect 7931 413 8132 436
rect 7943 411 8065 413
rect 8067 411 8132 413
rect 7943 409 8132 411
rect 8139 454 9353 510
rect 9441 530 9541 538
rect 9552 530 9567 545
rect 9421 498 9436 507
rect 9441 498 9567 530
rect 9421 494 9479 498
rect 9521 496 9567 498
rect 9487 494 9503 496
rect 9421 492 9503 494
rect 9421 473 9479 492
rect 9515 483 9567 496
rect 9574 483 9590 514
rect 9515 480 9590 483
rect 9515 473 9567 480
rect 9379 464 9567 473
rect 9379 454 9519 464
rect 8139 449 9519 454
rect 9521 449 9567 464
rect 9615 449 9978 584
rect 8139 432 9978 449
rect 10021 659 10092 674
rect 10941 665 10999 671
rect 10021 432 10091 659
rect 10941 631 10953 665
rect 10941 625 10999 631
rect 10203 591 10261 597
rect 10203 557 10215 591
rect 10373 568 10407 586
rect 10795 568 10829 586
rect 10203 551 10261 557
rect 10373 532 10443 568
rect 8139 415 10091 432
rect 8139 409 9390 415
rect 158 390 5861 402
rect 158 375 2320 390
rect 158 362 2312 375
rect 2340 374 5861 390
rect 158 348 644 362
rect 650 358 2312 362
rect 650 353 2310 358
rect 650 350 698 353
rect 704 350 2310 353
rect 650 348 704 350
rect 710 349 2310 350
rect 158 343 704 348
rect 712 347 2310 349
rect 2342 347 5861 374
rect 710 343 2310 347
rect 2338 343 5861 347
rect 5869 381 9390 409
rect 9407 405 9472 415
rect 9478 405 9547 415
rect 9407 387 9547 405
rect 9407 381 9548 387
rect 5869 347 9548 381
rect 5869 343 9390 347
rect 158 330 2298 343
rect 158 323 2322 330
rect 158 300 1382 323
rect 158 291 874 300
rect 875 291 1382 300
rect 158 243 1382 291
rect 1397 311 2322 323
rect 2326 323 5867 343
rect 2326 320 5125 323
rect 2326 311 5129 320
rect 1397 310 5129 311
rect 1397 306 1528 310
rect 1536 308 1584 310
rect 1604 308 5129 310
rect 5133 308 5867 323
rect 1536 306 2322 308
rect 1397 296 2322 306
rect 2326 296 5867 308
rect 5871 323 9390 343
rect 5871 318 8769 323
rect 8877 322 9390 323
rect 9407 322 9548 347
rect 5871 305 8763 318
rect 8877 313 9548 322
rect 5871 303 8800 305
rect 8877 303 9478 313
rect 5871 296 9478 303
rect 1397 288 9478 296
rect 1397 287 9353 288
rect 9379 287 9478 288
rect 9480 287 9548 313
rect 9581 353 9601 415
rect 9615 396 10091 415
rect 10390 498 10461 532
rect 9615 362 10103 396
rect 10159 362 10199 396
rect 9615 353 10091 362
rect 9581 287 10091 353
rect 10165 330 10199 362
rect 10177 300 10199 321
rect 1397 286 10091 287
rect 1397 268 9338 286
rect 1385 258 9338 268
rect 9379 266 10091 286
rect 1385 253 9333 258
rect 1385 243 2234 253
rect 158 226 2234 243
rect 2238 238 2322 253
rect 2326 238 5804 253
rect 2250 226 2322 238
rect 2338 226 5804 238
rect 158 209 5804 226
rect 5805 220 9333 253
rect 5805 209 9319 220
rect 9322 214 9333 220
rect 158 186 9319 209
rect 9326 186 9333 214
rect 158 184 9333 186
rect 158 170 9319 184
rect 158 167 9316 170
rect 9326 167 9333 184
rect 9367 253 10091 266
rect 9367 243 9514 253
rect 9367 214 9387 243
rect 9393 224 9514 243
rect 9393 214 9425 224
rect 9367 184 9425 214
rect 9367 176 9413 184
rect 9417 176 9419 184
rect 9427 176 9514 224
rect 9581 235 10091 253
rect 10165 299 10199 300
rect 10165 289 10223 299
rect 10165 283 10261 289
rect 10390 286 10460 498
rect 10572 430 10630 436
rect 10572 396 10584 430
rect 10572 390 10630 396
rect 10390 284 10493 286
rect 10165 250 10223 283
rect 10107 235 10151 250
rect 10165 239 10276 250
rect 10373 243 10493 284
rect 10165 235 10265 239
rect 9581 216 10373 235
rect 10390 216 10493 243
rect 9581 181 10141 216
rect 10165 181 10199 216
rect 9581 176 10119 181
rect 9367 167 10119 176
rect 158 164 10119 167
rect 158 160 6277 164
rect 158 130 630 160
rect 638 152 789 160
rect 798 159 2170 160
rect 814 152 2170 159
rect 650 148 798 152
rect 828 150 2170 152
rect 826 148 2170 150
rect 652 144 798 148
rect 663 142 798 144
rect 828 142 2170 148
rect 664 138 742 142
rect 167 116 630 130
rect 678 125 742 138
rect 678 120 692 125
rect 694 120 742 125
rect 708 116 742 120
rect 744 116 752 142
rect 764 138 786 142
rect 814 116 828 140
rect 840 138 2170 142
rect 2174 143 2234 160
rect 2250 159 2334 160
rect 2338 159 2436 160
rect 2174 141 2204 143
rect 2186 138 2204 141
rect 2216 141 2234 143
rect 2262 141 2334 159
rect 2216 138 2246 141
rect 2276 138 2334 141
rect 2342 138 2436 159
rect 852 122 2436 138
rect 835 120 2436 122
rect 835 116 2344 120
rect 2388 116 2436 120
rect 2441 157 6277 160
rect 2441 144 2603 157
rect 2631 144 2725 157
rect 2441 136 2496 144
rect 2505 141 2603 144
rect 2643 141 2725 144
rect 2748 141 2755 144
rect 2757 142 6277 157
rect 2757 141 6037 142
rect 2505 140 6037 141
rect 6048 141 6139 142
rect 6156 141 6277 142
rect 6295 162 9728 164
rect 6295 157 9316 162
rect 9326 157 9333 162
rect 9367 157 9728 162
rect 6295 142 9728 157
rect 6295 141 8407 142
rect 2441 116 2489 136
rect 167 92 2489 116
rect 144 84 2489 92
rect 2505 129 2539 140
rect 2543 136 6025 140
rect 2505 120 2538 129
rect 2543 122 5925 136
rect 5926 122 6018 136
rect 6048 131 8407 141
rect 8426 137 8428 142
rect 8430 131 9413 142
rect 6048 122 9413 131
rect 9427 122 9461 142
rect 9467 122 9514 142
rect 9581 122 9668 142
rect 2543 120 9668 122
rect 9670 120 9728 142
rect 2505 114 9668 120
rect 9682 114 9728 120
rect 2505 107 9728 114
rect 2505 84 2539 107
rect 2543 88 2703 107
rect 2555 84 2703 88
rect 2757 88 6144 107
rect 2757 84 6032 88
rect 144 82 6032 84
rect 144 14 630 82
rect 743 77 806 82
rect 834 80 835 82
rect 852 80 2278 82
rect 650 73 684 77
rect 738 74 806 77
rect 819 74 2278 80
rect 738 73 2278 74
rect 638 64 2278 73
rect 2344 74 6032 82
rect 6052 84 6144 88
rect 6156 84 6277 107
rect 6295 105 9728 107
rect 6295 97 9722 105
rect 6295 84 8407 97
rect 8420 93 9722 97
rect 8420 91 9728 93
rect 8408 85 8428 91
rect 6052 78 8407 84
rect 6052 74 6086 78
rect 6092 74 8407 78
rect 2344 72 8407 74
rect 638 63 698 64
rect 726 63 2278 64
rect 638 56 710 63
rect 727 62 2191 63
rect 727 56 2170 62
rect 2214 60 2228 63
rect 2230 60 2278 63
rect 2244 56 2278 60
rect 2348 68 8407 72
rect 2348 56 8306 68
rect 8310 56 8407 68
rect 638 52 8306 56
rect 8320 52 8354 56
rect 8360 53 8407 56
rect 8426 81 8428 85
rect 8430 88 9728 91
rect 8430 81 9514 88
rect 8426 74 9514 81
rect 9581 80 9728 88
rect 9736 80 9883 164
rect 9884 161 9904 164
rect 9929 161 9942 164
rect 9560 74 9573 80
rect 8426 62 9577 74
rect 8360 52 8422 53
rect 638 29 8296 52
rect 8320 29 8422 52
rect 8426 46 9464 62
rect 9467 54 9577 62
rect 8426 29 9461 46
rect 638 18 9461 29
rect 638 14 8279 18
rect 144 3 8279 14
rect 8296 6 9461 18
rect 8289 3 9461 6
rect 144 -5 9461 3
rect 144 -6 8296 -5
rect 144 -9 828 -6
rect 835 -9 8296 -6
rect 144 -20 8296 -9
rect 8300 -16 8422 -5
rect 144 -45 710 -20
rect 738 -45 798 -20
rect 835 -28 8296 -20
rect 8320 -28 8354 -16
rect 835 -31 8354 -28
rect 8364 -31 8422 -16
rect 8474 -30 8510 -5
rect 8515 -16 8561 -5
rect 8565 -16 9461 -5
rect 835 -34 8422 -31
rect 835 -35 8330 -34
rect 835 -37 6970 -35
rect 144 -58 711 -45
rect 738 -58 799 -45
rect 835 -48 6964 -37
rect 852 -52 6964 -48
rect 826 -54 6964 -52
rect 852 -56 6964 -54
rect 814 -58 6964 -56
rect 7015 -50 8330 -35
rect 8339 -37 8422 -34
rect 8470 -37 8510 -30
rect 8339 -46 8407 -37
rect 8354 -50 8407 -46
rect 7015 -58 8407 -50
rect 144 -68 732 -58
rect 738 -65 8407 -58
rect 738 -66 8322 -65
rect 8342 -66 8407 -65
rect 8474 -66 8508 -37
rect 8527 -66 8561 -16
rect 8567 -66 9461 -16
rect 738 -68 9461 -66
rect 144 -82 9461 -68
rect 144 -94 9413 -82
rect 144 -101 8723 -94
rect 144 -112 7891 -101
rect 7893 -102 8080 -101
rect 8092 -102 8723 -101
rect 7893 -112 8723 -102
rect 144 -113 8723 -112
rect 144 -150 7891 -113
rect 144 -172 6993 -150
rect 80 -176 6993 -172
rect 144 -177 6993 -176
rect 6998 -161 7891 -150
rect 7893 -118 8723 -113
rect 8742 -98 9413 -94
rect 7893 -137 8705 -118
rect 8742 -122 9403 -98
rect 9427 -117 9461 -82
rect 9467 -34 9514 54
rect 9527 40 9539 54
rect 9547 40 9577 54
rect 9560 34 9573 40
rect 9581 -7 9668 80
rect 9682 78 9883 80
rect 9670 46 9883 78
rect 9559 -22 9668 -7
rect 9467 -56 9517 -34
rect 9537 -56 9538 -28
rect 9559 -56 9578 -22
rect 9581 -48 9668 -22
rect 9682 34 9830 46
rect 9836 34 9883 46
rect 9682 -48 9883 34
rect 9581 -56 9883 -48
rect 9467 -92 9883 -56
rect 9467 -94 9830 -92
rect 9467 -98 9628 -94
rect 8742 -128 8776 -122
rect 8789 -128 9403 -122
rect 8742 -137 8757 -128
rect 8773 -137 8776 -128
rect 8796 -137 9403 -128
rect 9423 -135 9461 -117
rect 9471 -107 9624 -98
rect 9634 -107 9670 -94
rect 9471 -118 9670 -107
rect 9471 -125 9672 -118
rect 9678 -125 9830 -94
rect 9471 -134 9830 -125
rect 9836 -134 9883 -92
rect 9950 108 10018 164
rect 9950 91 9984 108
rect 9997 91 10018 108
rect 10054 154 10119 164
rect 10153 164 10311 181
rect 10153 158 10315 164
rect 10054 147 10122 154
rect 10153 147 10326 158
rect 10389 147 10493 216
rect 10572 230 10630 236
rect 10572 196 10584 230
rect 10572 190 10630 196
rect 10054 91 10141 147
rect 10165 91 10199 147
rect 10253 114 10265 147
rect 10253 108 10311 114
rect 10390 109 10493 147
rect 10390 94 10622 109
rect 10759 94 10829 568
rect 10941 177 10999 183
rect 10941 143 10953 177
rect 10941 137 10999 143
rect 10390 91 10493 94
rect 9950 55 10493 91
rect 10759 58 10812 94
rect 11130 58 11145 714
rect 9950 21 10534 55
rect 10795 41 10991 56
rect 11056 41 11145 58
rect 11164 680 11199 714
rect 11164 41 11198 680
rect 11310 612 11368 618
rect 11310 578 11322 612
rect 11310 572 11368 578
rect 11480 409 11514 427
rect 13324 415 13359 449
rect 11480 373 11550 409
rect 13325 396 13359 415
rect 11497 339 11568 373
rect 11848 339 11883 373
rect 11310 124 11368 130
rect 11310 90 11322 124
rect 11310 84 11368 90
rect 9950 2 10493 21
rect 10759 5 10973 38
rect 11164 7 11179 41
rect 11497 40 11567 339
rect 11849 320 11883 339
rect 11679 271 11737 277
rect 11679 237 11691 271
rect 11679 231 11737 237
rect 11679 71 11737 77
rect 11679 42 11691 71
rect 11679 40 11713 42
rect 11497 37 11713 40
rect 11497 31 11737 37
rect 11260 4 11418 22
rect 11206 3 11418 4
rect 9950 -7 10534 2
rect 9950 -13 10602 -7
rect 9950 -91 10493 -13
rect 10500 -32 10602 -13
rect 10687 -32 10903 2
rect 11144 -12 11418 3
rect 11421 -12 11452 4
rect 11144 -15 11364 -12
rect 11074 -30 11364 -15
rect 10534 -84 10545 -73
rect 10553 -84 10568 -32
rect 10534 -91 10568 -84
rect 10587 -84 10621 -32
rect 10688 -51 10722 -32
rect 10707 -53 10722 -51
rect 10587 -91 10602 -84
rect 10698 -91 10722 -53
rect 10741 -60 10903 -51
rect 10741 -85 10971 -60
rect 11074 -82 11359 -30
rect 11445 -64 11460 -60
rect 10741 -91 10775 -85
rect 9950 -125 10826 -91
rect 9950 -134 10510 -125
rect 10514 -134 10580 -125
rect 7893 -151 9403 -137
rect 9411 -141 9469 -135
rect 9471 -141 9719 -134
rect 9724 -135 9898 -134
rect 9724 -141 9794 -135
rect 9796 -141 9898 -135
rect 9407 -146 9724 -141
rect 9407 -150 9720 -146
rect 9736 -147 9898 -141
rect 9738 -150 9772 -147
rect 9407 -151 9776 -150
rect 7893 -156 9776 -151
rect 9792 -156 9898 -147
rect 7893 -158 9898 -156
rect 7897 -161 9898 -158
rect 6998 -164 9898 -161
rect 9928 -153 10510 -134
rect 10518 -140 10576 -134
rect 10534 -153 10568 -140
rect 9928 -164 10568 -153
rect 6998 -171 9830 -164
rect 6998 -177 8705 -171
rect 8780 -172 8798 -171
rect 8808 -172 8826 -171
rect 144 -200 8705 -177
rect 8773 -178 8839 -172
rect 8860 -175 9830 -171
rect 80 -204 8705 -200
rect 144 -211 8705 -204
rect 8780 -208 8798 -178
rect 8808 -208 8826 -178
rect 8860 -180 9668 -175
rect 8860 -181 9684 -180
rect 8860 -185 9668 -181
rect 8860 -190 9403 -185
rect 9427 -187 9523 -185
rect 9565 -187 9668 -185
rect 9427 -190 9495 -187
rect 8860 -191 9495 -190
rect 9581 -191 9668 -187
rect 8860 -208 9427 -191
rect 9432 -208 9461 -191
rect 9466 -208 9514 -191
rect 9581 -208 9624 -191
rect 9634 -204 9668 -191
rect 9685 -204 9719 -175
rect 9738 -204 9772 -175
rect 9782 -188 9830 -175
rect 9840 -170 9884 -164
rect 9782 -194 9838 -188
rect 9840 -194 9886 -170
rect 9950 -194 10568 -164
rect 10587 -168 10621 -125
rect 10688 -150 10722 -125
rect 10729 -134 10775 -125
rect 10733 -140 10791 -134
rect 9776 -204 10568 -194
rect 9634 -208 10568 -204
rect 144 -216 6993 -211
rect 6998 -216 8705 -211
rect 8860 -209 10568 -208
rect 8860 -212 9615 -209
rect 144 -220 8705 -216
rect 144 -222 2305 -220
rect 2326 -222 8705 -220
rect 144 -224 8705 -222
rect 144 -229 2308 -224
rect 144 -232 2298 -229
rect 2326 -230 8705 -224
rect 8756 -215 9615 -212
rect 8756 -222 9461 -215
rect 9466 -222 9514 -215
rect 9581 -222 9615 -215
rect 9634 -211 10568 -209
rect 10574 -211 10621 -168
rect 10667 -168 10722 -150
rect 10741 -153 10775 -140
rect 10792 -153 10826 -125
rect 10903 -137 10914 -126
rect 10922 -137 10937 -85
rect 10903 -144 10937 -137
rect 10956 -137 10990 -85
rect 10956 -144 10971 -137
rect 11074 -144 11352 -82
rect 11433 -103 11460 -64
rect 11497 -92 11711 31
rect 11868 -48 11883 320
rect 11794 -65 11883 -48
rect 11902 286 11937 320
rect 12217 286 12252 320
rect 12640 303 12675 321
rect 11902 -65 11936 286
rect 12218 267 12252 286
rect 12604 288 12675 303
rect 12048 218 12106 224
rect 12048 184 12060 218
rect 12048 178 12106 184
rect 12048 18 12106 24
rect 12048 -16 12060 18
rect 12048 -22 12106 -16
rect 11902 -66 11917 -65
rect 12237 -66 12252 267
rect 12271 233 12306 267
rect 12271 -66 12305 233
rect 12417 165 12475 171
rect 12417 131 12429 165
rect 12417 125 12475 131
rect 12417 -35 12475 -29
rect 12417 -64 12429 -35
rect 12417 -66 12451 -64
rect 11471 -98 11711 -92
rect 10667 -184 10735 -168
rect 10741 -172 10826 -153
rect 10845 -148 11352 -144
rect 11426 -121 11460 -103
rect 11467 -101 11711 -98
rect 11812 -69 12451 -66
rect 11812 -75 12475 -69
rect 11467 -121 11498 -101
rect 11812 -106 12449 -75
rect 11515 -121 11517 -110
rect 11645 -121 11675 -108
rect 11866 -121 12449 -106
rect 10845 -161 11359 -148
rect 11426 -154 12449 -121
rect 12604 -154 12674 288
rect 12786 220 12844 226
rect 12786 186 12798 220
rect 12786 180 12844 186
rect 12786 -88 12844 -82
rect 12786 -122 12798 -88
rect 12786 -128 12844 -122
rect 11426 -157 12097 -154
rect 11405 -161 12097 -157
rect 10741 -184 10835 -172
rect 10688 -187 10835 -184
rect 10845 -178 12097 -161
rect 12183 -170 12198 -166
rect 10845 -187 10879 -178
rect 10883 -187 10949 -178
rect 8756 -224 9519 -222
rect 8756 -230 9423 -224
rect 144 -236 2296 -232
rect 144 -244 644 -236
rect 650 -238 2296 -236
rect 650 -244 2298 -238
rect 144 -245 2298 -244
rect 144 -247 2211 -245
rect 144 -256 698 -247
rect 710 -251 2211 -247
rect 713 -252 2211 -251
rect 725 -253 732 -252
rect 710 -256 732 -253
rect 738 -256 786 -252
rect 790 -256 2211 -252
rect 2214 -256 2298 -245
rect 2326 -243 9423 -230
rect 9457 -243 9519 -224
rect 9527 -234 9561 -222
rect 9576 -234 9624 -222
rect 9547 -243 9624 -234
rect 9634 -238 10621 -211
rect 10622 -193 10680 -187
rect 10622 -227 10646 -193
rect 10654 -227 10684 -193
rect 10688 -211 10775 -187
rect 10789 -206 10879 -187
rect 10887 -193 10945 -187
rect 10903 -206 10937 -193
rect 10622 -233 10680 -227
rect 9634 -243 9734 -238
rect 9738 -243 9772 -238
rect 9782 -240 9949 -238
rect 9950 -240 10621 -238
rect 9782 -243 9914 -240
rect 2326 -244 9914 -243
rect 9928 -244 9934 -240
rect 2326 -252 8705 -244
rect 8727 -249 9914 -244
rect 9967 -249 10621 -240
rect 2326 -256 6993 -252
rect 144 -264 6993 -256
rect 6997 -256 8705 -252
rect 8722 -256 9914 -249
rect 6997 -264 9914 -256
rect 144 -268 9914 -264
rect 144 -290 6981 -268
rect 144 -300 1368 -290
rect 144 -344 630 -300
rect 638 -326 690 -300
rect 704 -326 1368 -300
rect 638 -344 684 -326
rect 710 -328 1368 -326
rect 710 -344 772 -328
rect 786 -342 1368 -328
rect 798 -344 1368 -342
rect 144 -357 1368 -344
rect 1383 -347 6981 -290
rect 6985 -271 9914 -268
rect 9950 -250 10621 -249
rect 9950 -266 10520 -250
rect 10524 -262 10621 -250
rect 6985 -277 9888 -271
rect 6985 -280 9500 -277
rect 9511 -280 9888 -277
rect 6985 -290 9888 -280
rect 6985 -333 8705 -290
rect 8722 -297 9386 -290
rect 9407 -291 9447 -290
rect 8756 -302 9386 -297
rect 9396 -302 9447 -291
rect 8756 -303 9407 -302
rect 8722 -330 9407 -303
rect 9413 -330 9447 -302
rect 8722 -331 9447 -330
rect 8756 -333 9447 -331
rect 6985 -334 9447 -333
rect 6989 -336 9447 -334
rect 9466 -336 9500 -290
rect 9581 -302 9615 -290
rect 9634 -296 9668 -290
rect 9685 -293 9702 -290
rect 9704 -293 9719 -290
rect 9685 -296 9719 -293
rect 9738 -296 9869 -290
rect 9880 -296 9883 -290
rect 9896 -296 9902 -287
rect 9916 -296 9946 -287
rect 9950 -296 10510 -266
rect 10534 -294 10568 -262
rect 10574 -265 10621 -262
rect 10688 -250 10777 -211
rect 10789 -250 10937 -206
rect 10956 -221 10990 -178
rect 11057 -188 12097 -178
rect 11057 -203 12090 -188
rect 10688 -262 10778 -250
rect 10789 -262 10829 -250
rect 10688 -265 10735 -262
rect 10574 -266 10630 -265
rect 10578 -290 10630 -266
rect 10672 -266 10735 -265
rect 10741 -266 10775 -262
rect 10789 -266 10826 -262
rect 10672 -290 10775 -266
rect 9634 -302 9685 -296
rect 9581 -320 9685 -302
rect 9580 -324 9702 -320
rect 9581 -330 9714 -324
rect 9719 -330 10510 -296
rect 10518 -300 10576 -294
rect 10578 -300 10621 -290
rect 9581 -336 9719 -330
rect 6989 -340 9719 -336
rect 1383 -353 2238 -347
rect 1383 -354 1443 -353
rect 1448 -354 2238 -353
rect 2240 -354 2250 -347
rect 2262 -354 2320 -347
rect 2328 -353 6981 -347
rect 2328 -354 5790 -353
rect 5807 -354 6981 -353
rect 6998 -346 9719 -340
rect 6998 -353 9513 -346
rect 6998 -354 9142 -353
rect 1383 -356 2238 -354
rect 1383 -357 1526 -356
rect 1531 -357 2238 -356
rect 2250 -357 9142 -354
rect 144 -368 2238 -357
rect 2262 -362 5790 -357
rect 2262 -368 2320 -362
rect 2328 -368 5790 -362
rect 144 -402 5790 -368
rect 5824 -367 9142 -357
rect 5824 -368 8722 -367
rect 5824 -402 6981 -368
rect 6998 -402 8722 -368
rect 144 -425 8722 -402
rect 144 -434 2106 -425
rect 2119 -434 8722 -425
rect 144 -436 8722 -434
rect 144 -460 630 -436
rect 638 -437 775 -436
rect 798 -437 806 -436
rect 638 -438 814 -437
rect 851 -438 2106 -436
rect 638 -442 2106 -438
rect 638 -448 2066 -442
rect 650 -452 664 -448
rect 676 -450 738 -448
rect 764 -450 772 -448
rect 676 -452 772 -450
rect 158 -470 630 -460
rect 678 -468 744 -452
rect 167 -506 174 -470
rect 193 -506 201 -470
rect 158 -508 201 -506
rect 216 -508 630 -470
rect 638 -475 744 -468
rect 638 -478 696 -475
rect 678 -482 696 -478
rect 704 -480 744 -475
rect 759 -478 770 -464
rect 814 -468 2066 -448
rect 2072 -468 2106 -442
rect 2174 -459 2232 -436
rect 2262 -442 2320 -436
rect 2240 -459 2320 -442
rect 2328 -450 2422 -436
rect 2436 -450 2494 -436
rect 2505 -449 2589 -436
rect 2624 -438 2677 -436
rect 2590 -449 2595 -442
rect 2618 -449 2623 -442
rect 2643 -449 2677 -438
rect 2757 -448 6176 -436
rect 2757 -449 5905 -448
rect 2505 -450 5905 -449
rect 2186 -463 2234 -459
rect 2187 -468 2206 -463
rect 2215 -468 2234 -463
rect 2240 -468 2265 -459
rect 2274 -463 2308 -459
rect 2328 -468 2382 -450
rect 814 -470 2382 -468
rect 2388 -470 2422 -450
rect 2441 -454 2482 -450
rect 2441 -456 2475 -454
rect 814 -480 2422 -470
rect 2436 -470 2475 -456
rect 2436 -480 2489 -470
rect 2494 -472 2524 -450
rect 2533 -468 5905 -450
rect 5924 -468 5984 -448
rect 6038 -468 6139 -448
rect 2533 -472 6139 -468
rect 2494 -478 6139 -472
rect 726 -482 738 -480
rect 678 -484 742 -482
rect 678 -486 788 -484
rect 678 -488 778 -486
rect 814 -488 2342 -480
rect 2354 -487 2382 -480
rect 678 -489 788 -488
rect 678 -492 804 -489
rect 678 -496 699 -492
rect 726 -496 804 -492
rect 685 -500 699 -496
rect 144 -586 630 -508
rect 646 -527 699 -500
rect 738 -505 804 -496
rect 638 -536 699 -527
rect 704 -518 804 -505
rect 635 -544 696 -536
rect 704 -539 806 -518
rect 821 -520 846 -488
rect 852 -495 2342 -488
rect 852 -512 1747 -495
rect 1762 -512 1814 -495
rect 713 -544 806 -539
rect 852 -544 1737 -512
rect 1768 -520 1814 -512
rect 1756 -521 1814 -520
rect 1844 -503 1902 -495
rect 1903 -503 1911 -495
rect 1918 -503 1948 -495
rect 1951 -497 2342 -495
rect 1951 -501 2305 -497
rect 1844 -520 1853 -503
rect 1856 -520 1902 -503
rect 1918 -520 1945 -503
rect 1951 -509 2316 -501
rect 2348 -509 2382 -487
rect 1951 -512 2382 -509
rect 1951 -518 2066 -512
rect 1951 -520 2013 -518
rect 1844 -521 1902 -520
rect 1756 -544 1823 -521
rect 1853 -544 1911 -521
rect 1962 -544 2013 -520
rect 2019 -536 2066 -518
rect 2072 -536 2106 -512
rect 2111 -527 2280 -512
rect 2111 -528 2191 -527
rect 2019 -544 2106 -536
rect 2125 -538 2191 -528
rect 2214 -540 2280 -527
rect 2348 -516 2382 -512
rect 2388 -508 2422 -480
rect 2441 -498 2475 -480
rect 2505 -483 6139 -478
rect 2441 -508 2456 -498
rect 2471 -501 2475 -498
rect 2464 -508 2475 -501
rect 2388 -512 2482 -508
rect 2543 -512 2601 -483
rect 2660 -498 2683 -496
rect 2649 -505 2689 -498
rect 2631 -512 2689 -505
rect 2757 -502 6139 -483
rect 2388 -516 2422 -512
rect 2441 -516 2475 -512
rect 2555 -516 2619 -512
rect 2757 -516 5984 -502
rect 2348 -528 6034 -516
rect 2348 -544 5896 -528
rect 635 -550 5896 -544
rect 635 -578 5884 -550
rect 635 -586 684 -578
rect 727 -586 784 -578
rect 852 -586 2328 -578
rect 144 -590 2328 -586
rect 2332 -590 5884 -578
rect 144 -608 2129 -590
rect 2130 -596 2180 -590
rect 2234 -596 2291 -590
rect 2130 -608 2192 -596
rect 2222 -608 2291 -596
rect 2305 -600 5884 -590
rect 2305 -606 4753 -600
rect 4757 -606 4899 -600
rect 2305 -608 3160 -606
rect 144 -613 2328 -608
rect 144 -625 570 -613
rect 596 -618 2328 -613
rect 596 -620 2331 -618
rect 607 -623 625 -620
rect 144 -635 604 -625
rect 607 -630 628 -623
rect 635 -630 696 -620
rect 607 -635 696 -630
rect 719 -632 732 -620
rect 738 -632 799 -620
rect 821 -624 2331 -620
rect 2332 -624 3160 -608
rect 144 -645 696 -635
rect 704 -636 719 -632
rect 732 -636 784 -632
rect 799 -636 806 -632
rect 144 -657 622 -645
rect 628 -657 696 -645
rect 144 -661 696 -657
rect 719 -654 732 -636
rect 738 -654 799 -636
rect 719 -658 799 -654
rect 821 -642 3160 -624
rect 821 -658 2075 -642
rect 711 -660 2075 -658
rect 144 -663 705 -661
rect 711 -662 793 -660
rect 799 -662 2075 -660
rect 2081 -646 2297 -642
rect 2305 -646 3160 -642
rect 2081 -652 3160 -646
rect 2081 -658 2192 -652
rect 2203 -658 3160 -652
rect 3179 -612 4753 -606
rect 4771 -612 4899 -606
rect 3179 -622 4899 -612
rect 3179 -625 4784 -622
rect 3179 -652 3213 -625
rect 3281 -627 3331 -625
rect 3369 -627 3427 -625
rect 3286 -631 3327 -627
rect 3339 -631 3358 -627
rect 3374 -631 3415 -627
rect 3286 -649 3405 -631
rect 3303 -652 3405 -649
rect 3179 -658 3405 -652
rect 3472 -658 4784 -625
rect 4821 -627 4899 -622
rect 4909 -604 4914 -600
rect 4921 -604 5884 -600
rect 4909 -615 5884 -604
rect 4833 -631 4879 -627
rect 4854 -632 4879 -631
rect 4796 -636 4826 -632
rect 4796 -640 4833 -636
rect 4854 -640 4868 -632
rect 4909 -634 4979 -615
rect 4787 -655 4845 -640
rect 2081 -662 2129 -658
rect 711 -663 845 -662
rect 144 -674 845 -663
rect 144 -680 705 -674
rect 711 -680 845 -674
rect 144 -691 845 -680
rect 144 -710 570 -691
rect 582 -698 845 -691
rect 852 -670 2066 -662
rect 2081 -668 2100 -662
rect 2112 -668 2129 -662
rect 2134 -668 2141 -658
rect 2146 -668 3156 -658
rect 2083 -670 3156 -668
rect 852 -674 3156 -670
rect 852 -698 2066 -674
rect 2095 -678 2100 -674
rect 2112 -678 2129 -674
rect 2134 -692 3156 -674
rect 3179 -665 3449 -658
rect 3179 -674 3274 -665
rect 3275 -669 3418 -665
rect 3286 -674 3418 -669
rect 3461 -674 4784 -658
rect 4793 -665 4845 -655
rect 4793 -668 4839 -665
rect 4854 -668 4867 -640
rect 4877 -665 4917 -650
rect 4877 -668 4927 -665
rect 4793 -674 4927 -668
rect 4931 -674 4979 -634
rect 3179 -676 4979 -674
rect 4984 -634 5884 -615
rect 5892 -634 5896 -550
rect 5924 -550 6034 -528
rect 5924 -597 5984 -550
rect 6038 -578 6086 -502
rect 6091 -578 6139 -502
rect 6142 -578 6176 -448
rect 6193 -520 6253 -436
rect 6293 -453 6598 -436
rect 6610 -443 6981 -436
rect 6293 -470 6353 -453
rect 6407 -466 6455 -453
rect 6397 -470 6455 -466
rect 6293 -520 6343 -470
rect 6353 -478 6355 -470
rect 6385 -478 6455 -470
rect 6397 -487 6455 -478
rect 6407 -499 6455 -487
rect 6511 -499 6545 -453
rect 6564 -476 6599 -453
rect 6633 -462 6981 -443
rect 6998 -462 8722 -436
rect 6633 -465 6964 -462
rect 6622 -476 6964 -465
rect 6564 -499 6598 -476
rect 6646 -499 6964 -476
rect 6979 -496 8722 -462
rect 6407 -506 6964 -499
rect 6407 -520 6968 -506
rect 6193 -550 6265 -520
rect 6293 -550 6355 -520
rect 6385 -529 6968 -520
rect 6385 -542 6950 -529
rect 6385 -550 6860 -542
rect 6193 -578 6253 -550
rect 6293 -556 6343 -550
rect 6287 -557 6343 -556
rect 6038 -580 6253 -578
rect 6028 -597 6253 -580
rect 6263 -584 6343 -557
rect 5924 -609 5972 -597
rect 6016 -604 6253 -597
rect 6259 -604 6343 -584
rect 5924 -634 5974 -609
rect 6016 -614 6343 -604
rect 6012 -618 6343 -614
rect 5995 -628 6343 -618
rect 4984 -646 5974 -634
rect 5984 -642 5995 -628
rect 5978 -646 5995 -642
rect 6012 -638 6343 -628
rect 6012 -646 6253 -638
rect 4984 -658 6139 -646
rect 6142 -658 6253 -646
rect 6259 -654 6279 -638
rect 3179 -680 4958 -676
rect 3179 -686 4979 -680
rect 2112 -698 2129 -694
rect 582 -701 622 -698
rect 144 -801 596 -710
rect 616 -713 622 -701
rect 638 -707 2066 -698
rect 2109 -700 2129 -698
rect 644 -710 650 -707
rect 671 -710 2066 -707
rect 644 -740 2066 -710
rect 2092 -736 2097 -720
rect 644 -741 2070 -740
rect 650 -766 2070 -741
rect 2088 -766 2097 -736
rect 2112 -735 2129 -700
rect 2134 -698 3173 -692
rect 2134 -717 2192 -698
rect 2200 -717 3173 -698
rect 2134 -724 3173 -717
rect 2140 -731 3173 -724
rect 2140 -734 2691 -731
rect 2112 -739 2131 -735
rect 2140 -739 2280 -734
rect 2126 -740 2131 -739
rect 2115 -751 2139 -740
rect 2144 -746 2280 -739
rect 2284 -746 2324 -734
rect 2144 -751 2324 -746
rect 650 -770 2097 -766
rect 644 -784 2097 -770
rect 2126 -754 2324 -751
rect 644 -788 2116 -784
rect 2126 -785 2185 -754
rect 2190 -770 2270 -754
rect 2278 -770 2324 -754
rect 2190 -785 2324 -770
rect 2126 -788 2324 -785
rect 644 -794 2270 -788
rect 644 -798 696 -794
rect 699 -798 2270 -794
rect 2278 -792 2324 -788
rect 2328 -792 2691 -734
rect 2717 -754 3173 -731
rect 3179 -754 3213 -686
rect 2717 -767 3213 -754
rect 3228 -692 4979 -686
rect 3228 -722 3267 -692
rect 3321 -699 3409 -692
rect 3321 -715 3374 -699
rect 3228 -767 3274 -722
rect 3328 -744 3362 -715
rect 3416 -733 3450 -692
rect 3281 -760 3286 -744
rect 3316 -760 3362 -744
rect 3281 -767 3362 -760
rect 3421 -767 3450 -733
rect 3455 -699 4979 -692
rect 3455 -701 4927 -699
rect 3455 -707 4346 -701
rect 4350 -702 4384 -701
rect 4348 -703 4384 -702
rect 4388 -703 4394 -701
rect 4400 -703 4544 -701
rect 3455 -767 4336 -707
rect 2717 -776 3227 -767
rect 2717 -784 3173 -776
rect 2717 -792 2932 -784
rect 2278 -798 2703 -792
rect 144 -812 602 -801
rect 607 -804 625 -798
rect 635 -804 2703 -798
rect 638 -810 2703 -804
rect 144 -856 618 -812
rect 638 -816 2284 -810
rect 2294 -812 2324 -810
rect 2290 -814 2324 -812
rect 2328 -814 2703 -810
rect 2717 -804 2804 -792
rect 638 -820 2260 -816
rect 2328 -820 2691 -814
rect 638 -822 2261 -820
rect 638 -834 696 -822
rect 639 -844 696 -834
rect 699 -835 2261 -822
rect 699 -842 2197 -835
rect 650 -846 684 -844
rect 703 -846 784 -842
rect 799 -846 806 -842
rect 814 -844 2197 -842
rect 826 -846 2197 -844
rect 2202 -846 2261 -835
rect 2291 -836 2691 -820
rect 2717 -836 2810 -804
rect 2291 -846 2810 -836
rect 650 -856 2810 -846
rect 144 -870 2810 -856
rect 2872 -848 2932 -792
rect 2942 -800 2952 -784
rect 2960 -800 3008 -784
rect 3096 -792 3173 -784
rect 2978 -845 3008 -800
rect 2872 -860 2910 -848
rect 2963 -860 3018 -845
rect 2910 -870 3002 -860
rect 144 -873 2691 -870
rect 181 -878 2691 -873
rect 181 -879 638 -878
rect 181 -880 649 -879
rect 679 -880 2691 -878
rect 195 -886 649 -880
rect 195 -890 667 -886
rect 685 -890 2691 -880
rect 216 -893 238 -890
rect 201 -908 238 -893
rect 621 -896 639 -890
rect 649 -896 667 -890
rect 737 -904 767 -890
rect 784 -904 814 -890
rect 446 -944 458 -913
rect 474 -944 486 -913
rect 869 -926 1324 -890
rect 635 -950 1324 -926
rect 1394 -908 1429 -890
rect 1432 -894 1455 -890
rect 1475 -906 1482 -890
rect 1486 -902 1516 -890
rect 1551 -892 2080 -890
rect 2088 -892 2185 -890
rect 1551 -896 2070 -892
rect 1590 -903 2070 -896
rect 2092 -903 2172 -892
rect 2180 -896 2185 -892
rect 2174 -903 2191 -896
rect 2202 -903 2260 -890
rect 2328 -903 2691 -890
rect 1590 -904 2691 -903
rect 1394 -910 1445 -908
rect 1475 -910 1482 -908
rect 1517 -910 1524 -906
rect 1551 -908 1583 -906
rect 1590 -908 2051 -904
rect 1394 -925 1429 -910
rect 1551 -922 2051 -908
rect 1517 -924 2051 -922
rect 1394 -932 1428 -925
rect 1533 -928 2051 -924
rect 1398 -935 1428 -932
rect 1517 -932 2051 -928
rect 2092 -908 2691 -904
rect 2092 -919 2328 -908
rect 2092 -924 2139 -919
rect 1398 -950 1429 -935
rect 144 -990 216 -960
rect 430 -961 464 -958
rect 635 -962 1341 -950
rect 1371 -958 1429 -950
rect 1517 -936 2047 -932
rect 1517 -956 1583 -936
rect 1590 -937 2047 -936
rect 1370 -962 1528 -958
rect 1590 -962 2046 -937
rect 2092 -944 2097 -924
rect 2109 -926 2139 -924
rect 2172 -926 2219 -919
rect 2248 -924 2328 -919
rect 2261 -926 2291 -924
rect 2098 -928 2150 -926
rect 2161 -928 2219 -926
rect 2098 -932 2242 -928
rect 2250 -932 2302 -926
rect 2098 -937 2302 -932
rect 2362 -937 2691 -908
rect 2172 -944 2181 -937
rect 2092 -947 2194 -944
rect 2236 -947 2282 -944
rect 2172 -950 2181 -947
rect 2328 -950 2339 -939
rect 2351 -950 2362 -939
rect 178 -996 216 -990
rect 272 -992 326 -966
rect 356 -992 414 -966
rect 556 -992 625 -966
rect 635 -979 2046 -962
rect 2170 -966 2204 -958
rect 2328 -966 2362 -950
rect 2365 -956 2691 -937
rect 2717 -881 2804 -870
rect 2890 -873 3002 -870
rect 2878 -881 3002 -873
rect 2717 -882 3002 -881
rect 2717 -956 2804 -882
rect 2878 -886 2898 -882
rect 2960 -891 3002 -882
rect 3086 -870 3097 -859
rect 3103 -870 3173 -792
rect 3179 -801 3227 -776
rect 3228 -770 4336 -767
rect 4348 -714 4544 -703
rect 4579 -713 4927 -701
rect 4939 -713 4979 -699
rect 4579 -714 4979 -713
rect 4348 -718 4979 -714
rect 4984 -684 6253 -658
rect 6287 -682 6343 -638
rect 4984 -692 5122 -684
rect 5140 -685 5198 -684
rect 5214 -685 6253 -684
rect 4348 -754 4790 -718
rect 4793 -730 4833 -718
rect 4799 -734 4833 -730
rect 4348 -758 4636 -754
rect 4348 -769 4534 -758
rect 4541 -769 4636 -758
rect 4348 -770 4636 -769
rect 3228 -779 4342 -770
rect 4348 -777 4440 -770
rect 4476 -777 4513 -770
rect 4348 -779 4416 -777
rect 3228 -780 4416 -779
rect 3228 -781 4303 -780
rect 4320 -781 4336 -780
rect 4602 -781 4636 -770
rect 3228 -801 4636 -781
rect 4683 -756 4790 -754
rect 4683 -767 4753 -756
rect 4765 -758 4790 -756
rect 4765 -767 4784 -758
rect 4838 -767 4884 -718
rect 4984 -727 5032 -692
rect 5035 -727 5122 -692
rect 5152 -727 5156 -685
rect 5164 -700 5198 -685
rect 5231 -694 6253 -685
rect 5231 -697 5880 -694
rect 5882 -697 5892 -694
rect 5231 -698 5892 -697
rect 5231 -700 5880 -698
rect 5882 -700 5892 -698
rect 5914 -700 6253 -694
rect 5164 -706 5186 -700
rect 5168 -718 5186 -706
rect 5231 -712 6253 -700
rect 5246 -718 6253 -712
rect 5253 -724 6253 -718
rect 5253 -727 6086 -724
rect 4984 -733 6086 -727
rect 4951 -734 6086 -733
rect 6091 -734 6139 -724
rect 6142 -734 6253 -724
rect 6293 -724 6343 -682
rect 6407 -552 6860 -550
rect 6880 -552 6950 -542
rect 6407 -588 6950 -552
rect 7015 -563 8722 -496
rect 7015 -565 8007 -563
rect 7015 -588 7229 -565
rect 6407 -595 7229 -588
rect 7280 -595 8007 -565
rect 8018 -595 8722 -563
rect 6407 -598 7083 -595
rect 7144 -598 7179 -595
rect 6407 -627 7097 -598
rect 7144 -627 7193 -598
rect 6407 -632 7193 -627
rect 6407 -681 6950 -632
rect 7145 -641 7193 -632
rect 7384 -601 8722 -595
rect 8728 -373 9142 -367
rect 9212 -364 9246 -353
rect 9265 -364 9323 -353
rect 9212 -369 9323 -364
rect 9212 -373 9327 -369
rect 9369 -370 9513 -353
rect 9546 -354 9719 -346
rect 9738 -354 9772 -330
rect 9776 -340 9869 -330
rect 9780 -346 9869 -340
rect 9782 -354 9816 -346
rect 9835 -354 9869 -346
rect 9950 -349 10510 -330
rect 10514 -334 10621 -300
rect 10518 -340 10576 -334
rect 10534 -349 10568 -340
rect 9546 -364 9880 -354
rect 9546 -370 9869 -364
rect 9373 -373 9407 -370
rect 9413 -373 9447 -370
rect 9466 -373 9501 -370
rect 9505 -373 9513 -370
rect 9530 -373 9567 -370
rect 8728 -388 9567 -373
rect 9568 -387 9869 -370
rect 9950 -383 10568 -349
rect 10578 -348 10580 -334
rect 10584 -348 10621 -334
rect 10688 -294 10775 -290
rect 10688 -300 10791 -294
rect 10792 -300 10826 -266
rect 10688 -348 10724 -300
rect 10729 -334 10775 -300
rect 10779 -334 10826 -300
rect 10843 -264 10937 -250
rect 10943 -264 10990 -221
rect 11036 -237 12090 -203
rect 12171 -209 12198 -170
rect 12235 -198 12449 -154
rect 12532 -171 12674 -154
rect 12604 -172 12657 -171
rect 12209 -204 12449 -198
rect 10843 -303 10990 -264
rect 10991 -246 11049 -240
rect 10991 -280 11015 -246
rect 11023 -280 11053 -246
rect 11057 -254 12090 -237
rect 12164 -227 12198 -209
rect 12205 -207 12449 -204
rect 12550 -194 12657 -172
rect 12205 -227 12236 -207
rect 12550 -208 12725 -194
rect 12736 -208 12894 -190
rect 12975 -208 12990 322
rect 13009 -208 13043 376
rect 13155 347 13213 353
rect 13155 313 13167 347
rect 13155 307 13213 313
rect 13187 -135 13342 -64
rect 13155 -141 13342 -135
rect 13155 -170 13167 -141
rect 13187 -170 13342 -141
rect 13155 -174 13342 -170
rect 13151 -175 13342 -174
rect 13155 -181 13342 -175
rect 12550 -212 12894 -208
rect 12253 -227 12255 -216
rect 12383 -227 12413 -214
rect 12620 -224 12894 -212
rect 12897 -224 12928 -208
rect 13043 -209 13151 -208
rect 12620 -227 12840 -224
rect 12164 -242 12840 -227
rect 13043 -242 13117 -209
rect 11057 -267 12097 -254
rect 12164 -263 12835 -242
rect 12143 -267 12835 -263
rect 10991 -286 11049 -280
rect 10843 -315 10889 -303
rect 10893 -315 10990 -303
rect 10733 -340 10791 -334
rect 10578 -350 10621 -348
rect 10578 -355 10622 -350
rect 10684 -355 10724 -348
rect 9568 -388 9880 -387
rect 8728 -601 9564 -388
rect 7384 -618 8007 -601
rect 7384 -630 7616 -618
rect 7384 -641 7615 -630
rect 7164 -681 7193 -641
rect 7198 -681 7247 -641
rect 7294 -648 7615 -641
rect 7294 -651 7452 -648
rect 7294 -675 7466 -651
rect 7308 -680 7466 -675
rect 6407 -692 7187 -681
rect 6407 -704 6968 -692
rect 6971 -694 7187 -692
rect 7248 -685 7514 -680
rect 6971 -704 7193 -694
rect 6407 -715 7193 -704
rect 7248 -715 7283 -685
rect 6407 -724 6967 -715
rect 6971 -724 7035 -715
rect 6293 -725 6355 -724
rect 4951 -741 5860 -734
rect 5864 -736 6181 -734
rect 6193 -735 6253 -734
rect 5864 -740 5993 -736
rect 5864 -741 5980 -740
rect 6016 -741 6035 -736
rect 6038 -741 6086 -736
rect 4951 -758 6086 -741
rect 4984 -761 6086 -758
rect 4964 -767 4985 -761
rect 4998 -767 5085 -761
rect 4683 -778 4902 -767
rect 4939 -770 5085 -767
rect 5094 -762 6086 -761
rect 6091 -762 6139 -736
rect 5094 -764 6139 -762
rect 4683 -780 4891 -778
rect 4683 -784 4826 -780
rect 4719 -790 4826 -784
rect 4861 -790 4891 -780
rect 4985 -790 5027 -770
rect 5094 -771 6086 -764
rect 5054 -774 5073 -771
rect 4719 -792 4837 -790
rect 4850 -792 4902 -790
rect 4985 -792 5038 -790
rect 5054 -792 5069 -774
rect 4719 -798 5069 -792
rect 3259 -806 3274 -801
rect 3240 -828 3274 -806
rect 3281 -810 3286 -801
rect 3316 -806 3347 -801
rect 3316 -828 3362 -806
rect 3240 -835 3287 -828
rect 3316 -832 3375 -828
rect 3240 -842 3274 -835
rect 3286 -844 3287 -835
rect 3328 -835 3375 -832
rect 3328 -842 3362 -835
rect 3374 -844 3375 -835
rect 2916 -907 2932 -901
rect 2912 -920 2928 -907
rect 2365 -966 2804 -956
rect 3086 -950 3173 -870
rect 3253 -854 3287 -844
rect 3341 -854 3375 -844
rect 3253 -880 3299 -854
rect 3341 -880 3387 -854
rect 3421 -858 3450 -801
rect 3455 -820 4636 -801
rect 4716 -801 5069 -798
rect 5088 -801 5122 -771
rect 5214 -772 6086 -771
rect 5237 -798 5255 -772
rect 5265 -798 5283 -772
rect 5299 -798 5306 -772
rect 5317 -775 6086 -772
rect 5317 -777 5980 -775
rect 6022 -777 6086 -775
rect 5317 -781 5944 -777
rect 5317 -791 5892 -781
rect 5922 -791 5944 -781
rect 5317 -798 5880 -791
rect 6038 -798 6086 -777
rect 4716 -808 4838 -801
rect 4861 -804 4868 -801
rect 5088 -804 5107 -801
rect 5111 -804 5122 -801
rect 5088 -820 5122 -804
rect 5317 -805 6086 -798
rect 5317 -809 5968 -805
rect 5317 -812 5860 -809
rect 5984 -812 6024 -809
rect 5317 -820 5880 -812
rect 3455 -846 4672 -820
rect 5088 -833 5880 -820
rect 5914 -824 6024 -812
rect 6038 -820 6086 -805
rect 6091 -794 6139 -764
rect 6142 -794 6176 -736
rect 6193 -737 6251 -735
rect 6295 -737 6355 -725
rect 6191 -747 6355 -737
rect 6191 -750 6232 -747
rect 6249 -750 6274 -747
rect 6191 -751 6274 -750
rect 6191 -764 6232 -751
rect 6249 -754 6274 -751
rect 6295 -754 6355 -747
rect 6385 -730 6967 -724
rect 6385 -743 6975 -730
rect 6985 -734 7051 -724
rect 6989 -740 7047 -734
rect 6385 -754 7001 -743
rect 6251 -760 6274 -754
rect 6297 -760 6343 -754
rect 6195 -794 6229 -764
rect 6249 -784 6343 -760
rect 6233 -792 6343 -784
rect 6407 -784 7001 -754
rect 7031 -762 7065 -758
rect 7019 -767 7077 -762
rect 7019 -768 7071 -767
rect 7019 -772 7048 -768
rect 7020 -774 7048 -772
rect 7075 -772 7077 -767
rect 7031 -784 7065 -774
rect 7075 -783 7091 -772
rect 7075 -784 7141 -783
rect 6233 -794 6385 -792
rect 6407 -794 6991 -784
rect 6091 -804 6173 -794
rect 6176 -804 6991 -794
rect 6091 -820 6991 -804
rect 5914 -833 6034 -824
rect 6038 -828 6991 -820
rect 6038 -830 6406 -828
rect 6407 -830 6991 -828
rect 6038 -833 6371 -830
rect 5088 -844 6371 -833
rect 6385 -834 6391 -830
rect 6421 -834 6991 -830
rect 6424 -839 6991 -834
rect 5088 -846 5099 -844
rect 5184 -846 6371 -844
rect 3374 -907 3387 -880
rect 3241 -922 3299 -907
rect 3329 -922 3387 -907
rect 3455 -862 6371 -846
rect 6407 -850 6991 -839
rect 7031 -817 7141 -784
rect 7031 -840 7091 -817
rect 7045 -850 7091 -840
rect 6407 -852 6968 -850
rect 6974 -852 6989 -850
rect 6407 -856 7059 -852
rect 7078 -855 7091 -850
rect 6407 -862 7071 -856
rect 3455 -877 6393 -862
rect 6407 -866 6991 -862
rect 3455 -880 6345 -877
rect 3455 -886 6139 -880
rect 6142 -886 6176 -880
rect 6195 -886 6323 -880
rect 6337 -886 6341 -880
rect 6353 -886 6359 -877
rect 6373 -886 6403 -877
rect 6407 -886 6967 -866
rect 7035 -867 7073 -862
rect 3455 -890 6144 -886
rect 3086 -966 3156 -950
rect 3297 -960 3331 -958
rect 635 -980 965 -979
rect 635 -992 879 -980
rect 891 -992 965 -980
rect 995 -992 1044 -979
rect 178 -1004 238 -996
rect 298 -1003 367 -992
rect 403 -995 567 -992
rect 403 -1003 480 -995
rect 298 -1015 322 -1003
rect 326 -1015 356 -1003
rect 414 -1011 480 -1003
rect 526 -1003 567 -995
rect 526 -1015 556 -1003
rect 625 -1014 925 -992
rect 954 -994 1006 -992
rect 1007 -994 1044 -992
rect 954 -996 1018 -994
rect 954 -1003 1045 -996
rect 158 -1024 174 -1018
rect 298 -1025 367 -1015
rect 515 -1025 567 -1015
rect 625 -1018 913 -1014
rect 625 -1025 879 -1018
rect 965 -1024 1045 -1003
rect 1007 -1025 1044 -1024
rect 298 -1026 1044 -1025
rect 635 -1048 879 -1026
rect 1098 -1038 1117 -979
rect 1126 -980 1253 -979
rect 1126 -992 1241 -980
rect 1274 -990 2046 -979
rect 1274 -992 1528 -990
rect 1607 -992 2046 -990
rect 2139 -971 2261 -966
rect 2139 -980 2154 -971
rect 2220 -980 2261 -971
rect 2139 -992 2181 -980
rect 2220 -992 2262 -980
rect 2291 -990 3156 -966
rect 2291 -992 2691 -990
rect 2734 -992 3156 -990
rect 3455 -966 3542 -890
rect 3659 -924 3662 -890
rect 3687 -896 3690 -890
rect 3698 -938 3708 -890
rect 3710 -928 3744 -890
rect 3610 -951 3708 -938
rect 3610 -966 3723 -951
rect 3455 -992 3682 -966
rect 1152 -996 2231 -992
rect 1152 -1009 1429 -996
rect 1445 -1009 1475 -996
rect 1607 -1003 2231 -996
rect 2250 -1003 2302 -992
rect 1607 -1006 2139 -1003
rect 1607 -1009 2069 -1006
rect 2154 -1009 2220 -1003
rect 2261 -1009 2291 -1003
rect 2328 -1009 2362 -992
rect 2365 -1009 2804 -992
rect 2832 -1009 3066 -992
rect 3074 -1009 3156 -992
rect 3270 -994 3542 -992
rect 3253 -1008 3542 -994
rect 3588 -997 3682 -992
rect 3588 -1004 3656 -997
rect 1152 -1026 3074 -1009
rect 1607 -1068 2046 -1026
rect 2328 -1068 2362 -1026
rect 2734 -1060 2945 -1026
rect 3090 -1032 3156 -1009
rect 3229 -1025 3542 -1008
rect 3616 -1013 3656 -1004
rect 3616 -1015 3648 -1013
rect 3650 -1015 3682 -1013
rect 3616 -1025 3682 -1015
rect 3229 -1026 3682 -1025
rect 3079 -1043 3156 -1032
rect 1607 -1079 2080 -1068
rect 2250 -1070 2475 -1068
rect 1607 -1085 2069 -1079
rect 188 -1128 238 -1090
rect 180 -1140 238 -1128
rect 268 -1140 326 -1090
rect 356 -1128 406 -1090
rect 2012 -1092 2069 -1085
rect 2111 -1091 2177 -1078
rect 2250 -1079 2291 -1070
rect 2261 -1091 2291 -1079
rect 2351 -1081 2362 -1070
rect 2734 -1079 2911 -1060
rect 3103 -1079 3156 -1043
rect 2111 -1092 2188 -1091
rect 1195 -1110 1210 -1095
rect 1414 -1110 1429 -1095
rect 2012 -1099 2188 -1092
rect 2250 -1099 2302 -1091
rect 3472 -1096 3542 -1026
rect 3650 -1047 3682 -1026
rect 2012 -1102 2362 -1099
rect 1195 -1128 1253 -1110
rect 356 -1140 414 -1128
rect 180 -1155 195 -1140
rect 180 -1164 196 -1160
rect 180 -1182 208 -1164
rect 280 -1182 314 -1140
rect 399 -1155 414 -1140
rect 399 -1182 414 -1167
rect 713 -1176 779 -1140
rect 1203 -1160 1253 -1128
rect 1283 -1160 1341 -1110
rect 1371 -1128 1429 -1110
rect 1371 -1160 1421 -1128
rect 1976 -1138 2195 -1106
rect 3472 -1132 3525 -1096
rect 3667 -1126 3719 -1115
rect 3678 -1138 3708 -1126
rect 3667 -1149 3719 -1138
rect 3843 -1149 3858 -890
rect 3877 -943 4672 -890
rect 4711 -904 4869 -890
rect 4930 -904 4965 -890
rect 4931 -923 4965 -904
rect 5041 -923 5054 -896
rect 5069 -923 5082 -896
rect 5317 -902 5388 -890
rect 5317 -923 5387 -902
rect 3877 -1149 3911 -943
rect 4210 -996 4672 -943
rect 4761 -972 4819 -966
rect 154 -1232 174 -1198
rect 180 -1212 238 -1182
rect 268 -1212 326 -1182
rect 356 -1212 414 -1182
rect 180 -1232 208 -1212
rect 180 -1263 189 -1232
rect 192 -1266 208 -1232
rect 280 -1224 314 -1212
rect 368 -1224 414 -1212
rect 446 -1224 636 -1191
rect 883 -1212 997 -1182
rect 3877 -1183 3892 -1149
rect 845 -1224 994 -1218
rect 1098 -1224 1117 -1212
rect 1341 -1220 1567 -1200
rect 1341 -1224 1677 -1220
rect 1729 -1224 1763 -1190
rect 1817 -1224 1851 -1190
rect 1905 -1224 1939 -1190
rect 1993 -1224 2027 -1190
rect 2081 -1224 2115 -1190
rect 2485 -1204 2519 -1190
rect 4210 -1202 4280 -996
rect 4392 -1119 4450 -1113
rect 4392 -1153 4404 -1119
rect 4392 -1159 4450 -1153
rect 4102 -1220 4128 -1202
rect 280 -1258 1034 -1224
rect 1055 -1252 1068 -1236
rect 1083 -1252 1101 -1240
rect 192 -1270 196 -1266
rect 280 -1274 314 -1258
rect 399 -1274 414 -1259
rect 216 -1293 238 -1274
rect 201 -1308 238 -1293
rect 268 -1304 326 -1274
rect 356 -1304 414 -1274
rect 468 -1274 483 -1259
rect 599 -1274 614 -1259
rect 468 -1303 526 -1274
rect 399 -1308 414 -1304
rect 476 -1304 526 -1303
rect 556 -1303 614 -1274
rect 667 -1280 717 -1258
rect 556 -1304 606 -1303
rect 476 -1306 606 -1304
rect 188 -1324 238 -1308
rect 268 -1324 326 -1308
rect 356 -1324 406 -1308
rect 446 -1344 458 -1306
rect 270 -1402 320 -1356
rect 262 -1406 320 -1402
rect 350 -1402 400 -1356
rect 440 -1398 458 -1344
rect 474 -1324 606 -1306
rect 659 -1304 717 -1280
rect 747 -1280 797 -1258
rect 867 -1274 882 -1259
rect 967 -1274 1001 -1258
rect 747 -1304 805 -1280
rect 867 -1304 925 -1274
rect 955 -1286 1013 -1274
rect 1055 -1286 1072 -1252
rect 1089 -1255 1101 -1252
rect 1098 -1286 1101 -1255
rect 1152 -1258 1158 -1224
rect 1242 -1235 1294 -1224
rect 1330 -1235 1341 -1224
rect 1253 -1242 1283 -1235
rect 1487 -1242 1555 -1224
rect 1567 -1242 1643 -1224
rect 1660 -1235 1712 -1224
rect 1176 -1254 1363 -1242
rect 1176 -1258 1367 -1254
rect 1487 -1258 1655 -1242
rect 1671 -1247 1701 -1235
rect 1660 -1258 1712 -1247
rect 1717 -1258 2127 -1224
rect 2250 -1235 2302 -1224
rect 2338 -1235 2390 -1224
rect 2458 -1235 2546 -1224
rect 2261 -1246 2291 -1235
rect 2349 -1246 2379 -1235
rect 1203 -1280 1253 -1258
rect 659 -1318 674 -1304
rect 790 -1318 805 -1304
rect 474 -1372 486 -1324
rect 526 -1329 556 -1324
rect 659 -1340 726 -1318
rect 747 -1340 805 -1318
rect 650 -1368 726 -1340
rect 659 -1370 726 -1368
rect 738 -1368 805 -1340
rect 667 -1372 717 -1370
rect 738 -1372 739 -1368
rect 747 -1370 805 -1368
rect 821 -1306 851 -1304
rect 867 -1306 882 -1304
rect 821 -1358 860 -1306
rect 867 -1318 888 -1306
rect 904 -1312 913 -1304
rect 904 -1318 919 -1312
rect 867 -1330 925 -1318
rect 955 -1330 1014 -1286
rect 1026 -1330 1035 -1306
rect 1043 -1330 1101 -1286
rect 1195 -1300 1253 -1280
rect 1283 -1280 1333 -1258
rect 1509 -1270 1524 -1258
rect 1684 -1270 1701 -1258
rect 1717 -1264 1775 -1258
rect 1805 -1264 1863 -1258
rect 1893 -1264 1951 -1258
rect 1981 -1264 2039 -1258
rect 2069 -1264 2127 -1258
rect 2203 -1258 2437 -1246
rect 2469 -1247 2535 -1235
rect 2469 -1254 2546 -1247
rect 4102 -1248 4142 -1230
rect 4210 -1236 4263 -1202
rect 4581 -1236 4596 -996
rect 4210 -1238 4596 -1236
rect 2494 -1258 2546 -1254
rect 4246 -1254 4596 -1238
rect 4615 -1254 4649 -996
rect 4761 -1006 4773 -972
rect 4761 -1012 4819 -1006
rect 4761 -1172 4819 -1166
rect 4761 -1206 4773 -1172
rect 4761 -1212 4819 -1206
rect 4246 -1255 4672 -1254
rect 2203 -1270 2218 -1258
rect 2422 -1270 2437 -1258
rect 1283 -1300 1341 -1280
rect 1195 -1306 1241 -1300
rect 1294 -1306 1324 -1300
rect 1110 -1318 1241 -1306
rect 1195 -1324 1241 -1318
rect 1261 -1324 1266 -1306
rect 1289 -1320 1324 -1306
rect 1326 -1315 1341 -1300
rect 1509 -1300 1567 -1270
rect 1597 -1280 1620 -1270
rect 1509 -1315 1524 -1300
rect 1597 -1320 1655 -1280
rect 1726 -1306 1743 -1270
rect 1756 -1300 1951 -1290
rect 2203 -1300 2261 -1270
rect 2291 -1300 2349 -1270
rect 2379 -1300 2437 -1270
rect 2535 -1300 2731 -1282
rect 4250 -1291 4672 -1255
rect 1726 -1312 1763 -1306
rect 1768 -1312 1791 -1306
rect 904 -1334 913 -1330
rect 967 -1334 1001 -1330
rect 1014 -1334 1089 -1330
rect 1173 -1334 1178 -1330
rect 1195 -1334 1266 -1324
rect 938 -1340 972 -1336
rect 984 -1340 997 -1334
rect 1014 -1340 1064 -1334
rect 926 -1358 978 -1340
rect 1014 -1356 1066 -1340
rect 1020 -1358 1066 -1356
rect 1132 -1346 1184 -1334
rect 1132 -1349 1162 -1346
rect 784 -1372 789 -1370
rect 468 -1398 486 -1372
rect 350 -1406 371 -1402
rect 262 -1412 277 -1406
rect 356 -1412 371 -1406
rect 262 -1421 308 -1412
rect 356 -1417 396 -1412
rect 274 -1446 308 -1421
rect 362 -1446 396 -1417
rect 474 -1446 508 -1412
rect 562 -1446 596 -1384
rect 644 -1398 690 -1372
rect 704 -1374 705 -1372
rect 726 -1384 762 -1372
rect 607 -1404 625 -1398
rect 635 -1404 653 -1398
rect 726 -1404 772 -1384
rect 792 -1398 793 -1370
rect 821 -1372 851 -1358
rect 926 -1368 972 -1358
rect 1026 -1368 1060 -1358
rect 814 -1384 866 -1372
rect 814 -1387 860 -1384
rect 820 -1398 851 -1387
rect 821 -1404 851 -1398
rect 857 -1404 872 -1389
rect 638 -1434 696 -1404
rect 726 -1434 784 -1404
rect 814 -1434 872 -1404
rect 926 -1392 955 -1368
rect 1057 -1392 1072 -1389
rect 926 -1430 984 -1392
rect 607 -1446 625 -1434
rect 181 -1457 257 -1446
rect 181 -1469 205 -1457
rect 216 -1469 246 -1457
rect 181 -1480 257 -1469
rect 262 -1480 408 -1446
rect 440 -1480 625 -1446
rect 440 -1580 458 -1486
rect 468 -1552 486 -1486
rect 562 -1540 596 -1480
rect 607 -1486 625 -1480
rect 635 -1446 684 -1434
rect 738 -1446 772 -1434
rect 826 -1446 872 -1434
rect 934 -1446 984 -1430
rect 1014 -1430 1072 -1392
rect 1132 -1392 1147 -1349
rect 1169 -1392 1184 -1346
rect 1195 -1358 1272 -1334
rect 1286 -1355 1341 -1320
rect 1509 -1332 1655 -1320
rect 1676 -1332 1806 -1312
rect 1676 -1334 1726 -1332
rect 1668 -1349 1726 -1334
rect 1195 -1370 1220 -1358
rect 1232 -1370 1272 -1358
rect 1283 -1370 1341 -1355
rect 1671 -1362 1726 -1349
rect 1729 -1334 1806 -1332
rect 1207 -1374 1212 -1370
rect 1232 -1392 1278 -1370
rect 1132 -1424 1190 -1392
rect 1220 -1424 1278 -1392
rect 1294 -1374 1329 -1370
rect 1294 -1404 1324 -1374
rect 1352 -1386 1363 -1370
rect 1352 -1389 1367 -1386
rect 1340 -1396 1367 -1389
rect 1340 -1404 1363 -1396
rect 1440 -1404 1474 -1386
rect 1559 -1404 1574 -1389
rect 1144 -1428 1178 -1424
rect 1232 -1428 1266 -1424
rect 1014 -1446 1064 -1430
rect 1253 -1434 1262 -1428
rect 1340 -1434 1398 -1404
rect 1428 -1434 1486 -1404
rect 1516 -1434 1574 -1404
rect 1668 -1392 1683 -1389
rect 1701 -1392 1720 -1362
rect 1668 -1424 1726 -1392
rect 1729 -1398 1748 -1334
rect 1756 -1362 1814 -1334
rect 1799 -1377 1814 -1362
rect 1966 -1370 1984 -1306
rect 1994 -1370 2012 -1306
rect 2203 -1315 2218 -1300
rect 2422 -1315 2437 -1300
rect 4286 -1307 4321 -1291
rect 4250 -1324 4321 -1307
rect 2203 -1336 2261 -1327
rect 2291 -1336 2349 -1327
rect 2379 -1336 2437 -1327
rect 2174 -1372 2349 -1362
rect 2379 -1372 2424 -1362
rect 2676 -1369 2704 -1368
rect 1982 -1377 1996 -1372
rect 3917 -1377 3952 -1343
rect 1799 -1392 1814 -1389
rect 1340 -1446 1386 -1434
rect 1440 -1446 1474 -1434
rect 1528 -1446 1574 -1434
rect 1676 -1446 1726 -1424
rect 1756 -1424 1814 -1392
rect 1982 -1404 1997 -1389
rect 2113 -1404 2128 -1389
rect 1756 -1446 1806 -1424
rect 1982 -1434 2040 -1404
rect 2070 -1434 2128 -1404
rect 1982 -1446 2028 -1434
rect 2082 -1446 2128 -1434
rect 2168 -1440 2577 -1418
rect 2168 -1446 2600 -1440
rect 635 -1480 872 -1446
rect 900 -1456 1098 -1446
rect 1106 -1450 1335 -1446
rect 904 -1468 1094 -1456
rect 1110 -1457 1335 -1450
rect 1110 -1462 1324 -1457
rect 984 -1469 1014 -1468
rect 1294 -1469 1324 -1462
rect 1340 -1464 1574 -1446
rect 1579 -1457 1631 -1446
rect 1642 -1450 1840 -1446
rect 1590 -1464 1620 -1457
rect 1646 -1462 1836 -1450
rect 1982 -1462 2128 -1446
rect 2133 -1452 2600 -1446
rect 2764 -1451 2822 -1448
rect 2133 -1457 2611 -1452
rect 1398 -1469 1428 -1464
rect 1486 -1469 1516 -1464
rect 1525 -1469 1674 -1464
rect 1726 -1466 1756 -1462
rect 2040 -1466 2070 -1462
rect 973 -1480 1025 -1469
rect 1283 -1480 1335 -1469
rect 1387 -1480 1439 -1469
rect 1475 -1480 1674 -1469
rect 635 -1486 684 -1480
rect 644 -1514 684 -1486
rect 665 -1518 684 -1514
rect 738 -1540 772 -1480
rect 1525 -1486 1674 -1480
rect 1714 -1486 1798 -1466
rect 1998 -1469 2082 -1466
rect 2144 -1469 2611 -1457
rect 2676 -1458 2822 -1451
rect 2852 -1458 2910 -1448
rect 3328 -1449 3362 -1392
rect 3548 -1401 3615 -1396
rect 3548 -1430 3662 -1401
rect 3667 -1407 3719 -1396
rect 3678 -1419 3708 -1407
rect 3667 -1430 3719 -1419
rect 1803 -1480 2082 -1469
rect 2133 -1480 2611 -1469
rect 1998 -1486 2082 -1480
rect 1784 -1490 1798 -1486
rect 1525 -1514 1646 -1492
rect 1714 -1514 1798 -1494
rect 1998 -1514 2082 -1494
rect 2290 -1504 2324 -1480
rect 2337 -1504 2600 -1480
rect 2942 -1500 3008 -1468
rect 3145 -1502 3162 -1474
rect 1756 -1518 1798 -1514
rect 2190 -1519 2600 -1504
rect 2810 -1513 2863 -1502
rect 2908 -1508 3162 -1502
rect 2810 -1519 2852 -1513
rect 2190 -1529 2405 -1519
rect 2454 -1529 2512 -1519
rect 2542 -1529 2668 -1519
rect 2190 -1530 2668 -1529
rect 2774 -1525 2852 -1519
rect 2908 -1516 3160 -1508
rect 2466 -1534 2500 -1530
rect 2554 -1534 2588 -1530
rect 2774 -1536 2863 -1525
rect 2908 -1534 3042 -1516
rect 3096 -1524 3160 -1516
rect 3110 -1525 3140 -1524
rect 3099 -1536 3140 -1525
rect 2774 -1555 2844 -1536
rect 2441 -1560 2622 -1555
rect 2441 -1568 2650 -1560
rect 2723 -1566 2844 -1555
rect 2441 -1589 2476 -1568
rect 2512 -1578 2542 -1568
rect 2501 -1582 2542 -1578
rect 2584 -1578 2650 -1568
rect 2734 -1578 2764 -1566
rect 2584 -1582 2661 -1578
rect 2501 -1589 2661 -1582
rect 2723 -1589 2764 -1578
rect 2072 -1619 2097 -1608
rect 2237 -1619 2289 -1608
rect 2321 -1619 2373 -1608
rect 2072 -1627 2086 -1619
rect 2248 -1624 2278 -1619
rect 1703 -1695 1902 -1661
rect 1907 -1672 2053 -1661
rect 1918 -1684 2053 -1672
rect 1907 -1690 2053 -1684
rect 1907 -1695 1959 -1690
rect 2038 -1695 2053 -1690
rect 1334 -1731 1386 -1714
rect 1427 -1721 1559 -1714
rect 1427 -1725 1479 -1721
rect 1579 -1725 1631 -1714
rect 929 -1746 1386 -1731
rect 1438 -1737 1468 -1725
rect 1590 -1737 1620 -1725
rect 1427 -1746 1479 -1737
rect 1579 -1743 1631 -1737
rect 1515 -1746 1631 -1743
rect 1668 -1746 1684 -1714
rect 929 -1748 1684 -1746
rect 440 -1798 458 -1774
rect 272 -1824 320 -1798
rect 350 -1824 462 -1798
rect 474 -1802 508 -1790
rect 468 -1818 508 -1802
rect 474 -1824 508 -1818
rect 562 -1820 596 -1790
rect 650 -1820 684 -1790
rect 692 -1798 738 -1790
rect 772 -1798 826 -1790
rect 692 -1814 826 -1798
rect 850 -1814 860 -1790
rect 692 -1820 860 -1814
rect 929 -1820 1368 -1748
rect 1392 -1800 1402 -1796
rect 1458 -1800 1514 -1782
rect 1568 -1800 1576 -1796
rect 562 -1824 872 -1820
rect 926 -1824 1368 -1820
rect 286 -1837 1368 -1824
rect 216 -1858 1368 -1837
rect 216 -1972 630 -1858
rect 650 -1874 664 -1858
rect 857 -1874 872 -1859
rect 638 -1904 696 -1874
rect 726 -1888 784 -1874
rect 814 -1875 872 -1874
rect 788 -1888 872 -1875
rect 720 -1904 872 -1888
rect 650 -1946 664 -1904
rect 720 -1906 738 -1904
rect 778 -1906 838 -1904
rect 720 -1916 784 -1906
rect 788 -1916 838 -1906
rect 720 -1922 838 -1916
rect 857 -1919 872 -1904
rect 738 -1946 838 -1922
rect 650 -1970 684 -1946
rect 650 -1972 664 -1970
rect 676 -1972 684 -1970
rect 738 -1956 860 -1946
rect 738 -1972 784 -1956
rect 792 -1962 800 -1956
rect 820 -1970 860 -1956
rect 820 -1972 838 -1970
rect 216 -1982 872 -1972
rect 912 -1982 1368 -1858
rect 1380 -1859 1422 -1800
rect 1458 -1812 1576 -1800
rect 1458 -1816 1602 -1812
rect 1476 -1850 1602 -1816
rect 1380 -1980 1426 -1859
rect 1476 -1866 1526 -1850
rect 1534 -1856 1538 -1850
rect 1480 -1869 1524 -1866
rect 1448 -1898 1460 -1893
rect 1438 -1909 1468 -1898
rect 1480 -1909 1525 -1869
rect 1562 -1884 1566 -1850
rect 1536 -1897 1548 -1893
rect 1448 -1968 1525 -1909
rect 1448 -1980 1482 -1968
rect 216 -2065 630 -1982
rect 181 -2233 185 -2065
rect 205 -2076 630 -2065
rect 214 -2088 630 -2076
rect 205 -2099 630 -2088
rect 193 -2100 630 -2099
rect 650 -1984 664 -1982
rect 676 -1984 690 -1982
rect 756 -1984 784 -1982
rect 820 -1984 866 -1982
rect 650 -2008 690 -1984
rect 710 -2003 718 -1999
rect 738 -2003 784 -1984
rect 798 -2003 806 -1999
rect 826 -2003 866 -1984
rect 650 -2100 664 -2008
rect 672 -2010 690 -2008
rect 672 -2044 684 -2010
rect 698 -2043 866 -2003
rect 872 -2043 1368 -1982
rect 1392 -1984 1402 -1980
rect 1414 -1984 1426 -1980
rect 672 -2072 690 -2044
rect 672 -2100 684 -2072
rect 698 -2100 1368 -2043
rect 1438 -2062 1482 -1980
rect 1502 -2008 1525 -1968
rect 1526 -1909 1556 -1897
rect 1568 -1909 1602 -1850
rect 1526 -1968 1602 -1909
rect 1526 -1991 1570 -1968
rect 1526 -2036 1582 -1991
rect 1536 -2044 1582 -2036
rect 1436 -2063 1482 -2062
rect 1502 -2063 1525 -2044
rect 1530 -2051 1582 -2044
rect 1530 -2063 1570 -2051
rect 1436 -2077 1494 -2063
rect 1502 -2072 1582 -2063
rect 1524 -2077 1582 -2072
rect 1494 -2078 1510 -2077
rect 193 -2140 876 -2100
rect 878 -2126 900 -2100
rect 912 -2113 1368 -2100
rect 1492 -2113 1526 -2092
rect 1650 -2094 1684 -1748
rect 1703 -1837 1737 -1695
rect 1768 -1837 1771 -1695
rect 1827 -1742 1856 -1729
rect 1895 -1732 1902 -1716
rect 1808 -1747 1856 -1742
rect 1887 -1747 1902 -1732
rect 1918 -1742 1948 -1705
rect 1962 -1742 1984 -1704
rect 1808 -1760 1902 -1747
rect 1907 -1760 1984 -1742
rect 1827 -1763 1902 -1760
rect 1918 -1763 1948 -1760
rect 1845 -1770 1948 -1763
rect 1990 -1770 2012 -1732
rect 1808 -1788 2012 -1770
rect 2019 -1748 2053 -1695
rect 2072 -1690 2087 -1627
rect 2130 -1631 2278 -1624
rect 2332 -1631 2362 -1619
rect 2119 -1642 2289 -1631
rect 2321 -1642 2373 -1631
rect 2172 -1654 2278 -1652
rect 2072 -1732 2106 -1690
rect 2019 -1782 2056 -1748
rect 2072 -1768 2090 -1732
rect 2095 -1768 2106 -1757
rect 1845 -1797 1948 -1788
rect 1783 -1818 1802 -1806
rect 1845 -1813 1902 -1797
rect 1918 -1813 1948 -1797
rect 1779 -1837 1802 -1818
rect 1856 -1828 1902 -1813
rect 1856 -1837 1893 -1828
rect 2019 -1837 2053 -1782
rect 2072 -1824 2106 -1768
rect 2190 -1778 2206 -1676
rect 2218 -1710 2276 -1704
rect 2407 -1710 2422 -1608
rect 2218 -1744 2234 -1710
rect 2218 -1750 2276 -1744
rect 2274 -1791 2308 -1786
rect 2174 -1820 2175 -1791
rect 2262 -1800 2320 -1791
rect 2406 -1800 2422 -1710
rect 2186 -1820 2220 -1803
rect 2262 -1806 2308 -1800
rect 2262 -1820 2264 -1806
rect 2274 -1820 2308 -1806
rect 2348 -1820 2374 -1800
rect 2388 -1820 2422 -1800
rect 2441 -1710 2475 -1589
rect 2541 -1612 2650 -1599
rect 2541 -1641 2542 -1612
rect 2584 -1626 2650 -1612
rect 2757 -1634 2764 -1589
rect 2774 -1604 2844 -1566
rect 2952 -1598 2990 -1592
rect 3126 -1598 3140 -1536
rect 3145 -1598 3160 -1524
rect 2952 -1604 3014 -1598
rect 3126 -1604 3160 -1598
rect 2774 -1634 3160 -1604
rect 2441 -1713 2456 -1710
rect 2441 -1796 2475 -1713
rect 2559 -1725 2570 -1676
rect 2583 -1698 2584 -1641
rect 2757 -1644 3160 -1634
rect 3179 -1524 3196 -1449
rect 3228 -1483 3462 -1449
rect 3516 -1458 3529 -1449
rect 3548 -1458 3582 -1430
rect 3516 -1479 3582 -1458
rect 3516 -1483 3529 -1479
rect 3548 -1480 3582 -1479
rect 3203 -1524 3213 -1483
rect 3179 -1625 3213 -1524
rect 3228 -1569 3267 -1483
rect 3495 -1491 3529 -1483
rect 3536 -1491 3582 -1480
rect 3495 -1495 3516 -1491
rect 3303 -1526 3328 -1517
rect 3299 -1530 3362 -1526
rect 3371 -1530 3409 -1513
rect 3299 -1564 3409 -1530
rect 3316 -1569 3409 -1564
rect 3416 -1569 3421 -1517
rect 3228 -1576 3286 -1569
rect 3316 -1576 3462 -1569
rect 3495 -1576 3529 -1495
rect 3240 -1580 3247 -1576
rect 3321 -1585 3374 -1576
rect 3382 -1585 3387 -1576
rect 3416 -1580 3421 -1576
rect 3321 -1601 3358 -1585
rect 3339 -1623 3358 -1601
rect 3374 -1623 3404 -1601
rect 3281 -1625 3331 -1623
rect 3369 -1625 3419 -1623
rect 3514 -1625 3529 -1576
rect 3548 -1625 3582 -1491
rect 3883 -1492 3898 -1396
rect 3628 -1608 3650 -1542
rect 3656 -1608 3708 -1570
rect 3727 -1608 3730 -1542
rect 3750 -1608 3784 -1574
rect 3864 -1608 3898 -1492
rect 3612 -1625 3616 -1608
rect 3628 -1625 3898 -1608
rect 3179 -1642 3898 -1625
rect 3179 -1644 3708 -1642
rect 3727 -1644 3730 -1642
rect 2587 -1657 2645 -1651
rect 2587 -1691 2599 -1657
rect 2757 -1668 3744 -1644
rect 2757 -1672 3766 -1668
rect 2587 -1697 2645 -1691
rect 2757 -1694 3778 -1672
rect 3781 -1694 3796 -1679
rect 2757 -1704 3796 -1694
rect 2757 -1710 3804 -1704
rect 2688 -1726 2711 -1710
rect 2643 -1738 2677 -1733
rect 2543 -1743 2601 -1738
rect 2567 -1750 2601 -1743
rect 2555 -1767 2601 -1750
rect 2643 -1754 2683 -1738
rect 2757 -1750 3796 -1710
rect 3804 -1738 3818 -1710
rect 2643 -1767 2677 -1754
rect 2757 -1767 3744 -1750
rect 3750 -1754 3798 -1750
rect 3754 -1760 3798 -1754
rect 2505 -1772 3744 -1767
rect 2441 -1820 2482 -1796
rect 2505 -1800 2529 -1772
rect 2543 -1778 3744 -1772
rect 3772 -1778 3798 -1760
rect 3864 -1778 3898 -1642
rect 3917 -1519 3951 -1377
rect 4250 -1519 4320 -1324
rect 4579 -1344 4672 -1291
rect 4950 -1308 4965 -923
rect 4984 -924 5387 -923
rect 4984 -957 5019 -924
rect 4984 -1308 5018 -957
rect 5041 -986 5054 -924
rect 5027 -1242 5054 -986
rect 5069 -1014 5082 -924
rect 5055 -1196 5082 -1014
rect 5102 -1196 5216 -1191
rect 5055 -1214 5255 -1196
rect 5130 -1224 5188 -1219
rect 4984 -1342 4999 -1308
rect 5041 -1342 5054 -1242
rect 5069 -1242 5269 -1224
rect 5069 -1342 5082 -1242
rect 5317 -1342 5387 -924
rect 5421 -920 5860 -890
rect 5421 -924 5870 -920
rect 5924 -924 5958 -920
rect 5421 -926 5860 -924
rect 6038 -926 6072 -890
rect 6091 -926 6126 -890
rect 6139 -914 6142 -890
rect 6176 -911 6967 -886
rect 6975 -890 7033 -884
rect 7035 -888 7081 -867
rect 7035 -890 7073 -888
rect 6176 -914 6403 -911
rect 6187 -920 6403 -914
rect 5421 -943 6080 -926
rect 5521 -1170 5527 -1023
rect 5549 -1198 5555 -1051
rect 5499 -1278 5557 -1272
rect 5499 -1296 5511 -1278
rect 5499 -1307 5545 -1296
rect 5688 -1307 5703 -943
rect 5722 -1307 5756 -943
rect 5826 -960 6080 -943
rect 6091 -960 6114 -926
rect 6139 -930 6195 -923
rect 6201 -925 6403 -920
rect 6407 -925 6967 -911
rect 6971 -924 7073 -890
rect 7145 -896 7193 -715
rect 7198 -896 7246 -715
rect 7145 -899 7246 -896
rect 6201 -930 6967 -925
rect 6139 -960 6176 -930
rect 5824 -1284 5882 -1236
rect 5912 -1278 5970 -1236
rect 5910 -1284 5970 -1278
rect 5836 -1288 5870 -1284
rect 5924 -1288 5958 -1284
rect 6038 -1290 6072 -960
rect 6091 -1290 6125 -960
rect 6195 -979 6229 -930
rect 6237 -936 6295 -930
rect 6407 -979 6967 -930
rect 6985 -934 7073 -924
rect 7135 -933 7246 -899
rect 7035 -938 7066 -934
rect 7145 -938 7193 -933
rect 7035 -945 7075 -938
rect 7141 -945 7193 -938
rect 7033 -950 7051 -945
rect 7091 -977 7131 -968
rect 6195 -992 6967 -979
rect 7079 -983 7137 -977
rect 7079 -992 7091 -983
rect 7111 -992 7141 -983
rect 7145 -992 7193 -945
rect 6195 -1013 7193 -992
rect 6407 -1017 7193 -1013
rect 6407 -1019 7141 -1017
rect 6407 -1099 6441 -1019
rect 6564 -1047 6579 -1019
rect 6793 -1031 7141 -1019
rect 7164 -1031 7193 -1017
rect 6793 -1036 7193 -1031
rect 6528 -1099 6731 -1049
rect 6793 -1062 6967 -1036
rect 6807 -1066 6967 -1062
rect 7198 -1045 7246 -933
rect 7249 -1045 7283 -715
rect 7531 -698 7615 -648
rect 7649 -631 8007 -618
rect 8018 -624 9564 -601
rect 8018 -629 8722 -624
rect 8728 -629 9564 -624
rect 8018 -631 9564 -629
rect 7649 -652 9564 -631
rect 7649 -665 8722 -652
rect 7649 -671 7967 -665
rect 7753 -688 7967 -671
rect 7531 -734 7688 -698
rect 7725 -701 7967 -688
rect 8018 -667 8722 -665
rect 8728 -667 9564 -652
rect 8018 -669 9564 -667
rect 8018 -685 8735 -669
rect 8018 -696 8705 -685
rect 8004 -701 8705 -696
rect 8709 -701 8728 -685
rect 8756 -701 9564 -669
rect 9568 -490 9668 -388
rect 9736 -389 9772 -388
rect 9782 -389 9816 -388
rect 9835 -389 9880 -388
rect 9950 -389 10510 -383
rect 9736 -399 10510 -389
rect 9736 -423 9882 -399
rect 9915 -402 10510 -399
rect 10587 -393 10621 -355
rect 10587 -402 10602 -393
rect 10618 -402 10621 -393
rect 10622 -393 10680 -387
rect 10622 -402 10634 -393
rect 10654 -402 10684 -393
rect 10688 -402 10722 -355
rect 10741 -402 10775 -340
rect 10792 -402 10826 -334
rect 10845 -319 10889 -315
rect 10845 -402 10879 -319
rect 10903 -347 10937 -315
rect 10943 -318 10990 -315
rect 11057 -294 12835 -267
rect 13043 -270 13117 -243
rect 12921 -276 12936 -272
rect 11057 -318 12828 -294
rect 10943 -319 10999 -318
rect 10947 -343 10999 -319
rect 11041 -343 12828 -318
rect 12909 -337 12936 -276
rect 13009 -276 13031 -272
rect 13043 -276 13185 -270
rect 13009 -277 13043 -276
rect 13105 -277 13185 -276
rect 12947 -310 13005 -304
rect 10887 -353 10945 -347
rect 10947 -353 10990 -343
rect 10883 -387 10990 -353
rect 10887 -393 10945 -387
rect 10903 -402 10937 -393
rect 9915 -419 10937 -402
rect 10947 -401 10949 -387
rect 10953 -401 10990 -387
rect 11057 -360 12828 -343
rect 11057 -373 12835 -360
rect 12907 -369 12936 -337
rect 12943 -344 12974 -310
rect 12993 -311 13009 -310
rect 13187 -313 13342 -181
rect 13344 -277 13359 396
rect 13378 362 13413 396
rect 13378 -277 13412 362
rect 13524 294 13582 300
rect 13524 260 13536 294
rect 13524 254 13582 260
rect 13694 91 13728 109
rect 13694 55 13764 91
rect 13711 21 13782 55
rect 14062 21 14097 55
rect 13524 -194 13582 -188
rect 13524 -228 13536 -194
rect 13524 -234 13582 -228
rect 13378 -300 13393 -277
rect 13378 -313 13463 -300
rect 13277 -318 13463 -313
rect 12947 -350 13005 -344
rect 13121 -354 13151 -320
rect 13378 -330 13463 -318
rect 13711 -330 13781 21
rect 14063 2 14097 21
rect 13893 -47 13951 -41
rect 13893 -81 13905 -47
rect 13893 -87 13951 -81
rect 13893 -247 13951 -241
rect 13893 -281 13905 -247
rect 13893 -287 13951 -281
rect 12881 -373 12936 -369
rect 13059 -373 13103 -354
rect 11057 -388 13103 -373
rect 13155 -388 13185 -354
rect 13344 -364 13409 -354
rect 13711 -366 13764 -330
rect 14082 -383 14097 2
rect 14116 -32 14151 2
rect 14431 -32 14466 0
rect 14116 -383 14150 -32
rect 14432 -51 14466 -32
rect 14262 -100 14320 -94
rect 14262 -134 14274 -100
rect 14262 -140 14320 -134
rect 14262 -300 14320 -294
rect 14262 -334 14274 -300
rect 14262 -340 14320 -334
rect 11057 -401 13093 -388
rect 10947 -403 10990 -401
rect 10947 -408 10991 -403
rect 11053 -408 13093 -401
rect 9915 -423 10088 -419
rect 9699 -440 9714 -425
rect 9672 -450 9714 -440
rect 9672 -456 9734 -450
rect 9736 -456 9816 -423
rect 9672 -490 9816 -456
rect 9568 -496 9734 -490
rect 9568 -537 9714 -496
rect 9736 -506 9738 -490
rect 9742 -506 9816 -490
rect 9736 -521 9816 -506
rect 9742 -524 9816 -521
rect 9732 -537 9736 -533
rect 9568 -672 9708 -537
rect 9568 -684 9620 -672
rect 9634 -684 9708 -672
rect 9726 -549 9736 -537
rect 9748 -549 9816 -524
rect 9580 -688 9615 -684
rect 7725 -722 7773 -701
rect 7739 -731 7773 -722
rect 7883 -711 7931 -701
rect 8004 -707 8709 -701
rect 8728 -707 9564 -701
rect 7723 -732 7789 -731
rect 7302 -745 7688 -734
rect 7302 -757 7337 -745
rect 7340 -751 7688 -745
rect 7883 -747 7967 -711
rect 8004 -737 8705 -707
rect 8709 -735 8728 -707
rect 8756 -722 9564 -707
rect 8756 -737 9114 -722
rect 7883 -751 7985 -747
rect 7340 -757 7985 -751
rect 7302 -768 7985 -757
rect 7302 -796 7336 -768
rect 7340 -777 7404 -768
rect 7354 -787 7420 -777
rect 7514 -787 7985 -768
rect 8004 -754 9114 -737
rect 9125 -754 9564 -722
rect 8004 -766 8336 -754
rect 8387 -760 9564 -754
rect 9581 -725 9615 -688
rect 9632 -705 9702 -684
rect 9726 -705 9816 -549
rect 9632 -717 9692 -705
rect 9726 -712 9736 -705
rect 9748 -706 9816 -705
rect 9835 -706 9880 -423
rect 9950 -509 10017 -423
rect 10082 -476 10083 -423
rect 10107 -442 10141 -419
rect 10151 -442 10185 -419
rect 10336 -436 10937 -419
rect 10107 -476 10137 -442
rect 10203 -476 10219 -442
rect 10336 -472 10510 -436
rect 10758 -441 10775 -436
rect 10440 -476 10510 -472
rect 10741 -455 10775 -441
rect 10792 -455 10826 -436
rect 10845 -455 10879 -436
rect 10956 -446 10990 -408
rect 10956 -455 10971 -446
rect 10987 -455 10990 -446
rect 10991 -446 11049 -440
rect 10991 -455 11003 -446
rect 11023 -455 11053 -446
rect 11057 -455 13093 -408
rect 10440 -481 10493 -476
rect 10151 -499 10185 -481
rect 10440 -495 10510 -481
rect 10741 -489 10792 -455
rect 10826 -470 13093 -455
rect 10837 -489 13093 -470
rect 10440 -499 10608 -495
rect 10151 -509 10608 -499
rect 9950 -512 10608 -509
rect 9950 -535 10221 -512
rect 10476 -529 10608 -512
rect 10707 -523 10792 -495
rect 10811 -529 10826 -489
rect 10845 -529 10879 -489
rect 10845 -534 10860 -529
rect 9950 -545 10239 -535
rect 10442 -544 10554 -535
rect 9950 -579 10221 -545
rect 10318 -569 10554 -544
rect 10318 -579 10353 -569
rect 9950 -691 10238 -579
rect 10319 -631 10353 -579
rect 10520 -588 10554 -569
rect 10845 -548 10879 -534
rect 11074 -548 13093 -489
rect 10845 -582 10977 -548
rect 11056 -582 13093 -548
rect 10539 -598 10554 -588
rect 10573 -598 10608 -588
rect 10811 -597 10923 -588
rect 10372 -603 10626 -598
rect 10372 -631 10446 -603
rect 10319 -632 10446 -631
rect 10468 -632 10626 -603
rect 10687 -622 10923 -597
rect 10687 -632 10722 -622
rect 10319 -637 10408 -632
rect 10346 -655 10362 -637
rect 9634 -725 9716 -717
rect 9581 -730 9716 -725
rect 9738 -730 9816 -706
rect 9581 -745 9816 -730
rect 9581 -747 9624 -745
rect 9634 -747 9816 -745
rect 9824 -747 9880 -706
rect 9949 -725 10238 -691
rect 9950 -737 10238 -725
rect 9967 -746 10238 -737
rect 9581 -751 9816 -747
rect 9581 -760 9756 -751
rect 9782 -760 9816 -751
rect 9835 -760 9880 -747
rect 8387 -766 9114 -760
rect 7358 -793 7416 -787
rect 7302 -815 7370 -796
rect 7400 -815 7434 -811
rect 7300 -837 7370 -815
rect 7388 -820 7446 -815
rect 7388 -821 7440 -820
rect 7388 -825 7417 -821
rect 7389 -827 7417 -825
rect 7444 -825 7446 -820
rect 7514 -821 7967 -787
rect 8004 -821 8353 -766
rect 7400 -837 7434 -827
rect 7444 -836 7460 -825
rect 7444 -837 7510 -836
rect 7300 -903 7360 -837
rect 7400 -870 7510 -837
rect 7400 -893 7460 -870
rect 7414 -903 7460 -893
rect 7300 -905 7337 -903
rect 7343 -905 7358 -903
rect 7302 -909 7428 -905
rect 7443 -908 7460 -903
rect 7471 -880 7482 -876
rect 7302 -915 7440 -909
rect 7302 -919 7360 -915
rect 7302 -1045 7336 -919
rect 7404 -920 7442 -915
rect 7443 -920 7456 -908
rect 7344 -943 7402 -937
rect 7404 -941 7456 -920
rect 7404 -943 7442 -941
rect 7340 -977 7442 -943
rect 7354 -987 7442 -977
rect 7404 -991 7435 -987
rect 7443 -991 7456 -941
rect 7404 -998 7456 -991
rect 7402 -1003 7420 -998
rect 7471 -1021 7484 -880
rect 7514 -952 7984 -821
rect 7504 -986 7984 -952
rect 7514 -991 7984 -986
rect 7510 -998 7984 -991
rect 7460 -1036 7500 -1021
rect 7480 -1045 7510 -1036
rect 7514 -1045 7984 -998
rect 6807 -1072 6950 -1066
rect 6846 -1077 6950 -1072
rect 7198 -1070 7227 -1045
rect 7294 -1070 7984 -1045
rect 7198 -1077 7212 -1070
rect 7294 -1077 7510 -1070
rect 6846 -1085 6967 -1077
rect 7198 -1078 7510 -1077
rect 7531 -1078 7984 -1070
rect 7198 -1079 7984 -1078
rect 7212 -1085 7984 -1079
rect 6846 -1089 7984 -1085
rect 6846 -1099 7283 -1089
rect 6407 -1135 6477 -1099
rect 6528 -1102 7283 -1099
rect 6933 -1119 7283 -1102
rect 7302 -1112 7984 -1089
rect 6407 -1169 6495 -1135
rect 6510 -1148 6776 -1135
rect 6933 -1148 7283 -1131
rect 6510 -1152 6846 -1148
rect 6897 -1152 7283 -1148
rect 6510 -1153 7283 -1152
rect 6510 -1165 7233 -1153
rect 6510 -1169 6967 -1165
rect 6407 -1201 6494 -1169
rect 6528 -1188 6967 -1169
rect 6528 -1193 6950 -1188
rect 6967 -1193 7179 -1188
rect 6528 -1199 7179 -1193
rect 6528 -1201 7001 -1199
rect 6407 -1222 7001 -1201
rect 7041 -1222 7179 -1199
rect 6407 -1237 6967 -1222
rect 7079 -1233 7137 -1227
rect 6193 -1271 6967 -1237
rect 5826 -1307 6080 -1290
rect 5034 -1360 5387 -1342
rect 5421 -1324 6080 -1307
rect 6091 -1324 6114 -1290
rect 6161 -1324 6176 -1290
rect 5421 -1360 5860 -1324
rect 5868 -1331 5926 -1325
rect 5034 -1361 5860 -1360
rect 5041 -1386 5054 -1361
rect 4432 -1392 4490 -1386
rect 4432 -1426 4444 -1392
rect 4432 -1432 4490 -1426
rect 4488 -1502 4522 -1468
rect 4602 -1502 4636 -1386
rect 5027 -1449 5054 -1386
rect 5069 -1414 5082 -1361
rect 5055 -1449 5082 -1414
rect 4719 -1466 4754 -1449
rect 3917 -1555 4320 -1519
rect 4350 -1536 4385 -1502
rect 4388 -1536 4636 -1502
rect 4683 -1483 4754 -1466
rect 4683 -1536 4753 -1483
rect 3917 -1725 4331 -1555
rect 3917 -1778 4339 -1725
rect 2543 -1800 4339 -1778
rect 2505 -1801 4339 -1800
rect 2505 -1812 2539 -1801
rect 2555 -1812 2589 -1801
rect 2072 -1837 2118 -1824
rect 2136 -1828 2171 -1820
rect 2174 -1828 2320 -1820
rect 2136 -1837 2320 -1828
rect 1703 -1854 2320 -1837
rect 2348 -1854 2486 -1820
rect 1703 -2094 2170 -1854
rect 2172 -1959 2220 -1854
rect 2262 -1888 2264 -1854
rect 2348 -1875 2374 -1854
rect 2348 -1888 2375 -1875
rect 2260 -1922 2274 -1888
rect 2305 -1906 2320 -1891
rect 2262 -1956 2264 -1922
rect 2278 -1956 2320 -1906
rect 2326 -1922 2340 -1916
rect 2322 -1956 2344 -1922
rect 2348 -1949 2378 -1888
rect 2388 -1949 2422 -1854
rect 2172 -1971 2206 -1959
rect 2262 -1971 2320 -1956
rect 2172 -2008 2218 -1971
rect 2274 -1975 2322 -1971
rect 2296 -1984 2322 -1975
rect 2348 -1980 2436 -1949
rect 2360 -1984 2422 -1980
rect 2250 -2003 2322 -1984
rect 2338 -2003 2372 -1999
rect 2172 -2012 2206 -2008
rect 2238 -2012 2298 -2003
rect 2332 -2008 2384 -2003
rect 2218 -2018 2298 -2012
rect 2338 -2018 2384 -2008
rect 2214 -2052 2298 -2018
rect 2214 -2058 2280 -2052
rect 2214 -2068 2234 -2058
rect 2238 -2068 2280 -2058
rect 2238 -2072 2264 -2068
rect 2190 -2078 2264 -2072
rect 2354 -2078 2384 -2018
rect 2190 -2086 2296 -2078
rect 1650 -2108 2170 -2094
rect 1650 -2113 1684 -2108
rect 1703 -2111 2170 -2108
rect 912 -2126 1694 -2113
rect 1731 -2120 2170 -2111
rect 2238 -2108 2296 -2086
rect 2326 -2108 2384 -2078
rect 2238 -2120 2253 -2108
rect 2338 -2120 2384 -2108
rect 2388 -2120 2422 -1984
rect 2441 -2067 2486 -1854
rect 2505 -1906 2589 -1812
rect 2505 -1931 2570 -1906
rect 2590 -1918 2595 -1801
rect 2613 -1812 2631 -1801
rect 2643 -1812 2677 -1801
rect 2757 -1804 4339 -1801
rect 4350 -1802 4384 -1536
rect 4388 -1653 4438 -1536
rect 4474 -1604 4488 -1570
rect 4519 -1588 4534 -1573
rect 4492 -1638 4534 -1588
rect 4542 -1638 4556 -1604
rect 4477 -1653 4534 -1638
rect 4400 -1657 4418 -1653
rect 4488 -1657 4536 -1653
rect 4510 -1666 4536 -1657
rect 4464 -1674 4536 -1666
rect 4444 -1685 4536 -1674
rect 4568 -1685 4586 -1681
rect 4444 -1700 4512 -1685
rect 4452 -1708 4512 -1700
rect 4568 -1708 4598 -1685
rect 4417 -1719 4598 -1708
rect 4428 -1731 4598 -1719
rect 4417 -1742 4598 -1731
rect 4602 -1740 4636 -1536
rect 4666 -1619 4753 -1536
rect 5027 -1566 5082 -1449
rect 5088 -1430 5123 -1396
rect 5088 -1566 5122 -1430
rect 5317 -1433 5860 -1361
rect 5864 -1358 5930 -1331
rect 5864 -1365 5898 -1358
rect 5926 -1365 5930 -1358
rect 5868 -1371 5930 -1365
rect 5926 -1376 5930 -1371
rect 5968 -1381 5972 -1376
rect 5972 -1392 6030 -1386
rect 5972 -1399 5984 -1392
rect 6004 -1399 6034 -1392
rect 5968 -1426 6034 -1399
rect 5972 -1432 6030 -1426
rect 6038 -1433 6072 -1324
rect 5317 -1450 6072 -1433
rect 5302 -1566 5327 -1542
rect 5423 -1566 5438 -1450
rect 4655 -1742 4753 -1619
rect 4833 -1655 4867 -1619
rect 4821 -1689 4967 -1655
rect 4833 -1717 4867 -1689
rect 5007 -1713 5021 -1689
rect 4452 -1765 4498 -1742
rect 4464 -1794 4498 -1765
rect 4552 -1776 4598 -1742
rect 4464 -1802 4510 -1794
rect 4546 -1802 4598 -1776
rect 4602 -1802 4636 -1742
rect 4350 -1804 4598 -1802
rect 2618 -1918 2623 -1812
rect 2624 -1838 2677 -1812
rect 2624 -1888 2689 -1838
rect 2697 -1888 2711 -1869
rect 2624 -1903 2711 -1888
rect 2624 -1909 2709 -1903
rect 2624 -1916 2689 -1909
rect 2734 -1916 2755 -1811
rect 2624 -1918 2755 -1916
rect 2505 -1968 2576 -1931
rect 2612 -1950 2670 -1918
rect 2683 -1919 2755 -1918
rect 2757 -1836 4598 -1804
rect 4604 -1836 4636 -1802
rect 4638 -1791 4753 -1742
rect 5024 -1751 5446 -1566
rect 4849 -1785 4911 -1751
rect 4849 -1791 4883 -1785
rect 2757 -1890 4384 -1836
rect 4464 -1844 4586 -1836
rect 4464 -1860 4510 -1844
rect 4518 -1850 4526 -1844
rect 4482 -1890 4510 -1860
rect 4546 -1878 4586 -1844
rect 4524 -1890 4532 -1887
rect 4552 -1890 4586 -1878
rect 2683 -1937 2737 -1919
rect 2734 -1946 2737 -1937
rect 2757 -1924 4598 -1890
rect 4604 -1924 4636 -1890
rect 2723 -1950 2741 -1946
rect 2612 -1951 2669 -1950
rect 2587 -1965 2604 -1959
rect 2608 -1962 2669 -1951
rect 2719 -1960 2753 -1950
rect 2612 -1965 2669 -1962
rect 2505 -2067 2539 -1968
rect 2549 -1980 2576 -1968
rect 2583 -1968 2669 -1965
rect 2692 -1962 2753 -1960
rect 2549 -1984 2570 -1980
rect 2583 -1999 2667 -1968
rect 2692 -1994 2707 -1962
rect 2719 -1965 2753 -1962
rect 2723 -1978 2753 -1965
rect 2587 -2005 2653 -1999
rect 2607 -2010 2653 -2005
rect 2559 -2015 2653 -2010
rect 2559 -2030 2622 -2015
rect 2559 -2033 2613 -2030
rect 2710 -2033 2753 -1978
rect 2707 -2067 2753 -2033
rect 2757 -2067 4384 -1924
rect 4424 -1958 4504 -1924
rect 4410 -1992 4512 -1958
rect 2441 -2072 2753 -2067
rect 2756 -2072 4384 -2067
rect 4424 -2026 4512 -1992
rect 4424 -2033 4504 -2026
rect 4424 -2035 4482 -2033
rect 4490 -2035 4504 -2033
rect 4424 -2045 4504 -2035
rect 4518 -2033 4598 -1924
rect 4518 -2045 4558 -2033
rect 4568 -2045 4598 -2033
rect 4424 -2049 4498 -2045
rect 4512 -2049 4586 -2045
rect 4424 -2058 4482 -2049
rect 4512 -2058 4570 -2049
rect 4424 -2069 4570 -2058
rect 2441 -2101 4384 -2072
rect 4400 -2071 4570 -2069
rect 4400 -2073 4434 -2071
rect 4436 -2073 4470 -2071
rect 1731 -2126 2384 -2120
rect 2407 -2126 2422 -2120
rect 2452 -2126 2486 -2101
rect 2505 -2126 2539 -2101
rect 2619 -2118 2653 -2101
rect 2707 -2118 2741 -2101
rect 2774 -2126 4384 -2101
rect 890 -2135 920 -2126
rect 929 -2132 4384 -2126
rect 4388 -2075 4470 -2073
rect 4474 -2073 4522 -2071
rect 4524 -2073 4558 -2071
rect 4474 -2075 4558 -2073
rect 4388 -2099 4440 -2075
rect 4474 -2086 4534 -2075
rect 4602 -2083 4636 -1924
rect 4474 -2092 4554 -2086
rect 4388 -2100 4438 -2099
rect 4388 -2109 4434 -2100
rect 4482 -2102 4558 -2092
rect 929 -2135 4356 -2132
rect 4388 -2134 4429 -2109
rect 4430 -2134 4434 -2109
rect 4476 -2109 4558 -2102
rect 193 -2152 872 -2140
rect 193 -2160 866 -2152
rect 883 -2158 4356 -2135
rect 883 -2160 4339 -2158
rect 193 -2178 630 -2160
rect 698 -2172 814 -2160
rect 829 -2172 844 -2160
rect 193 -2202 692 -2178
rect 698 -2183 844 -2172
rect 866 -2172 1694 -2160
rect 1731 -2161 2384 -2160
rect 1726 -2172 2384 -2161
rect 2385 -2172 2396 -2161
rect 866 -2181 2396 -2172
rect 706 -2202 756 -2183
rect 866 -2202 2170 -2181
rect 2238 -2183 2296 -2181
rect 2326 -2183 2396 -2181
rect 2250 -2187 2284 -2183
rect 2338 -2187 2396 -2183
rect 181 -2244 192 -2233
rect 193 -2244 630 -2202
rect 692 -2221 772 -2202
rect 708 -2222 756 -2221
rect 716 -2236 742 -2222
rect 758 -2230 772 -2221
rect 754 -2234 780 -2230
rect 754 -2238 788 -2234
rect 174 -2264 630 -2244
rect 738 -2264 804 -2238
rect 866 -2261 1711 -2202
rect 1731 -2208 2170 -2202
rect 2362 -2202 2396 -2187
rect 2362 -2208 2373 -2202
rect 1731 -2213 2373 -2208
rect 2385 -2208 2396 -2202
rect 2441 -2172 2486 -2160
rect 2505 -2172 2735 -2160
rect 2774 -2172 4339 -2160
rect 2441 -2189 4339 -2172
rect 2385 -2213 2422 -2208
rect 1731 -2233 2366 -2213
rect 1731 -2242 2373 -2233
rect 1731 -2261 2170 -2242
rect 2278 -2244 2296 -2242
rect 158 -2332 630 -2264
rect 784 -2272 820 -2264
rect 768 -2279 834 -2272
rect 752 -2283 834 -2279
rect 652 -2289 710 -2283
rect 652 -2332 653 -2289
rect 696 -2295 710 -2292
rect 664 -2298 710 -2295
rect 658 -2300 710 -2298
rect 740 -2298 834 -2283
rect 740 -2300 820 -2298
rect 832 -2300 834 -2298
rect 866 -2274 2170 -2261
rect 866 -2300 1712 -2274
rect 1731 -2300 2170 -2274
rect 2188 -2252 2254 -2249
rect 2278 -2252 2288 -2244
rect 2188 -2262 2322 -2252
rect 2328 -2262 2344 -2242
rect 2188 -2264 2344 -2262
rect 2362 -2243 2378 -2242
rect 2362 -2244 2396 -2243
rect 2407 -2244 2422 -2213
rect 2188 -2274 2322 -2264
rect 2188 -2276 2254 -2274
rect 2278 -2276 2322 -2274
rect 2188 -2280 2322 -2276
rect 2362 -2272 2422 -2244
rect 2441 -2272 2486 -2189
rect 2505 -2272 2539 -2189
rect 2663 -2198 2697 -2189
rect 2541 -2202 2691 -2199
rect 2647 -2227 2713 -2202
rect 2757 -2229 4339 -2189
rect 4361 -2194 4384 -2134
rect 4388 -2135 4438 -2134
rect 4464 -2135 4468 -2118
rect 4476 -2124 4534 -2109
rect 4542 -2124 4556 -2109
rect 4476 -2126 4556 -2124
rect 4476 -2135 4548 -2126
rect 4604 -2135 4636 -2083
rect 4638 -2129 4736 -1791
rect 4739 -1829 4753 -1791
rect 4781 -1829 4839 -1819
rect 4781 -1841 4845 -1829
rect 4781 -1853 4807 -1841
rect 4826 -1853 4845 -1841
rect 4854 -1853 4873 -1801
rect 4893 -1853 4927 -1819
rect 4793 -1887 4939 -1853
rect 5007 -1870 5446 -1751
rect 5457 -1747 5491 -1450
rect 5603 -1479 5615 -1450
rect 5686 -1467 6072 -1450
rect 5603 -1485 5661 -1479
rect 5686 -1503 5860 -1467
rect 5940 -1473 5974 -1469
rect 6028 -1473 6062 -1469
rect 5928 -1492 5986 -1473
rect 6016 -1492 6074 -1473
rect 5940 -1501 5974 -1492
rect 6028 -1501 6062 -1492
rect 5603 -1645 5661 -1639
rect 5603 -1679 5615 -1645
rect 5603 -1685 5661 -1679
rect 5457 -1781 5492 -1747
rect 5790 -1781 5860 -1503
rect 6057 -1554 6062 -1501
rect 6066 -1520 6074 -1492
rect 6091 -1486 6125 -1324
rect 6142 -1486 6176 -1324
rect 6193 -1299 6230 -1271
rect 6193 -1325 6239 -1299
rect 6306 -1305 6339 -1292
rect 6193 -1337 6230 -1325
rect 6303 -1337 6339 -1305
rect 6195 -1486 6229 -1337
rect 6303 -1341 6327 -1337
rect 6341 -1339 6399 -1333
rect 6337 -1363 6365 -1339
rect 6337 -1373 6361 -1363
rect 6373 -1373 6403 -1339
rect 6407 -1362 6967 -1271
rect 7075 -1256 7141 -1233
rect 7075 -1267 7091 -1256
rect 7111 -1267 7141 -1256
rect 7075 -1273 7137 -1267
rect 7075 -1283 7079 -1273
rect 7145 -1283 7179 -1222
rect 7268 -1227 7283 -1153
rect 7260 -1241 7283 -1227
rect 7302 -1138 7336 -1112
rect 7531 -1138 7984 -1112
rect 7302 -1146 7984 -1138
rect 7302 -1172 7337 -1146
rect 7410 -1151 7984 -1146
rect 7410 -1172 7971 -1151
rect 7302 -1241 7336 -1172
rect 7448 -1180 7506 -1174
rect 7444 -1206 7510 -1180
rect 7531 -1191 7971 -1172
rect 7448 -1207 7506 -1206
rect 7444 -1214 7510 -1207
rect 7448 -1220 7506 -1214
rect 7531 -1230 7953 -1191
rect 7382 -1241 7953 -1230
rect 7198 -1251 7233 -1241
rect 7294 -1248 7953 -1241
rect 7198 -1275 7235 -1251
rect 7294 -1252 7503 -1248
rect 7531 -1252 7953 -1248
rect 7294 -1275 7953 -1252
rect 7198 -1283 7232 -1275
rect 6975 -1290 7033 -1284
rect 6971 -1305 7037 -1290
rect 7047 -1305 7071 -1301
rect 6971 -1317 7071 -1305
rect 6971 -1324 7081 -1317
rect 6975 -1330 7033 -1324
rect 7035 -1340 7037 -1324
rect 7041 -1340 7081 -1324
rect 7035 -1349 7081 -1340
rect 7145 -1349 7232 -1283
rect 6237 -1384 6295 -1378
rect 6337 -1379 6399 -1373
rect 6233 -1418 6267 -1384
rect 6275 -1394 6299 -1384
rect 6337 -1389 6341 -1379
rect 6271 -1418 6299 -1394
rect 6237 -1424 6295 -1418
rect 6309 -1420 6333 -1416
rect 6297 -1449 6333 -1420
rect 6303 -1452 6333 -1449
rect 6407 -1452 6968 -1362
rect 7031 -1383 7081 -1349
rect 7135 -1383 7232 -1349
rect 7031 -1395 7065 -1383
rect 7145 -1395 7181 -1383
rect 7031 -1433 7077 -1395
rect 7079 -1433 7137 -1427
rect 7031 -1437 7071 -1433
rect 7075 -1437 7103 -1433
rect 7031 -1440 7103 -1437
rect 7041 -1452 7103 -1440
rect 6309 -1486 6343 -1452
rect 6407 -1486 6967 -1452
rect 7041 -1456 7065 -1452
rect 7075 -1467 7103 -1452
rect 7111 -1467 7141 -1433
rect 7075 -1473 7137 -1467
rect 7075 -1483 7079 -1473
rect 6091 -1520 6128 -1486
rect 6187 -1520 6967 -1486
rect 5972 -1700 6030 -1694
rect 5972 -1734 5984 -1700
rect 5972 -1740 6030 -1734
rect 5790 -1817 5843 -1781
rect 6161 -1836 6176 -1520
rect 6195 -1857 6229 -1520
rect 6424 -1535 6967 -1520
rect 6971 -1501 7014 -1490
rect 6971 -1524 7037 -1501
rect 7145 -1530 7179 -1395
rect 7164 -1535 7179 -1530
rect 7198 -1535 7232 -1383
rect 7249 -1535 7283 -1275
rect 7302 -1415 7336 -1275
rect 7404 -1309 7428 -1305
rect 7344 -1343 7402 -1337
rect 7404 -1342 7440 -1309
rect 7443 -1342 7456 -1275
rect 7340 -1377 7406 -1343
rect 7416 -1346 7440 -1342
rect 7344 -1383 7402 -1377
rect 7444 -1380 7448 -1364
rect 7471 -1370 7484 -1275
rect 7514 -1303 7953 -1275
rect 7504 -1330 7953 -1303
rect 7514 -1347 7953 -1330
rect 7987 -1204 8353 -821
rect 8356 -771 9114 -766
rect 8356 -777 8705 -771
rect 8356 -857 8390 -777
rect 8491 -794 8705 -777
rect 8463 -807 8705 -794
rect 8756 -777 9114 -771
rect 9125 -777 9565 -760
rect 8756 -779 9565 -777
rect 9581 -779 9880 -760
rect 8756 -781 9880 -779
rect 8756 -794 9581 -781
rect 9612 -794 9880 -781
rect 9955 -784 10238 -746
rect 10319 -671 10362 -655
rect 10372 -666 10412 -637
rect 10372 -671 10406 -666
rect 10319 -677 10408 -671
rect 10319 -687 10353 -677
rect 10372 -687 10406 -677
rect 10319 -753 10406 -687
rect 10520 -694 10554 -632
rect 10573 -694 10607 -632
rect 10688 -684 10722 -632
rect 10889 -641 10923 -622
rect 11074 -631 13093 -582
rect 10908 -651 10923 -641
rect 10942 -651 10977 -641
rect 10741 -656 10995 -651
rect 10741 -684 10815 -656
rect 10688 -685 10815 -684
rect 10837 -685 10995 -656
rect 11074 -654 11617 -631
rect 11627 -654 11661 -631
rect 11848 -648 11899 -631
rect 11916 -648 13093 -631
rect 11899 -654 13093 -648
rect 11074 -671 11600 -654
rect 11074 -682 11345 -671
rect 11431 -682 11460 -671
rect 10688 -690 10777 -685
rect 10518 -700 10607 -694
rect 8756 -802 9564 -794
rect 8463 -828 8511 -807
rect 8477 -837 8511 -828
rect 8621 -817 8669 -807
rect 8461 -838 8527 -837
rect 8621 -853 8705 -817
rect 8742 -824 9564 -802
rect 8742 -827 9060 -824
rect 8621 -857 8723 -853
rect 8356 -893 8723 -857
rect 8356 -949 8705 -893
rect 8742 -894 9074 -827
rect 9111 -833 9564 -824
rect 9581 -833 9615 -794
rect 9634 -833 9668 -794
rect 9672 -795 9706 -794
rect 9672 -798 9722 -795
rect 9676 -804 9734 -798
rect 9776 -828 9816 -794
rect 9832 -804 9880 -794
rect 9832 -824 9869 -804
rect 9832 -828 9864 -824
rect 9780 -833 9850 -828
rect 9111 -843 9547 -833
rect 9111 -877 9550 -843
rect 9562 -846 9720 -833
rect 9742 -834 9850 -833
rect 9742 -844 9816 -834
rect 9562 -866 9724 -846
rect 9742 -862 9782 -844
rect 9798 -866 9816 -844
rect 9832 -844 9850 -834
rect 9832 -866 9870 -844
rect 9562 -867 9784 -866
rect 9111 -890 9551 -877
rect 9626 -889 9784 -867
rect 9564 -890 9818 -889
rect 9832 -890 9866 -866
rect 8742 -900 9077 -894
rect 9111 -896 9866 -890
rect 9967 -881 10238 -784
rect 10318 -787 10406 -753
rect 10420 -772 10452 -721
rect 10518 -734 10554 -700
rect 10573 -734 10607 -700
rect 10715 -708 10731 -690
rect 10518 -740 10607 -734
rect 10319 -831 10353 -787
rect 10372 -803 10406 -787
rect 10474 -799 10506 -772
rect 10372 -831 10430 -803
rect 10319 -837 10430 -831
rect 10338 -871 10362 -837
rect 10372 -871 10430 -837
rect 10338 -877 10408 -871
rect 9111 -900 9888 -896
rect 8356 -953 8708 -949
rect 8742 -953 9091 -900
rect 7987 -1231 8342 -1204
rect 7987 -1244 8074 -1231
rect 8271 -1238 8276 -1231
rect 8280 -1238 8288 -1231
rect 8305 -1238 8342 -1231
rect 8356 -1238 8722 -953
rect 8271 -1244 8288 -1238
rect 8319 -1244 8722 -1238
rect 7987 -1278 8075 -1244
rect 8142 -1257 8722 -1244
rect 8142 -1278 8709 -1257
rect 8725 -1261 9091 -953
rect 7987 -1311 8074 -1278
rect 8154 -1293 8188 -1278
rect 8242 -1292 8288 -1278
rect 8356 -1292 8709 -1278
rect 8242 -1293 8276 -1292
rect 8280 -1293 8288 -1292
rect 8142 -1311 8200 -1293
rect 8230 -1311 8288 -1293
rect 8305 -1297 8709 -1292
rect 8305 -1311 8691 -1297
rect 7987 -1312 8691 -1311
rect 7987 -1326 8342 -1312
rect 7514 -1375 7971 -1347
rect 7987 -1367 8339 -1326
rect 7444 -1389 7468 -1380
rect 7410 -1415 7434 -1411
rect 7444 -1414 7472 -1389
rect 7480 -1414 7510 -1380
rect 7514 -1381 7987 -1375
rect 8004 -1381 8339 -1367
rect 7300 -1482 7337 -1415
rect 7410 -1445 7446 -1415
rect 7448 -1420 7468 -1414
rect 7514 -1429 7970 -1381
rect 7987 -1429 8339 -1381
rect 7514 -1443 7953 -1429
rect 7410 -1448 7440 -1445
rect 7422 -1452 7434 -1448
rect 7514 -1463 7959 -1443
rect 7514 -1482 7970 -1463
rect 7300 -1499 7970 -1482
rect 7300 -1505 7706 -1499
rect 7302 -1516 7706 -1505
rect 6424 -1538 7071 -1535
rect 6424 -1569 7145 -1538
rect 7198 -1569 7221 -1535
rect 7268 -1550 7283 -1535
rect 7344 -1543 7402 -1537
rect 7340 -1550 7406 -1543
rect 6424 -1592 6950 -1569
rect 6424 -1603 7145 -1592
rect 6424 -1609 6950 -1603
rect 5790 -1867 6229 -1857
rect 6341 -1827 6399 -1821
rect 6341 -1861 6353 -1827
rect 6341 -1867 6399 -1861
rect 4826 -1919 4845 -1887
rect 4854 -1947 4873 -1887
rect 5007 -1923 5105 -1870
rect 5007 -1996 5094 -1923
rect 5228 -1993 5255 -1870
rect 5256 -1965 5283 -1870
rect 5299 -1965 5302 -1870
rect 5327 -1970 5330 -1870
rect 5790 -1872 6215 -1867
rect 6530 -1944 6545 -1609
rect 6564 -1876 6598 -1609
rect 6793 -1662 6950 -1609
rect 7164 -1626 7179 -1569
rect 7198 -1626 7232 -1569
rect 7344 -1577 7356 -1550
rect 7514 -1552 7688 -1516
rect 7344 -1583 7402 -1577
rect 7514 -1583 7601 -1552
rect 7198 -1660 7213 -1626
rect 7531 -1679 7601 -1583
rect 7713 -1596 7771 -1590
rect 7713 -1630 7725 -1596
rect 7713 -1636 7771 -1630
rect 7531 -1715 7584 -1679
rect 7900 -1732 7970 -1499
rect 8004 -1484 8339 -1429
rect 8356 -1393 8691 -1312
rect 8742 -1310 9091 -1261
rect 9094 -913 9550 -900
rect 8742 -1337 9074 -1310
rect 9094 -1316 9443 -913
rect 8742 -1350 8812 -1337
rect 9043 -1344 9057 -1337
rect 8742 -1357 8813 -1350
rect 8742 -1393 8795 -1357
rect 8874 -1378 9057 -1350
rect 8874 -1393 9032 -1378
rect 8356 -1484 8390 -1393
rect 8451 -1394 8509 -1393
rect 8451 -1428 8463 -1394
rect 8742 -1399 9032 -1393
rect 9111 -1390 9443 -1316
rect 9463 -944 9550 -913
rect 9634 -930 9888 -900
rect 9967 -897 10221 -881
rect 9967 -920 10238 -897
rect 9630 -943 9664 -939
rect 9718 -943 9752 -939
rect 9630 -944 9676 -943
rect 9706 -944 9764 -943
rect 9832 -944 9866 -930
rect 9463 -978 9551 -944
rect 9600 -964 9866 -944
rect 9618 -978 9764 -964
rect 9463 -1272 9550 -978
rect 9636 -1030 9664 -1008
rect 9708 -1030 9755 -999
rect 9636 -1046 9676 -1030
rect 9706 -1046 9755 -1030
rect 9636 -1073 9755 -1046
rect 9618 -1123 9764 -1073
rect 9624 -1151 9670 -1127
rect 9708 -1151 9758 -1127
rect 9636 -1154 9664 -1151
rect 9708 -1154 9755 -1151
rect 9636 -1170 9676 -1154
rect 9706 -1170 9755 -1154
rect 9636 -1204 9755 -1170
rect 9636 -1220 9676 -1204
rect 9706 -1220 9746 -1204
rect 9636 -1238 9664 -1220
rect 9630 -1272 9664 -1238
rect 9718 -1238 9746 -1220
rect 9718 -1272 9752 -1238
rect 9463 -1306 9551 -1272
rect 9618 -1306 9764 -1272
rect 9770 -1295 9786 -1272
rect 9463 -1341 9550 -1306
rect 8621 -1417 8655 -1399
rect 8742 -1412 9078 -1399
rect 8742 -1417 8945 -1412
rect 9043 -1417 9078 -1412
rect 8451 -1434 8509 -1428
rect 8621 -1453 8691 -1417
rect 8742 -1432 9078 -1417
rect 8742 -1448 9077 -1432
rect 8419 -1475 8424 -1471
rect 8004 -1518 8328 -1484
rect 8382 -1518 8390 -1484
rect 8407 -1518 8444 -1475
rect 8638 -1487 8709 -1453
rect 8004 -1554 8339 -1518
rect 8419 -1552 8424 -1518
rect 8082 -1649 8140 -1643
rect 8082 -1683 8094 -1649
rect 8082 -1689 8140 -1683
rect 7900 -1768 7953 -1732
rect 6710 -1774 6768 -1768
rect 6710 -1808 6722 -1774
rect 6747 -1808 6768 -1774
rect 6710 -1814 6768 -1808
rect 6775 -1842 6796 -1776
rect 8269 -1785 8339 -1554
rect 8451 -1702 8509 -1696
rect 8451 -1736 8463 -1702
rect 8451 -1742 8509 -1736
rect 8269 -1821 8322 -1785
rect 8638 -1838 8708 -1487
rect 8820 -1555 8878 -1549
rect 8820 -1589 8832 -1555
rect 8820 -1595 8878 -1589
rect 8792 -1823 8798 -1721
rect 8820 -1755 8878 -1749
rect 8820 -1789 8832 -1755
rect 8820 -1795 8878 -1789
rect 8638 -1874 8691 -1838
rect 6564 -1910 6599 -1876
rect 6761 -1946 6950 -1889
rect 9007 -1891 9077 -1448
rect 9111 -1473 9429 -1390
rect 9480 -1437 9550 -1341
rect 9662 -1354 9720 -1348
rect 9662 -1388 9674 -1354
rect 9662 -1394 9720 -1388
rect 9832 -1394 9866 -964
rect 9967 -956 10221 -920
rect 10338 -939 10353 -877
rect 10372 -939 10406 -877
rect 10520 -894 10554 -740
rect 10573 -894 10607 -740
rect 10688 -724 10731 -708
rect 10741 -719 10781 -690
rect 10741 -724 10775 -719
rect 10688 -730 10777 -724
rect 10688 -740 10722 -730
rect 10741 -740 10775 -730
rect 10688 -806 10775 -740
rect 10889 -747 10923 -685
rect 10942 -747 10976 -685
rect 11074 -696 11340 -682
rect 11431 -688 11515 -682
rect 11679 -688 11695 -654
rect 11794 -688 13093 -654
rect 11057 -725 11340 -696
rect 11453 -715 11469 -688
rect 11426 -721 11469 -715
rect 11501 -721 11503 -710
rect 11627 -711 11661 -693
rect 11916 -702 13093 -688
rect 11848 -711 13093 -702
rect 11627 -720 13093 -711
rect 13117 -483 13147 -388
rect 14116 -417 14131 -383
rect 14451 -436 14466 -51
rect 14485 -85 14520 -51
rect 14485 -436 14519 -85
rect 14631 -153 14689 -147
rect 14631 -187 14643 -153
rect 14631 -193 14689 -187
rect 14631 -353 14689 -347
rect 14631 -387 14643 -353
rect 14631 -393 14689 -387
rect 13205 -456 13263 -450
rect 13117 -720 13151 -483
rect 13205 -490 13217 -456
rect 14485 -470 14500 -436
rect 13205 -496 13263 -490
rect 14818 -525 14871 -15
rect 13173 -537 13185 -533
rect 13161 -717 13205 -537
rect 15187 -578 15240 -121
rect 15556 -631 15609 -121
rect 15925 -684 15965 -227
rect 11627 -721 13089 -720
rect 11426 -724 13089 -721
rect 11057 -743 11345 -725
rect 10887 -753 10976 -747
rect 10687 -840 10775 -806
rect 10789 -825 10821 -774
rect 10887 -787 10923 -753
rect 10942 -787 10976 -753
rect 11074 -761 11345 -743
rect 10887 -793 10976 -787
rect 10688 -884 10722 -840
rect 10741 -856 10775 -840
rect 10843 -852 10875 -825
rect 10741 -884 10799 -856
rect 10688 -890 10799 -884
rect 10518 -900 10607 -894
rect 10518 -905 10554 -900
rect 10514 -934 10554 -905
rect 10573 -934 10607 -900
rect 10707 -924 10731 -890
rect 10741 -924 10799 -890
rect 10707 -930 10777 -924
rect 10518 -939 10588 -934
rect 10300 -948 10458 -939
rect 10480 -940 10588 -939
rect 10480 -948 10554 -940
rect 9967 -966 10020 -956
rect 10300 -973 10554 -948
rect 10573 -950 10588 -940
rect 10573 -973 10607 -950
rect 10338 -983 10353 -973
rect 10372 -983 10406 -973
rect 10372 -1017 10387 -983
rect 10573 -1002 10588 -973
rect 10707 -992 10722 -930
rect 10741 -992 10775 -930
rect 10889 -947 10923 -793
rect 10942 -947 10976 -793
rect 11057 -859 11345 -761
rect 11056 -893 11345 -859
rect 11057 -943 11345 -893
rect 11426 -747 11697 -724
rect 11812 -737 13089 -724
rect 11426 -757 11715 -747
rect 11426 -791 11697 -757
rect 11812 -760 12355 -737
rect 12365 -760 12399 -737
rect 12586 -754 12637 -737
rect 12654 -754 13089 -737
rect 13139 -744 13151 -720
rect 13173 -721 13185 -717
rect 13093 -754 13151 -744
rect 12637 -760 13093 -754
rect 11812 -777 12338 -760
rect 11812 -788 12083 -777
rect 12169 -788 12198 -777
rect 11426 -903 11714 -791
rect 11812 -802 12078 -788
rect 12169 -794 12253 -788
rect 12417 -794 12433 -760
rect 12532 -794 13093 -760
rect 11795 -831 12078 -802
rect 12191 -821 12207 -794
rect 12654 -798 13093 -794
rect 13205 -764 13263 -758
rect 13205 -798 13217 -764
rect 12164 -827 12207 -821
rect 12239 -827 12241 -816
rect 12365 -817 12399 -799
rect 12654 -808 13076 -798
rect 13205 -804 13263 -798
rect 12586 -817 13076 -808
rect 12365 -827 13076 -817
rect 12164 -830 13076 -827
rect 11795 -849 12083 -831
rect 11812 -867 12083 -849
rect 11425 -937 11714 -903
rect 10887 -953 10976 -947
rect 10887 -958 10923 -953
rect 10883 -987 10923 -958
rect 10942 -987 10976 -953
rect 11074 -959 11345 -943
rect 11426 -949 11714 -937
rect 11443 -958 11714 -949
rect 11074 -968 11328 -959
rect 10887 -992 10957 -987
rect 10406 -1007 10588 -1002
rect 10669 -1001 10827 -992
rect 10849 -993 10957 -992
rect 10849 -1001 10923 -993
rect 10669 -1026 10923 -1001
rect 10942 -1003 10957 -993
rect 10942 -1026 10976 -1003
rect 10707 -1036 10722 -1026
rect 10741 -1036 10775 -1026
rect 10741 -1070 10756 -1036
rect 10942 -1055 10957 -1026
rect 10775 -1060 10957 -1055
rect 11074 -1040 11340 -968
rect 11431 -996 11714 -958
rect 11795 -965 12083 -867
rect 11074 -1056 11328 -1040
rect 11074 -1079 11345 -1056
rect 11074 -1115 11328 -1079
rect 11443 -1093 11714 -996
rect 11794 -999 12083 -965
rect 11795 -1049 12083 -999
rect 12164 -853 12435 -830
rect 12550 -832 13076 -830
rect 13093 -832 13103 -812
rect 12164 -863 12453 -853
rect 12164 -897 12435 -863
rect 12550 -866 13093 -832
rect 13103 -866 13137 -832
rect 12550 -883 13076 -866
rect 12550 -894 12821 -883
rect 12907 -894 12936 -883
rect 12164 -1009 12452 -897
rect 12550 -908 12816 -894
rect 12907 -900 12991 -894
rect 13155 -900 13171 -866
rect 12533 -937 12816 -908
rect 12929 -927 12945 -900
rect 12902 -934 12945 -927
rect 12533 -955 12821 -937
rect 12550 -973 12821 -955
rect 12163 -1043 12452 -1009
rect 11812 -1065 12083 -1049
rect 12164 -1055 12452 -1043
rect 12181 -1064 12452 -1055
rect 11812 -1074 12066 -1065
rect 11443 -1109 11697 -1093
rect 11074 -1125 11127 -1115
rect 11443 -1132 11714 -1109
rect 11443 -1168 11697 -1132
rect 11812 -1146 12078 -1074
rect 12169 -1102 12452 -1064
rect 12533 -1071 12821 -973
rect 11812 -1162 12066 -1146
rect 11443 -1178 11496 -1168
rect 11812 -1185 12083 -1162
rect 11812 -1221 12066 -1185
rect 12181 -1199 12452 -1102
rect 12532 -1105 12821 -1071
rect 12533 -1155 12821 -1105
rect 12902 -940 12991 -934
rect 12902 -959 12936 -940
rect 12902 -1115 12969 -959
rect 12901 -1149 12969 -1115
rect 12550 -1171 12821 -1155
rect 12902 -1161 12936 -1149
rect 12550 -1180 12804 -1171
rect 12181 -1215 12435 -1199
rect 11812 -1231 11865 -1221
rect 12181 -1238 12452 -1215
rect 12181 -1274 12435 -1238
rect 12550 -1252 12816 -1180
rect 12907 -1202 12936 -1170
rect 12907 -1208 12991 -1202
rect 12929 -1242 12945 -1208
rect 12929 -1248 12991 -1242
rect 12550 -1268 12804 -1252
rect 12929 -1258 12936 -1248
rect 12181 -1284 12234 -1274
rect 12550 -1291 12821 -1268
rect 12925 -1269 12936 -1258
rect 12550 -1327 12804 -1291
rect 12550 -1337 12603 -1327
rect 9480 -1473 9533 -1437
rect 9189 -1500 9247 -1494
rect 9189 -1534 9201 -1500
rect 9480 -1526 9683 -1473
rect 9189 -1540 9247 -1534
rect 9189 -1808 9247 -1802
rect 9189 -1842 9201 -1808
rect 9189 -1848 9247 -1842
rect 9007 -1927 9060 -1891
rect 6159 -1963 6215 -1946
rect 5007 -1997 5206 -1996
rect 5024 -2014 5206 -1997
rect 6159 -1999 6581 -1963
rect 5024 -2024 5094 -2014
rect 5024 -2042 5206 -2024
rect 5024 -2093 5094 -2042
rect 5024 -2095 5082 -2093
rect 5024 -2113 5094 -2095
rect 5206 -2113 5241 -2095
rect 5024 -2114 5241 -2113
rect 5280 -2114 5460 -2094
rect 5024 -2128 5460 -2114
rect 5521 -2128 5556 -2094
rect 4638 -2132 4700 -2129
rect 4638 -2135 4690 -2132
rect 2567 -2257 2633 -2245
rect 2757 -2246 4381 -2229
rect 4388 -2246 4736 -2135
rect 5024 -2148 5314 -2128
rect 5522 -2147 5556 -2128
rect 4837 -2170 4852 -2149
rect 5024 -2152 5240 -2148
rect 4871 -2170 5240 -2152
rect 4781 -2171 5240 -2170
rect 4763 -2205 5240 -2171
rect 5541 -2190 5556 -2147
rect 4764 -2206 5240 -2205
rect 2757 -2254 4736 -2246
rect 2567 -2262 2599 -2257
rect 2757 -2261 4339 -2254
rect 2567 -2272 2633 -2262
rect 2757 -2272 4349 -2261
rect 2188 -2283 2298 -2280
rect 2196 -2300 2298 -2283
rect 2362 -2300 4349 -2272
rect 4395 -2264 4736 -2254
rect 4781 -2264 5240 -2206
rect 4395 -2300 5240 -2264
rect 5320 -2300 5354 -2266
rect 5408 -2300 5442 -2266
rect 5522 -2300 5556 -2190
rect 5575 -2181 5610 -2147
rect 5575 -2300 5609 -2181
rect 7366 -2213 7401 -2179
rect 5721 -2249 5779 -2243
rect 5721 -2262 5733 -2249
rect 5721 -2264 5767 -2262
rect 5721 -2266 5779 -2264
rect 5717 -2283 5783 -2266
rect 5891 -2272 5925 -2243
rect 6277 -2272 6488 -2217
rect 7367 -2232 7401 -2213
rect 5721 -2289 5779 -2283
rect 5693 -2300 5807 -2292
rect 5891 -2300 6234 -2272
rect 658 -2332 6234 -2300
rect 158 -2343 649 -2332
rect 652 -2334 6234 -2332
rect 158 -2346 638 -2343
rect 652 -2346 850 -2334
rect 158 -2347 639 -2346
rect 158 -2374 584 -2347
rect 596 -2348 639 -2347
rect 649 -2348 850 -2346
rect 866 -2340 4349 -2334
rect 866 -2346 4320 -2340
rect 866 -2347 3170 -2346
rect 866 -2348 2043 -2347
rect 596 -2352 2043 -2348
rect 2046 -2352 2106 -2347
rect 596 -2366 2106 -2352
rect 2136 -2366 3170 -2347
rect 621 -2374 639 -2366
rect 158 -2388 639 -2374
rect 649 -2374 710 -2366
rect 649 -2388 746 -2374
rect 158 -2398 584 -2388
rect 650 -2396 710 -2388
rect 752 -2396 798 -2366
rect 866 -2374 2106 -2366
rect 847 -2388 2106 -2374
rect 813 -2396 820 -2388
rect 650 -2398 738 -2396
rect 752 -2398 826 -2396
rect 158 -2400 596 -2398
rect 650 -2400 860 -2398
rect 158 -2402 584 -2400
rect 650 -2402 738 -2400
rect 158 -2416 602 -2402
rect 644 -2414 746 -2402
rect 752 -2414 826 -2400
rect 644 -2416 826 -2414
rect 158 -2437 584 -2416
rect 650 -2420 826 -2416
rect 832 -2402 860 -2400
rect 866 -2402 2106 -2388
rect 832 -2416 2106 -2402
rect 832 -2420 860 -2416
rect 866 -2420 2106 -2416
rect 596 -2437 2106 -2420
rect 158 -2454 2106 -2437
rect 158 -2526 630 -2454
rect 650 -2476 684 -2454
rect 691 -2463 704 -2454
rect 719 -2463 792 -2454
rect 691 -2467 698 -2463
rect 719 -2467 786 -2463
rect 719 -2476 772 -2467
rect 807 -2475 860 -2454
rect 158 -2558 643 -2526
rect 650 -2558 690 -2476
rect 719 -2491 776 -2476
rect 692 -2504 696 -2494
rect 692 -2510 718 -2504
rect 725 -2506 776 -2491
rect 725 -2510 784 -2506
rect 692 -2516 784 -2510
rect 788 -2516 860 -2475
rect 692 -2544 860 -2516
rect 692 -2550 718 -2544
rect 725 -2549 860 -2544
rect 866 -2476 2106 -2454
rect 2148 -2380 2194 -2366
rect 2200 -2380 2282 -2366
rect 2148 -2387 2282 -2380
rect 2288 -2387 3170 -2366
rect 2148 -2388 3170 -2387
rect 2148 -2391 2308 -2388
rect 2148 -2398 2314 -2391
rect 2317 -2398 2320 -2391
rect 2148 -2414 2335 -2398
rect 2148 -2439 2160 -2414
rect 2148 -2448 2163 -2439
rect 2168 -2448 2335 -2414
rect 2148 -2450 2220 -2448
rect 2248 -2450 2335 -2448
rect 2148 -2454 2230 -2450
rect 866 -2480 2111 -2476
rect 2148 -2480 2226 -2454
rect 2242 -2466 2335 -2450
rect 2242 -2480 2320 -2466
rect 866 -2549 2117 -2480
rect 2140 -2495 2145 -2491
rect 2134 -2496 2145 -2495
rect 2160 -2495 2226 -2480
rect 2228 -2482 2320 -2480
rect 2160 -2496 2220 -2495
rect 2228 -2496 2308 -2482
rect 2129 -2507 2153 -2496
rect 2160 -2498 2308 -2496
rect 2165 -2507 2262 -2498
rect 692 -2558 696 -2550
rect 725 -2556 2117 -2549
rect 158 -2582 698 -2558
rect 725 -2562 800 -2556
rect 725 -2568 786 -2562
rect 807 -2568 2117 -2556
rect 158 -2607 634 -2582
rect 158 -2612 630 -2607
rect 638 -2612 688 -2582
rect 710 -2598 786 -2568
rect 798 -2582 2117 -2568
rect 798 -2586 860 -2582
rect 798 -2598 859 -2586
rect 710 -2599 725 -2598
rect 710 -2603 718 -2599
rect 726 -2603 739 -2598
rect 744 -2602 772 -2598
rect 756 -2603 772 -2602
rect 798 -2599 813 -2598
rect 798 -2603 806 -2599
rect 832 -2602 847 -2598
rect 698 -2608 741 -2603
rect 698 -2610 725 -2608
rect 691 -2612 725 -2610
rect 726 -2612 741 -2608
rect 764 -2612 772 -2603
rect 786 -2612 829 -2603
rect 841 -2612 844 -2603
rect 866 -2612 2117 -2582
rect 158 -2620 2117 -2612
rect 158 -2636 630 -2620
rect 638 -2623 688 -2620
rect 691 -2623 2117 -2620
rect 646 -2636 664 -2623
rect 691 -2626 1377 -2623
rect 698 -2636 1377 -2626
rect 158 -2646 844 -2636
rect 864 -2646 1377 -2636
rect 158 -2690 630 -2646
rect 710 -2690 744 -2646
rect 751 -2690 756 -2646
rect 786 -2658 814 -2646
rect 829 -2658 844 -2646
rect 786 -2688 844 -2658
rect 798 -2690 844 -2688
rect 883 -2690 1377 -2646
rect 158 -2703 1377 -2690
rect 1397 -2703 1402 -2623
rect 1408 -2631 1525 -2623
rect 1530 -2631 1553 -2623
rect 1579 -2631 1582 -2623
rect 1408 -2650 1582 -2631
rect 1408 -2666 1494 -2650
rect 1408 -2688 1431 -2666
rect 1443 -2677 1494 -2666
rect 1500 -2677 1582 -2650
rect 1604 -2625 2117 -2623
rect 2134 -2510 2220 -2507
rect 2228 -2510 2262 -2507
rect 2274 -2510 2308 -2498
rect 2134 -2556 2308 -2510
rect 2317 -2556 2320 -2482
rect 2134 -2571 2320 -2556
rect 2342 -2500 3170 -2388
rect 3179 -2414 3213 -2346
rect 3215 -2361 3249 -2346
rect 3277 -2357 3303 -2346
rect 3277 -2360 3327 -2357
rect 3381 -2360 3415 -2346
rect 3277 -2361 3339 -2360
rect 3369 -2361 3427 -2360
rect 3486 -2361 4320 -2346
rect 3215 -2377 4320 -2361
rect 4395 -2352 5572 -2334
rect 5575 -2352 5609 -2334
rect 5651 -2346 5823 -2334
rect 3215 -2395 4327 -2377
rect 3281 -2403 3339 -2395
rect 3369 -2403 3427 -2395
rect 3486 -2402 4327 -2395
rect 3293 -2407 3327 -2403
rect 3381 -2407 3415 -2403
rect 3486 -2413 4341 -2402
rect 3486 -2414 4330 -2413
rect 3179 -2418 4330 -2414
rect 4342 -2418 4349 -2388
rect 4395 -2402 5609 -2352
rect 5689 -2372 5723 -2346
rect 5777 -2367 5811 -2346
rect 5747 -2372 5811 -2367
rect 5871 -2362 5877 -2346
rect 5891 -2362 6234 -2334
rect 5747 -2380 5794 -2372
rect 4382 -2418 5609 -2402
rect 5679 -2414 5689 -2380
rect 5729 -2388 5797 -2380
rect 5697 -2408 5735 -2398
rect 5747 -2408 5797 -2388
rect 3179 -2429 5609 -2418
rect 3179 -2476 3194 -2429
rect 3259 -2441 3449 -2429
rect 3486 -2436 5609 -2429
rect 3310 -2448 3398 -2441
rect 3486 -2451 4321 -2436
rect 3179 -2481 3213 -2476
rect 3321 -2491 3387 -2458
rect 3486 -2476 4303 -2451
rect 4308 -2463 4321 -2451
rect 4308 -2467 4315 -2463
rect 2134 -2575 2296 -2571
rect 2134 -2618 2274 -2575
rect 2342 -2597 3187 -2500
rect 3486 -2507 4305 -2476
rect 4336 -2489 4353 -2436
rect 4336 -2491 4349 -2489
rect 4342 -2501 4349 -2491
rect 3311 -2516 3345 -2509
rect 3201 -2577 3455 -2543
rect 3486 -2557 4113 -2507
rect 4203 -2510 4207 -2507
rect 4129 -2542 4139 -2526
rect 4124 -2557 4139 -2542
rect 4220 -2537 4241 -2507
rect 4242 -2537 4305 -2507
rect 4361 -2537 4388 -2436
rect 4395 -2537 5609 -2436
rect 5697 -2416 5797 -2408
rect 5808 -2416 5823 -2401
rect 5677 -2448 5692 -2439
rect 5697 -2448 5823 -2416
rect 5677 -2452 5735 -2448
rect 5777 -2450 5823 -2448
rect 5743 -2452 5759 -2450
rect 5677 -2454 5759 -2452
rect 5635 -2480 5640 -2476
rect 5677 -2480 5735 -2454
rect 5635 -2492 5646 -2480
rect 4220 -2544 5609 -2537
rect 3486 -2560 4139 -2557
rect 3267 -2588 3301 -2584
rect 3355 -2588 3389 -2584
rect 2134 -2625 2205 -2618
rect 1604 -2648 2205 -2625
rect 1604 -2659 2174 -2648
rect 2180 -2659 2205 -2648
rect 2214 -2652 2296 -2618
rect 2216 -2659 2274 -2652
rect 1604 -2660 2316 -2659
rect 1448 -2681 1465 -2677
rect 1410 -2703 1431 -2688
rect 1494 -2700 1525 -2677
rect 1531 -2678 1566 -2677
rect 1531 -2700 1597 -2678
rect 1494 -2703 1597 -2700
rect 1604 -2693 2067 -2660
rect 2106 -2666 2111 -2660
rect 2123 -2666 2316 -2660
rect 2342 -2666 2376 -2597
rect 2379 -2666 3187 -2597
rect 3255 -2602 3313 -2588
rect 3343 -2602 3401 -2588
rect 3267 -2611 3301 -2602
rect 3355 -2611 3389 -2602
rect 2106 -2675 2945 -2666
rect 2106 -2686 2168 -2675
rect 2180 -2682 2228 -2675
rect 2175 -2686 2228 -2682
rect 2234 -2686 2945 -2675
rect 2106 -2693 2945 -2686
rect 1604 -2703 2060 -2693
rect 158 -2724 2060 -2703
rect 158 -2726 630 -2724
rect 710 -2726 744 -2724
rect 751 -2726 756 -2724
rect 798 -2726 832 -2724
rect 839 -2726 2060 -2724
rect 158 -2737 2060 -2726
rect 2072 -2703 2111 -2693
rect 2072 -2720 2106 -2703
rect 2126 -2706 2252 -2693
rect 2150 -2720 2252 -2706
rect 2275 -2720 2276 -2693
rect 2342 -2720 2376 -2693
rect 2379 -2697 2945 -2693
rect 2379 -2703 2988 -2697
rect 2379 -2720 2945 -2703
rect 2072 -2727 2945 -2720
rect 2072 -2731 2326 -2727
rect 2072 -2732 2114 -2731
rect 2123 -2732 2153 -2731
rect 2072 -2737 2153 -2732
rect 2168 -2737 2326 -2731
rect 158 -2754 2326 -2737
rect 2342 -2754 2376 -2727
rect 2379 -2737 2945 -2727
rect 2379 -2754 2705 -2737
rect 158 -2760 2305 -2754
rect 158 -2816 630 -2760
rect 654 -2768 775 -2760
rect 698 -2783 775 -2768
rect 818 -2779 844 -2760
rect 786 -2783 844 -2779
rect 852 -2762 2316 -2760
rect 2342 -2762 2705 -2754
rect 852 -2770 2094 -2762
rect 2157 -2770 2316 -2762
rect 852 -2771 2316 -2770
rect 852 -2773 2066 -2771
rect 2275 -2772 2276 -2771
rect 852 -2783 2043 -2773
rect 710 -2786 744 -2783
rect 682 -2787 744 -2786
rect 682 -2792 725 -2787
rect 678 -2804 744 -2792
rect 676 -2811 744 -2804
rect 193 -2846 201 -2816
rect 172 -2854 201 -2846
rect 227 -2854 261 -2816
rect 281 -2829 295 -2825
rect 369 -2829 403 -2825
rect 269 -2844 297 -2829
rect 357 -2840 415 -2829
rect 269 -2854 295 -2844
rect 357 -2854 403 -2840
rect 500 -2843 630 -2816
rect 678 -2812 744 -2811
rect 751 -2812 786 -2783
rect 818 -2787 832 -2783
rect 852 -2786 866 -2783
rect 869 -2786 2043 -2783
rect 678 -2814 786 -2812
rect 852 -2804 2043 -2786
rect 852 -2805 1000 -2804
rect 1048 -2805 2043 -2804
rect 678 -2821 744 -2814
rect 678 -2842 696 -2824
rect 704 -2826 744 -2821
rect 759 -2824 770 -2814
rect 726 -2830 738 -2826
rect 726 -2835 778 -2830
rect 726 -2842 804 -2835
rect 483 -2854 630 -2843
rect 144 -2901 630 -2854
rect 646 -2866 696 -2846
rect 738 -2864 804 -2842
rect 738 -2866 806 -2864
rect 649 -2873 696 -2866
rect 743 -2869 806 -2866
rect 738 -2873 806 -2869
rect 638 -2878 806 -2873
rect 638 -2882 828 -2878
rect 835 -2880 846 -2824
rect 852 -2854 982 -2805
rect 1131 -2854 1155 -2805
rect 1157 -2807 2043 -2805
rect 2053 -2807 2066 -2773
rect 2376 -2776 2705 -2762
rect 2379 -2781 2705 -2776
rect 2342 -2792 2353 -2781
rect 2371 -2782 2705 -2781
rect 2371 -2792 2382 -2782
rect 1157 -2824 2066 -2807
rect 2275 -2824 2282 -2792
rect 2342 -2824 2382 -2792
rect 2480 -2807 2705 -2782
rect 2748 -2782 2945 -2737
rect 2748 -2789 2959 -2782
rect 3117 -2789 3187 -2666
rect 3486 -2613 3565 -2560
rect 3674 -2573 4139 -2560
rect 3674 -2607 4161 -2573
rect 4207 -2597 5609 -2544
rect 5631 -2597 5646 -2492
rect 5669 -2495 5674 -2491
rect 5663 -2496 5674 -2495
rect 5689 -2495 5735 -2480
rect 5771 -2463 5823 -2450
rect 5830 -2463 5846 -2432
rect 5771 -2466 5846 -2463
rect 5771 -2482 5823 -2466
rect 5757 -2495 5762 -2491
rect 5658 -2507 5682 -2496
rect 5689 -2498 5734 -2495
rect 5751 -2496 5762 -2495
rect 5746 -2497 5765 -2496
rect 5777 -2497 5823 -2482
rect 5871 -2497 6234 -2362
rect 5694 -2507 5734 -2498
rect 3674 -2612 4139 -2607
rect 4207 -2612 5646 -2597
rect 3299 -2716 3357 -2710
rect 3486 -2715 3556 -2613
rect 3674 -2623 5646 -2612
rect 3674 -2629 5015 -2623
rect 3724 -2652 3769 -2629
rect 3823 -2652 3945 -2629
rect 3999 -2652 4039 -2629
rect 4045 -2635 5015 -2629
rect 4079 -2641 5015 -2635
rect 4079 -2646 4139 -2641
rect 4175 -2643 5015 -2641
rect 5018 -2643 5025 -2623
rect 5027 -2643 5054 -2623
rect 5055 -2643 5082 -2623
rect 5133 -2624 5646 -2623
rect 5663 -2510 5734 -2507
rect 5736 -2510 6234 -2497
rect 5663 -2541 5728 -2510
rect 5735 -2520 5803 -2510
rect 5804 -2514 6234 -2510
rect 6277 -2287 6348 -2272
rect 7197 -2281 7255 -2275
rect 6277 -2514 6347 -2287
rect 7197 -2315 7209 -2281
rect 7197 -2321 7255 -2315
rect 6459 -2355 6517 -2349
rect 6459 -2389 6471 -2355
rect 6629 -2378 6663 -2360
rect 7051 -2378 7085 -2360
rect 6459 -2395 6517 -2389
rect 6629 -2414 6699 -2378
rect 5804 -2520 6347 -2514
rect 5735 -2523 6347 -2520
rect 5734 -2531 6347 -2523
rect 5734 -2541 5803 -2531
rect 5663 -2559 5803 -2541
rect 5871 -2550 6347 -2531
rect 6646 -2448 6717 -2414
rect 5663 -2607 5804 -2559
rect 5871 -2584 6359 -2550
rect 6415 -2584 6455 -2550
rect 5871 -2599 6347 -2584
rect 5663 -2624 5734 -2607
rect 5133 -2643 5734 -2624
rect 4175 -2646 5734 -2643
rect 3724 -2664 3758 -2652
rect 3838 -2664 3872 -2652
rect 3692 -2679 3758 -2664
rect 3766 -2679 3770 -2664
rect 3692 -2711 3770 -2679
rect 3299 -2738 3311 -2716
rect 3299 -2756 3357 -2738
rect 3271 -2784 3385 -2766
rect 3469 -2769 3556 -2715
rect 3624 -2722 3664 -2715
rect 3712 -2735 3773 -2711
rect 3712 -2746 3793 -2735
rect 3712 -2760 3762 -2746
rect 3668 -2769 3726 -2763
rect 3727 -2769 3754 -2760
rect 2748 -2799 3187 -2789
rect 2748 -2807 2959 -2799
rect 2671 -2816 2705 -2807
rect 2734 -2816 2959 -2807
rect 1157 -2835 2094 -2824
rect 2163 -2834 2251 -2824
rect 2125 -2835 2251 -2834
rect 2264 -2826 2382 -2824
rect 2264 -2835 2305 -2826
rect 2371 -2833 2382 -2826
rect 1157 -2836 2083 -2835
rect 2125 -2836 2240 -2835
rect 2275 -2836 2305 -2835
rect 2348 -2836 2382 -2833
rect 1157 -2841 2382 -2836
rect 1157 -2854 1697 -2841
rect 852 -2862 1697 -2854
rect 1743 -2862 1747 -2841
rect 635 -2890 696 -2882
rect 726 -2890 828 -2882
rect 852 -2890 1765 -2862
rect 1777 -2867 1811 -2856
rect 1823 -2867 1853 -2841
rect 1873 -2856 1895 -2841
rect 1865 -2867 1899 -2856
rect 1979 -2862 2013 -2841
rect 2026 -2858 2382 -2841
rect 1911 -2867 2013 -2862
rect 1771 -2868 1823 -2867
rect 1774 -2879 1823 -2868
rect 1777 -2882 1823 -2879
rect 1858 -2882 2013 -2867
rect 1777 -2890 1819 -2882
rect 1865 -2890 1907 -2882
rect 1911 -2890 2013 -2882
rect 2032 -2890 2066 -2858
rect 2125 -2873 2240 -2858
rect 2125 -2884 2191 -2873
rect 2275 -2889 2282 -2858
rect 2348 -2862 2382 -2858
rect 2734 -2862 2945 -2816
rect 3117 -2852 3174 -2799
rect 3472 -2803 3557 -2769
rect 3653 -2780 3827 -2769
rect 3664 -2792 3754 -2780
rect 3781 -2792 3811 -2780
rect 3857 -2788 3872 -2664
rect 3653 -2803 3754 -2792
rect 3770 -2803 3822 -2792
rect 3472 -2852 3556 -2803
rect 3668 -2809 3726 -2803
rect 3727 -2813 3754 -2803
rect 3664 -2819 3754 -2813
rect 3727 -2830 3754 -2819
rect 3843 -2816 3872 -2788
rect 3891 -2664 3925 -2652
rect 3843 -2822 3877 -2816
rect 3891 -2822 3906 -2664
rect 3923 -2785 3925 -2683
rect 3993 -2686 4002 -2664
rect 4005 -2670 4039 -2652
rect 4207 -2658 5734 -2646
rect 4207 -2659 5609 -2658
rect 5635 -2659 5734 -2658
rect 5736 -2659 5804 -2607
rect 5878 -2649 6347 -2599
rect 6421 -2616 6455 -2584
rect 6433 -2646 6455 -2625
rect 4207 -2660 5845 -2659
rect 4005 -2686 4052 -2670
rect 3957 -2751 3959 -2717
rect 3993 -2751 4052 -2686
rect 4207 -2688 5594 -2660
rect 5635 -2670 5845 -2660
rect 5635 -2682 5834 -2670
rect 5896 -2680 6347 -2649
rect 5838 -2682 6347 -2680
rect 4207 -2693 5590 -2688
rect 5635 -2692 6347 -2682
rect 3993 -2767 4023 -2751
rect 4081 -2760 4099 -2717
rect 4207 -2726 5589 -2693
rect 5635 -2703 5640 -2692
rect 5641 -2693 6347 -2692
rect 5679 -2720 5724 -2693
rect 5679 -2722 5693 -2720
rect 3993 -2768 4008 -2767
rect 4081 -2768 4114 -2760
rect 3993 -2775 4033 -2768
rect 4081 -2775 4139 -2768
rect 4207 -2776 5575 -2726
rect 5578 -2732 5589 -2726
rect 4207 -2779 5572 -2776
rect 5582 -2779 5589 -2732
rect 5683 -2756 5693 -2722
rect 5697 -2722 5724 -2720
rect 5736 -2722 5781 -2693
rect 5697 -2727 5781 -2722
rect 5697 -2756 5724 -2727
rect 5683 -2762 5724 -2756
rect 5736 -2756 5781 -2727
rect 4207 -2784 5637 -2779
rect 4207 -2804 5572 -2784
rect 3843 -2838 3906 -2822
rect 3925 -2822 4025 -2816
rect 4083 -2822 4095 -2820
rect 3925 -2833 4110 -2822
rect 3925 -2838 4025 -2833
rect 3843 -2842 4025 -2838
rect 2192 -2890 2222 -2889
rect 2348 -2890 2691 -2862
rect 635 -2901 2691 -2890
rect 144 -2924 2691 -2901
rect 144 -2932 696 -2924
rect 727 -2932 793 -2924
rect 852 -2930 2029 -2924
rect 2032 -2930 2083 -2924
rect 2108 -2925 2305 -2924
rect 2108 -2930 2316 -2925
rect 852 -2932 2316 -2930
rect 144 -2934 2316 -2932
rect 144 -2936 2328 -2934
rect 144 -2966 2075 -2936
rect 144 -2969 696 -2966
rect 144 -3000 570 -2969
rect 116 -3006 570 -3000
rect 144 -3058 570 -3006
rect 582 -3058 604 -2969
rect 607 -2978 625 -2969
rect 607 -3006 622 -2978
rect 612 -3047 622 -3006
rect 616 -3058 622 -3047
rect 628 -3032 696 -2969
rect 738 -2967 772 -2966
rect 738 -2978 784 -2967
rect 704 -3007 719 -2978
rect 732 -3007 784 -2978
rect 704 -3008 784 -3007
rect 799 -3008 806 -2978
rect 852 -3002 2075 -2966
rect 2095 -2942 2100 -2936
rect 2112 -2942 2129 -2936
rect 2095 -2962 2129 -2942
rect 711 -3009 778 -3008
rect 700 -3020 778 -3009
rect 711 -3025 778 -3020
rect 793 -3014 806 -3008
rect 818 -3008 833 -3004
rect 852 -3008 2083 -3002
rect 818 -3014 845 -3008
rect 793 -3025 845 -3014
rect 711 -3032 845 -3025
rect 628 -3058 845 -3032
rect 144 -3059 845 -3058
rect 144 -3164 570 -3059
rect 582 -3063 604 -3059
rect 673 -3066 674 -3059
rect 685 -3066 845 -3059
rect 660 -3100 845 -3066
rect 673 -3114 845 -3100
rect 673 -3126 833 -3114
rect 678 -3134 762 -3126
rect 597 -3160 602 -3147
rect 678 -3150 757 -3134
rect 699 -3154 714 -3150
rect 621 -3160 639 -3154
rect 649 -3160 714 -3154
rect 731 -3160 757 -3150
rect 773 -3154 779 -3126
rect 818 -3160 833 -3126
rect 835 -3160 845 -3114
rect 144 -3168 586 -3164
rect 639 -3168 757 -3160
rect 144 -3197 602 -3168
rect 639 -3190 667 -3168
rect 699 -3188 757 -3168
rect 787 -3188 845 -3160
rect 852 -3016 2066 -3008
rect 2067 -3016 2083 -3008
rect 2095 -3016 2100 -2962
rect 2108 -2978 2129 -2962
rect 2134 -2970 2141 -2936
rect 2146 -2962 2180 -2936
rect 2234 -2957 2268 -2936
rect 2204 -2962 2268 -2957
rect 2146 -2970 2167 -2962
rect 2204 -2970 2251 -2962
rect 2134 -2978 2167 -2970
rect 2186 -2978 2254 -2970
rect 2108 -2988 2167 -2978
rect 2204 -2980 2254 -2978
rect 2275 -2974 2328 -2936
rect 2275 -2978 2331 -2974
rect 2275 -2980 2328 -2978
rect 2348 -2980 2691 -2924
rect 2108 -2998 2192 -2988
rect 2204 -2998 2691 -2980
rect 2108 -3006 2691 -2998
rect 2108 -3008 2129 -3006
rect 2112 -3016 2129 -3008
rect 2134 -3016 2141 -3006
rect 852 -3020 2141 -3016
rect 852 -3160 2066 -3020
rect 2067 -3044 2083 -3020
rect 2095 -3024 2100 -3020
rect 2112 -3024 2129 -3020
rect 2146 -3029 2691 -3006
rect 2134 -3038 2691 -3029
rect 2112 -3044 2129 -3040
rect 2109 -3046 2129 -3044
rect 2092 -3082 2097 -3066
rect 2088 -3160 2097 -3082
rect 2112 -3081 2129 -3046
rect 2134 -3042 2192 -3038
rect 2195 -3042 2216 -3040
rect 2134 -3044 2216 -3042
rect 2134 -3070 2192 -3044
rect 2217 -3056 2691 -3038
rect 2217 -3070 2303 -3056
rect 2112 -3085 2131 -3081
rect 2140 -3085 2192 -3070
rect 2214 -3072 2303 -3070
rect 2214 -3080 2297 -3072
rect 2214 -3085 2280 -3080
rect 2126 -3086 2131 -3085
rect 2115 -3097 2139 -3086
rect 2146 -3088 2191 -3085
rect 2208 -3086 2280 -3085
rect 2151 -3097 2191 -3088
rect 2203 -3091 2280 -3086
rect 2311 -3091 2691 -3056
rect 2203 -3092 2691 -3091
rect 2203 -3097 2222 -3092
rect 2246 -3097 2280 -3092
rect 2126 -3100 2191 -3097
rect 2208 -3100 2280 -3097
rect 2317 -3100 2691 -3092
rect 2126 -3131 2185 -3100
rect 2192 -3113 2197 -3100
rect 2202 -3113 2260 -3100
rect 2191 -3126 2260 -3113
rect 2283 -3120 2317 -3100
rect 2191 -3131 2317 -3126
rect 2126 -3134 2317 -3131
rect 2126 -3141 2197 -3134
rect 2202 -3141 2260 -3134
rect 2126 -3154 2260 -3141
rect 144 -3202 570 -3197
rect 621 -3202 639 -3190
rect 144 -3219 639 -3202
rect 195 -3235 502 -3219
rect 514 -3235 639 -3219
rect 195 -3236 639 -3235
rect 621 -3242 639 -3236
rect 649 -3242 667 -3190
rect 711 -3192 745 -3188
rect 787 -3202 837 -3188
rect 852 -3190 2109 -3160
rect 2126 -3162 2317 -3154
rect 2126 -3176 2260 -3162
rect 2328 -3176 2691 -3100
rect 2126 -3181 2261 -3176
rect 852 -3202 2097 -3190
rect 2126 -3197 2197 -3181
rect 2202 -3197 2261 -3181
rect 2126 -3202 2185 -3197
rect 2214 -3202 2261 -3197
rect 2291 -3202 2691 -3176
rect 677 -3213 2691 -3202
rect 677 -3221 1513 -3213
rect 1556 -3221 2691 -3213
rect 677 -3226 2691 -3221
rect 693 -3236 2691 -3226
rect 869 -3272 1308 -3236
rect 635 -3308 1308 -3272
rect 1394 -3271 1429 -3236
rect 1432 -3240 1455 -3236
rect 1475 -3252 1482 -3236
rect 1551 -3238 2080 -3236
rect 2088 -3238 2185 -3236
rect 1551 -3242 2066 -3238
rect 1394 -3278 1417 -3271
rect 1489 -3308 1511 -3242
rect 1517 -3268 1539 -3242
rect 1590 -3249 2066 -3242
rect 2092 -3249 2160 -3238
rect 2180 -3242 2185 -3238
rect 2214 -3242 2260 -3236
rect 2180 -3249 2191 -3242
rect 2208 -3249 2260 -3242
rect 1590 -3250 2328 -3249
rect 1551 -3268 1583 -3252
rect 1517 -3302 1583 -3268
rect 1590 -3278 2051 -3250
rect 2092 -3265 2328 -3250
rect 2092 -3270 2139 -3265
rect 1590 -3283 2047 -3278
rect 1517 -3308 1539 -3302
rect 1590 -3308 2046 -3283
rect 2092 -3293 2097 -3270
rect 2109 -3272 2139 -3270
rect 2172 -3270 2214 -3265
rect 2248 -3270 2328 -3265
rect 2172 -3272 2202 -3270
rect 2261 -3272 2291 -3270
rect 2098 -3274 2150 -3272
rect 2161 -3274 2213 -3272
rect 2098 -3278 2242 -3274
rect 2250 -3278 2302 -3272
rect 2098 -3283 2302 -3278
rect 2362 -3283 2691 -3236
rect 2112 -3296 2139 -3283
rect 2172 -3296 2181 -3283
rect 635 -3325 1429 -3308
rect 1434 -3319 2046 -3308
rect 393 -3384 416 -3355
rect 421 -3356 444 -3355
rect 402 -3428 416 -3384
rect 398 -3432 416 -3428
rect 430 -3456 444 -3356
rect 635 -3394 879 -3325
rect 1240 -3376 1241 -3325
rect 1274 -3342 1429 -3325
rect 1445 -3331 1475 -3319
rect 1483 -3331 2046 -3319
rect 1434 -3336 2046 -3331
rect 1434 -3342 1486 -3336
rect 1489 -3346 1511 -3336
rect 1607 -3395 2046 -3336
rect 2154 -3312 2181 -3296
rect 2154 -3317 2220 -3312
rect 2154 -3352 2181 -3317
rect 2261 -3362 2262 -3283
rect 1607 -3431 2029 -3395
rect 2039 -3414 2046 -3395
rect 2328 -3382 2339 -3371
rect 2351 -3382 2362 -3371
rect 2365 -3372 2691 -3283
rect 2734 -2877 2805 -2862
rect 2734 -3336 2804 -2877
rect 3117 -2888 3156 -2852
rect 3472 -2888 3539 -2852
rect 3843 -2862 3906 -2842
rect 3701 -2865 3803 -2862
rect 3824 -2865 3906 -2862
rect 3654 -2871 3803 -2865
rect 3639 -2882 3769 -2871
rect 3770 -2882 3822 -2871
rect 3650 -2884 3769 -2882
rect 3776 -2884 3811 -2882
rect 3843 -2884 3906 -2865
rect 3925 -2845 4025 -2842
rect 4033 -2845 4099 -2833
rect 3925 -2856 4110 -2845
rect 3925 -2866 4025 -2856
rect 4083 -2862 4095 -2856
rect 3910 -2870 4025 -2866
rect 3925 -2884 4025 -2870
rect 4033 -2872 4069 -2866
rect 3650 -2890 3945 -2884
rect 3650 -2894 3925 -2890
rect 3639 -2898 3925 -2894
rect 3556 -2905 3925 -2898
rect 3957 -2901 4025 -2884
rect 4111 -2890 4123 -2820
rect 4167 -2856 4204 -2855
rect 4193 -2866 4204 -2856
rect 4207 -2862 4294 -2804
rect 4362 -2822 4394 -2804
rect 4362 -2825 4408 -2822
rect 4362 -2837 4409 -2825
rect 4364 -2859 4394 -2837
rect 4420 -2859 4436 -2837
rect 4222 -2866 4294 -2862
rect 4193 -2896 4294 -2866
rect 4193 -2901 4204 -2896
rect 4222 -2901 4294 -2896
rect 3654 -2911 3712 -2905
rect 3723 -2930 3752 -2905
rect 3823 -2924 3925 -2905
rect 3943 -2918 4025 -2901
rect 4069 -2918 4294 -2901
rect 4306 -2915 4328 -2882
rect 3943 -2924 4294 -2918
rect 2916 -2945 2974 -2939
rect 2916 -2979 2928 -2945
rect 3086 -2968 3120 -2950
rect 3508 -2968 3542 -2950
rect 2916 -2985 2974 -2979
rect 3086 -3004 3156 -2968
rect 3103 -3038 3174 -3004
rect 2916 -3253 2974 -3247
rect 2916 -3287 2928 -3253
rect 2916 -3293 2974 -3287
rect 2734 -3372 2787 -3336
rect 2328 -3414 2362 -3382
rect 2039 -3425 2080 -3414
rect 2250 -3416 2362 -3414
rect 2039 -3437 2069 -3425
rect 2028 -3438 2069 -3437
rect 2111 -3437 2177 -3424
rect 2250 -3425 2291 -3416
rect 2261 -3437 2291 -3425
rect 2351 -3427 2362 -3416
rect 2734 -3406 2945 -3372
rect 3103 -3389 3173 -3038
rect 3285 -3106 3343 -3100
rect 3285 -3140 3297 -3106
rect 3285 -3146 3343 -3140
rect 3285 -3306 3343 -3300
rect 3285 -3340 3297 -3306
rect 3285 -3346 3343 -3340
rect 2734 -3425 2911 -3406
rect 3103 -3425 3156 -3389
rect 2111 -3438 2188 -3437
rect 2028 -3448 2188 -3438
rect 2250 -3448 2302 -3437
rect 3472 -3442 3542 -2968
rect 3723 -3052 3778 -2930
rect 3823 -2958 4294 -2924
rect 4402 -2925 4436 -2859
rect 3823 -3052 3911 -2958
rect 3925 -2969 4281 -2958
rect 3925 -2974 4069 -2969
rect 3925 -3005 4067 -2974
rect 4105 -2981 4109 -2969
rect 4111 -2983 4145 -2969
rect 4157 -2982 4281 -2969
rect 4388 -2977 4514 -2974
rect 4576 -2977 4610 -2804
rect 4629 -2977 4644 -2804
rect 4353 -2982 4456 -2977
rect 4079 -3005 4091 -3001
rect 4111 -3005 4147 -2983
rect 3723 -3063 3756 -3052
rect 3824 -3063 3858 -3052
rect 3877 -3063 3911 -3052
rect 3957 -3047 4147 -3005
rect 4157 -2996 4456 -2982
rect 4457 -2988 4509 -2977
rect 4545 -2980 4644 -2977
rect 4660 -2980 4663 -2804
rect 4686 -2807 5572 -2804
rect 5582 -2807 5589 -2784
rect 4686 -2822 5615 -2807
rect 4686 -2824 5612 -2822
rect 5683 -2824 5717 -2762
rect 5736 -2824 5770 -2756
rect 5838 -2777 5849 -2693
rect 5838 -2792 5853 -2777
rect 5871 -2792 5905 -2693
rect 5908 -2765 6347 -2693
rect 6421 -2647 6455 -2646
rect 6421 -2657 6479 -2647
rect 6421 -2663 6517 -2657
rect 6421 -2697 6479 -2663
rect 6421 -2703 6517 -2697
rect 6421 -2713 6479 -2703
rect 6421 -2765 6455 -2713
rect 5908 -2782 6353 -2765
rect 5938 -2792 5984 -2782
rect 5838 -2824 5905 -2792
rect 4686 -2841 5615 -2824
rect 4686 -2856 5384 -2841
rect 4686 -2878 5192 -2856
rect 5214 -2868 5240 -2856
rect 5242 -2868 5268 -2856
rect 5234 -2878 5246 -2876
rect 4686 -2908 5246 -2878
rect 4686 -2928 5192 -2908
rect 4702 -2942 5032 -2928
rect 4702 -2946 5082 -2942
rect 5100 -2943 5155 -2935
rect 5158 -2936 5182 -2928
rect 4826 -2966 5082 -2946
rect 5116 -2966 5152 -2947
rect 5158 -2965 5186 -2936
rect 5194 -2943 5246 -2908
rect 5280 -2930 5306 -2926
rect 5260 -2943 5306 -2930
rect 4826 -2968 4833 -2966
rect 4945 -2970 4979 -2966
rect 4998 -2970 5032 -2966
rect 4545 -2988 4586 -2980
rect 4468 -2996 4498 -2988
rect 4556 -2996 4586 -2988
rect 4595 -2992 4663 -2980
rect 4629 -2996 4663 -2992
rect 4854 -2994 5054 -2970
rect 5166 -2971 5186 -2965
rect 5144 -2981 5152 -2975
rect 5214 -2976 5244 -2943
rect 5266 -2971 5268 -2943
rect 5156 -2981 5244 -2976
rect 4854 -2996 4861 -2994
rect 4157 -3011 4610 -2996
rect 4157 -3047 4263 -3011
rect 4302 -3045 4336 -3032
rect 3957 -3058 4125 -3047
rect 4157 -3048 4227 -3047
rect 4157 -3058 4261 -3048
rect 3957 -3059 4261 -3058
rect 3957 -3063 4025 -3059
rect 3723 -3064 4025 -3063
rect 3659 -3270 3662 -3126
rect 3698 -3132 3717 -3080
rect 3741 -3132 3756 -3117
rect 3687 -3242 3690 -3154
rect 3698 -3162 3756 -3132
rect 3741 -3164 3756 -3162
rect 3710 -3176 3756 -3164
rect 3824 -3176 3858 -3064
rect 3877 -3132 3911 -3064
rect 3877 -3162 3899 -3132
rect 3957 -3154 3959 -3064
rect 3985 -3154 3987 -3064
rect 4045 -3154 4057 -3059
rect 4069 -3085 4099 -3059
rect 4073 -3097 4091 -3085
rect 4073 -3154 4085 -3097
rect 4202 -3114 4261 -3059
rect 4202 -3125 4227 -3114
rect 4263 -3125 4331 -3047
rect 4510 -3074 4544 -3011
rect 4629 -3064 4644 -2996
rect 4660 -3030 4663 -2996
rect 4716 -3030 4906 -3014
rect 4660 -3041 4701 -3030
rect 4716 -3036 4784 -3030
rect 4785 -3036 4872 -3030
rect 4883 -3036 4906 -3030
rect 4660 -3053 4690 -3041
rect 4716 -3048 4906 -3036
rect 4649 -3064 4701 -3053
rect 4725 -3064 4906 -3048
rect 4964 -3064 4979 -2994
rect 4998 -2998 5054 -2994
rect 5064 -2998 5066 -2994
rect 4998 -3049 5086 -2998
rect 5140 -3014 5244 -2981
rect 5280 -2986 5306 -2943
rect 5140 -3015 5255 -3014
rect 5140 -3031 5198 -3015
rect 5214 -3031 5255 -3015
rect 5266 -3020 5306 -2986
rect 5183 -3046 5198 -3031
rect 5238 -3048 5255 -3031
rect 4998 -3064 5098 -3049
rect 4998 -3098 5013 -3064
rect 5027 -3076 5098 -3064
rect 5152 -3076 5186 -3049
rect 5027 -3083 5086 -3076
rect 5244 -3083 5255 -3048
rect 5027 -3088 5198 -3083
rect 5203 -3088 5255 -3083
rect 5272 -3024 5306 -3020
rect 5314 -2930 5384 -2856
rect 5391 -2862 5401 -2841
rect 5391 -2876 5469 -2862
rect 5391 -2923 5490 -2876
rect 5395 -2930 5490 -2923
rect 5494 -2930 5524 -2841
rect 5536 -2930 5549 -2841
rect 5555 -2848 5615 -2841
rect 5651 -2826 5905 -2824
rect 5926 -2826 5984 -2792
rect 5651 -2847 5834 -2826
rect 5838 -2847 5905 -2826
rect 5651 -2848 5905 -2847
rect 5555 -2858 5905 -2848
rect 5938 -2841 5984 -2826
rect 5938 -2853 5972 -2841
rect 5582 -2862 5615 -2858
rect 5683 -2862 5770 -2858
rect 5582 -2893 5770 -2862
rect 5582 -2930 5612 -2893
rect 5615 -2930 5770 -2893
rect 5314 -3008 5428 -2930
rect 5469 -2941 5615 -2930
rect 5448 -2987 5615 -2941
rect 5618 -2942 5637 -2930
rect 5448 -3008 5482 -2987
rect 5502 -2991 5515 -2987
rect 5527 -2996 5570 -2987
rect 5590 -2991 5603 -2987
rect 5494 -3008 5597 -2996
rect 5314 -3019 5401 -3008
rect 5475 -3019 5482 -3008
rect 5485 -3019 5597 -3008
rect 5618 -3008 5641 -2942
rect 5618 -3015 5637 -3008
rect 5624 -3019 5637 -3015
rect 5649 -3019 5658 -2930
rect 5670 -2934 5770 -2930
rect 5838 -2934 5849 -2858
rect 5938 -2868 5984 -2853
rect 5670 -2948 5849 -2934
rect 5670 -2980 5888 -2948
rect 5892 -2980 5896 -2868
rect 5926 -2900 5984 -2868
rect 5938 -2915 5984 -2900
rect 5938 -2980 5972 -2915
rect 5981 -2960 5984 -2915
rect 6052 -2926 6086 -2782
rect 6105 -2900 6120 -2782
rect 6313 -2799 6353 -2782
rect 6409 -2799 6567 -2765
rect 6646 -2799 6716 -2448
rect 6828 -2516 6886 -2510
rect 6828 -2550 6840 -2516
rect 6828 -2556 6886 -2550
rect 6828 -2716 6886 -2710
rect 6828 -2750 6840 -2716
rect 6828 -2756 6886 -2750
rect 6421 -2855 6455 -2799
rect 6646 -2835 6699 -2799
rect 6682 -2852 6878 -2837
rect 7015 -2852 7085 -2378
rect 7197 -2769 7255 -2763
rect 7197 -2803 7209 -2769
rect 7197 -2809 7255 -2803
rect 6421 -2891 6491 -2855
rect 7015 -2888 7068 -2852
rect 5670 -3002 5914 -2980
rect 5938 -3002 6002 -2980
rect 6028 -2994 6031 -2960
rect 6052 -2994 6096 -2926
rect 5670 -3014 5771 -3002
rect 5670 -3019 5804 -3014
rect 5314 -3020 5804 -3019
rect 5272 -3088 5283 -3024
rect 5314 -3083 5401 -3020
rect 5475 -3024 5482 -3020
rect 5524 -3028 5574 -3020
rect 5513 -3034 5574 -3028
rect 5509 -3058 5575 -3034
rect 5582 -3046 5612 -3020
rect 5624 -3024 5637 -3020
rect 5649 -3024 5658 -3020
rect 5683 -3033 5692 -3020
rect 5702 -3033 5717 -3020
rect 5513 -3068 5574 -3058
rect 5513 -3074 5571 -3068
rect 5331 -3088 5401 -3083
rect 5683 -3087 5717 -3033
rect 5736 -3080 5804 -3020
rect 5838 -3028 6002 -3002
rect 5838 -3033 5980 -3028
rect 5838 -3040 5984 -3033
rect 5846 -3071 5880 -3040
rect 5922 -3064 5926 -3040
rect 5934 -3053 5966 -3049
rect 5886 -3071 5910 -3064
rect 5846 -3080 5910 -3071
rect 5736 -3087 5771 -3080
rect 5878 -3081 5910 -3080
rect 5912 -3071 5928 -3064
rect 5934 -3071 5968 -3053
rect 5912 -3080 5968 -3071
rect 5912 -3081 5944 -3080
rect 5878 -3087 5892 -3081
rect 5922 -3087 5944 -3081
rect 5980 -3087 6048 -3040
rect 6052 -3087 6086 -2994
rect 4202 -3126 4331 -3125
rect 4193 -3154 4204 -3149
rect 4150 -3160 4168 -3154
rect 4178 -3160 4204 -3154
rect 4210 -3160 4263 -3127
rect 4302 -3130 4336 -3129
rect 5027 -3154 5054 -3088
rect 5055 -3154 5082 -3088
rect 5110 -3114 5140 -3088
rect 5203 -3094 5401 -3088
rect 5214 -3106 5401 -3094
rect 5203 -3117 5401 -3106
rect 5244 -3154 5255 -3117
rect 5272 -3154 5283 -3117
rect 5331 -3118 5401 -3117
rect 5331 -3148 5384 -3118
rect 5390 -3129 5401 -3118
rect 5688 -3148 5717 -3087
rect 5331 -3153 5717 -3148
rect 3877 -3176 3911 -3162
rect 4193 -3163 4263 -3160
rect 3710 -3177 3979 -3176
rect 3710 -3202 3744 -3177
rect 3756 -3202 3979 -3177
rect 3991 -3202 4025 -3168
rect 4079 -3202 4113 -3168
rect 4125 -3202 4177 -3176
rect 4193 -3190 4596 -3163
rect 5367 -3170 5717 -3153
rect 5722 -3092 5980 -3087
rect 5722 -3121 5771 -3092
rect 5804 -3118 5834 -3092
rect 5842 -3110 5944 -3092
rect 5842 -3121 5955 -3110
rect 6037 -3121 6086 -3087
rect 5722 -3176 5770 -3121
rect 5854 -3126 5908 -3121
rect 5922 -3126 5944 -3121
rect 5854 -3127 5944 -3126
rect 5854 -3137 5892 -3127
rect 5922 -3137 5944 -3127
rect 5854 -3154 5880 -3137
rect 6038 -3140 6086 -3121
rect 6105 -3140 6139 -2900
rect 6421 -2925 6509 -2891
rect 6789 -2925 6824 -2891
rect 7051 -2905 7247 -2890
rect 7386 -2905 7401 -2232
rect 7420 -2266 7455 -2232
rect 7420 -2905 7454 -2266
rect 7566 -2334 7624 -2328
rect 7566 -2368 7578 -2334
rect 7566 -2374 7624 -2368
rect 7736 -2537 7770 -2519
rect 9580 -2531 9615 -2497
rect 7736 -2573 7806 -2537
rect 9581 -2550 9615 -2531
rect 7753 -2607 7824 -2573
rect 8104 -2607 8139 -2573
rect 7566 -2822 7624 -2816
rect 7566 -2856 7578 -2822
rect 7566 -2862 7624 -2856
rect 6207 -3080 6222 -3065
rect 6232 -3080 6247 -3078
rect 6207 -3093 6247 -3080
rect 6313 -3093 6353 -3086
rect 6205 -3110 6232 -3093
rect 6265 -3110 6274 -3093
rect 6251 -3140 6309 -3134
rect 5854 -3155 5968 -3154
rect 6038 -3160 6049 -3149
rect 6057 -3160 6086 -3140
rect 5331 -3178 5770 -3176
rect 3710 -3235 3782 -3202
rect 3790 -3235 3911 -3202
rect 3957 -3235 4125 -3202
rect 4127 -3235 4147 -3202
rect 4150 -3235 4177 -3202
rect 3710 -3236 4177 -3235
rect 4178 -3197 4562 -3190
rect 4178 -3202 4280 -3197
rect 4585 -3201 4596 -3190
rect 5317 -3189 5770 -3178
rect 5832 -3189 5880 -3168
rect 5914 -3189 5990 -3168
rect 6038 -3176 6086 -3160
rect 6091 -3148 6140 -3140
rect 6091 -3160 6187 -3148
rect 6236 -3151 6324 -3140
rect 6091 -3163 6198 -3160
rect 6091 -3174 6201 -3163
rect 6091 -3176 6139 -3174
rect 6038 -3189 6170 -3176
rect 5317 -3190 6170 -3189
rect 5317 -3202 5756 -3190
rect 5832 -3202 5990 -3190
rect 6038 -3202 6170 -3190
rect 6223 -3202 6232 -3154
rect 6247 -3163 6313 -3151
rect 6236 -3174 6324 -3163
rect 6251 -3180 6309 -3174
rect 6421 -3180 6508 -2925
rect 6790 -2944 6824 -2925
rect 7015 -2941 7229 -2908
rect 7420 -2939 7435 -2905
rect 7753 -2906 7823 -2607
rect 8105 -2626 8139 -2607
rect 7935 -2675 7993 -2669
rect 7935 -2709 7947 -2675
rect 7935 -2715 7993 -2709
rect 7935 -2875 7993 -2869
rect 7935 -2904 7947 -2875
rect 7935 -2906 7969 -2904
rect 7753 -2909 7969 -2906
rect 7753 -2915 7993 -2909
rect 7643 -2942 7674 -2924
rect 6620 -2993 6678 -2987
rect 6620 -3027 6632 -2993
rect 6620 -3033 6678 -3027
rect 6247 -3190 6313 -3184
rect 4178 -3214 4263 -3202
rect 4280 -3214 4562 -3202
rect 5333 -3204 6086 -3202
rect 5415 -3214 5641 -3204
rect 5688 -3214 6086 -3204
rect 4178 -3223 6086 -3214
rect 4178 -3235 5756 -3223
rect 5770 -3235 6072 -3223
rect 6091 -3235 6170 -3202
rect 4178 -3236 6170 -3235
rect 3710 -3274 3744 -3236
rect 3654 -3359 3712 -3353
rect 3654 -3393 3666 -3359
rect 3699 -3393 3712 -3359
rect 3654 -3399 3712 -3393
rect 3727 -3427 3740 -3376
rect 2338 -3448 2362 -3447
rect 398 -3460 444 -3456
rect 1976 -3484 2195 -3452
rect 3472 -3478 3525 -3442
rect 3843 -3495 3858 -3236
rect 3877 -3495 3911 -3236
rect 4150 -3242 4168 -3236
rect 4178 -3242 4280 -3236
rect 4364 -3242 4478 -3236
rect 4196 -3270 4280 -3242
rect 4392 -3265 4450 -3259
rect 4388 -3270 4454 -3265
rect 4023 -3412 4081 -3406
rect 4023 -3446 4035 -3412
rect 4023 -3452 4081 -3446
rect 3877 -3529 3892 -3495
rect 1283 -3556 1325 -3532
rect 4210 -3548 4280 -3270
rect 4392 -3274 4438 -3270
rect 4392 -3299 4404 -3274
rect 4392 -3305 4450 -3299
rect 4392 -3465 4450 -3459
rect 4392 -3499 4404 -3465
rect 4392 -3505 4450 -3499
rect 605 -3626 614 -3572
rect 1311 -3584 1325 -3560
rect 1487 -3570 1525 -3560
rect 659 -3649 668 -3626
rect 1487 -3706 1511 -3570
rect 4210 -3584 4263 -3548
rect 1515 -3598 1553 -3588
rect 1515 -3678 1539 -3598
rect 4581 -3601 4596 -3236
rect 4615 -3250 4650 -3236
rect 4711 -3250 4869 -3236
rect 4930 -3250 4965 -3236
rect 4615 -3601 4649 -3250
rect 4931 -3269 4965 -3250
rect 5317 -3248 5388 -3236
rect 5317 -3269 5387 -3248
rect 4761 -3318 4819 -3312
rect 4761 -3352 4773 -3318
rect 4761 -3358 4819 -3352
rect 4761 -3518 4819 -3512
rect 4761 -3552 4773 -3518
rect 4761 -3558 4819 -3552
rect 4615 -3635 4630 -3601
rect 4950 -3654 4965 -3269
rect 4984 -3270 5387 -3269
rect 4984 -3303 5019 -3270
rect 4984 -3654 5018 -3303
rect 5130 -3371 5188 -3365
rect 5130 -3405 5142 -3371
rect 5130 -3411 5188 -3405
rect 5130 -3571 5188 -3565
rect 5130 -3605 5142 -3571
rect 5130 -3611 5188 -3605
rect 1493 -3744 1511 -3706
rect 1521 -3744 1539 -3678
rect 4984 -3688 4999 -3654
rect 5317 -3707 5387 -3270
rect 5499 -3316 5557 -3310
rect 5499 -3350 5511 -3316
rect 5499 -3356 5557 -3350
rect 5499 -3624 5557 -3618
rect 5499 -3658 5511 -3624
rect 5499 -3664 5557 -3658
rect 5317 -3743 5370 -3707
rect 607 -3750 625 -3744
rect 635 -3750 653 -3744
rect 5688 -3760 5703 -3236
rect 5722 -3760 5756 -3236
rect 5836 -3270 5870 -3266
rect 5924 -3270 5958 -3266
rect 5868 -3677 5926 -3671
rect 5868 -3711 5880 -3677
rect 5868 -3717 5926 -3711
rect 607 -3832 625 -3780
rect 635 -3832 653 -3780
rect 5722 -3794 5737 -3760
rect 6057 -3813 6072 -3236
rect 6091 -3276 6126 -3236
rect 6209 -3242 6232 -3208
rect 6237 -3242 6295 -3236
rect 6222 -3253 6310 -3242
rect 6233 -3265 6299 -3253
rect 6222 -3269 6310 -3265
rect 6139 -3276 6393 -3269
rect 6438 -3276 6508 -3180
rect 6620 -3193 6678 -3187
rect 6620 -3227 6632 -3193
rect 6620 -3233 6678 -3227
rect 6091 -3813 6125 -3276
rect 6237 -3282 6295 -3276
rect 6438 -3329 6495 -3276
rect 6809 -3329 6824 -2944
rect 6843 -2978 6878 -2944
rect 7158 -2978 7193 -2944
rect 7420 -2958 7616 -2943
rect 7677 -2958 7708 -2942
rect 7581 -2961 7616 -2958
rect 6843 -3329 6877 -2978
rect 7159 -2997 7193 -2978
rect 7384 -2976 7616 -2961
rect 7384 -2994 7615 -2976
rect 6989 -3046 7047 -3040
rect 6989 -3080 7001 -3046
rect 6989 -3086 7047 -3080
rect 6989 -3246 7047 -3240
rect 6989 -3280 7001 -3246
rect 6989 -3286 7047 -3280
rect 6438 -3365 6477 -3329
rect 6843 -3363 6858 -3329
rect 7178 -3382 7193 -2997
rect 7212 -3031 7247 -2997
rect 7212 -3382 7246 -3031
rect 7358 -3099 7416 -3093
rect 7358 -3133 7370 -3099
rect 7358 -3139 7416 -3133
rect 7358 -3299 7416 -3293
rect 7358 -3333 7370 -3299
rect 7358 -3339 7416 -3333
rect 7212 -3416 7227 -3382
rect 6407 -3445 6441 -3427
rect 7545 -3435 7615 -2994
rect 7753 -3038 7967 -2915
rect 8124 -3011 8139 -2626
rect 8158 -2660 8193 -2626
rect 8473 -2660 8508 -2626
rect 8896 -2643 8931 -2625
rect 8158 -3011 8192 -2660
rect 8474 -2679 8508 -2660
rect 8860 -2658 8931 -2643
rect 8304 -2728 8362 -2722
rect 8304 -2762 8316 -2728
rect 8304 -2768 8362 -2762
rect 8304 -2928 8362 -2922
rect 8304 -2962 8316 -2928
rect 8304 -2968 8362 -2962
rect 7727 -3044 7967 -3038
rect 7727 -3078 7739 -3044
rect 7753 -3047 7967 -3044
rect 8158 -3045 8173 -3011
rect 8493 -3012 8508 -2679
rect 8527 -2713 8562 -2679
rect 8527 -3012 8561 -2713
rect 8673 -2781 8731 -2775
rect 8673 -2815 8685 -2781
rect 8673 -2821 8731 -2815
rect 8673 -2981 8731 -2975
rect 8673 -3010 8685 -2981
rect 8673 -3012 8707 -3010
rect 8283 -3015 8707 -3012
rect 8283 -3021 8731 -3015
rect 8283 -3049 8705 -3021
rect 7897 -3067 7931 -3049
rect 8158 -3064 8705 -3049
rect 7727 -3084 7785 -3078
rect 7897 -3103 7967 -3067
rect 8283 -3100 8705 -3064
rect 7914 -3137 7985 -3103
rect 7727 -3352 7785 -3346
rect 7727 -3386 7739 -3352
rect 7727 -3392 7785 -3386
rect 6407 -3481 6477 -3445
rect 7545 -3471 7598 -3435
rect 7914 -3478 7984 -3137
rect 8096 -3205 8154 -3199
rect 8096 -3239 8108 -3205
rect 8096 -3245 8154 -3239
rect 8096 -3405 8154 -3399
rect 8096 -3439 8108 -3405
rect 8096 -3445 8154 -3439
rect 6424 -3515 6495 -3481
rect 6775 -3515 6810 -3481
rect 7581 -3488 7984 -3478
rect 6237 -3730 6295 -3724
rect 6237 -3764 6249 -3730
rect 6237 -3770 6295 -3764
rect 6091 -3847 6106 -3813
rect 6424 -3866 6494 -3515
rect 6776 -3534 6810 -3515
rect 6606 -3583 6664 -3577
rect 6606 -3617 6618 -3583
rect 6606 -3623 6664 -3617
rect 6606 -3783 6664 -3777
rect 6606 -3817 6618 -3783
rect 6606 -3823 6664 -3817
rect 6424 -3902 6477 -3866
rect 6795 -3919 6810 -3534
rect 6829 -3568 6864 -3534
rect 7144 -3568 7179 -3534
rect 7567 -3551 7602 -3533
rect 6829 -3919 6863 -3568
rect 7145 -3587 7179 -3568
rect 7531 -3566 7602 -3551
rect 7914 -3541 7971 -3488
rect 8283 -3541 8353 -3100
rect 8491 -3144 8705 -3100
rect 8465 -3150 8705 -3144
rect 8465 -3184 8477 -3150
rect 8491 -3153 8705 -3150
rect 8860 -3117 8930 -2658
rect 9042 -2726 9100 -2720
rect 9042 -2760 9054 -2726
rect 9042 -2766 9100 -2760
rect 9042 -3034 9100 -3028
rect 9042 -3068 9054 -3034
rect 9042 -3074 9100 -3068
rect 8860 -3153 8913 -3117
rect 8860 -3155 8959 -3153
rect 9119 -3154 9150 -3136
rect 9231 -3154 9246 -2624
rect 9265 -3154 9299 -2570
rect 9411 -2599 9469 -2593
rect 9411 -2633 9423 -2599
rect 9411 -2639 9469 -2633
rect 9411 -3087 9469 -3081
rect 9411 -3116 9423 -3087
rect 9411 -3120 9445 -3116
rect 9407 -3121 9445 -3120
rect 9411 -3127 9469 -3121
rect 8635 -3173 8669 -3155
rect 8860 -3170 9092 -3155
rect 9153 -3170 9184 -3154
rect 9299 -3155 9407 -3154
rect 8860 -3173 8959 -3170
rect 9057 -3173 9092 -3170
rect 8465 -3190 8523 -3184
rect 8635 -3209 8705 -3173
rect 8860 -3188 9092 -3173
rect 9299 -3188 9373 -3155
rect 8860 -3206 9091 -3188
rect 8652 -3243 8723 -3209
rect 8465 -3458 8523 -3452
rect 8465 -3492 8477 -3458
rect 8465 -3498 8523 -3492
rect 6975 -3636 7033 -3630
rect 6975 -3670 6987 -3636
rect 6975 -3676 7033 -3670
rect 6975 -3836 7033 -3830
rect 6975 -3870 6987 -3836
rect 6975 -3876 7033 -3870
rect 6829 -3953 6844 -3919
rect 7164 -3972 7179 -3587
rect 7198 -3621 7233 -3587
rect 7198 -3972 7232 -3621
rect 7344 -3689 7402 -3683
rect 7344 -3723 7356 -3689
rect 7344 -3729 7402 -3723
rect 7344 -3889 7402 -3883
rect 7344 -3923 7356 -3889
rect 7344 -3929 7402 -3923
rect 7198 -4006 7213 -3972
rect 7531 -4025 7601 -3566
rect 7914 -3577 7953 -3541
rect 8283 -3577 8336 -3541
rect 8652 -3584 8722 -3243
rect 8834 -3311 8892 -3305
rect 8834 -3345 8846 -3311
rect 8834 -3351 8892 -3345
rect 8834 -3511 8892 -3505
rect 8834 -3545 8846 -3511
rect 8834 -3551 8892 -3545
rect 8319 -3594 8722 -3584
rect 7713 -3634 7771 -3628
rect 7713 -3668 7725 -3634
rect 7883 -3657 7917 -3639
rect 8305 -3657 8340 -3639
rect 7713 -3674 7771 -3668
rect 7883 -3693 7953 -3657
rect 8269 -3672 8340 -3657
rect 8652 -3647 8709 -3594
rect 9021 -3647 9091 -3206
rect 9299 -3216 9373 -3189
rect 9265 -3222 9287 -3218
rect 9299 -3222 9441 -3216
rect 9265 -3223 9299 -3222
rect 9361 -3223 9441 -3222
rect 9600 -3223 9615 -2550
rect 9634 -2584 9669 -2550
rect 9634 -3223 9668 -2584
rect 9780 -2652 9838 -2646
rect 9780 -2686 9792 -2652
rect 9780 -2692 9838 -2686
rect 9950 -2855 9984 -2837
rect 9950 -2891 10020 -2855
rect 9967 -2925 10038 -2891
rect 10318 -2925 10353 -2891
rect 9780 -3140 9838 -3134
rect 9780 -3174 9792 -3140
rect 9780 -3180 9838 -3174
rect 9203 -3256 9261 -3250
rect 9203 -3290 9215 -3256
rect 9249 -3257 9265 -3256
rect 9634 -3257 9649 -3223
rect 9203 -3296 9261 -3290
rect 9598 -3312 9697 -3259
rect 9967 -3276 10037 -2925
rect 10319 -2944 10353 -2925
rect 10149 -2993 10207 -2987
rect 10149 -3027 10161 -2993
rect 10149 -3033 10207 -3027
rect 10149 -3193 10207 -3187
rect 10149 -3227 10161 -3193
rect 10149 -3233 10207 -3227
rect 9967 -3312 10020 -3276
rect 10338 -3329 10353 -2944
rect 10372 -2978 10407 -2944
rect 10687 -2978 10722 -2944
rect 11110 -2961 11145 -2943
rect 10372 -3329 10406 -2978
rect 10688 -2997 10722 -2978
rect 11074 -2976 11145 -2961
rect 10518 -3046 10576 -3040
rect 10518 -3080 10530 -3046
rect 10518 -3086 10576 -3080
rect 10518 -3246 10576 -3240
rect 10518 -3280 10530 -3246
rect 10518 -3286 10576 -3280
rect 10372 -3363 10387 -3329
rect 10707 -3382 10722 -2997
rect 10741 -3031 10776 -2997
rect 10741 -3382 10775 -3031
rect 10887 -3099 10945 -3093
rect 10887 -3133 10899 -3099
rect 10887 -3139 10945 -3133
rect 10887 -3299 10945 -3293
rect 10887 -3333 10899 -3299
rect 10887 -3339 10945 -3333
rect 10741 -3416 10756 -3382
rect 11074 -3435 11144 -2976
rect 11256 -3044 11314 -3038
rect 11256 -3078 11268 -3044
rect 11426 -3067 11460 -3049
rect 11848 -3067 11883 -3049
rect 11256 -3084 11314 -3078
rect 11426 -3103 11496 -3067
rect 11812 -3082 11883 -3067
rect 11443 -3137 11514 -3103
rect 11256 -3352 11314 -3346
rect 11256 -3386 11268 -3352
rect 11256 -3392 11314 -3386
rect 11074 -3471 11127 -3435
rect 11443 -3488 11513 -3137
rect 11625 -3205 11683 -3199
rect 11625 -3239 11637 -3205
rect 11625 -3245 11683 -3239
rect 11625 -3405 11683 -3399
rect 11625 -3439 11637 -3405
rect 11625 -3445 11683 -3439
rect 11443 -3524 11496 -3488
rect 11812 -3541 11882 -3082
rect 11994 -3150 12052 -3144
rect 11994 -3184 12006 -3150
rect 12164 -3173 12198 -3155
rect 12586 -3173 12621 -3155
rect 11994 -3190 12052 -3184
rect 12164 -3209 12234 -3173
rect 12550 -3188 12621 -3173
rect 12181 -3243 12252 -3209
rect 11994 -3458 12052 -3452
rect 11994 -3492 12006 -3458
rect 11994 -3498 12052 -3492
rect 9203 -3564 9261 -3558
rect 9203 -3598 9215 -3564
rect 11812 -3577 11865 -3541
rect 12181 -3594 12251 -3243
rect 12363 -3311 12421 -3305
rect 12363 -3345 12375 -3311
rect 12363 -3351 12421 -3345
rect 12363 -3511 12421 -3505
rect 12363 -3545 12375 -3511
rect 12363 -3551 12421 -3545
rect 9203 -3604 9261 -3598
rect 12181 -3630 12234 -3594
rect 12550 -3647 12620 -3188
rect 12732 -3256 12790 -3250
rect 12732 -3290 12744 -3256
rect 12732 -3296 12790 -3290
rect 12732 -3564 12790 -3558
rect 12732 -3598 12744 -3564
rect 12732 -3604 12790 -3598
rect 7900 -3727 7971 -3693
rect 7713 -3942 7771 -3936
rect 7713 -3976 7725 -3942
rect 7713 -3982 7771 -3976
rect 7531 -4061 7584 -4025
rect 7900 -4078 7970 -3727
rect 8082 -3795 8140 -3789
rect 8082 -3829 8094 -3795
rect 8082 -3835 8140 -3829
rect 8082 -3995 8140 -3989
rect 8082 -4029 8094 -3995
rect 8082 -4035 8140 -4029
rect 7900 -4114 7953 -4078
rect 8269 -4131 8339 -3672
rect 8652 -3683 8691 -3647
rect 9021 -3683 9074 -3647
rect 12550 -3683 12603 -3647
rect 9057 -3700 9407 -3690
rect 8451 -3740 8509 -3734
rect 8451 -3774 8463 -3740
rect 8621 -3763 8655 -3745
rect 9043 -3763 9078 -3745
rect 8451 -3780 8509 -3774
rect 8621 -3799 8691 -3763
rect 9007 -3778 9078 -3763
rect 8638 -3833 8709 -3799
rect 8451 -4048 8509 -4042
rect 8451 -4082 8463 -4048
rect 8451 -4088 8509 -4082
rect 358 -4166 384 -4148
rect 1311 -4160 1511 -4142
rect 8269 -4167 8322 -4131
rect 358 -4194 398 -4176
rect 1325 -4188 1525 -4170
rect 8638 -4184 8708 -3833
rect 8820 -3901 8878 -3895
rect 8820 -3935 8832 -3901
rect 8820 -3941 8878 -3935
rect 8820 -4101 8878 -4095
rect 8820 -4135 8832 -4101
rect 8820 -4141 8878 -4135
rect 8638 -4220 8691 -4184
rect 9007 -4237 9077 -3778
rect 9189 -3846 9247 -3840
rect 9189 -3880 9201 -3846
rect 9189 -3886 9247 -3880
rect 9189 -4154 9247 -4148
rect 9189 -4188 9201 -4154
rect 9189 -4194 9247 -4188
rect 9007 -4273 9060 -4237
rect 158 -4350 198 -4338
rect 184 -4378 198 -4366
rect 184 -4566 384 -4548
rect 1311 -4560 1511 -4542
rect 198 -4594 398 -4576
rect 1325 -4588 1525 -4570
rect 184 -4966 384 -4948
rect 1311 -4960 1511 -4942
rect 198 -4994 398 -4976
rect 1325 -4988 1525 -4970
<< nwell >>
rect 3696 2214 3718 2312
rect 3638 76 3662 174
rect 3652 -2270 3676 -2160
<< poly >>
rect 6 2346 26 2370
rect 78 2346 98 2370
rect 3694 2346 3716 2370
rect 3694 2344 3714 2346
rect 3694 -2062 3714 -2018
<< metal1 >>
rect -120 2168 220 2370
rect 3696 2214 3718 2312
rect -120 274 80 2168
rect 3772 1402 3972 2370
rect 3734 1276 3972 1402
rect 3716 1176 3972 1276
rect 3734 1040 3972 1176
rect -120 -176 260 274
rect 3638 76 3662 174
rect -120 -200 80 -176
rect -120 -400 200 -200
rect -120 -600 80 -400
rect -120 -800 200 -600
rect -120 -1000 80 -800
rect 3772 -944 3972 1040
rect -120 -1200 200 -1000
rect 3738 -1058 3972 -944
rect 3714 -1160 3972 -1058
rect -120 -1400 80 -1200
rect 3738 -1306 3972 -1160
rect -120 -1600 200 -1400
rect -120 -1800 80 -1600
rect -120 -2000 200 -1800
rect -120 -2070 80 -2000
rect -120 -2346 222 -2070
rect 3652 -2270 3676 -2160
rect 3772 -2346 3972 -1306
rect 0 -2400 200 -2346
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
<< metal2 >>
rect 3102 1558 3158 1614
rect 3102 828 3158 884
rect 3102 -788 3158 -732
rect 3102 -1518 3158 -1462
use c2b  c2b_0
timestamp 1624053917
transform 1 0 158 0 1 1196
box -158 -5010 13287 5060
use c2b  c2b_1
timestamp 1624053917
transform 1 0 158 0 1 -1150
box -158 -5010 13287 5060
use c2b  x1
timestamp 1624053917
transform 1 0 158 0 1 1796
box -158 -5010 13287 5060
use c2b  x2
timestamp 1624053917
transform 1 0 3902 0 1 1796
box -158 -5010 13287 5060
<< labels >>
rlabel poly 6 2346 26 2370 1 clr
rlabel poly 78 2346 98 2370 1 clk
rlabel poly 3694 2344 3714 2368 1 ce
rlabel metal2 3102 1558 3158 1614 1 b0
rlabel metal2 3102 828 3158 884 1 b1
rlabel metal2 3102 -788 3158 -732 1 b2
rlabel metal2 3102 -1518 3158 -1462 1 b3
rlabel metal1 -96 2302 -28 2348 1 vdd
rlabel metal1 3812 2272 3928 2344 1 vss
rlabel poly 3694 -2062 3714 -2018 1 out
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 ce
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 clr
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 b0
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 b1
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 b2
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 b3
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 out
port 10 nsew
<< end >>
