magic
tech sky130A
magscale 1 2
timestamp 1615997521
<< nwell >>
rect -3517 -919 3517 919
<< pmoslvt >>
rect -3321 -700 -3111 700
rect -3053 -700 -2843 700
rect -2785 -700 -2575 700
rect -2517 -700 -2307 700
rect -2249 -700 -2039 700
rect -1981 -700 -1771 700
rect -1713 -700 -1503 700
rect -1445 -700 -1235 700
rect -1177 -700 -967 700
rect -909 -700 -699 700
rect -641 -700 -431 700
rect -373 -700 -163 700
rect -105 -700 105 700
rect 163 -700 373 700
rect 431 -700 641 700
rect 699 -700 909 700
rect 967 -700 1177 700
rect 1235 -700 1445 700
rect 1503 -700 1713 700
rect 1771 -700 1981 700
rect 2039 -700 2249 700
rect 2307 -700 2517 700
rect 2575 -700 2785 700
rect 2843 -700 3053 700
rect 3111 -700 3321 700
<< pdiff >>
rect -3379 688 -3321 700
rect -3379 -688 -3367 688
rect -3333 -688 -3321 688
rect -3379 -700 -3321 -688
rect -3111 688 -3053 700
rect -3111 -688 -3099 688
rect -3065 -688 -3053 688
rect -3111 -700 -3053 -688
rect -2843 688 -2785 700
rect -2843 -688 -2831 688
rect -2797 -688 -2785 688
rect -2843 -700 -2785 -688
rect -2575 688 -2517 700
rect -2575 -688 -2563 688
rect -2529 -688 -2517 688
rect -2575 -700 -2517 -688
rect -2307 688 -2249 700
rect -2307 -688 -2295 688
rect -2261 -688 -2249 688
rect -2307 -700 -2249 -688
rect -2039 688 -1981 700
rect -2039 -688 -2027 688
rect -1993 -688 -1981 688
rect -2039 -700 -1981 -688
rect -1771 688 -1713 700
rect -1771 -688 -1759 688
rect -1725 -688 -1713 688
rect -1771 -700 -1713 -688
rect -1503 688 -1445 700
rect -1503 -688 -1491 688
rect -1457 -688 -1445 688
rect -1503 -700 -1445 -688
rect -1235 688 -1177 700
rect -1235 -688 -1223 688
rect -1189 -688 -1177 688
rect -1235 -700 -1177 -688
rect -967 688 -909 700
rect -967 -688 -955 688
rect -921 -688 -909 688
rect -967 -700 -909 -688
rect -699 688 -641 700
rect -699 -688 -687 688
rect -653 -688 -641 688
rect -699 -700 -641 -688
rect -431 688 -373 700
rect -431 -688 -419 688
rect -385 -688 -373 688
rect -431 -700 -373 -688
rect -163 688 -105 700
rect -163 -688 -151 688
rect -117 -688 -105 688
rect -163 -700 -105 -688
rect 105 688 163 700
rect 105 -688 117 688
rect 151 -688 163 688
rect 105 -700 163 -688
rect 373 688 431 700
rect 373 -688 385 688
rect 419 -688 431 688
rect 373 -700 431 -688
rect 641 688 699 700
rect 641 -688 653 688
rect 687 -688 699 688
rect 641 -700 699 -688
rect 909 688 967 700
rect 909 -688 921 688
rect 955 -688 967 688
rect 909 -700 967 -688
rect 1177 688 1235 700
rect 1177 -688 1189 688
rect 1223 -688 1235 688
rect 1177 -700 1235 -688
rect 1445 688 1503 700
rect 1445 -688 1457 688
rect 1491 -688 1503 688
rect 1445 -700 1503 -688
rect 1713 688 1771 700
rect 1713 -688 1725 688
rect 1759 -688 1771 688
rect 1713 -700 1771 -688
rect 1981 688 2039 700
rect 1981 -688 1993 688
rect 2027 -688 2039 688
rect 1981 -700 2039 -688
rect 2249 688 2307 700
rect 2249 -688 2261 688
rect 2295 -688 2307 688
rect 2249 -700 2307 -688
rect 2517 688 2575 700
rect 2517 -688 2529 688
rect 2563 -688 2575 688
rect 2517 -700 2575 -688
rect 2785 688 2843 700
rect 2785 -688 2797 688
rect 2831 -688 2843 688
rect 2785 -700 2843 -688
rect 3053 688 3111 700
rect 3053 -688 3065 688
rect 3099 -688 3111 688
rect 3053 -700 3111 -688
rect 3321 688 3379 700
rect 3321 -688 3333 688
rect 3367 -688 3379 688
rect 3321 -700 3379 -688
<< pdiffc >>
rect -3367 -688 -3333 688
rect -3099 -688 -3065 688
rect -2831 -688 -2797 688
rect -2563 -688 -2529 688
rect -2295 -688 -2261 688
rect -2027 -688 -1993 688
rect -1759 -688 -1725 688
rect -1491 -688 -1457 688
rect -1223 -688 -1189 688
rect -955 -688 -921 688
rect -687 -688 -653 688
rect -419 -688 -385 688
rect -151 -688 -117 688
rect 117 -688 151 688
rect 385 -688 419 688
rect 653 -688 687 688
rect 921 -688 955 688
rect 1189 -688 1223 688
rect 1457 -688 1491 688
rect 1725 -688 1759 688
rect 1993 -688 2027 688
rect 2261 -688 2295 688
rect 2529 -688 2563 688
rect 2797 -688 2831 688
rect 3065 -688 3099 688
rect 3333 -688 3367 688
<< nsubdiff >>
rect -3481 849 -3385 883
rect 3385 849 3481 883
rect -3481 787 -3447 849
rect 3447 787 3481 849
rect -3481 -849 -3447 -787
rect 3447 -849 3481 -787
rect -3481 -883 -3385 -849
rect 3385 -883 3481 -849
<< nsubdiffcont >>
rect -3385 849 3385 883
rect -3481 -787 -3447 787
rect 3447 -787 3481 787
rect -3385 -883 3385 -849
<< poly >>
rect -3321 781 -3111 797
rect -3321 747 -3305 781
rect -3127 747 -3111 781
rect -3321 700 -3111 747
rect -3053 781 -2843 797
rect -3053 747 -3037 781
rect -2859 747 -2843 781
rect -3053 700 -2843 747
rect -2785 781 -2575 797
rect -2785 747 -2769 781
rect -2591 747 -2575 781
rect -2785 700 -2575 747
rect -2517 781 -2307 797
rect -2517 747 -2501 781
rect -2323 747 -2307 781
rect -2517 700 -2307 747
rect -2249 781 -2039 797
rect -2249 747 -2233 781
rect -2055 747 -2039 781
rect -2249 700 -2039 747
rect -1981 781 -1771 797
rect -1981 747 -1965 781
rect -1787 747 -1771 781
rect -1981 700 -1771 747
rect -1713 781 -1503 797
rect -1713 747 -1697 781
rect -1519 747 -1503 781
rect -1713 700 -1503 747
rect -1445 781 -1235 797
rect -1445 747 -1429 781
rect -1251 747 -1235 781
rect -1445 700 -1235 747
rect -1177 781 -967 797
rect -1177 747 -1161 781
rect -983 747 -967 781
rect -1177 700 -967 747
rect -909 781 -699 797
rect -909 747 -893 781
rect -715 747 -699 781
rect -909 700 -699 747
rect -641 781 -431 797
rect -641 747 -625 781
rect -447 747 -431 781
rect -641 700 -431 747
rect -373 781 -163 797
rect -373 747 -357 781
rect -179 747 -163 781
rect -373 700 -163 747
rect -105 781 105 797
rect -105 747 -89 781
rect 89 747 105 781
rect -105 700 105 747
rect 163 781 373 797
rect 163 747 179 781
rect 357 747 373 781
rect 163 700 373 747
rect 431 781 641 797
rect 431 747 447 781
rect 625 747 641 781
rect 431 700 641 747
rect 699 781 909 797
rect 699 747 715 781
rect 893 747 909 781
rect 699 700 909 747
rect 967 781 1177 797
rect 967 747 983 781
rect 1161 747 1177 781
rect 967 700 1177 747
rect 1235 781 1445 797
rect 1235 747 1251 781
rect 1429 747 1445 781
rect 1235 700 1445 747
rect 1503 781 1713 797
rect 1503 747 1519 781
rect 1697 747 1713 781
rect 1503 700 1713 747
rect 1771 781 1981 797
rect 1771 747 1787 781
rect 1965 747 1981 781
rect 1771 700 1981 747
rect 2039 781 2249 797
rect 2039 747 2055 781
rect 2233 747 2249 781
rect 2039 700 2249 747
rect 2307 781 2517 797
rect 2307 747 2323 781
rect 2501 747 2517 781
rect 2307 700 2517 747
rect 2575 781 2785 797
rect 2575 747 2591 781
rect 2769 747 2785 781
rect 2575 700 2785 747
rect 2843 781 3053 797
rect 2843 747 2859 781
rect 3037 747 3053 781
rect 2843 700 3053 747
rect 3111 781 3321 797
rect 3111 747 3127 781
rect 3305 747 3321 781
rect 3111 700 3321 747
rect -3321 -747 -3111 -700
rect -3321 -781 -3305 -747
rect -3127 -781 -3111 -747
rect -3321 -797 -3111 -781
rect -3053 -747 -2843 -700
rect -3053 -781 -3037 -747
rect -2859 -781 -2843 -747
rect -3053 -797 -2843 -781
rect -2785 -747 -2575 -700
rect -2785 -781 -2769 -747
rect -2591 -781 -2575 -747
rect -2785 -797 -2575 -781
rect -2517 -747 -2307 -700
rect -2517 -781 -2501 -747
rect -2323 -781 -2307 -747
rect -2517 -797 -2307 -781
rect -2249 -747 -2039 -700
rect -2249 -781 -2233 -747
rect -2055 -781 -2039 -747
rect -2249 -797 -2039 -781
rect -1981 -747 -1771 -700
rect -1981 -781 -1965 -747
rect -1787 -781 -1771 -747
rect -1981 -797 -1771 -781
rect -1713 -747 -1503 -700
rect -1713 -781 -1697 -747
rect -1519 -781 -1503 -747
rect -1713 -797 -1503 -781
rect -1445 -747 -1235 -700
rect -1445 -781 -1429 -747
rect -1251 -781 -1235 -747
rect -1445 -797 -1235 -781
rect -1177 -747 -967 -700
rect -1177 -781 -1161 -747
rect -983 -781 -967 -747
rect -1177 -797 -967 -781
rect -909 -747 -699 -700
rect -909 -781 -893 -747
rect -715 -781 -699 -747
rect -909 -797 -699 -781
rect -641 -747 -431 -700
rect -641 -781 -625 -747
rect -447 -781 -431 -747
rect -641 -797 -431 -781
rect -373 -747 -163 -700
rect -373 -781 -357 -747
rect -179 -781 -163 -747
rect -373 -797 -163 -781
rect -105 -747 105 -700
rect -105 -781 -89 -747
rect 89 -781 105 -747
rect -105 -797 105 -781
rect 163 -747 373 -700
rect 163 -781 179 -747
rect 357 -781 373 -747
rect 163 -797 373 -781
rect 431 -747 641 -700
rect 431 -781 447 -747
rect 625 -781 641 -747
rect 431 -797 641 -781
rect 699 -747 909 -700
rect 699 -781 715 -747
rect 893 -781 909 -747
rect 699 -797 909 -781
rect 967 -747 1177 -700
rect 967 -781 983 -747
rect 1161 -781 1177 -747
rect 967 -797 1177 -781
rect 1235 -747 1445 -700
rect 1235 -781 1251 -747
rect 1429 -781 1445 -747
rect 1235 -797 1445 -781
rect 1503 -747 1713 -700
rect 1503 -781 1519 -747
rect 1697 -781 1713 -747
rect 1503 -797 1713 -781
rect 1771 -747 1981 -700
rect 1771 -781 1787 -747
rect 1965 -781 1981 -747
rect 1771 -797 1981 -781
rect 2039 -747 2249 -700
rect 2039 -781 2055 -747
rect 2233 -781 2249 -747
rect 2039 -797 2249 -781
rect 2307 -747 2517 -700
rect 2307 -781 2323 -747
rect 2501 -781 2517 -747
rect 2307 -797 2517 -781
rect 2575 -747 2785 -700
rect 2575 -781 2591 -747
rect 2769 -781 2785 -747
rect 2575 -797 2785 -781
rect 2843 -747 3053 -700
rect 2843 -781 2859 -747
rect 3037 -781 3053 -747
rect 2843 -797 3053 -781
rect 3111 -747 3321 -700
rect 3111 -781 3127 -747
rect 3305 -781 3321 -747
rect 3111 -797 3321 -781
<< polycont >>
rect -3305 747 -3127 781
rect -3037 747 -2859 781
rect -2769 747 -2591 781
rect -2501 747 -2323 781
rect -2233 747 -2055 781
rect -1965 747 -1787 781
rect -1697 747 -1519 781
rect -1429 747 -1251 781
rect -1161 747 -983 781
rect -893 747 -715 781
rect -625 747 -447 781
rect -357 747 -179 781
rect -89 747 89 781
rect 179 747 357 781
rect 447 747 625 781
rect 715 747 893 781
rect 983 747 1161 781
rect 1251 747 1429 781
rect 1519 747 1697 781
rect 1787 747 1965 781
rect 2055 747 2233 781
rect 2323 747 2501 781
rect 2591 747 2769 781
rect 2859 747 3037 781
rect 3127 747 3305 781
rect -3305 -781 -3127 -747
rect -3037 -781 -2859 -747
rect -2769 -781 -2591 -747
rect -2501 -781 -2323 -747
rect -2233 -781 -2055 -747
rect -1965 -781 -1787 -747
rect -1697 -781 -1519 -747
rect -1429 -781 -1251 -747
rect -1161 -781 -983 -747
rect -893 -781 -715 -747
rect -625 -781 -447 -747
rect -357 -781 -179 -747
rect -89 -781 89 -747
rect 179 -781 357 -747
rect 447 -781 625 -747
rect 715 -781 893 -747
rect 983 -781 1161 -747
rect 1251 -781 1429 -747
rect 1519 -781 1697 -747
rect 1787 -781 1965 -747
rect 2055 -781 2233 -747
rect 2323 -781 2501 -747
rect 2591 -781 2769 -747
rect 2859 -781 3037 -747
rect 3127 -781 3305 -747
<< locali >>
rect -3481 849 -3385 883
rect 3385 849 3481 883
rect -3481 787 -3447 849
rect 3447 787 3481 849
rect -3321 747 -3305 781
rect -3127 747 -3111 781
rect -3053 747 -3037 781
rect -2859 747 -2843 781
rect -2785 747 -2769 781
rect -2591 747 -2575 781
rect -2517 747 -2501 781
rect -2323 747 -2307 781
rect -2249 747 -2233 781
rect -2055 747 -2039 781
rect -1981 747 -1965 781
rect -1787 747 -1771 781
rect -1713 747 -1697 781
rect -1519 747 -1503 781
rect -1445 747 -1429 781
rect -1251 747 -1235 781
rect -1177 747 -1161 781
rect -983 747 -967 781
rect -909 747 -893 781
rect -715 747 -699 781
rect -641 747 -625 781
rect -447 747 -431 781
rect -373 747 -357 781
rect -179 747 -163 781
rect -105 747 -89 781
rect 89 747 105 781
rect 163 747 179 781
rect 357 747 373 781
rect 431 747 447 781
rect 625 747 641 781
rect 699 747 715 781
rect 893 747 909 781
rect 967 747 983 781
rect 1161 747 1177 781
rect 1235 747 1251 781
rect 1429 747 1445 781
rect 1503 747 1519 781
rect 1697 747 1713 781
rect 1771 747 1787 781
rect 1965 747 1981 781
rect 2039 747 2055 781
rect 2233 747 2249 781
rect 2307 747 2323 781
rect 2501 747 2517 781
rect 2575 747 2591 781
rect 2769 747 2785 781
rect 2843 747 2859 781
rect 3037 747 3053 781
rect 3111 747 3127 781
rect 3305 747 3321 781
rect -3367 688 -3333 704
rect -3367 -704 -3333 -688
rect -3099 688 -3065 704
rect -3099 -704 -3065 -688
rect -2831 688 -2797 704
rect -2831 -704 -2797 -688
rect -2563 688 -2529 704
rect -2563 -704 -2529 -688
rect -2295 688 -2261 704
rect -2295 -704 -2261 -688
rect -2027 688 -1993 704
rect -2027 -704 -1993 -688
rect -1759 688 -1725 704
rect -1759 -704 -1725 -688
rect -1491 688 -1457 704
rect -1491 -704 -1457 -688
rect -1223 688 -1189 704
rect -1223 -704 -1189 -688
rect -955 688 -921 704
rect -955 -704 -921 -688
rect -687 688 -653 704
rect -687 -704 -653 -688
rect -419 688 -385 704
rect -419 -704 -385 -688
rect -151 688 -117 704
rect -151 -704 -117 -688
rect 117 688 151 704
rect 117 -704 151 -688
rect 385 688 419 704
rect 385 -704 419 -688
rect 653 688 687 704
rect 653 -704 687 -688
rect 921 688 955 704
rect 921 -704 955 -688
rect 1189 688 1223 704
rect 1189 -704 1223 -688
rect 1457 688 1491 704
rect 1457 -704 1491 -688
rect 1725 688 1759 704
rect 1725 -704 1759 -688
rect 1993 688 2027 704
rect 1993 -704 2027 -688
rect 2261 688 2295 704
rect 2261 -704 2295 -688
rect 2529 688 2563 704
rect 2529 -704 2563 -688
rect 2797 688 2831 704
rect 2797 -704 2831 -688
rect 3065 688 3099 704
rect 3065 -704 3099 -688
rect 3333 688 3367 704
rect 3333 -704 3367 -688
rect -3321 -781 -3305 -747
rect -3127 -781 -3111 -747
rect -3053 -781 -3037 -747
rect -2859 -781 -2843 -747
rect -2785 -781 -2769 -747
rect -2591 -781 -2575 -747
rect -2517 -781 -2501 -747
rect -2323 -781 -2307 -747
rect -2249 -781 -2233 -747
rect -2055 -781 -2039 -747
rect -1981 -781 -1965 -747
rect -1787 -781 -1771 -747
rect -1713 -781 -1697 -747
rect -1519 -781 -1503 -747
rect -1445 -781 -1429 -747
rect -1251 -781 -1235 -747
rect -1177 -781 -1161 -747
rect -983 -781 -967 -747
rect -909 -781 -893 -747
rect -715 -781 -699 -747
rect -641 -781 -625 -747
rect -447 -781 -431 -747
rect -373 -781 -357 -747
rect -179 -781 -163 -747
rect -105 -781 -89 -747
rect 89 -781 105 -747
rect 163 -781 179 -747
rect 357 -781 373 -747
rect 431 -781 447 -747
rect 625 -781 641 -747
rect 699 -781 715 -747
rect 893 -781 909 -747
rect 967 -781 983 -747
rect 1161 -781 1177 -747
rect 1235 -781 1251 -747
rect 1429 -781 1445 -747
rect 1503 -781 1519 -747
rect 1697 -781 1713 -747
rect 1771 -781 1787 -747
rect 1965 -781 1981 -747
rect 2039 -781 2055 -747
rect 2233 -781 2249 -747
rect 2307 -781 2323 -747
rect 2501 -781 2517 -747
rect 2575 -781 2591 -747
rect 2769 -781 2785 -747
rect 2843 -781 2859 -747
rect 3037 -781 3053 -747
rect 3111 -781 3127 -747
rect 3305 -781 3321 -747
rect -3481 -849 -3447 -787
rect 3447 -849 3481 -787
rect -3481 -883 -3385 -849
rect 3385 -883 3481 -849
<< viali >>
rect -3305 747 -3127 781
rect -3037 747 -2859 781
rect -2769 747 -2591 781
rect -2501 747 -2323 781
rect -2233 747 -2055 781
rect -1965 747 -1787 781
rect -1697 747 -1519 781
rect -1429 747 -1251 781
rect -1161 747 -983 781
rect -893 747 -715 781
rect -625 747 -447 781
rect -357 747 -179 781
rect -89 747 89 781
rect 179 747 357 781
rect 447 747 625 781
rect 715 747 893 781
rect 983 747 1161 781
rect 1251 747 1429 781
rect 1519 747 1697 781
rect 1787 747 1965 781
rect 2055 747 2233 781
rect 2323 747 2501 781
rect 2591 747 2769 781
rect 2859 747 3037 781
rect 3127 747 3305 781
rect -3367 -688 -3333 688
rect -3099 -688 -3065 688
rect -2831 -688 -2797 688
rect -2563 -688 -2529 688
rect -2295 -688 -2261 688
rect -2027 -688 -1993 688
rect -1759 -688 -1725 688
rect -1491 -688 -1457 688
rect -1223 -688 -1189 688
rect -955 -688 -921 688
rect -687 -688 -653 688
rect -419 -688 -385 688
rect -151 -688 -117 688
rect 117 -688 151 688
rect 385 -688 419 688
rect 653 -688 687 688
rect 921 -688 955 688
rect 1189 -688 1223 688
rect 1457 -688 1491 688
rect 1725 -688 1759 688
rect 1993 -688 2027 688
rect 2261 -688 2295 688
rect 2529 -688 2563 688
rect 2797 -688 2831 688
rect 3065 -688 3099 688
rect 3333 -688 3367 688
rect -3305 -781 -3127 -747
rect -3037 -781 -2859 -747
rect -2769 -781 -2591 -747
rect -2501 -781 -2323 -747
rect -2233 -781 -2055 -747
rect -1965 -781 -1787 -747
rect -1697 -781 -1519 -747
rect -1429 -781 -1251 -747
rect -1161 -781 -983 -747
rect -893 -781 -715 -747
rect -625 -781 -447 -747
rect -357 -781 -179 -747
rect -89 -781 89 -747
rect 179 -781 357 -747
rect 447 -781 625 -747
rect 715 -781 893 -747
rect 983 -781 1161 -747
rect 1251 -781 1429 -747
rect 1519 -781 1697 -747
rect 1787 -781 1965 -747
rect 2055 -781 2233 -747
rect 2323 -781 2501 -747
rect 2591 -781 2769 -747
rect 2859 -781 3037 -747
rect 3127 -781 3305 -747
<< metal1 >>
rect -3317 781 -3115 787
rect -3317 747 -3305 781
rect -3127 747 -3115 781
rect -3317 741 -3115 747
rect -3049 781 -2847 787
rect -3049 747 -3037 781
rect -2859 747 -2847 781
rect -3049 741 -2847 747
rect -2781 781 -2579 787
rect -2781 747 -2769 781
rect -2591 747 -2579 781
rect -2781 741 -2579 747
rect -2513 781 -2311 787
rect -2513 747 -2501 781
rect -2323 747 -2311 781
rect -2513 741 -2311 747
rect -2245 781 -2043 787
rect -2245 747 -2233 781
rect -2055 747 -2043 781
rect -2245 741 -2043 747
rect -1977 781 -1775 787
rect -1977 747 -1965 781
rect -1787 747 -1775 781
rect -1977 741 -1775 747
rect -1709 781 -1507 787
rect -1709 747 -1697 781
rect -1519 747 -1507 781
rect -1709 741 -1507 747
rect -1441 781 -1239 787
rect -1441 747 -1429 781
rect -1251 747 -1239 781
rect -1441 741 -1239 747
rect -1173 781 -971 787
rect -1173 747 -1161 781
rect -983 747 -971 781
rect -1173 741 -971 747
rect -905 781 -703 787
rect -905 747 -893 781
rect -715 747 -703 781
rect -905 741 -703 747
rect -637 781 -435 787
rect -637 747 -625 781
rect -447 747 -435 781
rect -637 741 -435 747
rect -369 781 -167 787
rect -369 747 -357 781
rect -179 747 -167 781
rect -369 741 -167 747
rect -101 781 101 787
rect -101 747 -89 781
rect 89 747 101 781
rect -101 741 101 747
rect 167 781 369 787
rect 167 747 179 781
rect 357 747 369 781
rect 167 741 369 747
rect 435 781 637 787
rect 435 747 447 781
rect 625 747 637 781
rect 435 741 637 747
rect 703 781 905 787
rect 703 747 715 781
rect 893 747 905 781
rect 703 741 905 747
rect 971 781 1173 787
rect 971 747 983 781
rect 1161 747 1173 781
rect 971 741 1173 747
rect 1239 781 1441 787
rect 1239 747 1251 781
rect 1429 747 1441 781
rect 1239 741 1441 747
rect 1507 781 1709 787
rect 1507 747 1519 781
rect 1697 747 1709 781
rect 1507 741 1709 747
rect 1775 781 1977 787
rect 1775 747 1787 781
rect 1965 747 1977 781
rect 1775 741 1977 747
rect 2043 781 2245 787
rect 2043 747 2055 781
rect 2233 747 2245 781
rect 2043 741 2245 747
rect 2311 781 2513 787
rect 2311 747 2323 781
rect 2501 747 2513 781
rect 2311 741 2513 747
rect 2579 781 2781 787
rect 2579 747 2591 781
rect 2769 747 2781 781
rect 2579 741 2781 747
rect 2847 781 3049 787
rect 2847 747 2859 781
rect 3037 747 3049 781
rect 2847 741 3049 747
rect 3115 781 3317 787
rect 3115 747 3127 781
rect 3305 747 3317 781
rect 3115 741 3317 747
rect -3373 688 -3327 700
rect -3373 -688 -3367 688
rect -3333 -688 -3327 688
rect -3373 -700 -3327 -688
rect -3105 688 -3059 700
rect -3105 -688 -3099 688
rect -3065 -688 -3059 688
rect -3105 -700 -3059 -688
rect -2837 688 -2791 700
rect -2837 -688 -2831 688
rect -2797 -688 -2791 688
rect -2837 -700 -2791 -688
rect -2569 688 -2523 700
rect -2569 -688 -2563 688
rect -2529 -688 -2523 688
rect -2569 -700 -2523 -688
rect -2301 688 -2255 700
rect -2301 -688 -2295 688
rect -2261 -688 -2255 688
rect -2301 -700 -2255 -688
rect -2033 688 -1987 700
rect -2033 -688 -2027 688
rect -1993 -688 -1987 688
rect -2033 -700 -1987 -688
rect -1765 688 -1719 700
rect -1765 -688 -1759 688
rect -1725 -688 -1719 688
rect -1765 -700 -1719 -688
rect -1497 688 -1451 700
rect -1497 -688 -1491 688
rect -1457 -688 -1451 688
rect -1497 -700 -1451 -688
rect -1229 688 -1183 700
rect -1229 -688 -1223 688
rect -1189 -688 -1183 688
rect -1229 -700 -1183 -688
rect -961 688 -915 700
rect -961 -688 -955 688
rect -921 -688 -915 688
rect -961 -700 -915 -688
rect -693 688 -647 700
rect -693 -688 -687 688
rect -653 -688 -647 688
rect -693 -700 -647 -688
rect -425 688 -379 700
rect -425 -688 -419 688
rect -385 -688 -379 688
rect -425 -700 -379 -688
rect -157 688 -111 700
rect -157 -688 -151 688
rect -117 -688 -111 688
rect -157 -700 -111 -688
rect 111 688 157 700
rect 111 -688 117 688
rect 151 -688 157 688
rect 111 -700 157 -688
rect 379 688 425 700
rect 379 -688 385 688
rect 419 -688 425 688
rect 379 -700 425 -688
rect 647 688 693 700
rect 647 -688 653 688
rect 687 -688 693 688
rect 647 -700 693 -688
rect 915 688 961 700
rect 915 -688 921 688
rect 955 -688 961 688
rect 915 -700 961 -688
rect 1183 688 1229 700
rect 1183 -688 1189 688
rect 1223 -688 1229 688
rect 1183 -700 1229 -688
rect 1451 688 1497 700
rect 1451 -688 1457 688
rect 1491 -688 1497 688
rect 1451 -700 1497 -688
rect 1719 688 1765 700
rect 1719 -688 1725 688
rect 1759 -688 1765 688
rect 1719 -700 1765 -688
rect 1987 688 2033 700
rect 1987 -688 1993 688
rect 2027 -688 2033 688
rect 1987 -700 2033 -688
rect 2255 688 2301 700
rect 2255 -688 2261 688
rect 2295 -688 2301 688
rect 2255 -700 2301 -688
rect 2523 688 2569 700
rect 2523 -688 2529 688
rect 2563 -688 2569 688
rect 2523 -700 2569 -688
rect 2791 688 2837 700
rect 2791 -688 2797 688
rect 2831 -688 2837 688
rect 2791 -700 2837 -688
rect 3059 688 3105 700
rect 3059 -688 3065 688
rect 3099 -688 3105 688
rect 3059 -700 3105 -688
rect 3327 688 3373 700
rect 3327 -688 3333 688
rect 3367 -688 3373 688
rect 3327 -700 3373 -688
rect -3317 -747 -3115 -741
rect -3317 -781 -3305 -747
rect -3127 -781 -3115 -747
rect -3317 -787 -3115 -781
rect -3049 -747 -2847 -741
rect -3049 -781 -3037 -747
rect -2859 -781 -2847 -747
rect -3049 -787 -2847 -781
rect -2781 -747 -2579 -741
rect -2781 -781 -2769 -747
rect -2591 -781 -2579 -747
rect -2781 -787 -2579 -781
rect -2513 -747 -2311 -741
rect -2513 -781 -2501 -747
rect -2323 -781 -2311 -747
rect -2513 -787 -2311 -781
rect -2245 -747 -2043 -741
rect -2245 -781 -2233 -747
rect -2055 -781 -2043 -747
rect -2245 -787 -2043 -781
rect -1977 -747 -1775 -741
rect -1977 -781 -1965 -747
rect -1787 -781 -1775 -747
rect -1977 -787 -1775 -781
rect -1709 -747 -1507 -741
rect -1709 -781 -1697 -747
rect -1519 -781 -1507 -747
rect -1709 -787 -1507 -781
rect -1441 -747 -1239 -741
rect -1441 -781 -1429 -747
rect -1251 -781 -1239 -747
rect -1441 -787 -1239 -781
rect -1173 -747 -971 -741
rect -1173 -781 -1161 -747
rect -983 -781 -971 -747
rect -1173 -787 -971 -781
rect -905 -747 -703 -741
rect -905 -781 -893 -747
rect -715 -781 -703 -747
rect -905 -787 -703 -781
rect -637 -747 -435 -741
rect -637 -781 -625 -747
rect -447 -781 -435 -747
rect -637 -787 -435 -781
rect -369 -747 -167 -741
rect -369 -781 -357 -747
rect -179 -781 -167 -747
rect -369 -787 -167 -781
rect -101 -747 101 -741
rect -101 -781 -89 -747
rect 89 -781 101 -747
rect -101 -787 101 -781
rect 167 -747 369 -741
rect 167 -781 179 -747
rect 357 -781 369 -747
rect 167 -787 369 -781
rect 435 -747 637 -741
rect 435 -781 447 -747
rect 625 -781 637 -747
rect 435 -787 637 -781
rect 703 -747 905 -741
rect 703 -781 715 -747
rect 893 -781 905 -747
rect 703 -787 905 -781
rect 971 -747 1173 -741
rect 971 -781 983 -747
rect 1161 -781 1173 -747
rect 971 -787 1173 -781
rect 1239 -747 1441 -741
rect 1239 -781 1251 -747
rect 1429 -781 1441 -747
rect 1239 -787 1441 -781
rect 1507 -747 1709 -741
rect 1507 -781 1519 -747
rect 1697 -781 1709 -747
rect 1507 -787 1709 -781
rect 1775 -747 1977 -741
rect 1775 -781 1787 -747
rect 1965 -781 1977 -747
rect 1775 -787 1977 -781
rect 2043 -747 2245 -741
rect 2043 -781 2055 -747
rect 2233 -781 2245 -747
rect 2043 -787 2245 -781
rect 2311 -747 2513 -741
rect 2311 -781 2323 -747
rect 2501 -781 2513 -747
rect 2311 -787 2513 -781
rect 2579 -747 2781 -741
rect 2579 -781 2591 -747
rect 2769 -781 2781 -747
rect 2579 -787 2781 -781
rect 2847 -747 3049 -741
rect 2847 -781 2859 -747
rect 3037 -781 3049 -747
rect 2847 -787 3049 -781
rect 3115 -747 3317 -741
rect 3115 -781 3127 -747
rect 3305 -781 3317 -747
rect 3115 -787 3317 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -3464 -866 3464 866
string parameters w 7 l 1.05 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
