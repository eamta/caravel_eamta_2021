magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 334 1713 369 1747
rect 335 1694 369 1713
rect 165 1645 223 1651
rect 165 1611 177 1645
rect 165 1605 223 1611
rect 227 1400 267 1418
rect 354 1400 369 1694
rect 388 1660 423 1694
rect 388 1400 422 1660
rect 534 1592 592 1598
rect 534 1558 546 1592
rect 534 1552 592 1558
rect 704 1551 738 1605
rect 1126 1587 1161 1605
rect 1090 1572 1161 1587
rect 1441 1572 1476 1606
rect 0 1224 506 1400
rect 534 1302 592 1308
rect 534 1271 546 1302
rect 534 1268 580 1271
rect 534 1262 592 1268
rect 0 1200 531 1224
rect 0 1166 642 1200
rect 723 1166 738 1551
rect 757 1517 792 1551
rect 757 1166 791 1517
rect 1090 1455 1160 1572
rect 1442 1553 1476 1572
rect 1272 1504 1330 1510
rect 1272 1470 1284 1504
rect 1272 1464 1330 1470
rect 903 1449 961 1455
rect 903 1415 915 1449
rect 903 1409 961 1415
rect 1073 1348 1160 1455
rect 993 1312 1018 1317
rect 984 1287 1005 1312
rect 1073 1295 1370 1348
rect 1461 1295 1476 1553
rect 1495 1519 1530 1553
rect 1810 1519 1845 1553
rect 1495 1295 1529 1519
rect 1811 1500 1845 1519
rect 1641 1451 1699 1457
rect 1641 1417 1653 1451
rect 1641 1411 1699 1417
rect 984 1278 996 1287
rect 903 1249 961 1255
rect 903 1215 915 1249
rect 950 1215 965 1249
rect 984 1216 999 1278
rect 1073 1242 1739 1295
rect 1830 1242 1845 1500
rect 1864 1466 1899 1500
rect 1864 1242 1898 1466
rect 2010 1398 2068 1404
rect 2010 1364 2022 1398
rect 2010 1358 2068 1364
rect 903 1209 961 1215
rect -830 1049 -795 1083
rect -515 1064 -480 1082
rect -515 1049 -444 1064
rect -1199 996 -1164 1030
rect -1233 450 -1218 977
rect -1199 518 -1165 996
rect -1053 928 -995 934
rect -1053 894 -1041 928
rect -1053 888 -995 894
rect -1053 620 -995 626
rect -1053 586 -1041 620
rect -1053 580 -995 586
rect -1199 484 -1164 518
rect -864 503 -849 1030
rect -830 571 -796 1049
rect -514 1028 -444 1049
rect -497 994 -426 1028
rect -684 981 -626 987
rect -684 947 -672 981
rect -684 941 -626 947
rect -684 673 -626 679
rect -684 639 -672 673
rect -684 633 -626 639
rect -497 624 -427 994
rect -315 926 -257 932
rect -315 892 -303 926
rect -315 886 -257 892
rect -315 726 -257 732
rect -315 692 -303 726
rect -315 686 -257 692
rect -497 590 -426 624
rect -126 609 -111 1028
rect -92 677 -58 1082
rect 0 996 506 1166
rect 757 1132 772 1166
rect 984 1147 1018 1216
rect 1073 1209 2108 1242
rect 853 1113 1018 1147
rect 1090 1189 2108 1209
rect 1090 1138 2250 1189
rect 2424 1153 2477 1154
rect 1086 1113 2250 1138
rect 2406 1119 2477 1153
rect 2407 1118 2477 1119
rect 984 1022 1018 1113
rect 1090 1051 2250 1113
rect 2424 1084 2495 1118
rect 2775 1084 2810 1118
rect 1090 1024 2252 1051
rect 1300 1022 1334 1024
rect 1353 1022 1387 1024
rect 1459 1022 2252 1024
rect 2424 1022 2494 1084
rect 2776 1065 2810 1084
rect 2795 1022 2810 1065
rect 647 1021 663 1022
rect 22 980 60 984
rect 22 973 85 980
rect 10 912 85 973
rect 98 962 156 996
rect 224 990 311 996
rect 98 952 150 962
rect 98 924 144 952
rect 10 902 68 912
rect 10 887 56 902
rect 22 863 56 887
rect 98 886 150 924
rect 151 896 156 962
rect 166 928 178 970
rect 182 928 194 962
rect 166 914 178 924
rect 76 874 82 878
rect 98 877 144 886
rect 224 877 258 990
rect 274 956 311 990
rect 324 956 345 990
rect 277 877 311 956
rect 379 941 412 996
rect 382 895 412 941
rect 379 885 419 895
rect 379 882 425 885
rect 379 877 427 882
rect 646 877 663 1021
rect 948 986 2494 1022
rect 2618 1016 2652 1020
rect 2776 986 2810 1022
rect 2829 1040 2864 1065
rect 2829 1031 3053 1040
rect 3144 1031 3179 1065
rect 2829 986 2863 1031
rect 3145 1012 3179 1031
rect 728 963 2863 986
rect 2949 963 3021 986
rect 728 952 3021 963
rect 98 874 663 877
rect 76 873 88 874
rect 68 863 88 873
rect 22 836 88 863
rect 104 859 663 874
rect 98 851 663 859
rect 104 836 663 851
rect 22 829 82 836
rect 48 817 82 829
rect 110 829 663 836
rect 110 817 116 829
rect 136 817 663 829
rect 48 813 94 817
rect 32 779 94 813
rect 100 779 663 817
rect 50 745 663 779
rect 948 748 2494 952
rect 2540 941 2730 952
rect 2574 935 2608 939
rect 2662 935 2696 939
rect 2562 927 2620 935
rect 2650 927 2708 935
rect 2568 913 2614 927
rect 2656 913 2708 927
rect 2574 877 2614 913
rect 2624 895 2642 907
rect 2662 905 2708 913
rect 2650 895 2708 905
rect 50 731 94 745
rect 136 731 663 745
rect 36 694 94 731
rect 124 694 663 731
rect 1317 695 2494 748
rect 48 690 82 694
rect 136 690 663 694
rect 140 677 663 690
rect -92 643 -57 677
rect 0 660 663 677
rect 1686 660 2494 695
rect 2502 660 2528 802
rect 2540 727 2542 849
rect 2568 839 2570 849
rect 2574 839 2608 877
rect 2620 861 2708 895
rect 2650 855 2686 861
rect 2693 855 2708 861
rect 2650 851 2708 855
rect 2562 801 2608 839
rect 2562 798 2624 801
rect 2568 755 2570 798
rect 2574 767 2624 798
rect 2590 755 2624 767
rect 2628 755 2630 798
rect 2656 755 2658 826
rect 2660 801 2708 851
rect 2726 801 2730 805
rect 2742 801 2760 805
rect 2688 767 2702 801
rect 2692 755 2702 767
rect 2714 755 2762 801
rect 2590 742 2636 755
rect 2692 751 2696 755
rect 2584 708 2636 742
rect 2720 729 2734 755
rect 2720 727 2730 729
rect 2726 717 2730 727
rect 2602 660 2636 708
rect 2652 674 2658 708
rect 2742 660 2760 755
rect 0 659 316 660
rect 0 643 310 659
rect 140 641 310 643
rect 322 641 376 660
rect 382 659 422 660
rect 388 641 422 659
rect 476 641 510 660
rect 1686 642 2548 660
rect 53 606 510 641
rect -830 537 -795 571
rect -497 554 -444 590
rect 476 547 510 606
rect 2055 618 2548 642
rect 2578 618 2636 660
rect 2714 621 2772 660
rect 2055 606 2494 618
rect 2502 614 2536 618
rect 2590 614 2624 618
rect 2726 617 2760 621
rect 2776 606 2810 952
rect 2829 823 2863 952
rect 2987 941 3021 952
rect 2971 929 3037 941
rect 2971 919 2989 929
rect 2939 882 2989 919
rect 3019 913 3037 929
rect 3145 931 3156 942
rect 3164 935 3179 1012
rect 3198 978 3233 1012
rect 3513 978 3548 1012
rect 3198 935 3232 978
rect 3514 959 3548 978
rect 3164 931 3232 935
rect 3145 901 3232 931
rect 3316 941 3430 944
rect 3145 890 3156 901
rect 3164 887 3179 901
rect 2931 869 2989 882
rect 3019 870 3042 882
rect 2931 854 2977 869
rect 2829 805 2882 823
rect 2814 633 2882 805
rect 2943 821 2977 854
rect 3019 867 3065 870
rect 3019 833 3027 867
rect 2943 714 2985 821
rect 2951 671 2985 714
rect 2989 702 2996 832
rect 3031 821 3065 867
rect 3070 833 3077 882
rect 3145 855 3179 887
rect 3031 714 3073 821
rect 3039 702 3073 714
rect 2989 671 2997 702
rect 2951 655 2997 671
rect 3021 655 3073 702
rect 2814 621 2860 633
rect 2951 621 3073 655
rect 2814 617 2863 621
rect 2829 606 2863 617
rect 2055 603 2658 606
rect 2692 603 2863 606
rect 2055 589 2863 603
rect 2460 583 2863 589
rect 2460 580 2703 583
rect 2460 572 2501 580
rect 2548 573 2703 580
rect 2651 572 2703 573
rect 2761 574 2863 583
rect 2761 572 2810 574
rect 2829 553 2863 574
rect 2951 605 2997 621
rect 3027 605 3037 621
rect 2951 553 2985 605
rect 3039 553 3073 621
rect 3145 615 3195 855
rect 3145 553 3179 615
rect 2829 540 2887 553
rect 2829 530 2865 540
rect 2829 519 2840 530
rect 2925 519 3179 553
rect 3198 519 3232 901
rect 3241 867 3266 901
rect 3316 842 3331 941
rect 3344 910 3402 916
rect 3344 901 3359 910
rect 3340 880 3359 901
rect 3340 876 3372 880
rect 3388 876 3390 880
rect 3340 870 3402 876
rect 3340 860 3358 870
rect 3430 860 3448 901
rect 3533 871 3548 959
rect 3039 485 3073 519
rect 3198 473 3227 519
rect 3284 500 3286 833
rect 3372 829 3403 833
rect 3296 817 3330 821
rect 3342 817 3346 828
rect 3296 661 3346 817
rect 3296 636 3330 661
rect 3350 649 3352 829
rect 3373 821 3403 829
rect 3378 649 3380 821
rect 3384 817 3418 821
rect 3430 817 3434 828
rect 3384 661 3434 817
rect 3384 649 3418 661
rect 3438 649 3440 829
rect 3296 534 3336 636
rect 3340 602 3342 618
rect 3344 602 3364 608
rect 3372 602 3418 649
rect 3466 621 3468 833
rect 3340 568 3418 602
rect 3340 552 3342 568
rect 3344 562 3364 568
rect 3372 552 3418 568
rect 3296 500 3330 534
rect 3384 500 3418 552
rect 3480 534 3506 837
rect 3472 500 3506 534
rect 3514 500 3548 871
rect 3284 473 3518 500
rect 3331 466 3383 473
rect 3419 466 3471 473
rect 3533 466 3548 500
rect 3567 925 3602 959
rect 3882 925 3917 959
rect 3567 466 3601 925
rect 3883 906 3917 925
rect 3713 857 3771 863
rect 3713 823 3725 857
rect 3713 817 3771 823
rect 3713 549 3771 555
rect 3713 515 3725 549
rect 3713 509 3771 515
rect 3567 432 3582 466
rect 3902 413 3917 906
rect 3936 872 3971 906
rect 4251 872 4286 906
rect 3936 413 3970 872
rect 4252 853 4286 872
rect 4082 804 4140 810
rect 4082 770 4094 804
rect 4082 764 4140 770
rect 4082 496 4140 502
rect 4082 462 4094 496
rect 4082 456 4140 462
rect 3531 377 3586 411
rect 3936 379 3951 413
rect 4271 360 4286 853
rect 4305 819 4340 853
rect 4305 360 4339 819
rect 4451 751 4509 757
rect 4451 717 4463 751
rect 4621 728 4655 746
rect 4451 711 4509 717
rect 4621 692 4691 728
rect 4638 658 4709 692
rect 4451 443 4509 449
rect 4451 409 4463 443
rect 4451 403 4509 409
rect 4305 326 4320 360
rect 4638 307 4708 658
rect 4638 271 4691 307
rect 1025 201 1102 222
rect 1132 201 1201 222
rect 1025 173 1102 194
rect 1132 173 1229 194
rect 653 -1599 688 -1565
rect 654 -1618 688 -1599
rect 673 -1855 688 -1618
rect 707 -1652 742 -1618
rect 1022 -1652 1057 -1618
rect 707 -1855 741 -1652
rect 1023 -1671 1057 -1652
rect 853 -1720 911 -1714
rect 853 -1754 865 -1720
rect 853 -1760 911 -1754
rect 821 -1855 855 -1804
rect 909 -1855 943 -1804
rect 302 -1891 1002 -1855
rect 82 -1925 1002 -1891
rect 302 -2129 1002 -1925
rect 671 -2182 1002 -2129
rect 1042 -2146 1057 -1671
rect 1076 -1705 1111 -1671
rect 1391 -1705 1426 -1671
rect 1076 -2146 1110 -1705
rect 1392 -1724 1426 -1705
rect 1778 -1724 1831 -1723
rect 1194 -1799 1201 -1739
rect 1222 -1773 1280 -1767
rect 1222 -1807 1234 -1773
rect 1222 -1813 1280 -1807
rect 1222 -2063 1280 -2057
rect 1222 -2097 1234 -2063
rect 1222 -2103 1280 -2097
rect 1076 -2180 1091 -2146
rect 1411 -2199 1426 -1724
rect 1445 -1758 1480 -1724
rect 1760 -1758 1831 -1724
rect 1445 -2199 1479 -1758
rect 1761 -1759 1831 -1758
rect 1778 -1793 1849 -1759
rect 2129 -1793 2164 -1759
rect 1591 -1826 1649 -1820
rect 1591 -1860 1603 -1826
rect 1591 -1866 1649 -1860
rect 1591 -2116 1649 -2110
rect 1591 -2150 1603 -2116
rect 1591 -2156 1649 -2150
rect 1445 -2233 1460 -2199
rect 1778 -2252 1848 -1793
rect 2130 -1812 2164 -1793
rect 1960 -1861 2018 -1855
rect 1960 -1895 1972 -1861
rect 1960 -1901 2018 -1895
rect 1960 -2169 2018 -2163
rect 1960 -2203 1972 -2169
rect 1960 -2209 2018 -2203
rect 1778 -2288 1831 -2252
rect 2149 -2305 2164 -1812
rect 2183 -1846 2218 -1812
rect 2498 -1846 2533 -1812
rect 2183 -2305 2217 -1846
rect 2499 -1865 2533 -1846
rect 2329 -1914 2387 -1908
rect 2329 -1948 2341 -1914
rect 2329 -1954 2387 -1948
rect 2329 -2222 2387 -2216
rect 2329 -2256 2341 -2222
rect 2329 -2262 2387 -2256
rect 2183 -2339 2198 -2305
rect 2518 -2358 2533 -1865
rect 2552 -1899 2587 -1865
rect 2867 -1899 2902 -1865
rect 2552 -2358 2586 -1899
rect 2868 -1918 2902 -1899
rect 2698 -1967 2756 -1961
rect 2698 -2001 2710 -1967
rect 2698 -2007 2756 -2001
rect 2698 -2275 2756 -2269
rect 2698 -2309 2710 -2275
rect 2698 -2315 2756 -2309
rect 2552 -2392 2567 -2358
rect 2887 -2411 2902 -1918
rect 2921 -1952 2956 -1918
rect 3236 -1952 3271 -1918
rect 2921 -2411 2955 -1952
rect 3237 -1971 3271 -1952
rect 3067 -2020 3125 -2014
rect 3067 -2054 3079 -2020
rect 3067 -2060 3125 -2054
rect 3067 -2328 3125 -2322
rect 3067 -2362 3079 -2328
rect 3067 -2368 3125 -2362
rect 2921 -2445 2936 -2411
rect 3256 -2464 3271 -1971
rect 3290 -2005 3325 -1971
rect 3605 -2005 3640 -1971
rect 3290 -2464 3324 -2005
rect 3606 -2024 3640 -2005
rect 3436 -2073 3494 -2067
rect 3436 -2107 3448 -2073
rect 3436 -2113 3494 -2107
rect 3436 -2381 3494 -2375
rect 3436 -2415 3448 -2381
rect 3436 -2421 3494 -2415
rect 3290 -2498 3305 -2464
rect 3625 -2517 3640 -2024
rect 3659 -2058 3694 -2024
rect 3659 -2517 3693 -2058
rect 3805 -2126 3863 -2120
rect 3805 -2160 3817 -2126
rect 3975 -2149 4009 -2131
rect 3805 -2166 3863 -2160
rect 3975 -2185 4045 -2149
rect 3992 -2219 4063 -2185
rect 4343 -2219 4378 -2185
rect 3805 -2434 3863 -2428
rect 3805 -2468 3817 -2434
rect 3805 -2474 3863 -2468
rect 3659 -2551 3674 -2517
rect 3992 -2570 4062 -2219
rect 4344 -2238 4378 -2219
rect 4174 -2287 4232 -2281
rect 4174 -2321 4186 -2287
rect 4174 -2327 4232 -2321
rect 4174 -2487 4232 -2481
rect 4174 -2521 4186 -2487
rect 4174 -2527 4232 -2521
rect 3992 -2606 4045 -2570
rect 4363 -2623 4378 -2238
rect 4397 -2272 4432 -2238
rect 4397 -2623 4431 -2272
rect 4543 -2340 4601 -2334
rect 4543 -2374 4555 -2340
rect 4543 -2380 4601 -2374
rect 4543 -2540 4601 -2534
rect 4543 -2574 4555 -2540
rect 4543 -2580 4601 -2574
rect 379 -2676 456 -2655
rect 486 -2676 555 -2655
rect 4397 -2657 4412 -2623
rect 379 -2704 456 -2683
rect 486 -2704 583 -2683
<< metal1 >>
rect 602 971 3554 1022
rect 602 875 647 971
rect 140 349 228 483
rect 632 458 660 566
rect 638 378 648 430
rect 700 378 710 430
rect 1564 390 1574 442
rect 1626 390 1636 442
rect 1676 417 1742 475
rect 0 0 200 200
rect 646 77 647 78
rect 618 76 1648 77
rect 618 49 3524 76
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
<< via1 >>
rect 648 378 700 430
rect 1574 390 1626 442
<< metal2 >>
rect 3201 555 3253 607
rect 1086 514 2027 542
rect 1999 460 2027 514
rect 1574 442 1626 452
rect 648 430 700 440
rect 700 390 1574 409
rect 2834 409 2894 451
rect 1626 390 2895 409
rect 700 381 2895 390
rect 1574 380 1626 381
rect 648 368 700 378
use xor_lafe  xor_lafe_0
timestamp 1624053917
transform 1 0 1001 0 1 201
box -355 -2000 4428 1147
use xor_lafe  xor_lafe_1
timestamp 1624053917
transform 1 0 355 0 1 -2676
box -355 -2000 4428 1147
use and_lafe  and_lafe_0
timestamp 1624053917
transform -1 0 610 0 1 113
box -53 -2000 2214 1147
use and_lafe  and_lafe_1
timestamp 1624053917
transform 1 0 36 0 1 636
box -53 -2000 2214 1147
use dffc2  dffc2_0
timestamp 1624053917
transform 1 0 2672 0 1 457
box -1024 -425 882 565
<< labels >>
rlabel metal1 632 458 660 566 1 CE
rlabel metal1 1676 417 1742 475 1 CLK
rlabel metal2 3201 555 3253 607 1 CLR
rlabel metal1 602 971 3554 1022 1 vdd
rlabel metal1 646 49 3524 76 1 vss
rlabel metal2 2834 393 2894 451 1 Q
rlabel metal1 140 349 228 483 1 Sout
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Sout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLK
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 CLR
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 CE
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 vss
port 7 nsew
<< end >>
