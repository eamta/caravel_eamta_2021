magic
tech sky130A
magscale 1 2
timestamp 1617978432
<< nwell >>
rect 3414 1135 3477 1539
rect 2907 989 2908 991
rect 3983 989 3984 991
rect 3414 441 3485 845
<< poly >>
rect 1604 1863 1813 1893
rect 1782 1821 1813 1863
rect 5079 1863 5321 1893
rect 5079 1821 5109 1863
rect 1782 827 1812 1153
rect 5079 827 5109 1153
<< metal1 >>
rect 1876 1947 4986 1980
rect 2907 1935 3984 1947
rect 1546 1834 1556 1886
rect 1608 1834 1618 1886
rect 3414 1876 3478 1935
rect 6891 1921 6948 1980
rect 5253 1834 5263 1886
rect 5315 1834 5325 1886
rect 3326 1529 3414 1663
rect 3497 1533 3507 1585
rect 3559 1533 3569 1585
rect 2849 1417 2859 1469
rect 2911 1417 2921 1469
rect 4003 1433 4013 1485
rect 4065 1433 4075 1485
rect 3414 1135 3483 1255
rect -56 909 0 1071
rect 3414 725 3477 845
rect 1812 385 1878 443
rect 2894 426 2922 534
rect 3970 487 3980 539
rect 4032 487 4042 539
rect 3467 419 3477 471
rect 3529 419 3539 471
rect 3364 303 3416 336
rect 3344 251 3354 303
rect 3406 251 3416 303
rect 3414 47 3477 104
rect 6920 59 6948 1921
rect 1906 0 5172 47
rect 6891 0 6948 59
<< via1 >>
rect 1556 1834 1608 1886
rect 5263 1834 5315 1886
rect 3507 1533 3559 1585
rect 2859 1417 2911 1469
rect 4013 1433 4065 1485
rect 3980 487 4032 539
rect 3477 419 3529 471
rect 3354 251 3406 303
<< metal2 >>
rect 1556 1886 1608 1896
rect 5263 1886 5315 1896
rect 1608 1834 5263 1852
rect 1556 1824 5315 1834
rect 659 1556 721 1628
rect 3507 1585 3559 1595
rect 6170 1556 6232 1628
rect 3507 1523 3559 1533
rect 3529 1479 3557 1523
rect 2859 1469 3557 1479
rect 2911 1451 3557 1469
rect 4013 1485 4066 1495
rect 4065 1433 4066 1485
rect 4013 1423 4066 1433
rect 2859 1407 2911 1417
rect 316 577 344 1405
rect 4038 605 4066 1423
rect 3501 577 4066 605
rect 291 523 363 577
rect 316 122 344 523
rect 3501 481 3529 577
rect 6547 575 6575 1405
rect 3980 539 4032 549
rect 3477 471 3529 481
rect 659 349 721 424
rect 3477 409 3529 419
rect 3853 487 3980 508
rect 3853 480 4032 487
rect 3853 313 3881 480
rect 3980 477 4032 480
rect 6170 352 6232 424
rect 3354 303 3881 313
rect 3406 285 3881 303
rect 3354 241 3406 251
rect 6547 122 6575 572
rect 316 94 6575 122
use contador1bit  contador1bit_1 
timestamp 1617974880
transform 1 0 3337 0 1 -32
box 140 32 3554 1022
use contador1bit  contador1bit_0
timestamp 1617974880
transform -1 0 3554 0 1 -32
box 140 32 3554 1022
use contador1bit  contador1bit_2
timestamp 1617974880
transform 1 0 3337 0 -1 2012
box 140 32 3554 1022
use contador1bit  contador1bit_3
timestamp 1617974880
transform -1 0 3554 0 -1 2012
box 140 32 3554 1022
use contacto  contacto_0
timestamp 1616018980
transform 1 0 1558 0 1 1830
box 0 4 66 62
use contacto  contacto_1
timestamp 1616018980
transform 1 0 5263 0 1 1830
box 0 4 66 62
<< labels >>
rlabel metal1 1812 386 1878 442 1 CLK
rlabel metal2 291 523 363 577 1 CLR
rlabel metal2 659 1556 721 1628 1 Q3
rlabel metal2 6170 1556 6232 1628 1 Q2
rlabel metal2 6170 352 6232 424 1 Q1
rlabel metal2 659 349 721 424 1 Q0
rlabel metal1 2894 426 2922 534 1 CE
rlabel metal1 3326 1529 3414 1663 1 Sout
rlabel metal1 6920 0 6948 1980 1 vss
rlabel metal1 -56 909 0 1071 1 vdd
<< end >>
