magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -2381 481 -2323 487
rect -2189 481 -2131 487
rect -1997 481 -1939 487
rect -1805 481 -1747 487
rect -1613 481 -1555 487
rect -1421 481 -1363 487
rect -1229 481 -1171 487
rect -1037 481 -979 487
rect -845 481 -787 487
rect -653 481 -595 487
rect -461 481 -403 487
rect -269 481 -211 487
rect -77 481 -19 487
rect 115 481 173 487
rect 307 481 365 487
rect 499 481 557 487
rect 691 481 749 487
rect 883 481 941 487
rect 1075 481 1133 487
rect 1267 481 1325 487
rect 1459 481 1517 487
rect 1651 481 1709 487
rect 1843 481 1901 487
rect 2035 481 2093 487
rect 2227 481 2285 487
rect -2381 447 -2369 481
rect -2189 447 -2177 481
rect -1997 447 -1985 481
rect -1805 447 -1793 481
rect -1613 447 -1601 481
rect -1421 447 -1409 481
rect -1229 447 -1217 481
rect -1037 447 -1025 481
rect -845 447 -833 481
rect -653 447 -641 481
rect -461 447 -449 481
rect -269 447 -257 481
rect -77 447 -65 481
rect 115 447 127 481
rect 307 447 319 481
rect 499 447 511 481
rect 691 447 703 481
rect 883 447 895 481
rect 1075 447 1087 481
rect 1267 447 1279 481
rect 1459 447 1471 481
rect 1651 447 1663 481
rect 1843 447 1855 481
rect 2035 447 2047 481
rect 2227 447 2239 481
rect -2381 441 -2323 447
rect -2189 441 -2131 447
rect -1997 441 -1939 447
rect -1805 441 -1747 447
rect -1613 441 -1555 447
rect -1421 441 -1363 447
rect -1229 441 -1171 447
rect -1037 441 -979 447
rect -845 441 -787 447
rect -653 441 -595 447
rect -461 441 -403 447
rect -269 441 -211 447
rect -77 441 -19 447
rect 115 441 173 447
rect 307 441 365 447
rect 499 441 557 447
rect 691 441 749 447
rect 883 441 941 447
rect 1075 441 1133 447
rect 1267 441 1325 447
rect 1459 441 1517 447
rect 1651 441 1709 447
rect 1843 441 1901 447
rect 2035 441 2093 447
rect 2227 441 2285 447
rect -2285 71 -2227 77
rect -2093 71 -2035 77
rect -1901 71 -1843 77
rect -1709 71 -1651 77
rect -1517 71 -1459 77
rect -1325 71 -1267 77
rect -1133 71 -1075 77
rect -941 71 -883 77
rect -749 71 -691 77
rect -557 71 -499 77
rect -365 71 -307 77
rect -173 71 -115 77
rect 19 71 77 77
rect 211 71 269 77
rect 403 71 461 77
rect 595 71 653 77
rect 787 71 845 77
rect 979 71 1037 77
rect 1171 71 1229 77
rect 1363 71 1421 77
rect 1555 71 1613 77
rect 1747 71 1805 77
rect 1939 71 1997 77
rect 2131 71 2189 77
rect 2323 71 2381 77
rect -2285 37 -2273 71
rect -2093 37 -2081 71
rect -1901 37 -1889 71
rect -1709 37 -1697 71
rect -1517 37 -1505 71
rect -1325 37 -1313 71
rect -1133 37 -1121 71
rect -941 37 -929 71
rect -749 37 -737 71
rect -557 37 -545 71
rect -365 37 -353 71
rect -173 37 -161 71
rect 19 37 31 71
rect 211 37 223 71
rect 403 37 415 71
rect 595 37 607 71
rect 787 37 799 71
rect 979 37 991 71
rect 1171 37 1183 71
rect 1363 37 1375 71
rect 1555 37 1567 71
rect 1747 37 1759 71
rect 1939 37 1951 71
rect 2131 37 2143 71
rect 2323 37 2335 71
rect -2285 31 -2227 37
rect -2093 31 -2035 37
rect -1901 31 -1843 37
rect -1709 31 -1651 37
rect -1517 31 -1459 37
rect -1325 31 -1267 37
rect -1133 31 -1075 37
rect -941 31 -883 37
rect -749 31 -691 37
rect -557 31 -499 37
rect -365 31 -307 37
rect -173 31 -115 37
rect 19 31 77 37
rect 211 31 269 37
rect 403 31 461 37
rect 595 31 653 37
rect 787 31 845 37
rect 979 31 1037 37
rect 1171 31 1229 37
rect 1363 31 1421 37
rect 1555 31 1613 37
rect 1747 31 1805 37
rect 1939 31 1997 37
rect 2131 31 2189 37
rect 2323 31 2381 37
rect -2285 -37 -2227 -31
rect -2093 -37 -2035 -31
rect -1901 -37 -1843 -31
rect -1709 -37 -1651 -31
rect -1517 -37 -1459 -31
rect -1325 -37 -1267 -31
rect -1133 -37 -1075 -31
rect -941 -37 -883 -31
rect -749 -37 -691 -31
rect -557 -37 -499 -31
rect -365 -37 -307 -31
rect -173 -37 -115 -31
rect 19 -37 77 -31
rect 211 -37 269 -31
rect 403 -37 461 -31
rect 595 -37 653 -31
rect 787 -37 845 -31
rect 979 -37 1037 -31
rect 1171 -37 1229 -31
rect 1363 -37 1421 -31
rect 1555 -37 1613 -31
rect 1747 -37 1805 -31
rect 1939 -37 1997 -31
rect 2131 -37 2189 -31
rect 2323 -37 2381 -31
rect -2285 -71 -2273 -37
rect -2093 -71 -2081 -37
rect -1901 -71 -1889 -37
rect -1709 -71 -1697 -37
rect -1517 -71 -1505 -37
rect -1325 -71 -1313 -37
rect -1133 -71 -1121 -37
rect -941 -71 -929 -37
rect -749 -71 -737 -37
rect -557 -71 -545 -37
rect -365 -71 -353 -37
rect -173 -71 -161 -37
rect 19 -71 31 -37
rect 211 -71 223 -37
rect 403 -71 415 -37
rect 595 -71 607 -37
rect 787 -71 799 -37
rect 979 -71 991 -37
rect 1171 -71 1183 -37
rect 1363 -71 1375 -37
rect 1555 -71 1567 -37
rect 1747 -71 1759 -37
rect 1939 -71 1951 -37
rect 2131 -71 2143 -37
rect 2323 -71 2335 -37
rect -2285 -77 -2227 -71
rect -2093 -77 -2035 -71
rect -1901 -77 -1843 -71
rect -1709 -77 -1651 -71
rect -1517 -77 -1459 -71
rect -1325 -77 -1267 -71
rect -1133 -77 -1075 -71
rect -941 -77 -883 -71
rect -749 -77 -691 -71
rect -557 -77 -499 -71
rect -365 -77 -307 -71
rect -173 -77 -115 -71
rect 19 -77 77 -71
rect 211 -77 269 -71
rect 403 -77 461 -71
rect 595 -77 653 -71
rect 787 -77 845 -71
rect 979 -77 1037 -71
rect 1171 -77 1229 -71
rect 1363 -77 1421 -71
rect 1555 -77 1613 -71
rect 1747 -77 1805 -71
rect 1939 -77 1997 -71
rect 2131 -77 2189 -71
rect 2323 -77 2381 -71
rect -2381 -447 -2323 -441
rect -2189 -447 -2131 -441
rect -1997 -447 -1939 -441
rect -1805 -447 -1747 -441
rect -1613 -447 -1555 -441
rect -1421 -447 -1363 -441
rect -1229 -447 -1171 -441
rect -1037 -447 -979 -441
rect -845 -447 -787 -441
rect -653 -447 -595 -441
rect -461 -447 -403 -441
rect -269 -447 -211 -441
rect -77 -447 -19 -441
rect 115 -447 173 -441
rect 307 -447 365 -441
rect 499 -447 557 -441
rect 691 -447 749 -441
rect 883 -447 941 -441
rect 1075 -447 1133 -441
rect 1267 -447 1325 -441
rect 1459 -447 1517 -441
rect 1651 -447 1709 -441
rect 1843 -447 1901 -441
rect 2035 -447 2093 -441
rect 2227 -447 2285 -441
rect -2381 -481 -2369 -447
rect -2189 -481 -2177 -447
rect -1997 -481 -1985 -447
rect -1805 -481 -1793 -447
rect -1613 -481 -1601 -447
rect -1421 -481 -1409 -447
rect -1229 -481 -1217 -447
rect -1037 -481 -1025 -447
rect -845 -481 -833 -447
rect -653 -481 -641 -447
rect -461 -481 -449 -447
rect -269 -481 -257 -447
rect -77 -481 -65 -447
rect 115 -481 127 -447
rect 307 -481 319 -447
rect 499 -481 511 -447
rect 691 -481 703 -447
rect 883 -481 895 -447
rect 1075 -481 1087 -447
rect 1267 -481 1279 -447
rect 1459 -481 1471 -447
rect 1651 -481 1663 -447
rect 1843 -481 1855 -447
rect 2035 -481 2047 -447
rect 2227 -481 2239 -447
rect -2381 -487 -2323 -481
rect -2189 -487 -2131 -481
rect -1997 -487 -1939 -481
rect -1805 -487 -1747 -481
rect -1613 -487 -1555 -481
rect -1421 -487 -1363 -481
rect -1229 -487 -1171 -481
rect -1037 -487 -979 -481
rect -845 -487 -787 -481
rect -653 -487 -595 -481
rect -461 -487 -403 -481
rect -269 -487 -211 -481
rect -77 -487 -19 -481
rect 115 -487 173 -481
rect 307 -487 365 -481
rect 499 -487 557 -481
rect 691 -487 749 -481
rect 883 -487 941 -481
rect 1075 -487 1133 -481
rect 1267 -487 1325 -481
rect 1459 -487 1517 -481
rect 1651 -487 1709 -481
rect 1843 -487 1901 -481
rect 2035 -487 2093 -481
rect 2227 -487 2285 -481
<< pwell >>
rect -2567 -619 2567 619
<< nmos >>
rect -2367 109 -2337 409
rect -2271 109 -2241 409
rect -2175 109 -2145 409
rect -2079 109 -2049 409
rect -1983 109 -1953 409
rect -1887 109 -1857 409
rect -1791 109 -1761 409
rect -1695 109 -1665 409
rect -1599 109 -1569 409
rect -1503 109 -1473 409
rect -1407 109 -1377 409
rect -1311 109 -1281 409
rect -1215 109 -1185 409
rect -1119 109 -1089 409
rect -1023 109 -993 409
rect -927 109 -897 409
rect -831 109 -801 409
rect -735 109 -705 409
rect -639 109 -609 409
rect -543 109 -513 409
rect -447 109 -417 409
rect -351 109 -321 409
rect -255 109 -225 409
rect -159 109 -129 409
rect -63 109 -33 409
rect 33 109 63 409
rect 129 109 159 409
rect 225 109 255 409
rect 321 109 351 409
rect 417 109 447 409
rect 513 109 543 409
rect 609 109 639 409
rect 705 109 735 409
rect 801 109 831 409
rect 897 109 927 409
rect 993 109 1023 409
rect 1089 109 1119 409
rect 1185 109 1215 409
rect 1281 109 1311 409
rect 1377 109 1407 409
rect 1473 109 1503 409
rect 1569 109 1599 409
rect 1665 109 1695 409
rect 1761 109 1791 409
rect 1857 109 1887 409
rect 1953 109 1983 409
rect 2049 109 2079 409
rect 2145 109 2175 409
rect 2241 109 2271 409
rect 2337 109 2367 409
rect -2367 -409 -2337 -109
rect -2271 -409 -2241 -109
rect -2175 -409 -2145 -109
rect -2079 -409 -2049 -109
rect -1983 -409 -1953 -109
rect -1887 -409 -1857 -109
rect -1791 -409 -1761 -109
rect -1695 -409 -1665 -109
rect -1599 -409 -1569 -109
rect -1503 -409 -1473 -109
rect -1407 -409 -1377 -109
rect -1311 -409 -1281 -109
rect -1215 -409 -1185 -109
rect -1119 -409 -1089 -109
rect -1023 -409 -993 -109
rect -927 -409 -897 -109
rect -831 -409 -801 -109
rect -735 -409 -705 -109
rect -639 -409 -609 -109
rect -543 -409 -513 -109
rect -447 -409 -417 -109
rect -351 -409 -321 -109
rect -255 -409 -225 -109
rect -159 -409 -129 -109
rect -63 -409 -33 -109
rect 33 -409 63 -109
rect 129 -409 159 -109
rect 225 -409 255 -109
rect 321 -409 351 -109
rect 417 -409 447 -109
rect 513 -409 543 -109
rect 609 -409 639 -109
rect 705 -409 735 -109
rect 801 -409 831 -109
rect 897 -409 927 -109
rect 993 -409 1023 -109
rect 1089 -409 1119 -109
rect 1185 -409 1215 -109
rect 1281 -409 1311 -109
rect 1377 -409 1407 -109
rect 1473 -409 1503 -109
rect 1569 -409 1599 -109
rect 1665 -409 1695 -109
rect 1761 -409 1791 -109
rect 1857 -409 1887 -109
rect 1953 -409 1983 -109
rect 2049 -409 2079 -109
rect 2145 -409 2175 -109
rect 2241 -409 2271 -109
rect 2337 -409 2367 -109
<< ndiff >>
rect -2429 397 -2367 409
rect -2429 121 -2417 397
rect -2383 121 -2367 397
rect -2429 109 -2367 121
rect -2337 397 -2271 409
rect -2337 121 -2321 397
rect -2287 121 -2271 397
rect -2337 109 -2271 121
rect -2241 397 -2175 409
rect -2241 121 -2225 397
rect -2191 121 -2175 397
rect -2241 109 -2175 121
rect -2145 397 -2079 409
rect -2145 121 -2129 397
rect -2095 121 -2079 397
rect -2145 109 -2079 121
rect -2049 397 -1983 409
rect -2049 121 -2033 397
rect -1999 121 -1983 397
rect -2049 109 -1983 121
rect -1953 397 -1887 409
rect -1953 121 -1937 397
rect -1903 121 -1887 397
rect -1953 109 -1887 121
rect -1857 397 -1791 409
rect -1857 121 -1841 397
rect -1807 121 -1791 397
rect -1857 109 -1791 121
rect -1761 397 -1695 409
rect -1761 121 -1745 397
rect -1711 121 -1695 397
rect -1761 109 -1695 121
rect -1665 397 -1599 409
rect -1665 121 -1649 397
rect -1615 121 -1599 397
rect -1665 109 -1599 121
rect -1569 397 -1503 409
rect -1569 121 -1553 397
rect -1519 121 -1503 397
rect -1569 109 -1503 121
rect -1473 397 -1407 409
rect -1473 121 -1457 397
rect -1423 121 -1407 397
rect -1473 109 -1407 121
rect -1377 397 -1311 409
rect -1377 121 -1361 397
rect -1327 121 -1311 397
rect -1377 109 -1311 121
rect -1281 397 -1215 409
rect -1281 121 -1265 397
rect -1231 121 -1215 397
rect -1281 109 -1215 121
rect -1185 397 -1119 409
rect -1185 121 -1169 397
rect -1135 121 -1119 397
rect -1185 109 -1119 121
rect -1089 397 -1023 409
rect -1089 121 -1073 397
rect -1039 121 -1023 397
rect -1089 109 -1023 121
rect -993 397 -927 409
rect -993 121 -977 397
rect -943 121 -927 397
rect -993 109 -927 121
rect -897 397 -831 409
rect -897 121 -881 397
rect -847 121 -831 397
rect -897 109 -831 121
rect -801 397 -735 409
rect -801 121 -785 397
rect -751 121 -735 397
rect -801 109 -735 121
rect -705 397 -639 409
rect -705 121 -689 397
rect -655 121 -639 397
rect -705 109 -639 121
rect -609 397 -543 409
rect -609 121 -593 397
rect -559 121 -543 397
rect -609 109 -543 121
rect -513 397 -447 409
rect -513 121 -497 397
rect -463 121 -447 397
rect -513 109 -447 121
rect -417 397 -351 409
rect -417 121 -401 397
rect -367 121 -351 397
rect -417 109 -351 121
rect -321 397 -255 409
rect -321 121 -305 397
rect -271 121 -255 397
rect -321 109 -255 121
rect -225 397 -159 409
rect -225 121 -209 397
rect -175 121 -159 397
rect -225 109 -159 121
rect -129 397 -63 409
rect -129 121 -113 397
rect -79 121 -63 397
rect -129 109 -63 121
rect -33 397 33 409
rect -33 121 -17 397
rect 17 121 33 397
rect -33 109 33 121
rect 63 397 129 409
rect 63 121 79 397
rect 113 121 129 397
rect 63 109 129 121
rect 159 397 225 409
rect 159 121 175 397
rect 209 121 225 397
rect 159 109 225 121
rect 255 397 321 409
rect 255 121 271 397
rect 305 121 321 397
rect 255 109 321 121
rect 351 397 417 409
rect 351 121 367 397
rect 401 121 417 397
rect 351 109 417 121
rect 447 397 513 409
rect 447 121 463 397
rect 497 121 513 397
rect 447 109 513 121
rect 543 397 609 409
rect 543 121 559 397
rect 593 121 609 397
rect 543 109 609 121
rect 639 397 705 409
rect 639 121 655 397
rect 689 121 705 397
rect 639 109 705 121
rect 735 397 801 409
rect 735 121 751 397
rect 785 121 801 397
rect 735 109 801 121
rect 831 397 897 409
rect 831 121 847 397
rect 881 121 897 397
rect 831 109 897 121
rect 927 397 993 409
rect 927 121 943 397
rect 977 121 993 397
rect 927 109 993 121
rect 1023 397 1089 409
rect 1023 121 1039 397
rect 1073 121 1089 397
rect 1023 109 1089 121
rect 1119 397 1185 409
rect 1119 121 1135 397
rect 1169 121 1185 397
rect 1119 109 1185 121
rect 1215 397 1281 409
rect 1215 121 1231 397
rect 1265 121 1281 397
rect 1215 109 1281 121
rect 1311 397 1377 409
rect 1311 121 1327 397
rect 1361 121 1377 397
rect 1311 109 1377 121
rect 1407 397 1473 409
rect 1407 121 1423 397
rect 1457 121 1473 397
rect 1407 109 1473 121
rect 1503 397 1569 409
rect 1503 121 1519 397
rect 1553 121 1569 397
rect 1503 109 1569 121
rect 1599 397 1665 409
rect 1599 121 1615 397
rect 1649 121 1665 397
rect 1599 109 1665 121
rect 1695 397 1761 409
rect 1695 121 1711 397
rect 1745 121 1761 397
rect 1695 109 1761 121
rect 1791 397 1857 409
rect 1791 121 1807 397
rect 1841 121 1857 397
rect 1791 109 1857 121
rect 1887 397 1953 409
rect 1887 121 1903 397
rect 1937 121 1953 397
rect 1887 109 1953 121
rect 1983 397 2049 409
rect 1983 121 1999 397
rect 2033 121 2049 397
rect 1983 109 2049 121
rect 2079 397 2145 409
rect 2079 121 2095 397
rect 2129 121 2145 397
rect 2079 109 2145 121
rect 2175 397 2241 409
rect 2175 121 2191 397
rect 2225 121 2241 397
rect 2175 109 2241 121
rect 2271 397 2337 409
rect 2271 121 2287 397
rect 2321 121 2337 397
rect 2271 109 2337 121
rect 2367 397 2429 409
rect 2367 121 2383 397
rect 2417 121 2429 397
rect 2367 109 2429 121
rect -2429 -121 -2367 -109
rect -2429 -397 -2417 -121
rect -2383 -397 -2367 -121
rect -2429 -409 -2367 -397
rect -2337 -121 -2271 -109
rect -2337 -397 -2321 -121
rect -2287 -397 -2271 -121
rect -2337 -409 -2271 -397
rect -2241 -121 -2175 -109
rect -2241 -397 -2225 -121
rect -2191 -397 -2175 -121
rect -2241 -409 -2175 -397
rect -2145 -121 -2079 -109
rect -2145 -397 -2129 -121
rect -2095 -397 -2079 -121
rect -2145 -409 -2079 -397
rect -2049 -121 -1983 -109
rect -2049 -397 -2033 -121
rect -1999 -397 -1983 -121
rect -2049 -409 -1983 -397
rect -1953 -121 -1887 -109
rect -1953 -397 -1937 -121
rect -1903 -397 -1887 -121
rect -1953 -409 -1887 -397
rect -1857 -121 -1791 -109
rect -1857 -397 -1841 -121
rect -1807 -397 -1791 -121
rect -1857 -409 -1791 -397
rect -1761 -121 -1695 -109
rect -1761 -397 -1745 -121
rect -1711 -397 -1695 -121
rect -1761 -409 -1695 -397
rect -1665 -121 -1599 -109
rect -1665 -397 -1649 -121
rect -1615 -397 -1599 -121
rect -1665 -409 -1599 -397
rect -1569 -121 -1503 -109
rect -1569 -397 -1553 -121
rect -1519 -397 -1503 -121
rect -1569 -409 -1503 -397
rect -1473 -121 -1407 -109
rect -1473 -397 -1457 -121
rect -1423 -397 -1407 -121
rect -1473 -409 -1407 -397
rect -1377 -121 -1311 -109
rect -1377 -397 -1361 -121
rect -1327 -397 -1311 -121
rect -1377 -409 -1311 -397
rect -1281 -121 -1215 -109
rect -1281 -397 -1265 -121
rect -1231 -397 -1215 -121
rect -1281 -409 -1215 -397
rect -1185 -121 -1119 -109
rect -1185 -397 -1169 -121
rect -1135 -397 -1119 -121
rect -1185 -409 -1119 -397
rect -1089 -121 -1023 -109
rect -1089 -397 -1073 -121
rect -1039 -397 -1023 -121
rect -1089 -409 -1023 -397
rect -993 -121 -927 -109
rect -993 -397 -977 -121
rect -943 -397 -927 -121
rect -993 -409 -927 -397
rect -897 -121 -831 -109
rect -897 -397 -881 -121
rect -847 -397 -831 -121
rect -897 -409 -831 -397
rect -801 -121 -735 -109
rect -801 -397 -785 -121
rect -751 -397 -735 -121
rect -801 -409 -735 -397
rect -705 -121 -639 -109
rect -705 -397 -689 -121
rect -655 -397 -639 -121
rect -705 -409 -639 -397
rect -609 -121 -543 -109
rect -609 -397 -593 -121
rect -559 -397 -543 -121
rect -609 -409 -543 -397
rect -513 -121 -447 -109
rect -513 -397 -497 -121
rect -463 -397 -447 -121
rect -513 -409 -447 -397
rect -417 -121 -351 -109
rect -417 -397 -401 -121
rect -367 -397 -351 -121
rect -417 -409 -351 -397
rect -321 -121 -255 -109
rect -321 -397 -305 -121
rect -271 -397 -255 -121
rect -321 -409 -255 -397
rect -225 -121 -159 -109
rect -225 -397 -209 -121
rect -175 -397 -159 -121
rect -225 -409 -159 -397
rect -129 -121 -63 -109
rect -129 -397 -113 -121
rect -79 -397 -63 -121
rect -129 -409 -63 -397
rect -33 -121 33 -109
rect -33 -397 -17 -121
rect 17 -397 33 -121
rect -33 -409 33 -397
rect 63 -121 129 -109
rect 63 -397 79 -121
rect 113 -397 129 -121
rect 63 -409 129 -397
rect 159 -121 225 -109
rect 159 -397 175 -121
rect 209 -397 225 -121
rect 159 -409 225 -397
rect 255 -121 321 -109
rect 255 -397 271 -121
rect 305 -397 321 -121
rect 255 -409 321 -397
rect 351 -121 417 -109
rect 351 -397 367 -121
rect 401 -397 417 -121
rect 351 -409 417 -397
rect 447 -121 513 -109
rect 447 -397 463 -121
rect 497 -397 513 -121
rect 447 -409 513 -397
rect 543 -121 609 -109
rect 543 -397 559 -121
rect 593 -397 609 -121
rect 543 -409 609 -397
rect 639 -121 705 -109
rect 639 -397 655 -121
rect 689 -397 705 -121
rect 639 -409 705 -397
rect 735 -121 801 -109
rect 735 -397 751 -121
rect 785 -397 801 -121
rect 735 -409 801 -397
rect 831 -121 897 -109
rect 831 -397 847 -121
rect 881 -397 897 -121
rect 831 -409 897 -397
rect 927 -121 993 -109
rect 927 -397 943 -121
rect 977 -397 993 -121
rect 927 -409 993 -397
rect 1023 -121 1089 -109
rect 1023 -397 1039 -121
rect 1073 -397 1089 -121
rect 1023 -409 1089 -397
rect 1119 -121 1185 -109
rect 1119 -397 1135 -121
rect 1169 -397 1185 -121
rect 1119 -409 1185 -397
rect 1215 -121 1281 -109
rect 1215 -397 1231 -121
rect 1265 -397 1281 -121
rect 1215 -409 1281 -397
rect 1311 -121 1377 -109
rect 1311 -397 1327 -121
rect 1361 -397 1377 -121
rect 1311 -409 1377 -397
rect 1407 -121 1473 -109
rect 1407 -397 1423 -121
rect 1457 -397 1473 -121
rect 1407 -409 1473 -397
rect 1503 -121 1569 -109
rect 1503 -397 1519 -121
rect 1553 -397 1569 -121
rect 1503 -409 1569 -397
rect 1599 -121 1665 -109
rect 1599 -397 1615 -121
rect 1649 -397 1665 -121
rect 1599 -409 1665 -397
rect 1695 -121 1761 -109
rect 1695 -397 1711 -121
rect 1745 -397 1761 -121
rect 1695 -409 1761 -397
rect 1791 -121 1857 -109
rect 1791 -397 1807 -121
rect 1841 -397 1857 -121
rect 1791 -409 1857 -397
rect 1887 -121 1953 -109
rect 1887 -397 1903 -121
rect 1937 -397 1953 -121
rect 1887 -409 1953 -397
rect 1983 -121 2049 -109
rect 1983 -397 1999 -121
rect 2033 -397 2049 -121
rect 1983 -409 2049 -397
rect 2079 -121 2145 -109
rect 2079 -397 2095 -121
rect 2129 -397 2145 -121
rect 2079 -409 2145 -397
rect 2175 -121 2241 -109
rect 2175 -397 2191 -121
rect 2225 -397 2241 -121
rect 2175 -409 2241 -397
rect 2271 -121 2337 -109
rect 2271 -397 2287 -121
rect 2321 -397 2337 -121
rect 2271 -409 2337 -397
rect 2367 -121 2429 -109
rect 2367 -397 2383 -121
rect 2417 -397 2429 -121
rect 2367 -409 2429 -397
<< ndiffc >>
rect -2417 121 -2383 397
rect -2321 121 -2287 397
rect -2225 121 -2191 397
rect -2129 121 -2095 397
rect -2033 121 -1999 397
rect -1937 121 -1903 397
rect -1841 121 -1807 397
rect -1745 121 -1711 397
rect -1649 121 -1615 397
rect -1553 121 -1519 397
rect -1457 121 -1423 397
rect -1361 121 -1327 397
rect -1265 121 -1231 397
rect -1169 121 -1135 397
rect -1073 121 -1039 397
rect -977 121 -943 397
rect -881 121 -847 397
rect -785 121 -751 397
rect -689 121 -655 397
rect -593 121 -559 397
rect -497 121 -463 397
rect -401 121 -367 397
rect -305 121 -271 397
rect -209 121 -175 397
rect -113 121 -79 397
rect -17 121 17 397
rect 79 121 113 397
rect 175 121 209 397
rect 271 121 305 397
rect 367 121 401 397
rect 463 121 497 397
rect 559 121 593 397
rect 655 121 689 397
rect 751 121 785 397
rect 847 121 881 397
rect 943 121 977 397
rect 1039 121 1073 397
rect 1135 121 1169 397
rect 1231 121 1265 397
rect 1327 121 1361 397
rect 1423 121 1457 397
rect 1519 121 1553 397
rect 1615 121 1649 397
rect 1711 121 1745 397
rect 1807 121 1841 397
rect 1903 121 1937 397
rect 1999 121 2033 397
rect 2095 121 2129 397
rect 2191 121 2225 397
rect 2287 121 2321 397
rect 2383 121 2417 397
rect -2417 -397 -2383 -121
rect -2321 -397 -2287 -121
rect -2225 -397 -2191 -121
rect -2129 -397 -2095 -121
rect -2033 -397 -1999 -121
rect -1937 -397 -1903 -121
rect -1841 -397 -1807 -121
rect -1745 -397 -1711 -121
rect -1649 -397 -1615 -121
rect -1553 -397 -1519 -121
rect -1457 -397 -1423 -121
rect -1361 -397 -1327 -121
rect -1265 -397 -1231 -121
rect -1169 -397 -1135 -121
rect -1073 -397 -1039 -121
rect -977 -397 -943 -121
rect -881 -397 -847 -121
rect -785 -397 -751 -121
rect -689 -397 -655 -121
rect -593 -397 -559 -121
rect -497 -397 -463 -121
rect -401 -397 -367 -121
rect -305 -397 -271 -121
rect -209 -397 -175 -121
rect -113 -397 -79 -121
rect -17 -397 17 -121
rect 79 -397 113 -121
rect 175 -397 209 -121
rect 271 -397 305 -121
rect 367 -397 401 -121
rect 463 -397 497 -121
rect 559 -397 593 -121
rect 655 -397 689 -121
rect 751 -397 785 -121
rect 847 -397 881 -121
rect 943 -397 977 -121
rect 1039 -397 1073 -121
rect 1135 -397 1169 -121
rect 1231 -397 1265 -121
rect 1327 -397 1361 -121
rect 1423 -397 1457 -121
rect 1519 -397 1553 -121
rect 1615 -397 1649 -121
rect 1711 -397 1745 -121
rect 1807 -397 1841 -121
rect 1903 -397 1937 -121
rect 1999 -397 2033 -121
rect 2095 -397 2129 -121
rect 2191 -397 2225 -121
rect 2287 -397 2321 -121
rect 2383 -397 2417 -121
<< psubdiff >>
rect -2531 549 -2435 583
rect 2435 549 2531 583
rect -2531 487 -2497 549
rect 2497 487 2531 549
rect -2531 -549 -2497 -487
rect 2497 -549 2531 -487
rect -2531 -583 -2435 -549
rect 2435 -583 2531 -549
<< psubdiffcont >>
rect -2435 549 2435 583
rect -2531 -487 -2497 487
rect 2497 -487 2531 487
rect -2435 -583 2435 -549
<< poly >>
rect -2385 481 -2319 497
rect -2385 447 -2369 481
rect -2335 447 -2319 481
rect -2385 431 -2319 447
rect -2193 481 -2127 497
rect -2193 447 -2177 481
rect -2143 447 -2127 481
rect -2367 409 -2337 431
rect -2271 409 -2241 435
rect -2193 431 -2127 447
rect -2001 481 -1935 497
rect -2001 447 -1985 481
rect -1951 447 -1935 481
rect -2175 409 -2145 431
rect -2079 409 -2049 435
rect -2001 431 -1935 447
rect -1809 481 -1743 497
rect -1809 447 -1793 481
rect -1759 447 -1743 481
rect -1983 409 -1953 431
rect -1887 409 -1857 435
rect -1809 431 -1743 447
rect -1617 481 -1551 497
rect -1617 447 -1601 481
rect -1567 447 -1551 481
rect -1791 409 -1761 431
rect -1695 409 -1665 435
rect -1617 431 -1551 447
rect -1425 481 -1359 497
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1599 409 -1569 431
rect -1503 409 -1473 435
rect -1425 431 -1359 447
rect -1233 481 -1167 497
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1407 409 -1377 431
rect -1311 409 -1281 435
rect -1233 431 -1167 447
rect -1041 481 -975 497
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -1215 409 -1185 431
rect -1119 409 -1089 435
rect -1041 431 -975 447
rect -849 481 -783 497
rect -849 447 -833 481
rect -799 447 -783 481
rect -1023 409 -993 431
rect -927 409 -897 435
rect -849 431 -783 447
rect -657 481 -591 497
rect -657 447 -641 481
rect -607 447 -591 481
rect -831 409 -801 431
rect -735 409 -705 435
rect -657 431 -591 447
rect -465 481 -399 497
rect -465 447 -449 481
rect -415 447 -399 481
rect -639 409 -609 431
rect -543 409 -513 435
rect -465 431 -399 447
rect -273 481 -207 497
rect -273 447 -257 481
rect -223 447 -207 481
rect -447 409 -417 431
rect -351 409 -321 435
rect -273 431 -207 447
rect -81 481 -15 497
rect -81 447 -65 481
rect -31 447 -15 481
rect -255 409 -225 431
rect -159 409 -129 435
rect -81 431 -15 447
rect 111 481 177 497
rect 111 447 127 481
rect 161 447 177 481
rect -63 409 -33 431
rect 33 409 63 435
rect 111 431 177 447
rect 303 481 369 497
rect 303 447 319 481
rect 353 447 369 481
rect 129 409 159 431
rect 225 409 255 435
rect 303 431 369 447
rect 495 481 561 497
rect 495 447 511 481
rect 545 447 561 481
rect 321 409 351 431
rect 417 409 447 435
rect 495 431 561 447
rect 687 481 753 497
rect 687 447 703 481
rect 737 447 753 481
rect 513 409 543 431
rect 609 409 639 435
rect 687 431 753 447
rect 879 481 945 497
rect 879 447 895 481
rect 929 447 945 481
rect 705 409 735 431
rect 801 409 831 435
rect 879 431 945 447
rect 1071 481 1137 497
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 897 409 927 431
rect 993 409 1023 435
rect 1071 431 1137 447
rect 1263 481 1329 497
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1089 409 1119 431
rect 1185 409 1215 435
rect 1263 431 1329 447
rect 1455 481 1521 497
rect 1455 447 1471 481
rect 1505 447 1521 481
rect 1281 409 1311 431
rect 1377 409 1407 435
rect 1455 431 1521 447
rect 1647 481 1713 497
rect 1647 447 1663 481
rect 1697 447 1713 481
rect 1473 409 1503 431
rect 1569 409 1599 435
rect 1647 431 1713 447
rect 1839 481 1905 497
rect 1839 447 1855 481
rect 1889 447 1905 481
rect 1665 409 1695 431
rect 1761 409 1791 435
rect 1839 431 1905 447
rect 2031 481 2097 497
rect 2031 447 2047 481
rect 2081 447 2097 481
rect 1857 409 1887 431
rect 1953 409 1983 435
rect 2031 431 2097 447
rect 2223 481 2289 497
rect 2223 447 2239 481
rect 2273 447 2289 481
rect 2049 409 2079 431
rect 2145 409 2175 435
rect 2223 431 2289 447
rect 2241 409 2271 431
rect 2337 409 2367 435
rect -2367 83 -2337 109
rect -2271 87 -2241 109
rect -2289 71 -2223 87
rect -2175 83 -2145 109
rect -2079 87 -2049 109
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2289 21 -2223 37
rect -2097 71 -2031 87
rect -1983 83 -1953 109
rect -1887 87 -1857 109
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -2097 21 -2031 37
rect -1905 71 -1839 87
rect -1791 83 -1761 109
rect -1695 87 -1665 109
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1905 21 -1839 37
rect -1713 71 -1647 87
rect -1599 83 -1569 109
rect -1503 87 -1473 109
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1713 21 -1647 37
rect -1521 71 -1455 87
rect -1407 83 -1377 109
rect -1311 87 -1281 109
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1521 21 -1455 37
rect -1329 71 -1263 87
rect -1215 83 -1185 109
rect -1119 87 -1089 109
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1329 21 -1263 37
rect -1137 71 -1071 87
rect -1023 83 -993 109
rect -927 87 -897 109
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -1137 21 -1071 37
rect -945 71 -879 87
rect -831 83 -801 109
rect -735 87 -705 109
rect -945 37 -929 71
rect -895 37 -879 71
rect -945 21 -879 37
rect -753 71 -687 87
rect -639 83 -609 109
rect -543 87 -513 109
rect -753 37 -737 71
rect -703 37 -687 71
rect -753 21 -687 37
rect -561 71 -495 87
rect -447 83 -417 109
rect -351 87 -321 109
rect -561 37 -545 71
rect -511 37 -495 71
rect -561 21 -495 37
rect -369 71 -303 87
rect -255 83 -225 109
rect -159 87 -129 109
rect -369 37 -353 71
rect -319 37 -303 71
rect -369 21 -303 37
rect -177 71 -111 87
rect -63 83 -33 109
rect 33 87 63 109
rect -177 37 -161 71
rect -127 37 -111 71
rect -177 21 -111 37
rect 15 71 81 87
rect 129 83 159 109
rect 225 87 255 109
rect 15 37 31 71
rect 65 37 81 71
rect 15 21 81 37
rect 207 71 273 87
rect 321 83 351 109
rect 417 87 447 109
rect 207 37 223 71
rect 257 37 273 71
rect 207 21 273 37
rect 399 71 465 87
rect 513 83 543 109
rect 609 87 639 109
rect 399 37 415 71
rect 449 37 465 71
rect 399 21 465 37
rect 591 71 657 87
rect 705 83 735 109
rect 801 87 831 109
rect 591 37 607 71
rect 641 37 657 71
rect 591 21 657 37
rect 783 71 849 87
rect 897 83 927 109
rect 993 87 1023 109
rect 783 37 799 71
rect 833 37 849 71
rect 783 21 849 37
rect 975 71 1041 87
rect 1089 83 1119 109
rect 1185 87 1215 109
rect 975 37 991 71
rect 1025 37 1041 71
rect 975 21 1041 37
rect 1167 71 1233 87
rect 1281 83 1311 109
rect 1377 87 1407 109
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1167 21 1233 37
rect 1359 71 1425 87
rect 1473 83 1503 109
rect 1569 87 1599 109
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1359 21 1425 37
rect 1551 71 1617 87
rect 1665 83 1695 109
rect 1761 87 1791 109
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1551 21 1617 37
rect 1743 71 1809 87
rect 1857 83 1887 109
rect 1953 87 1983 109
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1743 21 1809 37
rect 1935 71 2001 87
rect 2049 83 2079 109
rect 2145 87 2175 109
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 1935 21 2001 37
rect 2127 71 2193 87
rect 2241 83 2271 109
rect 2337 87 2367 109
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2127 21 2193 37
rect 2319 71 2385 87
rect 2319 37 2335 71
rect 2369 37 2385 71
rect 2319 21 2385 37
rect -2289 -37 -2223 -21
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2367 -109 -2337 -83
rect -2289 -87 -2223 -71
rect -2097 -37 -2031 -21
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -2271 -109 -2241 -87
rect -2175 -109 -2145 -83
rect -2097 -87 -2031 -71
rect -1905 -37 -1839 -21
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -2079 -109 -2049 -87
rect -1983 -109 -1953 -83
rect -1905 -87 -1839 -71
rect -1713 -37 -1647 -21
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1887 -109 -1857 -87
rect -1791 -109 -1761 -83
rect -1713 -87 -1647 -71
rect -1521 -37 -1455 -21
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1695 -109 -1665 -87
rect -1599 -109 -1569 -83
rect -1521 -87 -1455 -71
rect -1329 -37 -1263 -21
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1503 -109 -1473 -87
rect -1407 -109 -1377 -83
rect -1329 -87 -1263 -71
rect -1137 -37 -1071 -21
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -1311 -109 -1281 -87
rect -1215 -109 -1185 -83
rect -1137 -87 -1071 -71
rect -945 -37 -879 -21
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -1119 -109 -1089 -87
rect -1023 -109 -993 -83
rect -945 -87 -879 -71
rect -753 -37 -687 -21
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -927 -109 -897 -87
rect -831 -109 -801 -83
rect -753 -87 -687 -71
rect -561 -37 -495 -21
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -735 -109 -705 -87
rect -639 -109 -609 -83
rect -561 -87 -495 -71
rect -369 -37 -303 -21
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -543 -109 -513 -87
rect -447 -109 -417 -83
rect -369 -87 -303 -71
rect -177 -37 -111 -21
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect -351 -109 -321 -87
rect -255 -109 -225 -83
rect -177 -87 -111 -71
rect 15 -37 81 -21
rect 15 -71 31 -37
rect 65 -71 81 -37
rect -159 -109 -129 -87
rect -63 -109 -33 -83
rect 15 -87 81 -71
rect 207 -37 273 -21
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 33 -109 63 -87
rect 129 -109 159 -83
rect 207 -87 273 -71
rect 399 -37 465 -21
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 225 -109 255 -87
rect 321 -109 351 -83
rect 399 -87 465 -71
rect 591 -37 657 -21
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 417 -109 447 -87
rect 513 -109 543 -83
rect 591 -87 657 -71
rect 783 -37 849 -21
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 609 -109 639 -87
rect 705 -109 735 -83
rect 783 -87 849 -71
rect 975 -37 1041 -21
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 801 -109 831 -87
rect 897 -109 927 -83
rect 975 -87 1041 -71
rect 1167 -37 1233 -21
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 993 -109 1023 -87
rect 1089 -109 1119 -83
rect 1167 -87 1233 -71
rect 1359 -37 1425 -21
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1185 -109 1215 -87
rect 1281 -109 1311 -83
rect 1359 -87 1425 -71
rect 1551 -37 1617 -21
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1377 -109 1407 -87
rect 1473 -109 1503 -83
rect 1551 -87 1617 -71
rect 1743 -37 1809 -21
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1569 -109 1599 -87
rect 1665 -109 1695 -83
rect 1743 -87 1809 -71
rect 1935 -37 2001 -21
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 1761 -109 1791 -87
rect 1857 -109 1887 -83
rect 1935 -87 2001 -71
rect 2127 -37 2193 -21
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 1953 -109 1983 -87
rect 2049 -109 2079 -83
rect 2127 -87 2193 -71
rect 2319 -37 2385 -21
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect 2145 -109 2175 -87
rect 2241 -109 2271 -83
rect 2319 -87 2385 -71
rect 2337 -109 2367 -87
rect -2367 -431 -2337 -409
rect -2385 -447 -2319 -431
rect -2271 -435 -2241 -409
rect -2175 -431 -2145 -409
rect -2385 -481 -2369 -447
rect -2335 -481 -2319 -447
rect -2385 -497 -2319 -481
rect -2193 -447 -2127 -431
rect -2079 -435 -2049 -409
rect -1983 -431 -1953 -409
rect -2193 -481 -2177 -447
rect -2143 -481 -2127 -447
rect -2193 -497 -2127 -481
rect -2001 -447 -1935 -431
rect -1887 -435 -1857 -409
rect -1791 -431 -1761 -409
rect -2001 -481 -1985 -447
rect -1951 -481 -1935 -447
rect -2001 -497 -1935 -481
rect -1809 -447 -1743 -431
rect -1695 -435 -1665 -409
rect -1599 -431 -1569 -409
rect -1809 -481 -1793 -447
rect -1759 -481 -1743 -447
rect -1809 -497 -1743 -481
rect -1617 -447 -1551 -431
rect -1503 -435 -1473 -409
rect -1407 -431 -1377 -409
rect -1617 -481 -1601 -447
rect -1567 -481 -1551 -447
rect -1617 -497 -1551 -481
rect -1425 -447 -1359 -431
rect -1311 -435 -1281 -409
rect -1215 -431 -1185 -409
rect -1425 -481 -1409 -447
rect -1375 -481 -1359 -447
rect -1425 -497 -1359 -481
rect -1233 -447 -1167 -431
rect -1119 -435 -1089 -409
rect -1023 -431 -993 -409
rect -1233 -481 -1217 -447
rect -1183 -481 -1167 -447
rect -1233 -497 -1167 -481
rect -1041 -447 -975 -431
rect -927 -435 -897 -409
rect -831 -431 -801 -409
rect -1041 -481 -1025 -447
rect -991 -481 -975 -447
rect -1041 -497 -975 -481
rect -849 -447 -783 -431
rect -735 -435 -705 -409
rect -639 -431 -609 -409
rect -849 -481 -833 -447
rect -799 -481 -783 -447
rect -849 -497 -783 -481
rect -657 -447 -591 -431
rect -543 -435 -513 -409
rect -447 -431 -417 -409
rect -657 -481 -641 -447
rect -607 -481 -591 -447
rect -657 -497 -591 -481
rect -465 -447 -399 -431
rect -351 -435 -321 -409
rect -255 -431 -225 -409
rect -465 -481 -449 -447
rect -415 -481 -399 -447
rect -465 -497 -399 -481
rect -273 -447 -207 -431
rect -159 -435 -129 -409
rect -63 -431 -33 -409
rect -273 -481 -257 -447
rect -223 -481 -207 -447
rect -273 -497 -207 -481
rect -81 -447 -15 -431
rect 33 -435 63 -409
rect 129 -431 159 -409
rect -81 -481 -65 -447
rect -31 -481 -15 -447
rect -81 -497 -15 -481
rect 111 -447 177 -431
rect 225 -435 255 -409
rect 321 -431 351 -409
rect 111 -481 127 -447
rect 161 -481 177 -447
rect 111 -497 177 -481
rect 303 -447 369 -431
rect 417 -435 447 -409
rect 513 -431 543 -409
rect 303 -481 319 -447
rect 353 -481 369 -447
rect 303 -497 369 -481
rect 495 -447 561 -431
rect 609 -435 639 -409
rect 705 -431 735 -409
rect 495 -481 511 -447
rect 545 -481 561 -447
rect 495 -497 561 -481
rect 687 -447 753 -431
rect 801 -435 831 -409
rect 897 -431 927 -409
rect 687 -481 703 -447
rect 737 -481 753 -447
rect 687 -497 753 -481
rect 879 -447 945 -431
rect 993 -435 1023 -409
rect 1089 -431 1119 -409
rect 879 -481 895 -447
rect 929 -481 945 -447
rect 879 -497 945 -481
rect 1071 -447 1137 -431
rect 1185 -435 1215 -409
rect 1281 -431 1311 -409
rect 1071 -481 1087 -447
rect 1121 -481 1137 -447
rect 1071 -497 1137 -481
rect 1263 -447 1329 -431
rect 1377 -435 1407 -409
rect 1473 -431 1503 -409
rect 1263 -481 1279 -447
rect 1313 -481 1329 -447
rect 1263 -497 1329 -481
rect 1455 -447 1521 -431
rect 1569 -435 1599 -409
rect 1665 -431 1695 -409
rect 1455 -481 1471 -447
rect 1505 -481 1521 -447
rect 1455 -497 1521 -481
rect 1647 -447 1713 -431
rect 1761 -435 1791 -409
rect 1857 -431 1887 -409
rect 1647 -481 1663 -447
rect 1697 -481 1713 -447
rect 1647 -497 1713 -481
rect 1839 -447 1905 -431
rect 1953 -435 1983 -409
rect 2049 -431 2079 -409
rect 1839 -481 1855 -447
rect 1889 -481 1905 -447
rect 1839 -497 1905 -481
rect 2031 -447 2097 -431
rect 2145 -435 2175 -409
rect 2241 -431 2271 -409
rect 2031 -481 2047 -447
rect 2081 -481 2097 -447
rect 2031 -497 2097 -481
rect 2223 -447 2289 -431
rect 2337 -435 2367 -409
rect 2223 -481 2239 -447
rect 2273 -481 2289 -447
rect 2223 -497 2289 -481
<< polycont >>
rect -2369 447 -2335 481
rect -2177 447 -2143 481
rect -1985 447 -1951 481
rect -1793 447 -1759 481
rect -1601 447 -1567 481
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect 1663 447 1697 481
rect 1855 447 1889 481
rect 2047 447 2081 481
rect 2239 447 2273 481
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect -2369 -481 -2335 -447
rect -2177 -481 -2143 -447
rect -1985 -481 -1951 -447
rect -1793 -481 -1759 -447
rect -1601 -481 -1567 -447
rect -1409 -481 -1375 -447
rect -1217 -481 -1183 -447
rect -1025 -481 -991 -447
rect -833 -481 -799 -447
rect -641 -481 -607 -447
rect -449 -481 -415 -447
rect -257 -481 -223 -447
rect -65 -481 -31 -447
rect 127 -481 161 -447
rect 319 -481 353 -447
rect 511 -481 545 -447
rect 703 -481 737 -447
rect 895 -481 929 -447
rect 1087 -481 1121 -447
rect 1279 -481 1313 -447
rect 1471 -481 1505 -447
rect 1663 -481 1697 -447
rect 1855 -481 1889 -447
rect 2047 -481 2081 -447
rect 2239 -481 2273 -447
<< locali >>
rect -2531 549 -2435 583
rect 2435 549 2531 583
rect -2531 487 -2497 549
rect 2497 487 2531 549
rect -2385 447 -2369 481
rect -2335 447 -2319 481
rect -2193 447 -2177 481
rect -2143 447 -2127 481
rect -2001 447 -1985 481
rect -1951 447 -1935 481
rect -1809 447 -1793 481
rect -1759 447 -1743 481
rect -1617 447 -1601 481
rect -1567 447 -1551 481
rect -1425 447 -1409 481
rect -1375 447 -1359 481
rect -1233 447 -1217 481
rect -1183 447 -1167 481
rect -1041 447 -1025 481
rect -991 447 -975 481
rect -849 447 -833 481
rect -799 447 -783 481
rect -657 447 -641 481
rect -607 447 -591 481
rect -465 447 -449 481
rect -415 447 -399 481
rect -273 447 -257 481
rect -223 447 -207 481
rect -81 447 -65 481
rect -31 447 -15 481
rect 111 447 127 481
rect 161 447 177 481
rect 303 447 319 481
rect 353 447 369 481
rect 495 447 511 481
rect 545 447 561 481
rect 687 447 703 481
rect 737 447 753 481
rect 879 447 895 481
rect 929 447 945 481
rect 1071 447 1087 481
rect 1121 447 1137 481
rect 1263 447 1279 481
rect 1313 447 1329 481
rect 1455 447 1471 481
rect 1505 447 1521 481
rect 1647 447 1663 481
rect 1697 447 1713 481
rect 1839 447 1855 481
rect 1889 447 1905 481
rect 2031 447 2047 481
rect 2081 447 2097 481
rect 2223 447 2239 481
rect 2273 447 2289 481
rect -2417 397 -2383 413
rect -2417 105 -2383 121
rect -2321 397 -2287 413
rect -2321 105 -2287 121
rect -2225 397 -2191 413
rect -2225 105 -2191 121
rect -2129 397 -2095 413
rect -2129 105 -2095 121
rect -2033 397 -1999 413
rect -2033 105 -1999 121
rect -1937 397 -1903 413
rect -1937 105 -1903 121
rect -1841 397 -1807 413
rect -1841 105 -1807 121
rect -1745 397 -1711 413
rect -1745 105 -1711 121
rect -1649 397 -1615 413
rect -1649 105 -1615 121
rect -1553 397 -1519 413
rect -1553 105 -1519 121
rect -1457 397 -1423 413
rect -1457 105 -1423 121
rect -1361 397 -1327 413
rect -1361 105 -1327 121
rect -1265 397 -1231 413
rect -1265 105 -1231 121
rect -1169 397 -1135 413
rect -1169 105 -1135 121
rect -1073 397 -1039 413
rect -1073 105 -1039 121
rect -977 397 -943 413
rect -977 105 -943 121
rect -881 397 -847 413
rect -881 105 -847 121
rect -785 397 -751 413
rect -785 105 -751 121
rect -689 397 -655 413
rect -689 105 -655 121
rect -593 397 -559 413
rect -593 105 -559 121
rect -497 397 -463 413
rect -497 105 -463 121
rect -401 397 -367 413
rect -401 105 -367 121
rect -305 397 -271 413
rect -305 105 -271 121
rect -209 397 -175 413
rect -209 105 -175 121
rect -113 397 -79 413
rect -113 105 -79 121
rect -17 397 17 413
rect -17 105 17 121
rect 79 397 113 413
rect 79 105 113 121
rect 175 397 209 413
rect 175 105 209 121
rect 271 397 305 413
rect 271 105 305 121
rect 367 397 401 413
rect 367 105 401 121
rect 463 397 497 413
rect 463 105 497 121
rect 559 397 593 413
rect 559 105 593 121
rect 655 397 689 413
rect 655 105 689 121
rect 751 397 785 413
rect 751 105 785 121
rect 847 397 881 413
rect 847 105 881 121
rect 943 397 977 413
rect 943 105 977 121
rect 1039 397 1073 413
rect 1039 105 1073 121
rect 1135 397 1169 413
rect 1135 105 1169 121
rect 1231 397 1265 413
rect 1231 105 1265 121
rect 1327 397 1361 413
rect 1327 105 1361 121
rect 1423 397 1457 413
rect 1423 105 1457 121
rect 1519 397 1553 413
rect 1519 105 1553 121
rect 1615 397 1649 413
rect 1615 105 1649 121
rect 1711 397 1745 413
rect 1711 105 1745 121
rect 1807 397 1841 413
rect 1807 105 1841 121
rect 1903 397 1937 413
rect 1903 105 1937 121
rect 1999 397 2033 413
rect 1999 105 2033 121
rect 2095 397 2129 413
rect 2095 105 2129 121
rect 2191 397 2225 413
rect 2191 105 2225 121
rect 2287 397 2321 413
rect 2287 105 2321 121
rect 2383 397 2417 413
rect 2383 105 2417 121
rect -2289 37 -2273 71
rect -2239 37 -2223 71
rect -2097 37 -2081 71
rect -2047 37 -2031 71
rect -1905 37 -1889 71
rect -1855 37 -1839 71
rect -1713 37 -1697 71
rect -1663 37 -1647 71
rect -1521 37 -1505 71
rect -1471 37 -1455 71
rect -1329 37 -1313 71
rect -1279 37 -1263 71
rect -1137 37 -1121 71
rect -1087 37 -1071 71
rect -945 37 -929 71
rect -895 37 -879 71
rect -753 37 -737 71
rect -703 37 -687 71
rect -561 37 -545 71
rect -511 37 -495 71
rect -369 37 -353 71
rect -319 37 -303 71
rect -177 37 -161 71
rect -127 37 -111 71
rect 15 37 31 71
rect 65 37 81 71
rect 207 37 223 71
rect 257 37 273 71
rect 399 37 415 71
rect 449 37 465 71
rect 591 37 607 71
rect 641 37 657 71
rect 783 37 799 71
rect 833 37 849 71
rect 975 37 991 71
rect 1025 37 1041 71
rect 1167 37 1183 71
rect 1217 37 1233 71
rect 1359 37 1375 71
rect 1409 37 1425 71
rect 1551 37 1567 71
rect 1601 37 1617 71
rect 1743 37 1759 71
rect 1793 37 1809 71
rect 1935 37 1951 71
rect 1985 37 2001 71
rect 2127 37 2143 71
rect 2177 37 2193 71
rect 2319 37 2335 71
rect 2369 37 2385 71
rect -2289 -71 -2273 -37
rect -2239 -71 -2223 -37
rect -2097 -71 -2081 -37
rect -2047 -71 -2031 -37
rect -1905 -71 -1889 -37
rect -1855 -71 -1839 -37
rect -1713 -71 -1697 -37
rect -1663 -71 -1647 -37
rect -1521 -71 -1505 -37
rect -1471 -71 -1455 -37
rect -1329 -71 -1313 -37
rect -1279 -71 -1263 -37
rect -1137 -71 -1121 -37
rect -1087 -71 -1071 -37
rect -945 -71 -929 -37
rect -895 -71 -879 -37
rect -753 -71 -737 -37
rect -703 -71 -687 -37
rect -561 -71 -545 -37
rect -511 -71 -495 -37
rect -369 -71 -353 -37
rect -319 -71 -303 -37
rect -177 -71 -161 -37
rect -127 -71 -111 -37
rect 15 -71 31 -37
rect 65 -71 81 -37
rect 207 -71 223 -37
rect 257 -71 273 -37
rect 399 -71 415 -37
rect 449 -71 465 -37
rect 591 -71 607 -37
rect 641 -71 657 -37
rect 783 -71 799 -37
rect 833 -71 849 -37
rect 975 -71 991 -37
rect 1025 -71 1041 -37
rect 1167 -71 1183 -37
rect 1217 -71 1233 -37
rect 1359 -71 1375 -37
rect 1409 -71 1425 -37
rect 1551 -71 1567 -37
rect 1601 -71 1617 -37
rect 1743 -71 1759 -37
rect 1793 -71 1809 -37
rect 1935 -71 1951 -37
rect 1985 -71 2001 -37
rect 2127 -71 2143 -37
rect 2177 -71 2193 -37
rect 2319 -71 2335 -37
rect 2369 -71 2385 -37
rect -2417 -121 -2383 -105
rect -2417 -413 -2383 -397
rect -2321 -121 -2287 -105
rect -2321 -413 -2287 -397
rect -2225 -121 -2191 -105
rect -2225 -413 -2191 -397
rect -2129 -121 -2095 -105
rect -2129 -413 -2095 -397
rect -2033 -121 -1999 -105
rect -2033 -413 -1999 -397
rect -1937 -121 -1903 -105
rect -1937 -413 -1903 -397
rect -1841 -121 -1807 -105
rect -1841 -413 -1807 -397
rect -1745 -121 -1711 -105
rect -1745 -413 -1711 -397
rect -1649 -121 -1615 -105
rect -1649 -413 -1615 -397
rect -1553 -121 -1519 -105
rect -1553 -413 -1519 -397
rect -1457 -121 -1423 -105
rect -1457 -413 -1423 -397
rect -1361 -121 -1327 -105
rect -1361 -413 -1327 -397
rect -1265 -121 -1231 -105
rect -1265 -413 -1231 -397
rect -1169 -121 -1135 -105
rect -1169 -413 -1135 -397
rect -1073 -121 -1039 -105
rect -1073 -413 -1039 -397
rect -977 -121 -943 -105
rect -977 -413 -943 -397
rect -881 -121 -847 -105
rect -881 -413 -847 -397
rect -785 -121 -751 -105
rect -785 -413 -751 -397
rect -689 -121 -655 -105
rect -689 -413 -655 -397
rect -593 -121 -559 -105
rect -593 -413 -559 -397
rect -497 -121 -463 -105
rect -497 -413 -463 -397
rect -401 -121 -367 -105
rect -401 -413 -367 -397
rect -305 -121 -271 -105
rect -305 -413 -271 -397
rect -209 -121 -175 -105
rect -209 -413 -175 -397
rect -113 -121 -79 -105
rect -113 -413 -79 -397
rect -17 -121 17 -105
rect -17 -413 17 -397
rect 79 -121 113 -105
rect 79 -413 113 -397
rect 175 -121 209 -105
rect 175 -413 209 -397
rect 271 -121 305 -105
rect 271 -413 305 -397
rect 367 -121 401 -105
rect 367 -413 401 -397
rect 463 -121 497 -105
rect 463 -413 497 -397
rect 559 -121 593 -105
rect 559 -413 593 -397
rect 655 -121 689 -105
rect 655 -413 689 -397
rect 751 -121 785 -105
rect 751 -413 785 -397
rect 847 -121 881 -105
rect 847 -413 881 -397
rect 943 -121 977 -105
rect 943 -413 977 -397
rect 1039 -121 1073 -105
rect 1039 -413 1073 -397
rect 1135 -121 1169 -105
rect 1135 -413 1169 -397
rect 1231 -121 1265 -105
rect 1231 -413 1265 -397
rect 1327 -121 1361 -105
rect 1327 -413 1361 -397
rect 1423 -121 1457 -105
rect 1423 -413 1457 -397
rect 1519 -121 1553 -105
rect 1519 -413 1553 -397
rect 1615 -121 1649 -105
rect 1615 -413 1649 -397
rect 1711 -121 1745 -105
rect 1711 -413 1745 -397
rect 1807 -121 1841 -105
rect 1807 -413 1841 -397
rect 1903 -121 1937 -105
rect 1903 -413 1937 -397
rect 1999 -121 2033 -105
rect 1999 -413 2033 -397
rect 2095 -121 2129 -105
rect 2095 -413 2129 -397
rect 2191 -121 2225 -105
rect 2191 -413 2225 -397
rect 2287 -121 2321 -105
rect 2287 -413 2321 -397
rect 2383 -121 2417 -105
rect 2383 -413 2417 -397
rect -2385 -481 -2369 -447
rect -2335 -481 -2319 -447
rect -2193 -481 -2177 -447
rect -2143 -481 -2127 -447
rect -2001 -481 -1985 -447
rect -1951 -481 -1935 -447
rect -1809 -481 -1793 -447
rect -1759 -481 -1743 -447
rect -1617 -481 -1601 -447
rect -1567 -481 -1551 -447
rect -1425 -481 -1409 -447
rect -1375 -481 -1359 -447
rect -1233 -481 -1217 -447
rect -1183 -481 -1167 -447
rect -1041 -481 -1025 -447
rect -991 -481 -975 -447
rect -849 -481 -833 -447
rect -799 -481 -783 -447
rect -657 -481 -641 -447
rect -607 -481 -591 -447
rect -465 -481 -449 -447
rect -415 -481 -399 -447
rect -273 -481 -257 -447
rect -223 -481 -207 -447
rect -81 -481 -65 -447
rect -31 -481 -15 -447
rect 111 -481 127 -447
rect 161 -481 177 -447
rect 303 -481 319 -447
rect 353 -481 369 -447
rect 495 -481 511 -447
rect 545 -481 561 -447
rect 687 -481 703 -447
rect 737 -481 753 -447
rect 879 -481 895 -447
rect 929 -481 945 -447
rect 1071 -481 1087 -447
rect 1121 -481 1137 -447
rect 1263 -481 1279 -447
rect 1313 -481 1329 -447
rect 1455 -481 1471 -447
rect 1505 -481 1521 -447
rect 1647 -481 1663 -447
rect 1697 -481 1713 -447
rect 1839 -481 1855 -447
rect 1889 -481 1905 -447
rect 2031 -481 2047 -447
rect 2081 -481 2097 -447
rect 2223 -481 2239 -447
rect 2273 -481 2289 -447
rect -2531 -549 -2497 -487
rect 2497 -549 2531 -487
rect -2531 -583 -2435 -549
rect 2435 -583 2531 -549
<< viali >>
rect -2369 447 -2335 481
rect -2177 447 -2143 481
rect -1985 447 -1951 481
rect -1793 447 -1759 481
rect -1601 447 -1567 481
rect -1409 447 -1375 481
rect -1217 447 -1183 481
rect -1025 447 -991 481
rect -833 447 -799 481
rect -641 447 -607 481
rect -449 447 -415 481
rect -257 447 -223 481
rect -65 447 -31 481
rect 127 447 161 481
rect 319 447 353 481
rect 511 447 545 481
rect 703 447 737 481
rect 895 447 929 481
rect 1087 447 1121 481
rect 1279 447 1313 481
rect 1471 447 1505 481
rect 1663 447 1697 481
rect 1855 447 1889 481
rect 2047 447 2081 481
rect 2239 447 2273 481
rect -2417 121 -2383 397
rect -2321 121 -2287 397
rect -2225 121 -2191 397
rect -2129 121 -2095 397
rect -2033 121 -1999 397
rect -1937 121 -1903 397
rect -1841 121 -1807 397
rect -1745 121 -1711 397
rect -1649 121 -1615 397
rect -1553 121 -1519 397
rect -1457 121 -1423 397
rect -1361 121 -1327 397
rect -1265 121 -1231 397
rect -1169 121 -1135 397
rect -1073 121 -1039 397
rect -977 121 -943 397
rect -881 121 -847 397
rect -785 121 -751 397
rect -689 121 -655 397
rect -593 121 -559 397
rect -497 121 -463 397
rect -401 121 -367 397
rect -305 121 -271 397
rect -209 121 -175 397
rect -113 121 -79 397
rect -17 121 17 397
rect 79 121 113 397
rect 175 121 209 397
rect 271 121 305 397
rect 367 121 401 397
rect 463 121 497 397
rect 559 121 593 397
rect 655 121 689 397
rect 751 121 785 397
rect 847 121 881 397
rect 943 121 977 397
rect 1039 121 1073 397
rect 1135 121 1169 397
rect 1231 121 1265 397
rect 1327 121 1361 397
rect 1423 121 1457 397
rect 1519 121 1553 397
rect 1615 121 1649 397
rect 1711 121 1745 397
rect 1807 121 1841 397
rect 1903 121 1937 397
rect 1999 121 2033 397
rect 2095 121 2129 397
rect 2191 121 2225 397
rect 2287 121 2321 397
rect 2383 121 2417 397
rect -2273 37 -2239 71
rect -2081 37 -2047 71
rect -1889 37 -1855 71
rect -1697 37 -1663 71
rect -1505 37 -1471 71
rect -1313 37 -1279 71
rect -1121 37 -1087 71
rect -929 37 -895 71
rect -737 37 -703 71
rect -545 37 -511 71
rect -353 37 -319 71
rect -161 37 -127 71
rect 31 37 65 71
rect 223 37 257 71
rect 415 37 449 71
rect 607 37 641 71
rect 799 37 833 71
rect 991 37 1025 71
rect 1183 37 1217 71
rect 1375 37 1409 71
rect 1567 37 1601 71
rect 1759 37 1793 71
rect 1951 37 1985 71
rect 2143 37 2177 71
rect 2335 37 2369 71
rect -2273 -71 -2239 -37
rect -2081 -71 -2047 -37
rect -1889 -71 -1855 -37
rect -1697 -71 -1663 -37
rect -1505 -71 -1471 -37
rect -1313 -71 -1279 -37
rect -1121 -71 -1087 -37
rect -929 -71 -895 -37
rect -737 -71 -703 -37
rect -545 -71 -511 -37
rect -353 -71 -319 -37
rect -161 -71 -127 -37
rect 31 -71 65 -37
rect 223 -71 257 -37
rect 415 -71 449 -37
rect 607 -71 641 -37
rect 799 -71 833 -37
rect 991 -71 1025 -37
rect 1183 -71 1217 -37
rect 1375 -71 1409 -37
rect 1567 -71 1601 -37
rect 1759 -71 1793 -37
rect 1951 -71 1985 -37
rect 2143 -71 2177 -37
rect 2335 -71 2369 -37
rect -2417 -397 -2383 -121
rect -2321 -397 -2287 -121
rect -2225 -397 -2191 -121
rect -2129 -397 -2095 -121
rect -2033 -397 -1999 -121
rect -1937 -397 -1903 -121
rect -1841 -397 -1807 -121
rect -1745 -397 -1711 -121
rect -1649 -397 -1615 -121
rect -1553 -397 -1519 -121
rect -1457 -397 -1423 -121
rect -1361 -397 -1327 -121
rect -1265 -397 -1231 -121
rect -1169 -397 -1135 -121
rect -1073 -397 -1039 -121
rect -977 -397 -943 -121
rect -881 -397 -847 -121
rect -785 -397 -751 -121
rect -689 -397 -655 -121
rect -593 -397 -559 -121
rect -497 -397 -463 -121
rect -401 -397 -367 -121
rect -305 -397 -271 -121
rect -209 -397 -175 -121
rect -113 -397 -79 -121
rect -17 -397 17 -121
rect 79 -397 113 -121
rect 175 -397 209 -121
rect 271 -397 305 -121
rect 367 -397 401 -121
rect 463 -397 497 -121
rect 559 -397 593 -121
rect 655 -397 689 -121
rect 751 -397 785 -121
rect 847 -397 881 -121
rect 943 -397 977 -121
rect 1039 -397 1073 -121
rect 1135 -397 1169 -121
rect 1231 -397 1265 -121
rect 1327 -397 1361 -121
rect 1423 -397 1457 -121
rect 1519 -397 1553 -121
rect 1615 -397 1649 -121
rect 1711 -397 1745 -121
rect 1807 -397 1841 -121
rect 1903 -397 1937 -121
rect 1999 -397 2033 -121
rect 2095 -397 2129 -121
rect 2191 -397 2225 -121
rect 2287 -397 2321 -121
rect 2383 -397 2417 -121
rect -2369 -481 -2335 -447
rect -2177 -481 -2143 -447
rect -1985 -481 -1951 -447
rect -1793 -481 -1759 -447
rect -1601 -481 -1567 -447
rect -1409 -481 -1375 -447
rect -1217 -481 -1183 -447
rect -1025 -481 -991 -447
rect -833 -481 -799 -447
rect -641 -481 -607 -447
rect -449 -481 -415 -447
rect -257 -481 -223 -447
rect -65 -481 -31 -447
rect 127 -481 161 -447
rect 319 -481 353 -447
rect 511 -481 545 -447
rect 703 -481 737 -447
rect 895 -481 929 -447
rect 1087 -481 1121 -447
rect 1279 -481 1313 -447
rect 1471 -481 1505 -447
rect 1663 -481 1697 -447
rect 1855 -481 1889 -447
rect 2047 -481 2081 -447
rect 2239 -481 2273 -447
<< metal1 >>
rect -2381 481 -2323 487
rect -2381 447 -2369 481
rect -2335 447 -2323 481
rect -2381 441 -2323 447
rect -2189 481 -2131 487
rect -2189 447 -2177 481
rect -2143 447 -2131 481
rect -2189 441 -2131 447
rect -1997 481 -1939 487
rect -1997 447 -1985 481
rect -1951 447 -1939 481
rect -1997 441 -1939 447
rect -1805 481 -1747 487
rect -1805 447 -1793 481
rect -1759 447 -1747 481
rect -1805 441 -1747 447
rect -1613 481 -1555 487
rect -1613 447 -1601 481
rect -1567 447 -1555 481
rect -1613 441 -1555 447
rect -1421 481 -1363 487
rect -1421 447 -1409 481
rect -1375 447 -1363 481
rect -1421 441 -1363 447
rect -1229 481 -1171 487
rect -1229 447 -1217 481
rect -1183 447 -1171 481
rect -1229 441 -1171 447
rect -1037 481 -979 487
rect -1037 447 -1025 481
rect -991 447 -979 481
rect -1037 441 -979 447
rect -845 481 -787 487
rect -845 447 -833 481
rect -799 447 -787 481
rect -845 441 -787 447
rect -653 481 -595 487
rect -653 447 -641 481
rect -607 447 -595 481
rect -653 441 -595 447
rect -461 481 -403 487
rect -461 447 -449 481
rect -415 447 -403 481
rect -461 441 -403 447
rect -269 481 -211 487
rect -269 447 -257 481
rect -223 447 -211 481
rect -269 441 -211 447
rect -77 481 -19 487
rect -77 447 -65 481
rect -31 447 -19 481
rect -77 441 -19 447
rect 115 481 173 487
rect 115 447 127 481
rect 161 447 173 481
rect 115 441 173 447
rect 307 481 365 487
rect 307 447 319 481
rect 353 447 365 481
rect 307 441 365 447
rect 499 481 557 487
rect 499 447 511 481
rect 545 447 557 481
rect 499 441 557 447
rect 691 481 749 487
rect 691 447 703 481
rect 737 447 749 481
rect 691 441 749 447
rect 883 481 941 487
rect 883 447 895 481
rect 929 447 941 481
rect 883 441 941 447
rect 1075 481 1133 487
rect 1075 447 1087 481
rect 1121 447 1133 481
rect 1075 441 1133 447
rect 1267 481 1325 487
rect 1267 447 1279 481
rect 1313 447 1325 481
rect 1267 441 1325 447
rect 1459 481 1517 487
rect 1459 447 1471 481
rect 1505 447 1517 481
rect 1459 441 1517 447
rect 1651 481 1709 487
rect 1651 447 1663 481
rect 1697 447 1709 481
rect 1651 441 1709 447
rect 1843 481 1901 487
rect 1843 447 1855 481
rect 1889 447 1901 481
rect 1843 441 1901 447
rect 2035 481 2093 487
rect 2035 447 2047 481
rect 2081 447 2093 481
rect 2035 441 2093 447
rect 2227 481 2285 487
rect 2227 447 2239 481
rect 2273 447 2285 481
rect 2227 441 2285 447
rect -2423 397 -2377 409
rect -2423 121 -2417 397
rect -2383 121 -2377 397
rect -2423 109 -2377 121
rect -2327 397 -2281 409
rect -2327 121 -2321 397
rect -2287 121 -2281 397
rect -2327 109 -2281 121
rect -2231 397 -2185 409
rect -2231 121 -2225 397
rect -2191 121 -2185 397
rect -2231 109 -2185 121
rect -2135 397 -2089 409
rect -2135 121 -2129 397
rect -2095 121 -2089 397
rect -2135 109 -2089 121
rect -2039 397 -1993 409
rect -2039 121 -2033 397
rect -1999 121 -1993 397
rect -2039 109 -1993 121
rect -1943 397 -1897 409
rect -1943 121 -1937 397
rect -1903 121 -1897 397
rect -1943 109 -1897 121
rect -1847 397 -1801 409
rect -1847 121 -1841 397
rect -1807 121 -1801 397
rect -1847 109 -1801 121
rect -1751 397 -1705 409
rect -1751 121 -1745 397
rect -1711 121 -1705 397
rect -1751 109 -1705 121
rect -1655 397 -1609 409
rect -1655 121 -1649 397
rect -1615 121 -1609 397
rect -1655 109 -1609 121
rect -1559 397 -1513 409
rect -1559 121 -1553 397
rect -1519 121 -1513 397
rect -1559 109 -1513 121
rect -1463 397 -1417 409
rect -1463 121 -1457 397
rect -1423 121 -1417 397
rect -1463 109 -1417 121
rect -1367 397 -1321 409
rect -1367 121 -1361 397
rect -1327 121 -1321 397
rect -1367 109 -1321 121
rect -1271 397 -1225 409
rect -1271 121 -1265 397
rect -1231 121 -1225 397
rect -1271 109 -1225 121
rect -1175 397 -1129 409
rect -1175 121 -1169 397
rect -1135 121 -1129 397
rect -1175 109 -1129 121
rect -1079 397 -1033 409
rect -1079 121 -1073 397
rect -1039 121 -1033 397
rect -1079 109 -1033 121
rect -983 397 -937 409
rect -983 121 -977 397
rect -943 121 -937 397
rect -983 109 -937 121
rect -887 397 -841 409
rect -887 121 -881 397
rect -847 121 -841 397
rect -887 109 -841 121
rect -791 397 -745 409
rect -791 121 -785 397
rect -751 121 -745 397
rect -791 109 -745 121
rect -695 397 -649 409
rect -695 121 -689 397
rect -655 121 -649 397
rect -695 109 -649 121
rect -599 397 -553 409
rect -599 121 -593 397
rect -559 121 -553 397
rect -599 109 -553 121
rect -503 397 -457 409
rect -503 121 -497 397
rect -463 121 -457 397
rect -503 109 -457 121
rect -407 397 -361 409
rect -407 121 -401 397
rect -367 121 -361 397
rect -407 109 -361 121
rect -311 397 -265 409
rect -311 121 -305 397
rect -271 121 -265 397
rect -311 109 -265 121
rect -215 397 -169 409
rect -215 121 -209 397
rect -175 121 -169 397
rect -215 109 -169 121
rect -119 397 -73 409
rect -119 121 -113 397
rect -79 121 -73 397
rect -119 109 -73 121
rect -23 397 23 409
rect -23 121 -17 397
rect 17 121 23 397
rect -23 109 23 121
rect 73 397 119 409
rect 73 121 79 397
rect 113 121 119 397
rect 73 109 119 121
rect 169 397 215 409
rect 169 121 175 397
rect 209 121 215 397
rect 169 109 215 121
rect 265 397 311 409
rect 265 121 271 397
rect 305 121 311 397
rect 265 109 311 121
rect 361 397 407 409
rect 361 121 367 397
rect 401 121 407 397
rect 361 109 407 121
rect 457 397 503 409
rect 457 121 463 397
rect 497 121 503 397
rect 457 109 503 121
rect 553 397 599 409
rect 553 121 559 397
rect 593 121 599 397
rect 553 109 599 121
rect 649 397 695 409
rect 649 121 655 397
rect 689 121 695 397
rect 649 109 695 121
rect 745 397 791 409
rect 745 121 751 397
rect 785 121 791 397
rect 745 109 791 121
rect 841 397 887 409
rect 841 121 847 397
rect 881 121 887 397
rect 841 109 887 121
rect 937 397 983 409
rect 937 121 943 397
rect 977 121 983 397
rect 937 109 983 121
rect 1033 397 1079 409
rect 1033 121 1039 397
rect 1073 121 1079 397
rect 1033 109 1079 121
rect 1129 397 1175 409
rect 1129 121 1135 397
rect 1169 121 1175 397
rect 1129 109 1175 121
rect 1225 397 1271 409
rect 1225 121 1231 397
rect 1265 121 1271 397
rect 1225 109 1271 121
rect 1321 397 1367 409
rect 1321 121 1327 397
rect 1361 121 1367 397
rect 1321 109 1367 121
rect 1417 397 1463 409
rect 1417 121 1423 397
rect 1457 121 1463 397
rect 1417 109 1463 121
rect 1513 397 1559 409
rect 1513 121 1519 397
rect 1553 121 1559 397
rect 1513 109 1559 121
rect 1609 397 1655 409
rect 1609 121 1615 397
rect 1649 121 1655 397
rect 1609 109 1655 121
rect 1705 397 1751 409
rect 1705 121 1711 397
rect 1745 121 1751 397
rect 1705 109 1751 121
rect 1801 397 1847 409
rect 1801 121 1807 397
rect 1841 121 1847 397
rect 1801 109 1847 121
rect 1897 397 1943 409
rect 1897 121 1903 397
rect 1937 121 1943 397
rect 1897 109 1943 121
rect 1993 397 2039 409
rect 1993 121 1999 397
rect 2033 121 2039 397
rect 1993 109 2039 121
rect 2089 397 2135 409
rect 2089 121 2095 397
rect 2129 121 2135 397
rect 2089 109 2135 121
rect 2185 397 2231 409
rect 2185 121 2191 397
rect 2225 121 2231 397
rect 2185 109 2231 121
rect 2281 397 2327 409
rect 2281 121 2287 397
rect 2321 121 2327 397
rect 2281 109 2327 121
rect 2377 397 2423 409
rect 2377 121 2383 397
rect 2417 121 2423 397
rect 2377 109 2423 121
rect -2285 71 -2227 77
rect -2285 37 -2273 71
rect -2239 37 -2227 71
rect -2285 31 -2227 37
rect -2093 71 -2035 77
rect -2093 37 -2081 71
rect -2047 37 -2035 71
rect -2093 31 -2035 37
rect -1901 71 -1843 77
rect -1901 37 -1889 71
rect -1855 37 -1843 71
rect -1901 31 -1843 37
rect -1709 71 -1651 77
rect -1709 37 -1697 71
rect -1663 37 -1651 71
rect -1709 31 -1651 37
rect -1517 71 -1459 77
rect -1517 37 -1505 71
rect -1471 37 -1459 71
rect -1517 31 -1459 37
rect -1325 71 -1267 77
rect -1325 37 -1313 71
rect -1279 37 -1267 71
rect -1325 31 -1267 37
rect -1133 71 -1075 77
rect -1133 37 -1121 71
rect -1087 37 -1075 71
rect -1133 31 -1075 37
rect -941 71 -883 77
rect -941 37 -929 71
rect -895 37 -883 71
rect -941 31 -883 37
rect -749 71 -691 77
rect -749 37 -737 71
rect -703 37 -691 71
rect -749 31 -691 37
rect -557 71 -499 77
rect -557 37 -545 71
rect -511 37 -499 71
rect -557 31 -499 37
rect -365 71 -307 77
rect -365 37 -353 71
rect -319 37 -307 71
rect -365 31 -307 37
rect -173 71 -115 77
rect -173 37 -161 71
rect -127 37 -115 71
rect -173 31 -115 37
rect 19 71 77 77
rect 19 37 31 71
rect 65 37 77 71
rect 19 31 77 37
rect 211 71 269 77
rect 211 37 223 71
rect 257 37 269 71
rect 211 31 269 37
rect 403 71 461 77
rect 403 37 415 71
rect 449 37 461 71
rect 403 31 461 37
rect 595 71 653 77
rect 595 37 607 71
rect 641 37 653 71
rect 595 31 653 37
rect 787 71 845 77
rect 787 37 799 71
rect 833 37 845 71
rect 787 31 845 37
rect 979 71 1037 77
rect 979 37 991 71
rect 1025 37 1037 71
rect 979 31 1037 37
rect 1171 71 1229 77
rect 1171 37 1183 71
rect 1217 37 1229 71
rect 1171 31 1229 37
rect 1363 71 1421 77
rect 1363 37 1375 71
rect 1409 37 1421 71
rect 1363 31 1421 37
rect 1555 71 1613 77
rect 1555 37 1567 71
rect 1601 37 1613 71
rect 1555 31 1613 37
rect 1747 71 1805 77
rect 1747 37 1759 71
rect 1793 37 1805 71
rect 1747 31 1805 37
rect 1939 71 1997 77
rect 1939 37 1951 71
rect 1985 37 1997 71
rect 1939 31 1997 37
rect 2131 71 2189 77
rect 2131 37 2143 71
rect 2177 37 2189 71
rect 2131 31 2189 37
rect 2323 71 2381 77
rect 2323 37 2335 71
rect 2369 37 2381 71
rect 2323 31 2381 37
rect -2285 -37 -2227 -31
rect -2285 -71 -2273 -37
rect -2239 -71 -2227 -37
rect -2285 -77 -2227 -71
rect -2093 -37 -2035 -31
rect -2093 -71 -2081 -37
rect -2047 -71 -2035 -37
rect -2093 -77 -2035 -71
rect -1901 -37 -1843 -31
rect -1901 -71 -1889 -37
rect -1855 -71 -1843 -37
rect -1901 -77 -1843 -71
rect -1709 -37 -1651 -31
rect -1709 -71 -1697 -37
rect -1663 -71 -1651 -37
rect -1709 -77 -1651 -71
rect -1517 -37 -1459 -31
rect -1517 -71 -1505 -37
rect -1471 -71 -1459 -37
rect -1517 -77 -1459 -71
rect -1325 -37 -1267 -31
rect -1325 -71 -1313 -37
rect -1279 -71 -1267 -37
rect -1325 -77 -1267 -71
rect -1133 -37 -1075 -31
rect -1133 -71 -1121 -37
rect -1087 -71 -1075 -37
rect -1133 -77 -1075 -71
rect -941 -37 -883 -31
rect -941 -71 -929 -37
rect -895 -71 -883 -37
rect -941 -77 -883 -71
rect -749 -37 -691 -31
rect -749 -71 -737 -37
rect -703 -71 -691 -37
rect -749 -77 -691 -71
rect -557 -37 -499 -31
rect -557 -71 -545 -37
rect -511 -71 -499 -37
rect -557 -77 -499 -71
rect -365 -37 -307 -31
rect -365 -71 -353 -37
rect -319 -71 -307 -37
rect -365 -77 -307 -71
rect -173 -37 -115 -31
rect -173 -71 -161 -37
rect -127 -71 -115 -37
rect -173 -77 -115 -71
rect 19 -37 77 -31
rect 19 -71 31 -37
rect 65 -71 77 -37
rect 19 -77 77 -71
rect 211 -37 269 -31
rect 211 -71 223 -37
rect 257 -71 269 -37
rect 211 -77 269 -71
rect 403 -37 461 -31
rect 403 -71 415 -37
rect 449 -71 461 -37
rect 403 -77 461 -71
rect 595 -37 653 -31
rect 595 -71 607 -37
rect 641 -71 653 -37
rect 595 -77 653 -71
rect 787 -37 845 -31
rect 787 -71 799 -37
rect 833 -71 845 -37
rect 787 -77 845 -71
rect 979 -37 1037 -31
rect 979 -71 991 -37
rect 1025 -71 1037 -37
rect 979 -77 1037 -71
rect 1171 -37 1229 -31
rect 1171 -71 1183 -37
rect 1217 -71 1229 -37
rect 1171 -77 1229 -71
rect 1363 -37 1421 -31
rect 1363 -71 1375 -37
rect 1409 -71 1421 -37
rect 1363 -77 1421 -71
rect 1555 -37 1613 -31
rect 1555 -71 1567 -37
rect 1601 -71 1613 -37
rect 1555 -77 1613 -71
rect 1747 -37 1805 -31
rect 1747 -71 1759 -37
rect 1793 -71 1805 -37
rect 1747 -77 1805 -71
rect 1939 -37 1997 -31
rect 1939 -71 1951 -37
rect 1985 -71 1997 -37
rect 1939 -77 1997 -71
rect 2131 -37 2189 -31
rect 2131 -71 2143 -37
rect 2177 -71 2189 -37
rect 2131 -77 2189 -71
rect 2323 -37 2381 -31
rect 2323 -71 2335 -37
rect 2369 -71 2381 -37
rect 2323 -77 2381 -71
rect -2423 -121 -2377 -109
rect -2423 -397 -2417 -121
rect -2383 -397 -2377 -121
rect -2423 -409 -2377 -397
rect -2327 -121 -2281 -109
rect -2327 -397 -2321 -121
rect -2287 -397 -2281 -121
rect -2327 -409 -2281 -397
rect -2231 -121 -2185 -109
rect -2231 -397 -2225 -121
rect -2191 -397 -2185 -121
rect -2231 -409 -2185 -397
rect -2135 -121 -2089 -109
rect -2135 -397 -2129 -121
rect -2095 -397 -2089 -121
rect -2135 -409 -2089 -397
rect -2039 -121 -1993 -109
rect -2039 -397 -2033 -121
rect -1999 -397 -1993 -121
rect -2039 -409 -1993 -397
rect -1943 -121 -1897 -109
rect -1943 -397 -1937 -121
rect -1903 -397 -1897 -121
rect -1943 -409 -1897 -397
rect -1847 -121 -1801 -109
rect -1847 -397 -1841 -121
rect -1807 -397 -1801 -121
rect -1847 -409 -1801 -397
rect -1751 -121 -1705 -109
rect -1751 -397 -1745 -121
rect -1711 -397 -1705 -121
rect -1751 -409 -1705 -397
rect -1655 -121 -1609 -109
rect -1655 -397 -1649 -121
rect -1615 -397 -1609 -121
rect -1655 -409 -1609 -397
rect -1559 -121 -1513 -109
rect -1559 -397 -1553 -121
rect -1519 -397 -1513 -121
rect -1559 -409 -1513 -397
rect -1463 -121 -1417 -109
rect -1463 -397 -1457 -121
rect -1423 -397 -1417 -121
rect -1463 -409 -1417 -397
rect -1367 -121 -1321 -109
rect -1367 -397 -1361 -121
rect -1327 -397 -1321 -121
rect -1367 -409 -1321 -397
rect -1271 -121 -1225 -109
rect -1271 -397 -1265 -121
rect -1231 -397 -1225 -121
rect -1271 -409 -1225 -397
rect -1175 -121 -1129 -109
rect -1175 -397 -1169 -121
rect -1135 -397 -1129 -121
rect -1175 -409 -1129 -397
rect -1079 -121 -1033 -109
rect -1079 -397 -1073 -121
rect -1039 -397 -1033 -121
rect -1079 -409 -1033 -397
rect -983 -121 -937 -109
rect -983 -397 -977 -121
rect -943 -397 -937 -121
rect -983 -409 -937 -397
rect -887 -121 -841 -109
rect -887 -397 -881 -121
rect -847 -397 -841 -121
rect -887 -409 -841 -397
rect -791 -121 -745 -109
rect -791 -397 -785 -121
rect -751 -397 -745 -121
rect -791 -409 -745 -397
rect -695 -121 -649 -109
rect -695 -397 -689 -121
rect -655 -397 -649 -121
rect -695 -409 -649 -397
rect -599 -121 -553 -109
rect -599 -397 -593 -121
rect -559 -397 -553 -121
rect -599 -409 -553 -397
rect -503 -121 -457 -109
rect -503 -397 -497 -121
rect -463 -397 -457 -121
rect -503 -409 -457 -397
rect -407 -121 -361 -109
rect -407 -397 -401 -121
rect -367 -397 -361 -121
rect -407 -409 -361 -397
rect -311 -121 -265 -109
rect -311 -397 -305 -121
rect -271 -397 -265 -121
rect -311 -409 -265 -397
rect -215 -121 -169 -109
rect -215 -397 -209 -121
rect -175 -397 -169 -121
rect -215 -409 -169 -397
rect -119 -121 -73 -109
rect -119 -397 -113 -121
rect -79 -397 -73 -121
rect -119 -409 -73 -397
rect -23 -121 23 -109
rect -23 -397 -17 -121
rect 17 -397 23 -121
rect -23 -409 23 -397
rect 73 -121 119 -109
rect 73 -397 79 -121
rect 113 -397 119 -121
rect 73 -409 119 -397
rect 169 -121 215 -109
rect 169 -397 175 -121
rect 209 -397 215 -121
rect 169 -409 215 -397
rect 265 -121 311 -109
rect 265 -397 271 -121
rect 305 -397 311 -121
rect 265 -409 311 -397
rect 361 -121 407 -109
rect 361 -397 367 -121
rect 401 -397 407 -121
rect 361 -409 407 -397
rect 457 -121 503 -109
rect 457 -397 463 -121
rect 497 -397 503 -121
rect 457 -409 503 -397
rect 553 -121 599 -109
rect 553 -397 559 -121
rect 593 -397 599 -121
rect 553 -409 599 -397
rect 649 -121 695 -109
rect 649 -397 655 -121
rect 689 -397 695 -121
rect 649 -409 695 -397
rect 745 -121 791 -109
rect 745 -397 751 -121
rect 785 -397 791 -121
rect 745 -409 791 -397
rect 841 -121 887 -109
rect 841 -397 847 -121
rect 881 -397 887 -121
rect 841 -409 887 -397
rect 937 -121 983 -109
rect 937 -397 943 -121
rect 977 -397 983 -121
rect 937 -409 983 -397
rect 1033 -121 1079 -109
rect 1033 -397 1039 -121
rect 1073 -397 1079 -121
rect 1033 -409 1079 -397
rect 1129 -121 1175 -109
rect 1129 -397 1135 -121
rect 1169 -397 1175 -121
rect 1129 -409 1175 -397
rect 1225 -121 1271 -109
rect 1225 -397 1231 -121
rect 1265 -397 1271 -121
rect 1225 -409 1271 -397
rect 1321 -121 1367 -109
rect 1321 -397 1327 -121
rect 1361 -397 1367 -121
rect 1321 -409 1367 -397
rect 1417 -121 1463 -109
rect 1417 -397 1423 -121
rect 1457 -397 1463 -121
rect 1417 -409 1463 -397
rect 1513 -121 1559 -109
rect 1513 -397 1519 -121
rect 1553 -397 1559 -121
rect 1513 -409 1559 -397
rect 1609 -121 1655 -109
rect 1609 -397 1615 -121
rect 1649 -397 1655 -121
rect 1609 -409 1655 -397
rect 1705 -121 1751 -109
rect 1705 -397 1711 -121
rect 1745 -397 1751 -121
rect 1705 -409 1751 -397
rect 1801 -121 1847 -109
rect 1801 -397 1807 -121
rect 1841 -397 1847 -121
rect 1801 -409 1847 -397
rect 1897 -121 1943 -109
rect 1897 -397 1903 -121
rect 1937 -397 1943 -121
rect 1897 -409 1943 -397
rect 1993 -121 2039 -109
rect 1993 -397 1999 -121
rect 2033 -397 2039 -121
rect 1993 -409 2039 -397
rect 2089 -121 2135 -109
rect 2089 -397 2095 -121
rect 2129 -397 2135 -121
rect 2089 -409 2135 -397
rect 2185 -121 2231 -109
rect 2185 -397 2191 -121
rect 2225 -397 2231 -121
rect 2185 -409 2231 -397
rect 2281 -121 2327 -109
rect 2281 -397 2287 -121
rect 2321 -397 2327 -121
rect 2281 -409 2327 -397
rect 2377 -121 2423 -109
rect 2377 -397 2383 -121
rect 2417 -397 2423 -121
rect 2377 -409 2423 -397
rect -2381 -447 -2323 -441
rect -2381 -481 -2369 -447
rect -2335 -481 -2323 -447
rect -2381 -487 -2323 -481
rect -2189 -447 -2131 -441
rect -2189 -481 -2177 -447
rect -2143 -481 -2131 -447
rect -2189 -487 -2131 -481
rect -1997 -447 -1939 -441
rect -1997 -481 -1985 -447
rect -1951 -481 -1939 -447
rect -1997 -487 -1939 -481
rect -1805 -447 -1747 -441
rect -1805 -481 -1793 -447
rect -1759 -481 -1747 -447
rect -1805 -487 -1747 -481
rect -1613 -447 -1555 -441
rect -1613 -481 -1601 -447
rect -1567 -481 -1555 -447
rect -1613 -487 -1555 -481
rect -1421 -447 -1363 -441
rect -1421 -481 -1409 -447
rect -1375 -481 -1363 -447
rect -1421 -487 -1363 -481
rect -1229 -447 -1171 -441
rect -1229 -481 -1217 -447
rect -1183 -481 -1171 -447
rect -1229 -487 -1171 -481
rect -1037 -447 -979 -441
rect -1037 -481 -1025 -447
rect -991 -481 -979 -447
rect -1037 -487 -979 -481
rect -845 -447 -787 -441
rect -845 -481 -833 -447
rect -799 -481 -787 -447
rect -845 -487 -787 -481
rect -653 -447 -595 -441
rect -653 -481 -641 -447
rect -607 -481 -595 -447
rect -653 -487 -595 -481
rect -461 -447 -403 -441
rect -461 -481 -449 -447
rect -415 -481 -403 -447
rect -461 -487 -403 -481
rect -269 -447 -211 -441
rect -269 -481 -257 -447
rect -223 -481 -211 -447
rect -269 -487 -211 -481
rect -77 -447 -19 -441
rect -77 -481 -65 -447
rect -31 -481 -19 -447
rect -77 -487 -19 -481
rect 115 -447 173 -441
rect 115 -481 127 -447
rect 161 -481 173 -447
rect 115 -487 173 -481
rect 307 -447 365 -441
rect 307 -481 319 -447
rect 353 -481 365 -447
rect 307 -487 365 -481
rect 499 -447 557 -441
rect 499 -481 511 -447
rect 545 -481 557 -447
rect 499 -487 557 -481
rect 691 -447 749 -441
rect 691 -481 703 -447
rect 737 -481 749 -447
rect 691 -487 749 -481
rect 883 -447 941 -441
rect 883 -481 895 -447
rect 929 -481 941 -447
rect 883 -487 941 -481
rect 1075 -447 1133 -441
rect 1075 -481 1087 -447
rect 1121 -481 1133 -447
rect 1075 -487 1133 -481
rect 1267 -447 1325 -441
rect 1267 -481 1279 -447
rect 1313 -481 1325 -447
rect 1267 -487 1325 -481
rect 1459 -447 1517 -441
rect 1459 -481 1471 -447
rect 1505 -481 1517 -447
rect 1459 -487 1517 -481
rect 1651 -447 1709 -441
rect 1651 -481 1663 -447
rect 1697 -481 1709 -447
rect 1651 -487 1709 -481
rect 1843 -447 1901 -441
rect 1843 -481 1855 -447
rect 1889 -481 1901 -447
rect 1843 -487 1901 -481
rect 2035 -447 2093 -441
rect 2035 -481 2047 -447
rect 2081 -481 2093 -447
rect 2035 -487 2093 -481
rect 2227 -447 2285 -441
rect 2227 -481 2239 -447
rect 2273 -481 2285 -447
rect 2227 -487 2285 -481
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2514 -566 2514 566
string parameters w 1.5 l 0.150 m 2 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
