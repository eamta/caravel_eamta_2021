magic
tech sky130A
magscale 1 2
timestamp 1615923543
<< error_p >>
rect -5870 -307 -5812 -301
rect -5752 -307 -5694 -301
rect -5634 -307 -5576 -301
rect -5516 -307 -5458 -301
rect -5398 -307 -5340 -301
rect -5280 -307 -5222 -301
rect -5162 -307 -5104 -301
rect -5044 -307 -4986 -301
rect -4926 -307 -4868 -301
rect -4808 -307 -4750 -301
rect -4690 -307 -4632 -301
rect -4572 -307 -4514 -301
rect -4454 -307 -4396 -301
rect -4336 -307 -4278 -301
rect -4218 -307 -4160 -301
rect -4100 -307 -4042 -301
rect -3982 -307 -3924 -301
rect -3864 -307 -3806 -301
rect -3746 -307 -3688 -301
rect -3628 -307 -3570 -301
rect -3510 -307 -3452 -301
rect -3392 -307 -3334 -301
rect -3274 -307 -3216 -301
rect -3156 -307 -3098 -301
rect -3038 -307 -2980 -301
rect -2920 -307 -2862 -301
rect -2802 -307 -2744 -301
rect -2684 -307 -2626 -301
rect -2566 -307 -2508 -301
rect -2448 -307 -2390 -301
rect -2330 -307 -2272 -301
rect -2212 -307 -2154 -301
rect -2094 -307 -2036 -301
rect -1976 -307 -1918 -301
rect -1858 -307 -1800 -301
rect -1740 -307 -1682 -301
rect -1622 -307 -1564 -301
rect -1504 -307 -1446 -301
rect -1386 -307 -1328 -301
rect -1268 -307 -1210 -301
rect -1150 -307 -1092 -301
rect -1032 -307 -974 -301
rect -914 -307 -856 -301
rect -796 -307 -738 -301
rect -678 -307 -620 -301
rect -560 -307 -502 -301
rect -442 -307 -384 -301
rect -324 -307 -266 -301
rect -206 -307 -148 -301
rect -88 -307 -30 -301
rect 30 -307 88 -301
rect 148 -307 206 -301
rect 266 -307 324 -301
rect 384 -307 442 -301
rect 502 -307 560 -301
rect 620 -307 678 -301
rect 738 -307 796 -301
rect 856 -307 914 -301
rect 974 -307 1032 -301
rect 1092 -307 1150 -301
rect 1210 -307 1268 -301
rect 1328 -307 1386 -301
rect 1446 -307 1504 -301
rect 1564 -307 1622 -301
rect 1682 -307 1740 -301
rect 1800 -307 1858 -301
rect 1918 -307 1976 -301
rect 2036 -307 2094 -301
rect 2154 -307 2212 -301
rect 2272 -307 2330 -301
rect 2390 -307 2448 -301
rect 2508 -307 2566 -301
rect 2626 -307 2684 -301
rect 2744 -307 2802 -301
rect 2862 -307 2920 -301
rect 2980 -307 3038 -301
rect 3098 -307 3156 -301
rect 3216 -307 3274 -301
rect 3334 -307 3392 -301
rect 3452 -307 3510 -301
rect 3570 -307 3628 -301
rect 3688 -307 3746 -301
rect 3806 -307 3864 -301
rect 3924 -307 3982 -301
rect 4042 -307 4100 -301
rect 4160 -307 4218 -301
rect 4278 -307 4336 -301
rect 4396 -307 4454 -301
rect 4514 -307 4572 -301
rect 4632 -307 4690 -301
rect 4750 -307 4808 -301
rect 4868 -307 4926 -301
rect 4986 -307 5044 -301
rect 5104 -307 5162 -301
rect 5222 -307 5280 -301
rect 5340 -307 5398 -301
rect 5458 -307 5516 -301
rect 5576 -307 5634 -301
rect 5694 -307 5752 -301
rect 5812 -307 5870 -301
rect -5870 -341 -5858 -307
rect -5752 -341 -5740 -307
rect -5634 -341 -5622 -307
rect -5516 -341 -5504 -307
rect -5398 -341 -5386 -307
rect -5280 -341 -5268 -307
rect -5162 -341 -5150 -307
rect -5044 -341 -5032 -307
rect -4926 -341 -4914 -307
rect -4808 -341 -4796 -307
rect -4690 -341 -4678 -307
rect -4572 -341 -4560 -307
rect -4454 -341 -4442 -307
rect -4336 -341 -4324 -307
rect -4218 -341 -4206 -307
rect -4100 -341 -4088 -307
rect -3982 -341 -3970 -307
rect -3864 -341 -3852 -307
rect -3746 -341 -3734 -307
rect -3628 -341 -3616 -307
rect -3510 -341 -3498 -307
rect -3392 -341 -3380 -307
rect -3274 -341 -3262 -307
rect -3156 -341 -3144 -307
rect -3038 -341 -3026 -307
rect -2920 -341 -2908 -307
rect -2802 -341 -2790 -307
rect -2684 -341 -2672 -307
rect -2566 -341 -2554 -307
rect -2448 -341 -2436 -307
rect -2330 -341 -2318 -307
rect -2212 -341 -2200 -307
rect -2094 -341 -2082 -307
rect -1976 -341 -1964 -307
rect -1858 -341 -1846 -307
rect -1740 -341 -1728 -307
rect -1622 -341 -1610 -307
rect -1504 -341 -1492 -307
rect -1386 -341 -1374 -307
rect -1268 -341 -1256 -307
rect -1150 -341 -1138 -307
rect -1032 -341 -1020 -307
rect -914 -341 -902 -307
rect -796 -341 -784 -307
rect -678 -341 -666 -307
rect -560 -341 -548 -307
rect -442 -341 -430 -307
rect -324 -341 -312 -307
rect -206 -341 -194 -307
rect -88 -341 -76 -307
rect 30 -341 42 -307
rect 148 -341 160 -307
rect 266 -341 278 -307
rect 384 -341 396 -307
rect 502 -341 514 -307
rect 620 -341 632 -307
rect 738 -341 750 -307
rect 856 -341 868 -307
rect 974 -341 986 -307
rect 1092 -341 1104 -307
rect 1210 -341 1222 -307
rect 1328 -341 1340 -307
rect 1446 -341 1458 -307
rect 1564 -341 1576 -307
rect 1682 -341 1694 -307
rect 1800 -341 1812 -307
rect 1918 -341 1930 -307
rect 2036 -341 2048 -307
rect 2154 -341 2166 -307
rect 2272 -341 2284 -307
rect 2390 -341 2402 -307
rect 2508 -341 2520 -307
rect 2626 -341 2638 -307
rect 2744 -341 2756 -307
rect 2862 -341 2874 -307
rect 2980 -341 2992 -307
rect 3098 -341 3110 -307
rect 3216 -341 3228 -307
rect 3334 -341 3346 -307
rect 3452 -341 3464 -307
rect 3570 -341 3582 -307
rect 3688 -341 3700 -307
rect 3806 -341 3818 -307
rect 3924 -341 3936 -307
rect 4042 -341 4054 -307
rect 4160 -341 4172 -307
rect 4278 -341 4290 -307
rect 4396 -341 4408 -307
rect 4514 -341 4526 -307
rect 4632 -341 4644 -307
rect 4750 -341 4762 -307
rect 4868 -341 4880 -307
rect 4986 -341 4998 -307
rect 5104 -341 5116 -307
rect 5222 -341 5234 -307
rect 5340 -341 5352 -307
rect 5458 -341 5470 -307
rect 5576 -341 5588 -307
rect 5694 -341 5706 -307
rect 5812 -341 5824 -307
rect -5870 -347 -5812 -341
rect -5752 -347 -5694 -341
rect -5634 -347 -5576 -341
rect -5516 -347 -5458 -341
rect -5398 -347 -5340 -341
rect -5280 -347 -5222 -341
rect -5162 -347 -5104 -341
rect -5044 -347 -4986 -341
rect -4926 -347 -4868 -341
rect -4808 -347 -4750 -341
rect -4690 -347 -4632 -341
rect -4572 -347 -4514 -341
rect -4454 -347 -4396 -341
rect -4336 -347 -4278 -341
rect -4218 -347 -4160 -341
rect -4100 -347 -4042 -341
rect -3982 -347 -3924 -341
rect -3864 -347 -3806 -341
rect -3746 -347 -3688 -341
rect -3628 -347 -3570 -341
rect -3510 -347 -3452 -341
rect -3392 -347 -3334 -341
rect -3274 -347 -3216 -341
rect -3156 -347 -3098 -341
rect -3038 -347 -2980 -341
rect -2920 -347 -2862 -341
rect -2802 -347 -2744 -341
rect -2684 -347 -2626 -341
rect -2566 -347 -2508 -341
rect -2448 -347 -2390 -341
rect -2330 -347 -2272 -341
rect -2212 -347 -2154 -341
rect -2094 -347 -2036 -341
rect -1976 -347 -1918 -341
rect -1858 -347 -1800 -341
rect -1740 -347 -1682 -341
rect -1622 -347 -1564 -341
rect -1504 -347 -1446 -341
rect -1386 -347 -1328 -341
rect -1268 -347 -1210 -341
rect -1150 -347 -1092 -341
rect -1032 -347 -974 -341
rect -914 -347 -856 -341
rect -796 -347 -738 -341
rect -678 -347 -620 -341
rect -560 -347 -502 -341
rect -442 -347 -384 -341
rect -324 -347 -266 -341
rect -206 -347 -148 -341
rect -88 -347 -30 -341
rect 30 -347 88 -341
rect 148 -347 206 -341
rect 266 -347 324 -341
rect 384 -347 442 -341
rect 502 -347 560 -341
rect 620 -347 678 -341
rect 738 -347 796 -341
rect 856 -347 914 -341
rect 974 -347 1032 -341
rect 1092 -347 1150 -341
rect 1210 -347 1268 -341
rect 1328 -347 1386 -341
rect 1446 -347 1504 -341
rect 1564 -347 1622 -341
rect 1682 -347 1740 -341
rect 1800 -347 1858 -341
rect 1918 -347 1976 -341
rect 2036 -347 2094 -341
rect 2154 -347 2212 -341
rect 2272 -347 2330 -341
rect 2390 -347 2448 -341
rect 2508 -347 2566 -341
rect 2626 -347 2684 -341
rect 2744 -347 2802 -341
rect 2862 -347 2920 -341
rect 2980 -347 3038 -341
rect 3098 -347 3156 -341
rect 3216 -347 3274 -341
rect 3334 -347 3392 -341
rect 3452 -347 3510 -341
rect 3570 -347 3628 -341
rect 3688 -347 3746 -341
rect 3806 -347 3864 -341
rect 3924 -347 3982 -341
rect 4042 -347 4100 -341
rect 4160 -347 4218 -341
rect 4278 -347 4336 -341
rect 4396 -347 4454 -341
rect 4514 -347 4572 -341
rect 4632 -347 4690 -341
rect 4750 -347 4808 -341
rect 4868 -347 4926 -341
rect 4986 -347 5044 -341
rect 5104 -347 5162 -341
rect 5222 -347 5280 -341
rect 5340 -347 5398 -341
rect 5458 -347 5516 -341
rect 5576 -347 5634 -341
rect 5694 -347 5752 -341
rect 5812 -347 5870 -341
<< nmos >>
rect -5871 -269 -5811 331
rect -5753 -269 -5693 331
rect -5635 -269 -5575 331
rect -5517 -269 -5457 331
rect -5399 -269 -5339 331
rect -5281 -269 -5221 331
rect -5163 -269 -5103 331
rect -5045 -269 -4985 331
rect -4927 -269 -4867 331
rect -4809 -269 -4749 331
rect -4691 -269 -4631 331
rect -4573 -269 -4513 331
rect -4455 -269 -4395 331
rect -4337 -269 -4277 331
rect -4219 -269 -4159 331
rect -4101 -269 -4041 331
rect -3983 -269 -3923 331
rect -3865 -269 -3805 331
rect -3747 -269 -3687 331
rect -3629 -269 -3569 331
rect -3511 -269 -3451 331
rect -3393 -269 -3333 331
rect -3275 -269 -3215 331
rect -3157 -269 -3097 331
rect -3039 -269 -2979 331
rect -2921 -269 -2861 331
rect -2803 -269 -2743 331
rect -2685 -269 -2625 331
rect -2567 -269 -2507 331
rect -2449 -269 -2389 331
rect -2331 -269 -2271 331
rect -2213 -269 -2153 331
rect -2095 -269 -2035 331
rect -1977 -269 -1917 331
rect -1859 -269 -1799 331
rect -1741 -269 -1681 331
rect -1623 -269 -1563 331
rect -1505 -269 -1445 331
rect -1387 -269 -1327 331
rect -1269 -269 -1209 331
rect -1151 -269 -1091 331
rect -1033 -269 -973 331
rect -915 -269 -855 331
rect -797 -269 -737 331
rect -679 -269 -619 331
rect -561 -269 -501 331
rect -443 -269 -383 331
rect -325 -269 -265 331
rect -207 -269 -147 331
rect -89 -269 -29 331
rect 29 -269 89 331
rect 147 -269 207 331
rect 265 -269 325 331
rect 383 -269 443 331
rect 501 -269 561 331
rect 619 -269 679 331
rect 737 -269 797 331
rect 855 -269 915 331
rect 973 -269 1033 331
rect 1091 -269 1151 331
rect 1209 -269 1269 331
rect 1327 -269 1387 331
rect 1445 -269 1505 331
rect 1563 -269 1623 331
rect 1681 -269 1741 331
rect 1799 -269 1859 331
rect 1917 -269 1977 331
rect 2035 -269 2095 331
rect 2153 -269 2213 331
rect 2271 -269 2331 331
rect 2389 -269 2449 331
rect 2507 -269 2567 331
rect 2625 -269 2685 331
rect 2743 -269 2803 331
rect 2861 -269 2921 331
rect 2979 -269 3039 331
rect 3097 -269 3157 331
rect 3215 -269 3275 331
rect 3333 -269 3393 331
rect 3451 -269 3511 331
rect 3569 -269 3629 331
rect 3687 -269 3747 331
rect 3805 -269 3865 331
rect 3923 -269 3983 331
rect 4041 -269 4101 331
rect 4159 -269 4219 331
rect 4277 -269 4337 331
rect 4395 -269 4455 331
rect 4513 -269 4573 331
rect 4631 -269 4691 331
rect 4749 -269 4809 331
rect 4867 -269 4927 331
rect 4985 -269 5045 331
rect 5103 -269 5163 331
rect 5221 -269 5281 331
rect 5339 -269 5399 331
rect 5457 -269 5517 331
rect 5575 -269 5635 331
rect 5693 -269 5753 331
rect 5811 -269 5871 331
<< ndiff >>
rect -5929 319 -5871 331
rect -5929 -257 -5917 319
rect -5883 -257 -5871 319
rect -5929 -269 -5871 -257
rect -5811 319 -5753 331
rect -5811 -257 -5799 319
rect -5765 -257 -5753 319
rect -5811 -269 -5753 -257
rect -5693 319 -5635 331
rect -5693 -257 -5681 319
rect -5647 -257 -5635 319
rect -5693 -269 -5635 -257
rect -5575 319 -5517 331
rect -5575 -257 -5563 319
rect -5529 -257 -5517 319
rect -5575 -269 -5517 -257
rect -5457 319 -5399 331
rect -5457 -257 -5445 319
rect -5411 -257 -5399 319
rect -5457 -269 -5399 -257
rect -5339 319 -5281 331
rect -5339 -257 -5327 319
rect -5293 -257 -5281 319
rect -5339 -269 -5281 -257
rect -5221 319 -5163 331
rect -5221 -257 -5209 319
rect -5175 -257 -5163 319
rect -5221 -269 -5163 -257
rect -5103 319 -5045 331
rect -5103 -257 -5091 319
rect -5057 -257 -5045 319
rect -5103 -269 -5045 -257
rect -4985 319 -4927 331
rect -4985 -257 -4973 319
rect -4939 -257 -4927 319
rect -4985 -269 -4927 -257
rect -4867 319 -4809 331
rect -4867 -257 -4855 319
rect -4821 -257 -4809 319
rect -4867 -269 -4809 -257
rect -4749 319 -4691 331
rect -4749 -257 -4737 319
rect -4703 -257 -4691 319
rect -4749 -269 -4691 -257
rect -4631 319 -4573 331
rect -4631 -257 -4619 319
rect -4585 -257 -4573 319
rect -4631 -269 -4573 -257
rect -4513 319 -4455 331
rect -4513 -257 -4501 319
rect -4467 -257 -4455 319
rect -4513 -269 -4455 -257
rect -4395 319 -4337 331
rect -4395 -257 -4383 319
rect -4349 -257 -4337 319
rect -4395 -269 -4337 -257
rect -4277 319 -4219 331
rect -4277 -257 -4265 319
rect -4231 -257 -4219 319
rect -4277 -269 -4219 -257
rect -4159 319 -4101 331
rect -4159 -257 -4147 319
rect -4113 -257 -4101 319
rect -4159 -269 -4101 -257
rect -4041 319 -3983 331
rect -4041 -257 -4029 319
rect -3995 -257 -3983 319
rect -4041 -269 -3983 -257
rect -3923 319 -3865 331
rect -3923 -257 -3911 319
rect -3877 -257 -3865 319
rect -3923 -269 -3865 -257
rect -3805 319 -3747 331
rect -3805 -257 -3793 319
rect -3759 -257 -3747 319
rect -3805 -269 -3747 -257
rect -3687 319 -3629 331
rect -3687 -257 -3675 319
rect -3641 -257 -3629 319
rect -3687 -269 -3629 -257
rect -3569 319 -3511 331
rect -3569 -257 -3557 319
rect -3523 -257 -3511 319
rect -3569 -269 -3511 -257
rect -3451 319 -3393 331
rect -3451 -257 -3439 319
rect -3405 -257 -3393 319
rect -3451 -269 -3393 -257
rect -3333 319 -3275 331
rect -3333 -257 -3321 319
rect -3287 -257 -3275 319
rect -3333 -269 -3275 -257
rect -3215 319 -3157 331
rect -3215 -257 -3203 319
rect -3169 -257 -3157 319
rect -3215 -269 -3157 -257
rect -3097 319 -3039 331
rect -3097 -257 -3085 319
rect -3051 -257 -3039 319
rect -3097 -269 -3039 -257
rect -2979 319 -2921 331
rect -2979 -257 -2967 319
rect -2933 -257 -2921 319
rect -2979 -269 -2921 -257
rect -2861 319 -2803 331
rect -2861 -257 -2849 319
rect -2815 -257 -2803 319
rect -2861 -269 -2803 -257
rect -2743 319 -2685 331
rect -2743 -257 -2731 319
rect -2697 -257 -2685 319
rect -2743 -269 -2685 -257
rect -2625 319 -2567 331
rect -2625 -257 -2613 319
rect -2579 -257 -2567 319
rect -2625 -269 -2567 -257
rect -2507 319 -2449 331
rect -2507 -257 -2495 319
rect -2461 -257 -2449 319
rect -2507 -269 -2449 -257
rect -2389 319 -2331 331
rect -2389 -257 -2377 319
rect -2343 -257 -2331 319
rect -2389 -269 -2331 -257
rect -2271 319 -2213 331
rect -2271 -257 -2259 319
rect -2225 -257 -2213 319
rect -2271 -269 -2213 -257
rect -2153 319 -2095 331
rect -2153 -257 -2141 319
rect -2107 -257 -2095 319
rect -2153 -269 -2095 -257
rect -2035 319 -1977 331
rect -2035 -257 -2023 319
rect -1989 -257 -1977 319
rect -2035 -269 -1977 -257
rect -1917 319 -1859 331
rect -1917 -257 -1905 319
rect -1871 -257 -1859 319
rect -1917 -269 -1859 -257
rect -1799 319 -1741 331
rect -1799 -257 -1787 319
rect -1753 -257 -1741 319
rect -1799 -269 -1741 -257
rect -1681 319 -1623 331
rect -1681 -257 -1669 319
rect -1635 -257 -1623 319
rect -1681 -269 -1623 -257
rect -1563 319 -1505 331
rect -1563 -257 -1551 319
rect -1517 -257 -1505 319
rect -1563 -269 -1505 -257
rect -1445 319 -1387 331
rect -1445 -257 -1433 319
rect -1399 -257 -1387 319
rect -1445 -269 -1387 -257
rect -1327 319 -1269 331
rect -1327 -257 -1315 319
rect -1281 -257 -1269 319
rect -1327 -269 -1269 -257
rect -1209 319 -1151 331
rect -1209 -257 -1197 319
rect -1163 -257 -1151 319
rect -1209 -269 -1151 -257
rect -1091 319 -1033 331
rect -1091 -257 -1079 319
rect -1045 -257 -1033 319
rect -1091 -269 -1033 -257
rect -973 319 -915 331
rect -973 -257 -961 319
rect -927 -257 -915 319
rect -973 -269 -915 -257
rect -855 319 -797 331
rect -855 -257 -843 319
rect -809 -257 -797 319
rect -855 -269 -797 -257
rect -737 319 -679 331
rect -737 -257 -725 319
rect -691 -257 -679 319
rect -737 -269 -679 -257
rect -619 319 -561 331
rect -619 -257 -607 319
rect -573 -257 -561 319
rect -619 -269 -561 -257
rect -501 319 -443 331
rect -501 -257 -489 319
rect -455 -257 -443 319
rect -501 -269 -443 -257
rect -383 319 -325 331
rect -383 -257 -371 319
rect -337 -257 -325 319
rect -383 -269 -325 -257
rect -265 319 -207 331
rect -265 -257 -253 319
rect -219 -257 -207 319
rect -265 -269 -207 -257
rect -147 319 -89 331
rect -147 -257 -135 319
rect -101 -257 -89 319
rect -147 -269 -89 -257
rect -29 319 29 331
rect -29 -257 -17 319
rect 17 -257 29 319
rect -29 -269 29 -257
rect 89 319 147 331
rect 89 -257 101 319
rect 135 -257 147 319
rect 89 -269 147 -257
rect 207 319 265 331
rect 207 -257 219 319
rect 253 -257 265 319
rect 207 -269 265 -257
rect 325 319 383 331
rect 325 -257 337 319
rect 371 -257 383 319
rect 325 -269 383 -257
rect 443 319 501 331
rect 443 -257 455 319
rect 489 -257 501 319
rect 443 -269 501 -257
rect 561 319 619 331
rect 561 -257 573 319
rect 607 -257 619 319
rect 561 -269 619 -257
rect 679 319 737 331
rect 679 -257 691 319
rect 725 -257 737 319
rect 679 -269 737 -257
rect 797 319 855 331
rect 797 -257 809 319
rect 843 -257 855 319
rect 797 -269 855 -257
rect 915 319 973 331
rect 915 -257 927 319
rect 961 -257 973 319
rect 915 -269 973 -257
rect 1033 319 1091 331
rect 1033 -257 1045 319
rect 1079 -257 1091 319
rect 1033 -269 1091 -257
rect 1151 319 1209 331
rect 1151 -257 1163 319
rect 1197 -257 1209 319
rect 1151 -269 1209 -257
rect 1269 319 1327 331
rect 1269 -257 1281 319
rect 1315 -257 1327 319
rect 1269 -269 1327 -257
rect 1387 319 1445 331
rect 1387 -257 1399 319
rect 1433 -257 1445 319
rect 1387 -269 1445 -257
rect 1505 319 1563 331
rect 1505 -257 1517 319
rect 1551 -257 1563 319
rect 1505 -269 1563 -257
rect 1623 319 1681 331
rect 1623 -257 1635 319
rect 1669 -257 1681 319
rect 1623 -269 1681 -257
rect 1741 319 1799 331
rect 1741 -257 1753 319
rect 1787 -257 1799 319
rect 1741 -269 1799 -257
rect 1859 319 1917 331
rect 1859 -257 1871 319
rect 1905 -257 1917 319
rect 1859 -269 1917 -257
rect 1977 319 2035 331
rect 1977 -257 1989 319
rect 2023 -257 2035 319
rect 1977 -269 2035 -257
rect 2095 319 2153 331
rect 2095 -257 2107 319
rect 2141 -257 2153 319
rect 2095 -269 2153 -257
rect 2213 319 2271 331
rect 2213 -257 2225 319
rect 2259 -257 2271 319
rect 2213 -269 2271 -257
rect 2331 319 2389 331
rect 2331 -257 2343 319
rect 2377 -257 2389 319
rect 2331 -269 2389 -257
rect 2449 319 2507 331
rect 2449 -257 2461 319
rect 2495 -257 2507 319
rect 2449 -269 2507 -257
rect 2567 319 2625 331
rect 2567 -257 2579 319
rect 2613 -257 2625 319
rect 2567 -269 2625 -257
rect 2685 319 2743 331
rect 2685 -257 2697 319
rect 2731 -257 2743 319
rect 2685 -269 2743 -257
rect 2803 319 2861 331
rect 2803 -257 2815 319
rect 2849 -257 2861 319
rect 2803 -269 2861 -257
rect 2921 319 2979 331
rect 2921 -257 2933 319
rect 2967 -257 2979 319
rect 2921 -269 2979 -257
rect 3039 319 3097 331
rect 3039 -257 3051 319
rect 3085 -257 3097 319
rect 3039 -269 3097 -257
rect 3157 319 3215 331
rect 3157 -257 3169 319
rect 3203 -257 3215 319
rect 3157 -269 3215 -257
rect 3275 319 3333 331
rect 3275 -257 3287 319
rect 3321 -257 3333 319
rect 3275 -269 3333 -257
rect 3393 319 3451 331
rect 3393 -257 3405 319
rect 3439 -257 3451 319
rect 3393 -269 3451 -257
rect 3511 319 3569 331
rect 3511 -257 3523 319
rect 3557 -257 3569 319
rect 3511 -269 3569 -257
rect 3629 319 3687 331
rect 3629 -257 3641 319
rect 3675 -257 3687 319
rect 3629 -269 3687 -257
rect 3747 319 3805 331
rect 3747 -257 3759 319
rect 3793 -257 3805 319
rect 3747 -269 3805 -257
rect 3865 319 3923 331
rect 3865 -257 3877 319
rect 3911 -257 3923 319
rect 3865 -269 3923 -257
rect 3983 319 4041 331
rect 3983 -257 3995 319
rect 4029 -257 4041 319
rect 3983 -269 4041 -257
rect 4101 319 4159 331
rect 4101 -257 4113 319
rect 4147 -257 4159 319
rect 4101 -269 4159 -257
rect 4219 319 4277 331
rect 4219 -257 4231 319
rect 4265 -257 4277 319
rect 4219 -269 4277 -257
rect 4337 319 4395 331
rect 4337 -257 4349 319
rect 4383 -257 4395 319
rect 4337 -269 4395 -257
rect 4455 319 4513 331
rect 4455 -257 4467 319
rect 4501 -257 4513 319
rect 4455 -269 4513 -257
rect 4573 319 4631 331
rect 4573 -257 4585 319
rect 4619 -257 4631 319
rect 4573 -269 4631 -257
rect 4691 319 4749 331
rect 4691 -257 4703 319
rect 4737 -257 4749 319
rect 4691 -269 4749 -257
rect 4809 319 4867 331
rect 4809 -257 4821 319
rect 4855 -257 4867 319
rect 4809 -269 4867 -257
rect 4927 319 4985 331
rect 4927 -257 4939 319
rect 4973 -257 4985 319
rect 4927 -269 4985 -257
rect 5045 319 5103 331
rect 5045 -257 5057 319
rect 5091 -257 5103 319
rect 5045 -269 5103 -257
rect 5163 319 5221 331
rect 5163 -257 5175 319
rect 5209 -257 5221 319
rect 5163 -269 5221 -257
rect 5281 319 5339 331
rect 5281 -257 5293 319
rect 5327 -257 5339 319
rect 5281 -269 5339 -257
rect 5399 319 5457 331
rect 5399 -257 5411 319
rect 5445 -257 5457 319
rect 5399 -269 5457 -257
rect 5517 319 5575 331
rect 5517 -257 5529 319
rect 5563 -257 5575 319
rect 5517 -269 5575 -257
rect 5635 319 5693 331
rect 5635 -257 5647 319
rect 5681 -257 5693 319
rect 5635 -269 5693 -257
rect 5753 319 5811 331
rect 5753 -257 5765 319
rect 5799 -257 5811 319
rect 5753 -269 5811 -257
rect 5871 319 5929 331
rect 5871 -257 5883 319
rect 5917 -257 5929 319
rect 5871 -269 5929 -257
<< ndiffc >>
rect -5917 -257 -5883 319
rect -5799 -257 -5765 319
rect -5681 -257 -5647 319
rect -5563 -257 -5529 319
rect -5445 -257 -5411 319
rect -5327 -257 -5293 319
rect -5209 -257 -5175 319
rect -5091 -257 -5057 319
rect -4973 -257 -4939 319
rect -4855 -257 -4821 319
rect -4737 -257 -4703 319
rect -4619 -257 -4585 319
rect -4501 -257 -4467 319
rect -4383 -257 -4349 319
rect -4265 -257 -4231 319
rect -4147 -257 -4113 319
rect -4029 -257 -3995 319
rect -3911 -257 -3877 319
rect -3793 -257 -3759 319
rect -3675 -257 -3641 319
rect -3557 -257 -3523 319
rect -3439 -257 -3405 319
rect -3321 -257 -3287 319
rect -3203 -257 -3169 319
rect -3085 -257 -3051 319
rect -2967 -257 -2933 319
rect -2849 -257 -2815 319
rect -2731 -257 -2697 319
rect -2613 -257 -2579 319
rect -2495 -257 -2461 319
rect -2377 -257 -2343 319
rect -2259 -257 -2225 319
rect -2141 -257 -2107 319
rect -2023 -257 -1989 319
rect -1905 -257 -1871 319
rect -1787 -257 -1753 319
rect -1669 -257 -1635 319
rect -1551 -257 -1517 319
rect -1433 -257 -1399 319
rect -1315 -257 -1281 319
rect -1197 -257 -1163 319
rect -1079 -257 -1045 319
rect -961 -257 -927 319
rect -843 -257 -809 319
rect -725 -257 -691 319
rect -607 -257 -573 319
rect -489 -257 -455 319
rect -371 -257 -337 319
rect -253 -257 -219 319
rect -135 -257 -101 319
rect -17 -257 17 319
rect 101 -257 135 319
rect 219 -257 253 319
rect 337 -257 371 319
rect 455 -257 489 319
rect 573 -257 607 319
rect 691 -257 725 319
rect 809 -257 843 319
rect 927 -257 961 319
rect 1045 -257 1079 319
rect 1163 -257 1197 319
rect 1281 -257 1315 319
rect 1399 -257 1433 319
rect 1517 -257 1551 319
rect 1635 -257 1669 319
rect 1753 -257 1787 319
rect 1871 -257 1905 319
rect 1989 -257 2023 319
rect 2107 -257 2141 319
rect 2225 -257 2259 319
rect 2343 -257 2377 319
rect 2461 -257 2495 319
rect 2579 -257 2613 319
rect 2697 -257 2731 319
rect 2815 -257 2849 319
rect 2933 -257 2967 319
rect 3051 -257 3085 319
rect 3169 -257 3203 319
rect 3287 -257 3321 319
rect 3405 -257 3439 319
rect 3523 -257 3557 319
rect 3641 -257 3675 319
rect 3759 -257 3793 319
rect 3877 -257 3911 319
rect 3995 -257 4029 319
rect 4113 -257 4147 319
rect 4231 -257 4265 319
rect 4349 -257 4383 319
rect 4467 -257 4501 319
rect 4585 -257 4619 319
rect 4703 -257 4737 319
rect 4821 -257 4855 319
rect 4939 -257 4973 319
rect 5057 -257 5091 319
rect 5175 -257 5209 319
rect 5293 -257 5327 319
rect 5411 -257 5445 319
rect 5529 -257 5563 319
rect 5647 -257 5681 319
rect 5765 -257 5799 319
rect 5883 -257 5917 319
<< poly >>
rect -5871 331 -5811 357
rect -5753 331 -5693 357
rect -5635 331 -5575 357
rect -5517 331 -5457 357
rect -5399 331 -5339 357
rect -5281 331 -5221 357
rect -5163 331 -5103 357
rect -5045 331 -4985 357
rect -4927 331 -4867 357
rect -4809 331 -4749 357
rect -4691 331 -4631 357
rect -4573 331 -4513 357
rect -4455 331 -4395 357
rect -4337 331 -4277 357
rect -4219 331 -4159 357
rect -4101 331 -4041 357
rect -3983 331 -3923 357
rect -3865 331 -3805 357
rect -3747 331 -3687 357
rect -3629 331 -3569 357
rect -3511 331 -3451 357
rect -3393 331 -3333 357
rect -3275 331 -3215 357
rect -3157 331 -3097 357
rect -3039 331 -2979 357
rect -2921 331 -2861 357
rect -2803 331 -2743 357
rect -2685 331 -2625 357
rect -2567 331 -2507 357
rect -2449 331 -2389 357
rect -2331 331 -2271 357
rect -2213 331 -2153 357
rect -2095 331 -2035 357
rect -1977 331 -1917 357
rect -1859 331 -1799 357
rect -1741 331 -1681 357
rect -1623 331 -1563 357
rect -1505 331 -1445 357
rect -1387 331 -1327 357
rect -1269 331 -1209 357
rect -1151 331 -1091 357
rect -1033 331 -973 357
rect -915 331 -855 357
rect -797 331 -737 357
rect -679 331 -619 357
rect -561 331 -501 357
rect -443 331 -383 357
rect -325 331 -265 357
rect -207 331 -147 357
rect -89 331 -29 357
rect 29 331 89 357
rect 147 331 207 357
rect 265 331 325 357
rect 383 331 443 357
rect 501 331 561 357
rect 619 331 679 357
rect 737 331 797 357
rect 855 331 915 357
rect 973 331 1033 357
rect 1091 331 1151 357
rect 1209 331 1269 357
rect 1327 331 1387 357
rect 1445 331 1505 357
rect 1563 331 1623 357
rect 1681 331 1741 357
rect 1799 331 1859 357
rect 1917 331 1977 357
rect 2035 331 2095 357
rect 2153 331 2213 357
rect 2271 331 2331 357
rect 2389 331 2449 357
rect 2507 331 2567 357
rect 2625 331 2685 357
rect 2743 331 2803 357
rect 2861 331 2921 357
rect 2979 331 3039 357
rect 3097 331 3157 357
rect 3215 331 3275 357
rect 3333 331 3393 357
rect 3451 331 3511 357
rect 3569 331 3629 357
rect 3687 331 3747 357
rect 3805 331 3865 357
rect 3923 331 3983 357
rect 4041 331 4101 357
rect 4159 331 4219 357
rect 4277 331 4337 357
rect 4395 331 4455 357
rect 4513 331 4573 357
rect 4631 331 4691 357
rect 4749 331 4809 357
rect 4867 331 4927 357
rect 4985 331 5045 357
rect 5103 331 5163 357
rect 5221 331 5281 357
rect 5339 331 5399 357
rect 5457 331 5517 357
rect 5575 331 5635 357
rect 5693 331 5753 357
rect 5811 331 5871 357
rect -5871 -291 -5811 -269
rect -5753 -291 -5693 -269
rect -5635 -291 -5575 -269
rect -5517 -291 -5457 -269
rect -5399 -291 -5339 -269
rect -5281 -291 -5221 -269
rect -5163 -291 -5103 -269
rect -5045 -291 -4985 -269
rect -4927 -291 -4867 -269
rect -4809 -291 -4749 -269
rect -4691 -291 -4631 -269
rect -4573 -291 -4513 -269
rect -4455 -291 -4395 -269
rect -4337 -291 -4277 -269
rect -4219 -291 -4159 -269
rect -4101 -291 -4041 -269
rect -3983 -291 -3923 -269
rect -3865 -291 -3805 -269
rect -3747 -291 -3687 -269
rect -3629 -291 -3569 -269
rect -3511 -291 -3451 -269
rect -3393 -291 -3333 -269
rect -3275 -291 -3215 -269
rect -3157 -291 -3097 -269
rect -3039 -291 -2979 -269
rect -2921 -291 -2861 -269
rect -2803 -291 -2743 -269
rect -2685 -291 -2625 -269
rect -2567 -291 -2507 -269
rect -2449 -291 -2389 -269
rect -2331 -291 -2271 -269
rect -2213 -291 -2153 -269
rect -2095 -291 -2035 -269
rect -1977 -291 -1917 -269
rect -1859 -291 -1799 -269
rect -1741 -291 -1681 -269
rect -1623 -291 -1563 -269
rect -1505 -291 -1445 -269
rect -1387 -291 -1327 -269
rect -1269 -291 -1209 -269
rect -1151 -291 -1091 -269
rect -1033 -291 -973 -269
rect -915 -291 -855 -269
rect -797 -291 -737 -269
rect -679 -291 -619 -269
rect -561 -291 -501 -269
rect -443 -291 -383 -269
rect -325 -291 -265 -269
rect -207 -291 -147 -269
rect -89 -291 -29 -269
rect 29 -291 89 -269
rect 147 -291 207 -269
rect 265 -291 325 -269
rect 383 -291 443 -269
rect 501 -291 561 -269
rect 619 -291 679 -269
rect 737 -291 797 -269
rect 855 -291 915 -269
rect 973 -291 1033 -269
rect 1091 -291 1151 -269
rect 1209 -291 1269 -269
rect 1327 -291 1387 -269
rect 1445 -291 1505 -269
rect 1563 -291 1623 -269
rect 1681 -291 1741 -269
rect 1799 -291 1859 -269
rect 1917 -291 1977 -269
rect 2035 -291 2095 -269
rect 2153 -291 2213 -269
rect 2271 -291 2331 -269
rect 2389 -291 2449 -269
rect 2507 -291 2567 -269
rect 2625 -291 2685 -269
rect 2743 -291 2803 -269
rect 2861 -291 2921 -269
rect 2979 -291 3039 -269
rect 3097 -291 3157 -269
rect 3215 -291 3275 -269
rect 3333 -291 3393 -269
rect 3451 -291 3511 -269
rect 3569 -291 3629 -269
rect 3687 -291 3747 -269
rect 3805 -291 3865 -269
rect 3923 -291 3983 -269
rect 4041 -291 4101 -269
rect 4159 -291 4219 -269
rect 4277 -291 4337 -269
rect 4395 -291 4455 -269
rect 4513 -291 4573 -269
rect 4631 -291 4691 -269
rect 4749 -291 4809 -269
rect 4867 -291 4927 -269
rect 4985 -291 5045 -269
rect 5103 -291 5163 -269
rect 5221 -291 5281 -269
rect 5339 -291 5399 -269
rect 5457 -291 5517 -269
rect 5575 -291 5635 -269
rect 5693 -291 5753 -269
rect 5811 -291 5871 -269
rect -5874 -307 -5808 -291
rect -5874 -341 -5858 -307
rect -5824 -341 -5808 -307
rect -5874 -357 -5808 -341
rect -5756 -307 -5690 -291
rect -5756 -341 -5740 -307
rect -5706 -341 -5690 -307
rect -5756 -357 -5690 -341
rect -5638 -307 -5572 -291
rect -5638 -341 -5622 -307
rect -5588 -341 -5572 -307
rect -5638 -357 -5572 -341
rect -5520 -307 -5454 -291
rect -5520 -341 -5504 -307
rect -5470 -341 -5454 -307
rect -5520 -357 -5454 -341
rect -5402 -307 -5336 -291
rect -5402 -341 -5386 -307
rect -5352 -341 -5336 -307
rect -5402 -357 -5336 -341
rect -5284 -307 -5218 -291
rect -5284 -341 -5268 -307
rect -5234 -341 -5218 -307
rect -5284 -357 -5218 -341
rect -5166 -307 -5100 -291
rect -5166 -341 -5150 -307
rect -5116 -341 -5100 -307
rect -5166 -357 -5100 -341
rect -5048 -307 -4982 -291
rect -5048 -341 -5032 -307
rect -4998 -341 -4982 -307
rect -5048 -357 -4982 -341
rect -4930 -307 -4864 -291
rect -4930 -341 -4914 -307
rect -4880 -341 -4864 -307
rect -4930 -357 -4864 -341
rect -4812 -307 -4746 -291
rect -4812 -341 -4796 -307
rect -4762 -341 -4746 -307
rect -4812 -357 -4746 -341
rect -4694 -307 -4628 -291
rect -4694 -341 -4678 -307
rect -4644 -341 -4628 -307
rect -4694 -357 -4628 -341
rect -4576 -307 -4510 -291
rect -4576 -341 -4560 -307
rect -4526 -341 -4510 -307
rect -4576 -357 -4510 -341
rect -4458 -307 -4392 -291
rect -4458 -341 -4442 -307
rect -4408 -341 -4392 -307
rect -4458 -357 -4392 -341
rect -4340 -307 -4274 -291
rect -4340 -341 -4324 -307
rect -4290 -341 -4274 -307
rect -4340 -357 -4274 -341
rect -4222 -307 -4156 -291
rect -4222 -341 -4206 -307
rect -4172 -341 -4156 -307
rect -4222 -357 -4156 -341
rect -4104 -307 -4038 -291
rect -4104 -341 -4088 -307
rect -4054 -341 -4038 -307
rect -4104 -357 -4038 -341
rect -3986 -307 -3920 -291
rect -3986 -341 -3970 -307
rect -3936 -341 -3920 -307
rect -3986 -357 -3920 -341
rect -3868 -307 -3802 -291
rect -3868 -341 -3852 -307
rect -3818 -341 -3802 -307
rect -3868 -357 -3802 -341
rect -3750 -307 -3684 -291
rect -3750 -341 -3734 -307
rect -3700 -341 -3684 -307
rect -3750 -357 -3684 -341
rect -3632 -307 -3566 -291
rect -3632 -341 -3616 -307
rect -3582 -341 -3566 -307
rect -3632 -357 -3566 -341
rect -3514 -307 -3448 -291
rect -3514 -341 -3498 -307
rect -3464 -341 -3448 -307
rect -3514 -357 -3448 -341
rect -3396 -307 -3330 -291
rect -3396 -341 -3380 -307
rect -3346 -341 -3330 -307
rect -3396 -357 -3330 -341
rect -3278 -307 -3212 -291
rect -3278 -341 -3262 -307
rect -3228 -341 -3212 -307
rect -3278 -357 -3212 -341
rect -3160 -307 -3094 -291
rect -3160 -341 -3144 -307
rect -3110 -341 -3094 -307
rect -3160 -357 -3094 -341
rect -3042 -307 -2976 -291
rect -3042 -341 -3026 -307
rect -2992 -341 -2976 -307
rect -3042 -357 -2976 -341
rect -2924 -307 -2858 -291
rect -2924 -341 -2908 -307
rect -2874 -341 -2858 -307
rect -2924 -357 -2858 -341
rect -2806 -307 -2740 -291
rect -2806 -341 -2790 -307
rect -2756 -341 -2740 -307
rect -2806 -357 -2740 -341
rect -2688 -307 -2622 -291
rect -2688 -341 -2672 -307
rect -2638 -341 -2622 -307
rect -2688 -357 -2622 -341
rect -2570 -307 -2504 -291
rect -2570 -341 -2554 -307
rect -2520 -341 -2504 -307
rect -2570 -357 -2504 -341
rect -2452 -307 -2386 -291
rect -2452 -341 -2436 -307
rect -2402 -341 -2386 -307
rect -2452 -357 -2386 -341
rect -2334 -307 -2268 -291
rect -2334 -341 -2318 -307
rect -2284 -341 -2268 -307
rect -2334 -357 -2268 -341
rect -2216 -307 -2150 -291
rect -2216 -341 -2200 -307
rect -2166 -341 -2150 -307
rect -2216 -357 -2150 -341
rect -2098 -307 -2032 -291
rect -2098 -341 -2082 -307
rect -2048 -341 -2032 -307
rect -2098 -357 -2032 -341
rect -1980 -307 -1914 -291
rect -1980 -341 -1964 -307
rect -1930 -341 -1914 -307
rect -1980 -357 -1914 -341
rect -1862 -307 -1796 -291
rect -1862 -341 -1846 -307
rect -1812 -341 -1796 -307
rect -1862 -357 -1796 -341
rect -1744 -307 -1678 -291
rect -1744 -341 -1728 -307
rect -1694 -341 -1678 -307
rect -1744 -357 -1678 -341
rect -1626 -307 -1560 -291
rect -1626 -341 -1610 -307
rect -1576 -341 -1560 -307
rect -1626 -357 -1560 -341
rect -1508 -307 -1442 -291
rect -1508 -341 -1492 -307
rect -1458 -341 -1442 -307
rect -1508 -357 -1442 -341
rect -1390 -307 -1324 -291
rect -1390 -341 -1374 -307
rect -1340 -341 -1324 -307
rect -1390 -357 -1324 -341
rect -1272 -307 -1206 -291
rect -1272 -341 -1256 -307
rect -1222 -341 -1206 -307
rect -1272 -357 -1206 -341
rect -1154 -307 -1088 -291
rect -1154 -341 -1138 -307
rect -1104 -341 -1088 -307
rect -1154 -357 -1088 -341
rect -1036 -307 -970 -291
rect -1036 -341 -1020 -307
rect -986 -341 -970 -307
rect -1036 -357 -970 -341
rect -918 -307 -852 -291
rect -918 -341 -902 -307
rect -868 -341 -852 -307
rect -918 -357 -852 -341
rect -800 -307 -734 -291
rect -800 -341 -784 -307
rect -750 -341 -734 -307
rect -800 -357 -734 -341
rect -682 -307 -616 -291
rect -682 -341 -666 -307
rect -632 -341 -616 -307
rect -682 -357 -616 -341
rect -564 -307 -498 -291
rect -564 -341 -548 -307
rect -514 -341 -498 -307
rect -564 -357 -498 -341
rect -446 -307 -380 -291
rect -446 -341 -430 -307
rect -396 -341 -380 -307
rect -446 -357 -380 -341
rect -328 -307 -262 -291
rect -328 -341 -312 -307
rect -278 -341 -262 -307
rect -328 -357 -262 -341
rect -210 -307 -144 -291
rect -210 -341 -194 -307
rect -160 -341 -144 -307
rect -210 -357 -144 -341
rect -92 -307 -26 -291
rect -92 -341 -76 -307
rect -42 -341 -26 -307
rect -92 -357 -26 -341
rect 26 -307 92 -291
rect 26 -341 42 -307
rect 76 -341 92 -307
rect 26 -357 92 -341
rect 144 -307 210 -291
rect 144 -341 160 -307
rect 194 -341 210 -307
rect 144 -357 210 -341
rect 262 -307 328 -291
rect 262 -341 278 -307
rect 312 -341 328 -307
rect 262 -357 328 -341
rect 380 -307 446 -291
rect 380 -341 396 -307
rect 430 -341 446 -307
rect 380 -357 446 -341
rect 498 -307 564 -291
rect 498 -341 514 -307
rect 548 -341 564 -307
rect 498 -357 564 -341
rect 616 -307 682 -291
rect 616 -341 632 -307
rect 666 -341 682 -307
rect 616 -357 682 -341
rect 734 -307 800 -291
rect 734 -341 750 -307
rect 784 -341 800 -307
rect 734 -357 800 -341
rect 852 -307 918 -291
rect 852 -341 868 -307
rect 902 -341 918 -307
rect 852 -357 918 -341
rect 970 -307 1036 -291
rect 970 -341 986 -307
rect 1020 -341 1036 -307
rect 970 -357 1036 -341
rect 1088 -307 1154 -291
rect 1088 -341 1104 -307
rect 1138 -341 1154 -307
rect 1088 -357 1154 -341
rect 1206 -307 1272 -291
rect 1206 -341 1222 -307
rect 1256 -341 1272 -307
rect 1206 -357 1272 -341
rect 1324 -307 1390 -291
rect 1324 -341 1340 -307
rect 1374 -341 1390 -307
rect 1324 -357 1390 -341
rect 1442 -307 1508 -291
rect 1442 -341 1458 -307
rect 1492 -341 1508 -307
rect 1442 -357 1508 -341
rect 1560 -307 1626 -291
rect 1560 -341 1576 -307
rect 1610 -341 1626 -307
rect 1560 -357 1626 -341
rect 1678 -307 1744 -291
rect 1678 -341 1694 -307
rect 1728 -341 1744 -307
rect 1678 -357 1744 -341
rect 1796 -307 1862 -291
rect 1796 -341 1812 -307
rect 1846 -341 1862 -307
rect 1796 -357 1862 -341
rect 1914 -307 1980 -291
rect 1914 -341 1930 -307
rect 1964 -341 1980 -307
rect 1914 -357 1980 -341
rect 2032 -307 2098 -291
rect 2032 -341 2048 -307
rect 2082 -341 2098 -307
rect 2032 -357 2098 -341
rect 2150 -307 2216 -291
rect 2150 -341 2166 -307
rect 2200 -341 2216 -307
rect 2150 -357 2216 -341
rect 2268 -307 2334 -291
rect 2268 -341 2284 -307
rect 2318 -341 2334 -307
rect 2268 -357 2334 -341
rect 2386 -307 2452 -291
rect 2386 -341 2402 -307
rect 2436 -341 2452 -307
rect 2386 -357 2452 -341
rect 2504 -307 2570 -291
rect 2504 -341 2520 -307
rect 2554 -341 2570 -307
rect 2504 -357 2570 -341
rect 2622 -307 2688 -291
rect 2622 -341 2638 -307
rect 2672 -341 2688 -307
rect 2622 -357 2688 -341
rect 2740 -307 2806 -291
rect 2740 -341 2756 -307
rect 2790 -341 2806 -307
rect 2740 -357 2806 -341
rect 2858 -307 2924 -291
rect 2858 -341 2874 -307
rect 2908 -341 2924 -307
rect 2858 -357 2924 -341
rect 2976 -307 3042 -291
rect 2976 -341 2992 -307
rect 3026 -341 3042 -307
rect 2976 -357 3042 -341
rect 3094 -307 3160 -291
rect 3094 -341 3110 -307
rect 3144 -341 3160 -307
rect 3094 -357 3160 -341
rect 3212 -307 3278 -291
rect 3212 -341 3228 -307
rect 3262 -341 3278 -307
rect 3212 -357 3278 -341
rect 3330 -307 3396 -291
rect 3330 -341 3346 -307
rect 3380 -341 3396 -307
rect 3330 -357 3396 -341
rect 3448 -307 3514 -291
rect 3448 -341 3464 -307
rect 3498 -341 3514 -307
rect 3448 -357 3514 -341
rect 3566 -307 3632 -291
rect 3566 -341 3582 -307
rect 3616 -341 3632 -307
rect 3566 -357 3632 -341
rect 3684 -307 3750 -291
rect 3684 -341 3700 -307
rect 3734 -341 3750 -307
rect 3684 -357 3750 -341
rect 3802 -307 3868 -291
rect 3802 -341 3818 -307
rect 3852 -341 3868 -307
rect 3802 -357 3868 -341
rect 3920 -307 3986 -291
rect 3920 -341 3936 -307
rect 3970 -341 3986 -307
rect 3920 -357 3986 -341
rect 4038 -307 4104 -291
rect 4038 -341 4054 -307
rect 4088 -341 4104 -307
rect 4038 -357 4104 -341
rect 4156 -307 4222 -291
rect 4156 -341 4172 -307
rect 4206 -341 4222 -307
rect 4156 -357 4222 -341
rect 4274 -307 4340 -291
rect 4274 -341 4290 -307
rect 4324 -341 4340 -307
rect 4274 -357 4340 -341
rect 4392 -307 4458 -291
rect 4392 -341 4408 -307
rect 4442 -341 4458 -307
rect 4392 -357 4458 -341
rect 4510 -307 4576 -291
rect 4510 -341 4526 -307
rect 4560 -341 4576 -307
rect 4510 -357 4576 -341
rect 4628 -307 4694 -291
rect 4628 -341 4644 -307
rect 4678 -341 4694 -307
rect 4628 -357 4694 -341
rect 4746 -307 4812 -291
rect 4746 -341 4762 -307
rect 4796 -341 4812 -307
rect 4746 -357 4812 -341
rect 4864 -307 4930 -291
rect 4864 -341 4880 -307
rect 4914 -341 4930 -307
rect 4864 -357 4930 -341
rect 4982 -307 5048 -291
rect 4982 -341 4998 -307
rect 5032 -341 5048 -307
rect 4982 -357 5048 -341
rect 5100 -307 5166 -291
rect 5100 -341 5116 -307
rect 5150 -341 5166 -307
rect 5100 -357 5166 -341
rect 5218 -307 5284 -291
rect 5218 -341 5234 -307
rect 5268 -341 5284 -307
rect 5218 -357 5284 -341
rect 5336 -307 5402 -291
rect 5336 -341 5352 -307
rect 5386 -341 5402 -307
rect 5336 -357 5402 -341
rect 5454 -307 5520 -291
rect 5454 -341 5470 -307
rect 5504 -341 5520 -307
rect 5454 -357 5520 -341
rect 5572 -307 5638 -291
rect 5572 -341 5588 -307
rect 5622 -341 5638 -307
rect 5572 -357 5638 -341
rect 5690 -307 5756 -291
rect 5690 -341 5706 -307
rect 5740 -341 5756 -307
rect 5690 -357 5756 -341
rect 5808 -307 5874 -291
rect 5808 -341 5824 -307
rect 5858 -341 5874 -307
rect 5808 -357 5874 -341
<< polycont >>
rect -5858 -341 -5824 -307
rect -5740 -341 -5706 -307
rect -5622 -341 -5588 -307
rect -5504 -341 -5470 -307
rect -5386 -341 -5352 -307
rect -5268 -341 -5234 -307
rect -5150 -341 -5116 -307
rect -5032 -341 -4998 -307
rect -4914 -341 -4880 -307
rect -4796 -341 -4762 -307
rect -4678 -341 -4644 -307
rect -4560 -341 -4526 -307
rect -4442 -341 -4408 -307
rect -4324 -341 -4290 -307
rect -4206 -341 -4172 -307
rect -4088 -341 -4054 -307
rect -3970 -341 -3936 -307
rect -3852 -341 -3818 -307
rect -3734 -341 -3700 -307
rect -3616 -341 -3582 -307
rect -3498 -341 -3464 -307
rect -3380 -341 -3346 -307
rect -3262 -341 -3228 -307
rect -3144 -341 -3110 -307
rect -3026 -341 -2992 -307
rect -2908 -341 -2874 -307
rect -2790 -341 -2756 -307
rect -2672 -341 -2638 -307
rect -2554 -341 -2520 -307
rect -2436 -341 -2402 -307
rect -2318 -341 -2284 -307
rect -2200 -341 -2166 -307
rect -2082 -341 -2048 -307
rect -1964 -341 -1930 -307
rect -1846 -341 -1812 -307
rect -1728 -341 -1694 -307
rect -1610 -341 -1576 -307
rect -1492 -341 -1458 -307
rect -1374 -341 -1340 -307
rect -1256 -341 -1222 -307
rect -1138 -341 -1104 -307
rect -1020 -341 -986 -307
rect -902 -341 -868 -307
rect -784 -341 -750 -307
rect -666 -341 -632 -307
rect -548 -341 -514 -307
rect -430 -341 -396 -307
rect -312 -341 -278 -307
rect -194 -341 -160 -307
rect -76 -341 -42 -307
rect 42 -341 76 -307
rect 160 -341 194 -307
rect 278 -341 312 -307
rect 396 -341 430 -307
rect 514 -341 548 -307
rect 632 -341 666 -307
rect 750 -341 784 -307
rect 868 -341 902 -307
rect 986 -341 1020 -307
rect 1104 -341 1138 -307
rect 1222 -341 1256 -307
rect 1340 -341 1374 -307
rect 1458 -341 1492 -307
rect 1576 -341 1610 -307
rect 1694 -341 1728 -307
rect 1812 -341 1846 -307
rect 1930 -341 1964 -307
rect 2048 -341 2082 -307
rect 2166 -341 2200 -307
rect 2284 -341 2318 -307
rect 2402 -341 2436 -307
rect 2520 -341 2554 -307
rect 2638 -341 2672 -307
rect 2756 -341 2790 -307
rect 2874 -341 2908 -307
rect 2992 -341 3026 -307
rect 3110 -341 3144 -307
rect 3228 -341 3262 -307
rect 3346 -341 3380 -307
rect 3464 -341 3498 -307
rect 3582 -341 3616 -307
rect 3700 -341 3734 -307
rect 3818 -341 3852 -307
rect 3936 -341 3970 -307
rect 4054 -341 4088 -307
rect 4172 -341 4206 -307
rect 4290 -341 4324 -307
rect 4408 -341 4442 -307
rect 4526 -341 4560 -307
rect 4644 -341 4678 -307
rect 4762 -341 4796 -307
rect 4880 -341 4914 -307
rect 4998 -341 5032 -307
rect 5116 -341 5150 -307
rect 5234 -341 5268 -307
rect 5352 -341 5386 -307
rect 5470 -341 5504 -307
rect 5588 -341 5622 -307
rect 5706 -341 5740 -307
rect 5824 -341 5858 -307
<< locali >>
rect -5917 319 -5883 335
rect -5917 -273 -5883 -257
rect -5799 319 -5765 335
rect -5799 -273 -5765 -257
rect -5681 319 -5647 335
rect -5681 -273 -5647 -257
rect -5563 319 -5529 335
rect -5563 -273 -5529 -257
rect -5445 319 -5411 335
rect -5445 -273 -5411 -257
rect -5327 319 -5293 335
rect -5327 -273 -5293 -257
rect -5209 319 -5175 335
rect -5209 -273 -5175 -257
rect -5091 319 -5057 335
rect -5091 -273 -5057 -257
rect -4973 319 -4939 335
rect -4973 -273 -4939 -257
rect -4855 319 -4821 335
rect -4855 -273 -4821 -257
rect -4737 319 -4703 335
rect -4737 -273 -4703 -257
rect -4619 319 -4585 335
rect -4619 -273 -4585 -257
rect -4501 319 -4467 335
rect -4501 -273 -4467 -257
rect -4383 319 -4349 335
rect -4383 -273 -4349 -257
rect -4265 319 -4231 335
rect -4265 -273 -4231 -257
rect -4147 319 -4113 335
rect -4147 -273 -4113 -257
rect -4029 319 -3995 335
rect -4029 -273 -3995 -257
rect -3911 319 -3877 335
rect -3911 -273 -3877 -257
rect -3793 319 -3759 335
rect -3793 -273 -3759 -257
rect -3675 319 -3641 335
rect -3675 -273 -3641 -257
rect -3557 319 -3523 335
rect -3557 -273 -3523 -257
rect -3439 319 -3405 335
rect -3439 -273 -3405 -257
rect -3321 319 -3287 335
rect -3321 -273 -3287 -257
rect -3203 319 -3169 335
rect -3203 -273 -3169 -257
rect -3085 319 -3051 335
rect -3085 -273 -3051 -257
rect -2967 319 -2933 335
rect -2967 -273 -2933 -257
rect -2849 319 -2815 335
rect -2849 -273 -2815 -257
rect -2731 319 -2697 335
rect -2731 -273 -2697 -257
rect -2613 319 -2579 335
rect -2613 -273 -2579 -257
rect -2495 319 -2461 335
rect -2495 -273 -2461 -257
rect -2377 319 -2343 335
rect -2377 -273 -2343 -257
rect -2259 319 -2225 335
rect -2259 -273 -2225 -257
rect -2141 319 -2107 335
rect -2141 -273 -2107 -257
rect -2023 319 -1989 335
rect -2023 -273 -1989 -257
rect -1905 319 -1871 335
rect -1905 -273 -1871 -257
rect -1787 319 -1753 335
rect -1787 -273 -1753 -257
rect -1669 319 -1635 335
rect -1669 -273 -1635 -257
rect -1551 319 -1517 335
rect -1551 -273 -1517 -257
rect -1433 319 -1399 335
rect -1433 -273 -1399 -257
rect -1315 319 -1281 335
rect -1315 -273 -1281 -257
rect -1197 319 -1163 335
rect -1197 -273 -1163 -257
rect -1079 319 -1045 335
rect -1079 -273 -1045 -257
rect -961 319 -927 335
rect -961 -273 -927 -257
rect -843 319 -809 335
rect -843 -273 -809 -257
rect -725 319 -691 335
rect -725 -273 -691 -257
rect -607 319 -573 335
rect -607 -273 -573 -257
rect -489 319 -455 335
rect -489 -273 -455 -257
rect -371 319 -337 335
rect -371 -273 -337 -257
rect -253 319 -219 335
rect -253 -273 -219 -257
rect -135 319 -101 335
rect -135 -273 -101 -257
rect -17 319 17 335
rect -17 -273 17 -257
rect 101 319 135 335
rect 101 -273 135 -257
rect 219 319 253 335
rect 219 -273 253 -257
rect 337 319 371 335
rect 337 -273 371 -257
rect 455 319 489 335
rect 455 -273 489 -257
rect 573 319 607 335
rect 573 -273 607 -257
rect 691 319 725 335
rect 691 -273 725 -257
rect 809 319 843 335
rect 809 -273 843 -257
rect 927 319 961 335
rect 927 -273 961 -257
rect 1045 319 1079 335
rect 1045 -273 1079 -257
rect 1163 319 1197 335
rect 1163 -273 1197 -257
rect 1281 319 1315 335
rect 1281 -273 1315 -257
rect 1399 319 1433 335
rect 1399 -273 1433 -257
rect 1517 319 1551 335
rect 1517 -273 1551 -257
rect 1635 319 1669 335
rect 1635 -273 1669 -257
rect 1753 319 1787 335
rect 1753 -273 1787 -257
rect 1871 319 1905 335
rect 1871 -273 1905 -257
rect 1989 319 2023 335
rect 1989 -273 2023 -257
rect 2107 319 2141 335
rect 2107 -273 2141 -257
rect 2225 319 2259 335
rect 2225 -273 2259 -257
rect 2343 319 2377 335
rect 2343 -273 2377 -257
rect 2461 319 2495 335
rect 2461 -273 2495 -257
rect 2579 319 2613 335
rect 2579 -273 2613 -257
rect 2697 319 2731 335
rect 2697 -273 2731 -257
rect 2815 319 2849 335
rect 2815 -273 2849 -257
rect 2933 319 2967 335
rect 2933 -273 2967 -257
rect 3051 319 3085 335
rect 3051 -273 3085 -257
rect 3169 319 3203 335
rect 3169 -273 3203 -257
rect 3287 319 3321 335
rect 3287 -273 3321 -257
rect 3405 319 3439 335
rect 3405 -273 3439 -257
rect 3523 319 3557 335
rect 3523 -273 3557 -257
rect 3641 319 3675 335
rect 3641 -273 3675 -257
rect 3759 319 3793 335
rect 3759 -273 3793 -257
rect 3877 319 3911 335
rect 3877 -273 3911 -257
rect 3995 319 4029 335
rect 3995 -273 4029 -257
rect 4113 319 4147 335
rect 4113 -273 4147 -257
rect 4231 319 4265 335
rect 4231 -273 4265 -257
rect 4349 319 4383 335
rect 4349 -273 4383 -257
rect 4467 319 4501 335
rect 4467 -273 4501 -257
rect 4585 319 4619 335
rect 4585 -273 4619 -257
rect 4703 319 4737 335
rect 4703 -273 4737 -257
rect 4821 319 4855 335
rect 4821 -273 4855 -257
rect 4939 319 4973 335
rect 4939 -273 4973 -257
rect 5057 319 5091 335
rect 5057 -273 5091 -257
rect 5175 319 5209 335
rect 5175 -273 5209 -257
rect 5293 319 5327 335
rect 5293 -273 5327 -257
rect 5411 319 5445 335
rect 5411 -273 5445 -257
rect 5529 319 5563 335
rect 5529 -273 5563 -257
rect 5647 319 5681 335
rect 5647 -273 5681 -257
rect 5765 319 5799 335
rect 5765 -273 5799 -257
rect 5883 319 5917 335
rect 5883 -273 5917 -257
rect -5874 -341 -5858 -307
rect -5824 -341 -5808 -307
rect -5756 -341 -5740 -307
rect -5706 -341 -5690 -307
rect -5638 -341 -5622 -307
rect -5588 -341 -5572 -307
rect -5520 -341 -5504 -307
rect -5470 -341 -5454 -307
rect -5402 -341 -5386 -307
rect -5352 -341 -5336 -307
rect -5284 -341 -5268 -307
rect -5234 -341 -5218 -307
rect -5166 -341 -5150 -307
rect -5116 -341 -5100 -307
rect -5048 -341 -5032 -307
rect -4998 -341 -4982 -307
rect -4930 -341 -4914 -307
rect -4880 -341 -4864 -307
rect -4812 -341 -4796 -307
rect -4762 -341 -4746 -307
rect -4694 -341 -4678 -307
rect -4644 -341 -4628 -307
rect -4576 -341 -4560 -307
rect -4526 -341 -4510 -307
rect -4458 -341 -4442 -307
rect -4408 -341 -4392 -307
rect -4340 -341 -4324 -307
rect -4290 -341 -4274 -307
rect -4222 -341 -4206 -307
rect -4172 -341 -4156 -307
rect -4104 -341 -4088 -307
rect -4054 -341 -4038 -307
rect -3986 -341 -3970 -307
rect -3936 -341 -3920 -307
rect -3868 -341 -3852 -307
rect -3818 -341 -3802 -307
rect -3750 -341 -3734 -307
rect -3700 -341 -3684 -307
rect -3632 -341 -3616 -307
rect -3582 -341 -3566 -307
rect -3514 -341 -3498 -307
rect -3464 -341 -3448 -307
rect -3396 -341 -3380 -307
rect -3346 -341 -3330 -307
rect -3278 -341 -3262 -307
rect -3228 -341 -3212 -307
rect -3160 -341 -3144 -307
rect -3110 -341 -3094 -307
rect -3042 -341 -3026 -307
rect -2992 -341 -2976 -307
rect -2924 -341 -2908 -307
rect -2874 -341 -2858 -307
rect -2806 -341 -2790 -307
rect -2756 -341 -2740 -307
rect -2688 -341 -2672 -307
rect -2638 -341 -2622 -307
rect -2570 -341 -2554 -307
rect -2520 -341 -2504 -307
rect -2452 -341 -2436 -307
rect -2402 -341 -2386 -307
rect -2334 -341 -2318 -307
rect -2284 -341 -2268 -307
rect -2216 -341 -2200 -307
rect -2166 -341 -2150 -307
rect -2098 -341 -2082 -307
rect -2048 -341 -2032 -307
rect -1980 -341 -1964 -307
rect -1930 -341 -1914 -307
rect -1862 -341 -1846 -307
rect -1812 -341 -1796 -307
rect -1744 -341 -1728 -307
rect -1694 -341 -1678 -307
rect -1626 -341 -1610 -307
rect -1576 -341 -1560 -307
rect -1508 -341 -1492 -307
rect -1458 -341 -1442 -307
rect -1390 -341 -1374 -307
rect -1340 -341 -1324 -307
rect -1272 -341 -1256 -307
rect -1222 -341 -1206 -307
rect -1154 -341 -1138 -307
rect -1104 -341 -1088 -307
rect -1036 -341 -1020 -307
rect -986 -341 -970 -307
rect -918 -341 -902 -307
rect -868 -341 -852 -307
rect -800 -341 -784 -307
rect -750 -341 -734 -307
rect -682 -341 -666 -307
rect -632 -341 -616 -307
rect -564 -341 -548 -307
rect -514 -341 -498 -307
rect -446 -341 -430 -307
rect -396 -341 -380 -307
rect -328 -341 -312 -307
rect -278 -341 -262 -307
rect -210 -341 -194 -307
rect -160 -341 -144 -307
rect -92 -341 -76 -307
rect -42 -341 -26 -307
rect 26 -341 42 -307
rect 76 -341 92 -307
rect 144 -341 160 -307
rect 194 -341 210 -307
rect 262 -341 278 -307
rect 312 -341 328 -307
rect 380 -341 396 -307
rect 430 -341 446 -307
rect 498 -341 514 -307
rect 548 -341 564 -307
rect 616 -341 632 -307
rect 666 -341 682 -307
rect 734 -341 750 -307
rect 784 -341 800 -307
rect 852 -341 868 -307
rect 902 -341 918 -307
rect 970 -341 986 -307
rect 1020 -341 1036 -307
rect 1088 -341 1104 -307
rect 1138 -341 1154 -307
rect 1206 -341 1222 -307
rect 1256 -341 1272 -307
rect 1324 -341 1340 -307
rect 1374 -341 1390 -307
rect 1442 -341 1458 -307
rect 1492 -341 1508 -307
rect 1560 -341 1576 -307
rect 1610 -341 1626 -307
rect 1678 -341 1694 -307
rect 1728 -341 1744 -307
rect 1796 -341 1812 -307
rect 1846 -341 1862 -307
rect 1914 -341 1930 -307
rect 1964 -341 1980 -307
rect 2032 -341 2048 -307
rect 2082 -341 2098 -307
rect 2150 -341 2166 -307
rect 2200 -341 2216 -307
rect 2268 -341 2284 -307
rect 2318 -341 2334 -307
rect 2386 -341 2402 -307
rect 2436 -341 2452 -307
rect 2504 -341 2520 -307
rect 2554 -341 2570 -307
rect 2622 -341 2638 -307
rect 2672 -341 2688 -307
rect 2740 -341 2756 -307
rect 2790 -341 2806 -307
rect 2858 -341 2874 -307
rect 2908 -341 2924 -307
rect 2976 -341 2992 -307
rect 3026 -341 3042 -307
rect 3094 -341 3110 -307
rect 3144 -341 3160 -307
rect 3212 -341 3228 -307
rect 3262 -341 3278 -307
rect 3330 -341 3346 -307
rect 3380 -341 3396 -307
rect 3448 -341 3464 -307
rect 3498 -341 3514 -307
rect 3566 -341 3582 -307
rect 3616 -341 3632 -307
rect 3684 -341 3700 -307
rect 3734 -341 3750 -307
rect 3802 -341 3818 -307
rect 3852 -341 3868 -307
rect 3920 -341 3936 -307
rect 3970 -341 3986 -307
rect 4038 -341 4054 -307
rect 4088 -341 4104 -307
rect 4156 -341 4172 -307
rect 4206 -341 4222 -307
rect 4274 -341 4290 -307
rect 4324 -341 4340 -307
rect 4392 -341 4408 -307
rect 4442 -341 4458 -307
rect 4510 -341 4526 -307
rect 4560 -341 4576 -307
rect 4628 -341 4644 -307
rect 4678 -341 4694 -307
rect 4746 -341 4762 -307
rect 4796 -341 4812 -307
rect 4864 -341 4880 -307
rect 4914 -341 4930 -307
rect 4982 -341 4998 -307
rect 5032 -341 5048 -307
rect 5100 -341 5116 -307
rect 5150 -341 5166 -307
rect 5218 -341 5234 -307
rect 5268 -341 5284 -307
rect 5336 -341 5352 -307
rect 5386 -341 5402 -307
rect 5454 -341 5470 -307
rect 5504 -341 5520 -307
rect 5572 -341 5588 -307
rect 5622 -341 5638 -307
rect 5690 -341 5706 -307
rect 5740 -341 5756 -307
rect 5808 -341 5824 -307
rect 5858 -341 5874 -307
<< viali >>
rect -5917 -257 -5883 319
rect -5799 -257 -5765 319
rect -5681 -257 -5647 319
rect -5563 -257 -5529 319
rect -5445 -257 -5411 319
rect -5327 -257 -5293 319
rect -5209 -257 -5175 319
rect -5091 -257 -5057 319
rect -4973 -257 -4939 319
rect -4855 -257 -4821 319
rect -4737 -257 -4703 319
rect -4619 -257 -4585 319
rect -4501 -257 -4467 319
rect -4383 -257 -4349 319
rect -4265 -257 -4231 319
rect -4147 -257 -4113 319
rect -4029 -257 -3995 319
rect -3911 -257 -3877 319
rect -3793 -257 -3759 319
rect -3675 -257 -3641 319
rect -3557 -257 -3523 319
rect -3439 -257 -3405 319
rect -3321 -257 -3287 319
rect -3203 -257 -3169 319
rect -3085 -257 -3051 319
rect -2967 -257 -2933 319
rect -2849 -257 -2815 319
rect -2731 -257 -2697 319
rect -2613 -257 -2579 319
rect -2495 -257 -2461 319
rect -2377 -257 -2343 319
rect -2259 -257 -2225 319
rect -2141 -257 -2107 319
rect -2023 -257 -1989 319
rect -1905 -257 -1871 319
rect -1787 -257 -1753 319
rect -1669 -257 -1635 319
rect -1551 -257 -1517 319
rect -1433 -257 -1399 319
rect -1315 -257 -1281 319
rect -1197 -257 -1163 319
rect -1079 -257 -1045 319
rect -961 -257 -927 319
rect -843 -257 -809 319
rect -725 -257 -691 319
rect -607 -257 -573 319
rect -489 -257 -455 319
rect -371 -257 -337 319
rect -253 -257 -219 319
rect -135 -257 -101 319
rect -17 -257 17 319
rect 101 -257 135 319
rect 219 -257 253 319
rect 337 -257 371 319
rect 455 -257 489 319
rect 573 -257 607 319
rect 691 -257 725 319
rect 809 -257 843 319
rect 927 -257 961 319
rect 1045 -257 1079 319
rect 1163 -257 1197 319
rect 1281 -257 1315 319
rect 1399 -257 1433 319
rect 1517 -257 1551 319
rect 1635 -257 1669 319
rect 1753 -257 1787 319
rect 1871 -257 1905 319
rect 1989 -257 2023 319
rect 2107 -257 2141 319
rect 2225 -257 2259 319
rect 2343 -257 2377 319
rect 2461 -257 2495 319
rect 2579 -257 2613 319
rect 2697 -257 2731 319
rect 2815 -257 2849 319
rect 2933 -257 2967 319
rect 3051 -257 3085 319
rect 3169 -257 3203 319
rect 3287 -257 3321 319
rect 3405 -257 3439 319
rect 3523 -257 3557 319
rect 3641 -257 3675 319
rect 3759 -257 3793 319
rect 3877 -257 3911 319
rect 3995 -257 4029 319
rect 4113 -257 4147 319
rect 4231 -257 4265 319
rect 4349 -257 4383 319
rect 4467 -257 4501 319
rect 4585 -257 4619 319
rect 4703 -257 4737 319
rect 4821 -257 4855 319
rect 4939 -257 4973 319
rect 5057 -257 5091 319
rect 5175 -257 5209 319
rect 5293 -257 5327 319
rect 5411 -257 5445 319
rect 5529 -257 5563 319
rect 5647 -257 5681 319
rect 5765 -257 5799 319
rect 5883 -257 5917 319
rect -5858 -341 -5824 -307
rect -5740 -341 -5706 -307
rect -5622 -341 -5588 -307
rect -5504 -341 -5470 -307
rect -5386 -341 -5352 -307
rect -5268 -341 -5234 -307
rect -5150 -341 -5116 -307
rect -5032 -341 -4998 -307
rect -4914 -341 -4880 -307
rect -4796 -341 -4762 -307
rect -4678 -341 -4644 -307
rect -4560 -341 -4526 -307
rect -4442 -341 -4408 -307
rect -4324 -341 -4290 -307
rect -4206 -341 -4172 -307
rect -4088 -341 -4054 -307
rect -3970 -341 -3936 -307
rect -3852 -341 -3818 -307
rect -3734 -341 -3700 -307
rect -3616 -341 -3582 -307
rect -3498 -341 -3464 -307
rect -3380 -341 -3346 -307
rect -3262 -341 -3228 -307
rect -3144 -341 -3110 -307
rect -3026 -341 -2992 -307
rect -2908 -341 -2874 -307
rect -2790 -341 -2756 -307
rect -2672 -341 -2638 -307
rect -2554 -341 -2520 -307
rect -2436 -341 -2402 -307
rect -2318 -341 -2284 -307
rect -2200 -341 -2166 -307
rect -2082 -341 -2048 -307
rect -1964 -341 -1930 -307
rect -1846 -341 -1812 -307
rect -1728 -341 -1694 -307
rect -1610 -341 -1576 -307
rect -1492 -341 -1458 -307
rect -1374 -341 -1340 -307
rect -1256 -341 -1222 -307
rect -1138 -341 -1104 -307
rect -1020 -341 -986 -307
rect -902 -341 -868 -307
rect -784 -341 -750 -307
rect -666 -341 -632 -307
rect -548 -341 -514 -307
rect -430 -341 -396 -307
rect -312 -341 -278 -307
rect -194 -341 -160 -307
rect -76 -341 -42 -307
rect 42 -341 76 -307
rect 160 -341 194 -307
rect 278 -341 312 -307
rect 396 -341 430 -307
rect 514 -341 548 -307
rect 632 -341 666 -307
rect 750 -341 784 -307
rect 868 -341 902 -307
rect 986 -341 1020 -307
rect 1104 -341 1138 -307
rect 1222 -341 1256 -307
rect 1340 -341 1374 -307
rect 1458 -341 1492 -307
rect 1576 -341 1610 -307
rect 1694 -341 1728 -307
rect 1812 -341 1846 -307
rect 1930 -341 1964 -307
rect 2048 -341 2082 -307
rect 2166 -341 2200 -307
rect 2284 -341 2318 -307
rect 2402 -341 2436 -307
rect 2520 -341 2554 -307
rect 2638 -341 2672 -307
rect 2756 -341 2790 -307
rect 2874 -341 2908 -307
rect 2992 -341 3026 -307
rect 3110 -341 3144 -307
rect 3228 -341 3262 -307
rect 3346 -341 3380 -307
rect 3464 -341 3498 -307
rect 3582 -341 3616 -307
rect 3700 -341 3734 -307
rect 3818 -341 3852 -307
rect 3936 -341 3970 -307
rect 4054 -341 4088 -307
rect 4172 -341 4206 -307
rect 4290 -341 4324 -307
rect 4408 -341 4442 -307
rect 4526 -341 4560 -307
rect 4644 -341 4678 -307
rect 4762 -341 4796 -307
rect 4880 -341 4914 -307
rect 4998 -341 5032 -307
rect 5116 -341 5150 -307
rect 5234 -341 5268 -307
rect 5352 -341 5386 -307
rect 5470 -341 5504 -307
rect 5588 -341 5622 -307
rect 5706 -341 5740 -307
rect 5824 -341 5858 -307
<< metal1 >>
rect -5923 319 -5877 331
rect -5923 -257 -5917 319
rect -5883 -257 -5877 319
rect -5923 -269 -5877 -257
rect -5805 319 -5759 331
rect -5805 -257 -5799 319
rect -5765 -257 -5759 319
rect -5805 -269 -5759 -257
rect -5687 319 -5641 331
rect -5687 -257 -5681 319
rect -5647 -257 -5641 319
rect -5687 -269 -5641 -257
rect -5569 319 -5523 331
rect -5569 -257 -5563 319
rect -5529 -257 -5523 319
rect -5569 -269 -5523 -257
rect -5451 319 -5405 331
rect -5451 -257 -5445 319
rect -5411 -257 -5405 319
rect -5451 -269 -5405 -257
rect -5333 319 -5287 331
rect -5333 -257 -5327 319
rect -5293 -257 -5287 319
rect -5333 -269 -5287 -257
rect -5215 319 -5169 331
rect -5215 -257 -5209 319
rect -5175 -257 -5169 319
rect -5215 -269 -5169 -257
rect -5097 319 -5051 331
rect -5097 -257 -5091 319
rect -5057 -257 -5051 319
rect -5097 -269 -5051 -257
rect -4979 319 -4933 331
rect -4979 -257 -4973 319
rect -4939 -257 -4933 319
rect -4979 -269 -4933 -257
rect -4861 319 -4815 331
rect -4861 -257 -4855 319
rect -4821 -257 -4815 319
rect -4861 -269 -4815 -257
rect -4743 319 -4697 331
rect -4743 -257 -4737 319
rect -4703 -257 -4697 319
rect -4743 -269 -4697 -257
rect -4625 319 -4579 331
rect -4625 -257 -4619 319
rect -4585 -257 -4579 319
rect -4625 -269 -4579 -257
rect -4507 319 -4461 331
rect -4507 -257 -4501 319
rect -4467 -257 -4461 319
rect -4507 -269 -4461 -257
rect -4389 319 -4343 331
rect -4389 -257 -4383 319
rect -4349 -257 -4343 319
rect -4389 -269 -4343 -257
rect -4271 319 -4225 331
rect -4271 -257 -4265 319
rect -4231 -257 -4225 319
rect -4271 -269 -4225 -257
rect -4153 319 -4107 331
rect -4153 -257 -4147 319
rect -4113 -257 -4107 319
rect -4153 -269 -4107 -257
rect -4035 319 -3989 331
rect -4035 -257 -4029 319
rect -3995 -257 -3989 319
rect -4035 -269 -3989 -257
rect -3917 319 -3871 331
rect -3917 -257 -3911 319
rect -3877 -257 -3871 319
rect -3917 -269 -3871 -257
rect -3799 319 -3753 331
rect -3799 -257 -3793 319
rect -3759 -257 -3753 319
rect -3799 -269 -3753 -257
rect -3681 319 -3635 331
rect -3681 -257 -3675 319
rect -3641 -257 -3635 319
rect -3681 -269 -3635 -257
rect -3563 319 -3517 331
rect -3563 -257 -3557 319
rect -3523 -257 -3517 319
rect -3563 -269 -3517 -257
rect -3445 319 -3399 331
rect -3445 -257 -3439 319
rect -3405 -257 -3399 319
rect -3445 -269 -3399 -257
rect -3327 319 -3281 331
rect -3327 -257 -3321 319
rect -3287 -257 -3281 319
rect -3327 -269 -3281 -257
rect -3209 319 -3163 331
rect -3209 -257 -3203 319
rect -3169 -257 -3163 319
rect -3209 -269 -3163 -257
rect -3091 319 -3045 331
rect -3091 -257 -3085 319
rect -3051 -257 -3045 319
rect -3091 -269 -3045 -257
rect -2973 319 -2927 331
rect -2973 -257 -2967 319
rect -2933 -257 -2927 319
rect -2973 -269 -2927 -257
rect -2855 319 -2809 331
rect -2855 -257 -2849 319
rect -2815 -257 -2809 319
rect -2855 -269 -2809 -257
rect -2737 319 -2691 331
rect -2737 -257 -2731 319
rect -2697 -257 -2691 319
rect -2737 -269 -2691 -257
rect -2619 319 -2573 331
rect -2619 -257 -2613 319
rect -2579 -257 -2573 319
rect -2619 -269 -2573 -257
rect -2501 319 -2455 331
rect -2501 -257 -2495 319
rect -2461 -257 -2455 319
rect -2501 -269 -2455 -257
rect -2383 319 -2337 331
rect -2383 -257 -2377 319
rect -2343 -257 -2337 319
rect -2383 -269 -2337 -257
rect -2265 319 -2219 331
rect -2265 -257 -2259 319
rect -2225 -257 -2219 319
rect -2265 -269 -2219 -257
rect -2147 319 -2101 331
rect -2147 -257 -2141 319
rect -2107 -257 -2101 319
rect -2147 -269 -2101 -257
rect -2029 319 -1983 331
rect -2029 -257 -2023 319
rect -1989 -257 -1983 319
rect -2029 -269 -1983 -257
rect -1911 319 -1865 331
rect -1911 -257 -1905 319
rect -1871 -257 -1865 319
rect -1911 -269 -1865 -257
rect -1793 319 -1747 331
rect -1793 -257 -1787 319
rect -1753 -257 -1747 319
rect -1793 -269 -1747 -257
rect -1675 319 -1629 331
rect -1675 -257 -1669 319
rect -1635 -257 -1629 319
rect -1675 -269 -1629 -257
rect -1557 319 -1511 331
rect -1557 -257 -1551 319
rect -1517 -257 -1511 319
rect -1557 -269 -1511 -257
rect -1439 319 -1393 331
rect -1439 -257 -1433 319
rect -1399 -257 -1393 319
rect -1439 -269 -1393 -257
rect -1321 319 -1275 331
rect -1321 -257 -1315 319
rect -1281 -257 -1275 319
rect -1321 -269 -1275 -257
rect -1203 319 -1157 331
rect -1203 -257 -1197 319
rect -1163 -257 -1157 319
rect -1203 -269 -1157 -257
rect -1085 319 -1039 331
rect -1085 -257 -1079 319
rect -1045 -257 -1039 319
rect -1085 -269 -1039 -257
rect -967 319 -921 331
rect -967 -257 -961 319
rect -927 -257 -921 319
rect -967 -269 -921 -257
rect -849 319 -803 331
rect -849 -257 -843 319
rect -809 -257 -803 319
rect -849 -269 -803 -257
rect -731 319 -685 331
rect -731 -257 -725 319
rect -691 -257 -685 319
rect -731 -269 -685 -257
rect -613 319 -567 331
rect -613 -257 -607 319
rect -573 -257 -567 319
rect -613 -269 -567 -257
rect -495 319 -449 331
rect -495 -257 -489 319
rect -455 -257 -449 319
rect -495 -269 -449 -257
rect -377 319 -331 331
rect -377 -257 -371 319
rect -337 -257 -331 319
rect -377 -269 -331 -257
rect -259 319 -213 331
rect -259 -257 -253 319
rect -219 -257 -213 319
rect -259 -269 -213 -257
rect -141 319 -95 331
rect -141 -257 -135 319
rect -101 -257 -95 319
rect -141 -269 -95 -257
rect -23 319 23 331
rect -23 -257 -17 319
rect 17 -257 23 319
rect -23 -269 23 -257
rect 95 319 141 331
rect 95 -257 101 319
rect 135 -257 141 319
rect 95 -269 141 -257
rect 213 319 259 331
rect 213 -257 219 319
rect 253 -257 259 319
rect 213 -269 259 -257
rect 331 319 377 331
rect 331 -257 337 319
rect 371 -257 377 319
rect 331 -269 377 -257
rect 449 319 495 331
rect 449 -257 455 319
rect 489 -257 495 319
rect 449 -269 495 -257
rect 567 319 613 331
rect 567 -257 573 319
rect 607 -257 613 319
rect 567 -269 613 -257
rect 685 319 731 331
rect 685 -257 691 319
rect 725 -257 731 319
rect 685 -269 731 -257
rect 803 319 849 331
rect 803 -257 809 319
rect 843 -257 849 319
rect 803 -269 849 -257
rect 921 319 967 331
rect 921 -257 927 319
rect 961 -257 967 319
rect 921 -269 967 -257
rect 1039 319 1085 331
rect 1039 -257 1045 319
rect 1079 -257 1085 319
rect 1039 -269 1085 -257
rect 1157 319 1203 331
rect 1157 -257 1163 319
rect 1197 -257 1203 319
rect 1157 -269 1203 -257
rect 1275 319 1321 331
rect 1275 -257 1281 319
rect 1315 -257 1321 319
rect 1275 -269 1321 -257
rect 1393 319 1439 331
rect 1393 -257 1399 319
rect 1433 -257 1439 319
rect 1393 -269 1439 -257
rect 1511 319 1557 331
rect 1511 -257 1517 319
rect 1551 -257 1557 319
rect 1511 -269 1557 -257
rect 1629 319 1675 331
rect 1629 -257 1635 319
rect 1669 -257 1675 319
rect 1629 -269 1675 -257
rect 1747 319 1793 331
rect 1747 -257 1753 319
rect 1787 -257 1793 319
rect 1747 -269 1793 -257
rect 1865 319 1911 331
rect 1865 -257 1871 319
rect 1905 -257 1911 319
rect 1865 -269 1911 -257
rect 1983 319 2029 331
rect 1983 -257 1989 319
rect 2023 -257 2029 319
rect 1983 -269 2029 -257
rect 2101 319 2147 331
rect 2101 -257 2107 319
rect 2141 -257 2147 319
rect 2101 -269 2147 -257
rect 2219 319 2265 331
rect 2219 -257 2225 319
rect 2259 -257 2265 319
rect 2219 -269 2265 -257
rect 2337 319 2383 331
rect 2337 -257 2343 319
rect 2377 -257 2383 319
rect 2337 -269 2383 -257
rect 2455 319 2501 331
rect 2455 -257 2461 319
rect 2495 -257 2501 319
rect 2455 -269 2501 -257
rect 2573 319 2619 331
rect 2573 -257 2579 319
rect 2613 -257 2619 319
rect 2573 -269 2619 -257
rect 2691 319 2737 331
rect 2691 -257 2697 319
rect 2731 -257 2737 319
rect 2691 -269 2737 -257
rect 2809 319 2855 331
rect 2809 -257 2815 319
rect 2849 -257 2855 319
rect 2809 -269 2855 -257
rect 2927 319 2973 331
rect 2927 -257 2933 319
rect 2967 -257 2973 319
rect 2927 -269 2973 -257
rect 3045 319 3091 331
rect 3045 -257 3051 319
rect 3085 -257 3091 319
rect 3045 -269 3091 -257
rect 3163 319 3209 331
rect 3163 -257 3169 319
rect 3203 -257 3209 319
rect 3163 -269 3209 -257
rect 3281 319 3327 331
rect 3281 -257 3287 319
rect 3321 -257 3327 319
rect 3281 -269 3327 -257
rect 3399 319 3445 331
rect 3399 -257 3405 319
rect 3439 -257 3445 319
rect 3399 -269 3445 -257
rect 3517 319 3563 331
rect 3517 -257 3523 319
rect 3557 -257 3563 319
rect 3517 -269 3563 -257
rect 3635 319 3681 331
rect 3635 -257 3641 319
rect 3675 -257 3681 319
rect 3635 -269 3681 -257
rect 3753 319 3799 331
rect 3753 -257 3759 319
rect 3793 -257 3799 319
rect 3753 -269 3799 -257
rect 3871 319 3917 331
rect 3871 -257 3877 319
rect 3911 -257 3917 319
rect 3871 -269 3917 -257
rect 3989 319 4035 331
rect 3989 -257 3995 319
rect 4029 -257 4035 319
rect 3989 -269 4035 -257
rect 4107 319 4153 331
rect 4107 -257 4113 319
rect 4147 -257 4153 319
rect 4107 -269 4153 -257
rect 4225 319 4271 331
rect 4225 -257 4231 319
rect 4265 -257 4271 319
rect 4225 -269 4271 -257
rect 4343 319 4389 331
rect 4343 -257 4349 319
rect 4383 -257 4389 319
rect 4343 -269 4389 -257
rect 4461 319 4507 331
rect 4461 -257 4467 319
rect 4501 -257 4507 319
rect 4461 -269 4507 -257
rect 4579 319 4625 331
rect 4579 -257 4585 319
rect 4619 -257 4625 319
rect 4579 -269 4625 -257
rect 4697 319 4743 331
rect 4697 -257 4703 319
rect 4737 -257 4743 319
rect 4697 -269 4743 -257
rect 4815 319 4861 331
rect 4815 -257 4821 319
rect 4855 -257 4861 319
rect 4815 -269 4861 -257
rect 4933 319 4979 331
rect 4933 -257 4939 319
rect 4973 -257 4979 319
rect 4933 -269 4979 -257
rect 5051 319 5097 331
rect 5051 -257 5057 319
rect 5091 -257 5097 319
rect 5051 -269 5097 -257
rect 5169 319 5215 331
rect 5169 -257 5175 319
rect 5209 -257 5215 319
rect 5169 -269 5215 -257
rect 5287 319 5333 331
rect 5287 -257 5293 319
rect 5327 -257 5333 319
rect 5287 -269 5333 -257
rect 5405 319 5451 331
rect 5405 -257 5411 319
rect 5445 -257 5451 319
rect 5405 -269 5451 -257
rect 5523 319 5569 331
rect 5523 -257 5529 319
rect 5563 -257 5569 319
rect 5523 -269 5569 -257
rect 5641 319 5687 331
rect 5641 -257 5647 319
rect 5681 -257 5687 319
rect 5641 -269 5687 -257
rect 5759 319 5805 331
rect 5759 -257 5765 319
rect 5799 -257 5805 319
rect 5759 -269 5805 -257
rect 5877 319 5923 331
rect 5877 -257 5883 319
rect 5917 -257 5923 319
rect 5877 -269 5923 -257
rect -5870 -307 -5812 -301
rect -5870 -341 -5858 -307
rect -5824 -341 -5812 -307
rect -5870 -347 -5812 -341
rect -5752 -307 -5694 -301
rect -5752 -341 -5740 -307
rect -5706 -341 -5694 -307
rect -5752 -347 -5694 -341
rect -5634 -307 -5576 -301
rect -5634 -341 -5622 -307
rect -5588 -341 -5576 -307
rect -5634 -347 -5576 -341
rect -5516 -307 -5458 -301
rect -5516 -341 -5504 -307
rect -5470 -341 -5458 -307
rect -5516 -347 -5458 -341
rect -5398 -307 -5340 -301
rect -5398 -341 -5386 -307
rect -5352 -341 -5340 -307
rect -5398 -347 -5340 -341
rect -5280 -307 -5222 -301
rect -5280 -341 -5268 -307
rect -5234 -341 -5222 -307
rect -5280 -347 -5222 -341
rect -5162 -307 -5104 -301
rect -5162 -341 -5150 -307
rect -5116 -341 -5104 -307
rect -5162 -347 -5104 -341
rect -5044 -307 -4986 -301
rect -5044 -341 -5032 -307
rect -4998 -341 -4986 -307
rect -5044 -347 -4986 -341
rect -4926 -307 -4868 -301
rect -4926 -341 -4914 -307
rect -4880 -341 -4868 -307
rect -4926 -347 -4868 -341
rect -4808 -307 -4750 -301
rect -4808 -341 -4796 -307
rect -4762 -341 -4750 -307
rect -4808 -347 -4750 -341
rect -4690 -307 -4632 -301
rect -4690 -341 -4678 -307
rect -4644 -341 -4632 -307
rect -4690 -347 -4632 -341
rect -4572 -307 -4514 -301
rect -4572 -341 -4560 -307
rect -4526 -341 -4514 -307
rect -4572 -347 -4514 -341
rect -4454 -307 -4396 -301
rect -4454 -341 -4442 -307
rect -4408 -341 -4396 -307
rect -4454 -347 -4396 -341
rect -4336 -307 -4278 -301
rect -4336 -341 -4324 -307
rect -4290 -341 -4278 -307
rect -4336 -347 -4278 -341
rect -4218 -307 -4160 -301
rect -4218 -341 -4206 -307
rect -4172 -341 -4160 -307
rect -4218 -347 -4160 -341
rect -4100 -307 -4042 -301
rect -4100 -341 -4088 -307
rect -4054 -341 -4042 -307
rect -4100 -347 -4042 -341
rect -3982 -307 -3924 -301
rect -3982 -341 -3970 -307
rect -3936 -341 -3924 -307
rect -3982 -347 -3924 -341
rect -3864 -307 -3806 -301
rect -3864 -341 -3852 -307
rect -3818 -341 -3806 -307
rect -3864 -347 -3806 -341
rect -3746 -307 -3688 -301
rect -3746 -341 -3734 -307
rect -3700 -341 -3688 -307
rect -3746 -347 -3688 -341
rect -3628 -307 -3570 -301
rect -3628 -341 -3616 -307
rect -3582 -341 -3570 -307
rect -3628 -347 -3570 -341
rect -3510 -307 -3452 -301
rect -3510 -341 -3498 -307
rect -3464 -341 -3452 -307
rect -3510 -347 -3452 -341
rect -3392 -307 -3334 -301
rect -3392 -341 -3380 -307
rect -3346 -341 -3334 -307
rect -3392 -347 -3334 -341
rect -3274 -307 -3216 -301
rect -3274 -341 -3262 -307
rect -3228 -341 -3216 -307
rect -3274 -347 -3216 -341
rect -3156 -307 -3098 -301
rect -3156 -341 -3144 -307
rect -3110 -341 -3098 -307
rect -3156 -347 -3098 -341
rect -3038 -307 -2980 -301
rect -3038 -341 -3026 -307
rect -2992 -341 -2980 -307
rect -3038 -347 -2980 -341
rect -2920 -307 -2862 -301
rect -2920 -341 -2908 -307
rect -2874 -341 -2862 -307
rect -2920 -347 -2862 -341
rect -2802 -307 -2744 -301
rect -2802 -341 -2790 -307
rect -2756 -341 -2744 -307
rect -2802 -347 -2744 -341
rect -2684 -307 -2626 -301
rect -2684 -341 -2672 -307
rect -2638 -341 -2626 -307
rect -2684 -347 -2626 -341
rect -2566 -307 -2508 -301
rect -2566 -341 -2554 -307
rect -2520 -341 -2508 -307
rect -2566 -347 -2508 -341
rect -2448 -307 -2390 -301
rect -2448 -341 -2436 -307
rect -2402 -341 -2390 -307
rect -2448 -347 -2390 -341
rect -2330 -307 -2272 -301
rect -2330 -341 -2318 -307
rect -2284 -341 -2272 -307
rect -2330 -347 -2272 -341
rect -2212 -307 -2154 -301
rect -2212 -341 -2200 -307
rect -2166 -341 -2154 -307
rect -2212 -347 -2154 -341
rect -2094 -307 -2036 -301
rect -2094 -341 -2082 -307
rect -2048 -341 -2036 -307
rect -2094 -347 -2036 -341
rect -1976 -307 -1918 -301
rect -1976 -341 -1964 -307
rect -1930 -341 -1918 -307
rect -1976 -347 -1918 -341
rect -1858 -307 -1800 -301
rect -1858 -341 -1846 -307
rect -1812 -341 -1800 -307
rect -1858 -347 -1800 -341
rect -1740 -307 -1682 -301
rect -1740 -341 -1728 -307
rect -1694 -341 -1682 -307
rect -1740 -347 -1682 -341
rect -1622 -307 -1564 -301
rect -1622 -341 -1610 -307
rect -1576 -341 -1564 -307
rect -1622 -347 -1564 -341
rect -1504 -307 -1446 -301
rect -1504 -341 -1492 -307
rect -1458 -341 -1446 -307
rect -1504 -347 -1446 -341
rect -1386 -307 -1328 -301
rect -1386 -341 -1374 -307
rect -1340 -341 -1328 -307
rect -1386 -347 -1328 -341
rect -1268 -307 -1210 -301
rect -1268 -341 -1256 -307
rect -1222 -341 -1210 -307
rect -1268 -347 -1210 -341
rect -1150 -307 -1092 -301
rect -1150 -341 -1138 -307
rect -1104 -341 -1092 -307
rect -1150 -347 -1092 -341
rect -1032 -307 -974 -301
rect -1032 -341 -1020 -307
rect -986 -341 -974 -307
rect -1032 -347 -974 -341
rect -914 -307 -856 -301
rect -914 -341 -902 -307
rect -868 -341 -856 -307
rect -914 -347 -856 -341
rect -796 -307 -738 -301
rect -796 -341 -784 -307
rect -750 -341 -738 -307
rect -796 -347 -738 -341
rect -678 -307 -620 -301
rect -678 -341 -666 -307
rect -632 -341 -620 -307
rect -678 -347 -620 -341
rect -560 -307 -502 -301
rect -560 -341 -548 -307
rect -514 -341 -502 -307
rect -560 -347 -502 -341
rect -442 -307 -384 -301
rect -442 -341 -430 -307
rect -396 -341 -384 -307
rect -442 -347 -384 -341
rect -324 -307 -266 -301
rect -324 -341 -312 -307
rect -278 -341 -266 -307
rect -324 -347 -266 -341
rect -206 -307 -148 -301
rect -206 -341 -194 -307
rect -160 -341 -148 -307
rect -206 -347 -148 -341
rect -88 -307 -30 -301
rect -88 -341 -76 -307
rect -42 -341 -30 -307
rect -88 -347 -30 -341
rect 30 -307 88 -301
rect 30 -341 42 -307
rect 76 -341 88 -307
rect 30 -347 88 -341
rect 148 -307 206 -301
rect 148 -341 160 -307
rect 194 -341 206 -307
rect 148 -347 206 -341
rect 266 -307 324 -301
rect 266 -341 278 -307
rect 312 -341 324 -307
rect 266 -347 324 -341
rect 384 -307 442 -301
rect 384 -341 396 -307
rect 430 -341 442 -307
rect 384 -347 442 -341
rect 502 -307 560 -301
rect 502 -341 514 -307
rect 548 -341 560 -307
rect 502 -347 560 -341
rect 620 -307 678 -301
rect 620 -341 632 -307
rect 666 -341 678 -307
rect 620 -347 678 -341
rect 738 -307 796 -301
rect 738 -341 750 -307
rect 784 -341 796 -307
rect 738 -347 796 -341
rect 856 -307 914 -301
rect 856 -341 868 -307
rect 902 -341 914 -307
rect 856 -347 914 -341
rect 974 -307 1032 -301
rect 974 -341 986 -307
rect 1020 -341 1032 -307
rect 974 -347 1032 -341
rect 1092 -307 1150 -301
rect 1092 -341 1104 -307
rect 1138 -341 1150 -307
rect 1092 -347 1150 -341
rect 1210 -307 1268 -301
rect 1210 -341 1222 -307
rect 1256 -341 1268 -307
rect 1210 -347 1268 -341
rect 1328 -307 1386 -301
rect 1328 -341 1340 -307
rect 1374 -341 1386 -307
rect 1328 -347 1386 -341
rect 1446 -307 1504 -301
rect 1446 -341 1458 -307
rect 1492 -341 1504 -307
rect 1446 -347 1504 -341
rect 1564 -307 1622 -301
rect 1564 -341 1576 -307
rect 1610 -341 1622 -307
rect 1564 -347 1622 -341
rect 1682 -307 1740 -301
rect 1682 -341 1694 -307
rect 1728 -341 1740 -307
rect 1682 -347 1740 -341
rect 1800 -307 1858 -301
rect 1800 -341 1812 -307
rect 1846 -341 1858 -307
rect 1800 -347 1858 -341
rect 1918 -307 1976 -301
rect 1918 -341 1930 -307
rect 1964 -341 1976 -307
rect 1918 -347 1976 -341
rect 2036 -307 2094 -301
rect 2036 -341 2048 -307
rect 2082 -341 2094 -307
rect 2036 -347 2094 -341
rect 2154 -307 2212 -301
rect 2154 -341 2166 -307
rect 2200 -341 2212 -307
rect 2154 -347 2212 -341
rect 2272 -307 2330 -301
rect 2272 -341 2284 -307
rect 2318 -341 2330 -307
rect 2272 -347 2330 -341
rect 2390 -307 2448 -301
rect 2390 -341 2402 -307
rect 2436 -341 2448 -307
rect 2390 -347 2448 -341
rect 2508 -307 2566 -301
rect 2508 -341 2520 -307
rect 2554 -341 2566 -307
rect 2508 -347 2566 -341
rect 2626 -307 2684 -301
rect 2626 -341 2638 -307
rect 2672 -341 2684 -307
rect 2626 -347 2684 -341
rect 2744 -307 2802 -301
rect 2744 -341 2756 -307
rect 2790 -341 2802 -307
rect 2744 -347 2802 -341
rect 2862 -307 2920 -301
rect 2862 -341 2874 -307
rect 2908 -341 2920 -307
rect 2862 -347 2920 -341
rect 2980 -307 3038 -301
rect 2980 -341 2992 -307
rect 3026 -341 3038 -307
rect 2980 -347 3038 -341
rect 3098 -307 3156 -301
rect 3098 -341 3110 -307
rect 3144 -341 3156 -307
rect 3098 -347 3156 -341
rect 3216 -307 3274 -301
rect 3216 -341 3228 -307
rect 3262 -341 3274 -307
rect 3216 -347 3274 -341
rect 3334 -307 3392 -301
rect 3334 -341 3346 -307
rect 3380 -341 3392 -307
rect 3334 -347 3392 -341
rect 3452 -307 3510 -301
rect 3452 -341 3464 -307
rect 3498 -341 3510 -307
rect 3452 -347 3510 -341
rect 3570 -307 3628 -301
rect 3570 -341 3582 -307
rect 3616 -341 3628 -307
rect 3570 -347 3628 -341
rect 3688 -307 3746 -301
rect 3688 -341 3700 -307
rect 3734 -341 3746 -307
rect 3688 -347 3746 -341
rect 3806 -307 3864 -301
rect 3806 -341 3818 -307
rect 3852 -341 3864 -307
rect 3806 -347 3864 -341
rect 3924 -307 3982 -301
rect 3924 -341 3936 -307
rect 3970 -341 3982 -307
rect 3924 -347 3982 -341
rect 4042 -307 4100 -301
rect 4042 -341 4054 -307
rect 4088 -341 4100 -307
rect 4042 -347 4100 -341
rect 4160 -307 4218 -301
rect 4160 -341 4172 -307
rect 4206 -341 4218 -307
rect 4160 -347 4218 -341
rect 4278 -307 4336 -301
rect 4278 -341 4290 -307
rect 4324 -341 4336 -307
rect 4278 -347 4336 -341
rect 4396 -307 4454 -301
rect 4396 -341 4408 -307
rect 4442 -341 4454 -307
rect 4396 -347 4454 -341
rect 4514 -307 4572 -301
rect 4514 -341 4526 -307
rect 4560 -341 4572 -307
rect 4514 -347 4572 -341
rect 4632 -307 4690 -301
rect 4632 -341 4644 -307
rect 4678 -341 4690 -307
rect 4632 -347 4690 -341
rect 4750 -307 4808 -301
rect 4750 -341 4762 -307
rect 4796 -341 4808 -307
rect 4750 -347 4808 -341
rect 4868 -307 4926 -301
rect 4868 -341 4880 -307
rect 4914 -341 4926 -307
rect 4868 -347 4926 -341
rect 4986 -307 5044 -301
rect 4986 -341 4998 -307
rect 5032 -341 5044 -307
rect 4986 -347 5044 -341
rect 5104 -307 5162 -301
rect 5104 -341 5116 -307
rect 5150 -341 5162 -307
rect 5104 -347 5162 -341
rect 5222 -307 5280 -301
rect 5222 -341 5234 -307
rect 5268 -341 5280 -307
rect 5222 -347 5280 -341
rect 5340 -307 5398 -301
rect 5340 -341 5352 -307
rect 5386 -341 5398 -307
rect 5340 -347 5398 -341
rect 5458 -307 5516 -301
rect 5458 -341 5470 -307
rect 5504 -341 5516 -307
rect 5458 -347 5516 -341
rect 5576 -307 5634 -301
rect 5576 -341 5588 -307
rect 5622 -341 5634 -307
rect 5576 -347 5634 -341
rect 5694 -307 5752 -301
rect 5694 -341 5706 -307
rect 5740 -341 5752 -307
rect 5694 -347 5752 -341
rect 5812 -307 5870 -301
rect 5812 -341 5824 -307
rect 5858 -341 5870 -307
rect 5812 -347 5870 -341
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 3 l 0.3 m 1 nf 100 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
