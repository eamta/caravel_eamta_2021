magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 79 1084 237 1143
rect 17 1083 299 1084
rect 17 1049 299 1050
rect 141 981 175 1015
rect -17 617 17 627
rect 299 617 333 627
rect -17 609 333 617
rect -53 547 369 609
rect 109 257 129 265
<< nwell >>
rect -53 1083 369 1179
<< pwell >>
rect -53 112 355 124
rect -53 16 369 112
<< psubdiff >>
rect 55 53 79 87
rect 237 53 261 87
<< nsubdiff >>
rect 55 1109 79 1143
rect 237 1109 261 1143
<< psubdiffcont >>
rect 79 53 237 87
<< nsubdiffcont >>
rect 79 1109 237 1143
<< viali >>
rect -20 1143 336 1146
rect -20 1109 79 1143
rect 79 1109 237 1143
rect 237 1109 336 1143
rect -20 1106 336 1109
rect -20 1010 336 1050
rect -20 138 336 178
rect -20 87 336 90
rect -20 53 79 87
rect 79 53 237 87
rect 237 53 336 87
rect -20 50 336 53
<< metal1 >>
rect -53 1146 369 1152
rect -53 1106 -20 1146
rect 336 1106 369 1146
rect -53 1050 369 1106
rect -53 1010 -20 1050
rect 336 1010 369 1050
rect -53 1004 369 1010
rect 91 918 137 1004
rect 179 922 285 939
rect 125 573 191 729
rect 119 521 129 573
rect 181 521 191 573
rect 125 366 191 521
rect 219 573 285 922
rect 219 521 229 573
rect 281 521 291 573
rect 219 337 285 521
rect 91 200 137 257
rect 179 249 285 337
rect 0 184 200 200
rect -53 178 369 184
rect -53 138 -20 178
rect 336 138 369 178
rect -53 90 369 138
rect -53 50 -20 90
rect 336 50 369 90
rect -53 44 369 50
rect 0 0 200 44
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
<< via1 >>
rect 129 521 181 573
rect 229 521 281 573
<< metal2 >>
rect 129 573 181 583
rect -53 521 129 573
rect 129 511 181 521
rect 229 573 281 583
rect 281 521 369 573
rect 229 511 281 521
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 1624053917
transform 1 0 158 0 1 357
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_MQX2PY  XM2
timestamp 1624053917
transform 1 0 158 0 1 850
box -211 -303 211 303
<< labels >>
rlabel metal2 281 521 369 573 1 out
port 2 n
rlabel metal2 -53 521 129 573 1 in
port 3 n
rlabel metal1 -53 90 369 138 1 vss
port 4 n
rlabel metal1 -53 1050 369 1106 1 vdd
port 1 n
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 in
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vss
<< end >>
