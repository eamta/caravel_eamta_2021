magic
tech sky130A
magscale 1 2
timestamp 1624067212
<< nwell >>
rect -107 1050 1084 1271
rect 1090 1272 2550 1351
rect 3799 1272 5354 1352
rect 1090 1050 5354 1272
rect -107 767 5354 1050
rect -107 366 1147 767
rect 1090 339 1147 366
rect 1148 367 5354 767
rect 1148 339 2550 367
rect 3805 340 5354 367
rect 1090 -327 2550 -248
rect 3800 -327 5354 -247
rect 1090 -328 5354 -327
rect -107 -803 5354 -328
rect -107 -804 3800 -803
rect 3806 -804 5354 -803
rect -107 -1232 5354 -804
rect -107 -1233 2550 -1232
rect 1090 -1260 2550 -1233
rect 3806 -1259 5354 -1232
<< pwell >>
rect 1084 1698 5353 1735
rect -107 1666 5353 1698
rect -107 1624 3277 1666
rect 3580 1624 5353 1666
rect -107 1352 5353 1624
rect -107 1351 3799 1352
rect -107 1271 1084 1351
rect 2550 1272 3799 1351
rect -107 339 1084 366
rect 2550 340 3800 367
rect 2550 339 5354 340
rect -107 259 5354 339
rect -107 256 2684 259
rect 3509 256 5354 259
rect -107 167 5354 256
rect -107 164 1905 167
rect 1957 164 5354 167
rect -107 -247 5354 164
rect -107 -248 3800 -247
rect -107 -328 1084 -248
rect 2550 -327 3800 -248
rect -107 -1260 1090 -1233
rect 2550 -1259 3806 -1232
rect 2550 -1260 5353 -1259
rect -107 -1605 5353 -1260
<< psubdiff >>
rect 319 1628 343 1663
rect 1201 1628 1225 1663
rect 1827 1626 1851 1661
rect 1976 1626 2000 1661
rect 2397 1629 2421 1664
rect 2558 1629 2582 1664
rect 3043 1629 3067 1664
rect 3923 1629 3947 1664
rect 4565 1629 4589 1663
rect 4672 1629 4696 1663
rect 5115 1630 5139 1664
rect 5321 1630 5345 1664
rect 557 29 581 63
rect 900 29 924 63
rect 3139 30 3163 64
rect 3253 30 3277 64
rect 3644 30 3668 64
rect 36 -1570 60 -1536
rect 292 -1570 316 -1536
rect 552 -1571 576 -1536
rect 1397 -1571 1421 -1536
rect 2405 -1571 2429 -1535
rect 2981 -1571 3005 -1535
rect 3268 -1570 3292 -1536
rect 3605 -1570 3629 -1536
rect 3741 -1570 3765 -1536
rect 3877 -1570 3901 -1536
<< nsubdiff >>
rect 564 826 603 860
rect 690 826 724 860
<< psubdiffcont >>
rect 343 1628 1201 1663
rect 1851 1626 1976 1661
rect 2421 1629 2558 1664
rect 3067 1629 3923 1664
rect 4589 1629 4672 1663
rect 5139 1630 5321 1664
rect 581 29 900 63
rect 3277 30 3644 64
rect 60 -1570 292 -1536
rect 576 -1571 1397 -1536
rect 2429 -1571 2981 -1535
rect 3292 -1570 3605 -1536
rect 3765 -1570 3877 -1536
<< nsubdiffcont >>
rect 603 826 690 860
<< poly >>
rect 1118 808 1148 1311
rect 640 381 706 397
rect 640 347 656 381
rect 690 366 706 381
rect 690 347 1006 366
rect 640 336 1006 347
rect 640 331 676 336
rect 976 -80 1006 336
rect 1118 339 1147 808
rect 3356 382 3422 398
rect 3356 348 3372 382
rect 3406 367 3422 382
rect 3406 348 3722 367
rect 1118 -294 1148 339
rect 3356 337 3722 348
rect 3356 332 3392 337
rect 3692 -21 3722 337
rect 3833 323 3863 325
rect 3833 307 3899 323
rect 3833 273 3849 307
rect 3883 273 3899 307
rect 3833 257 3899 273
rect 3833 -240 3863 257
<< polycont >>
rect 656 347 690 381
rect 3372 348 3406 382
rect 3849 273 3883 307
<< locali >>
rect 640 381 706 397
rect 640 347 656 381
rect 690 347 706 381
rect 640 331 706 347
rect 3356 382 3422 398
rect 3356 348 3372 382
rect 3406 348 3422 382
rect 3356 332 3422 348
rect 3833 307 3899 323
rect 3833 273 3849 307
rect 3883 273 3899 307
rect 3833 257 3899 273
<< viali >>
rect 319 1628 343 1663
rect 343 1628 1201 1663
rect 1201 1628 1225 1663
rect 1827 1626 1851 1661
rect 1851 1626 1976 1661
rect 1976 1626 2000 1661
rect 2397 1629 2421 1664
rect 2421 1629 2558 1664
rect 2558 1629 2582 1664
rect 3043 1629 3067 1664
rect 3067 1629 3923 1664
rect 3923 1629 3947 1664
rect 4565 1629 4589 1663
rect 4589 1629 4672 1663
rect 4672 1629 4696 1663
rect 5115 1630 5139 1664
rect 5139 1630 5321 1664
rect 5321 1630 5345 1664
rect 564 826 603 860
rect 603 826 690 860
rect 690 826 724 860
rect 656 347 690 381
rect 3372 348 3406 382
rect 3849 273 3883 307
rect 557 29 581 63
rect 581 29 900 63
rect 900 29 924 63
rect 3253 30 3277 64
rect 3277 30 3644 64
rect 3644 30 3668 64
rect 36 -1570 60 -1536
rect 60 -1570 292 -1536
rect 292 -1570 316 -1536
rect 552 -1571 576 -1536
rect 576 -1571 1397 -1536
rect 1397 -1571 1421 -1536
rect 2405 -1571 2429 -1535
rect 2429 -1571 2981 -1535
rect 2981 -1571 3005 -1535
rect 3268 -1570 3292 -1536
rect 3292 -1570 3605 -1536
rect 3605 -1570 3629 -1536
rect 3741 -1570 3765 -1536
rect 3765 -1570 3877 -1536
rect 3877 -1570 3901 -1536
<< metal1 >>
rect 307 1668 1237 1669
rect 53 1667 2011 1668
rect 53 1663 2012 1667
rect 53 1662 319 1663
rect 53 1628 65 1662
rect 307 1628 319 1662
rect 1225 1662 2012 1663
rect 1225 1628 1237 1662
rect 1815 1661 2012 1662
rect 1815 1628 1827 1661
rect 53 1626 1827 1628
rect 2000 1626 2012 1661
rect 53 1622 2012 1626
rect 2385 1664 2594 1670
rect 3031 1669 3959 1670
rect 2385 1629 2397 1664
rect 2582 1629 2594 1664
rect 2385 1623 2594 1629
rect 1815 1620 2012 1622
rect 2599 1617 2609 1669
rect 2661 1664 3959 1669
rect 2661 1663 3043 1664
rect 2661 1629 2742 1663
rect 2768 1629 2780 1663
rect 3031 1629 3043 1663
rect 3947 1629 3959 1664
rect 2661 1623 3959 1629
rect 3969 1664 5357 1670
rect 3969 1630 3981 1664
rect 4553 1663 4708 1664
rect 4553 1630 4565 1663
rect 3969 1629 4565 1630
rect 4696 1630 4708 1663
rect 5103 1630 5115 1664
rect 5345 1630 5357 1664
rect 4696 1629 5357 1630
rect 3969 1624 5357 1629
rect 4553 1623 4708 1624
rect 2661 1622 2768 1623
rect 2661 1617 2671 1622
rect 2551 1403 2556 1437
rect 5270 1404 5271 1438
rect -62 816 -52 868
rect 0 816 10 868
rect 480 866 665 868
rect 480 862 736 866
rect 480 826 492 862
rect 552 860 736 862
rect 552 826 564 860
rect 724 826 736 860
rect 480 820 736 826
rect 2546 821 2723 869
rect 3190 863 3377 869
rect 3190 827 3202 863
rect 3365 827 3377 863
rect 3190 821 3377 827
rect 4456 863 4582 869
rect 4456 829 4468 863
rect 4570 829 4582 863
rect 4456 823 4582 829
rect 4949 824 4959 869
rect 604 381 706 397
rect 565 367 571 373
rect 604 367 656 381
rect 565 365 656 367
rect 640 347 656 365
rect 690 347 706 381
rect 3320 382 3422 398
rect 3320 367 3372 382
rect 640 331 706 347
rect 2431 323 2718 358
rect 3356 348 3372 367
rect 3406 348 3422 382
rect 3356 332 3422 348
rect 2674 318 2718 323
rect 1918 157 1952 306
rect 2674 266 2684 318
rect 2736 266 2746 318
rect 3833 307 3899 323
rect 3833 304 3849 307
rect 3353 273 3849 304
rect 3883 273 3899 307
rect 3353 270 3899 273
rect 3353 221 3387 270
rect 3833 257 3899 270
rect 2685 169 2695 221
rect 2747 169 2757 221
rect 3332 169 3342 221
rect 3394 169 3404 221
rect 3447 186 3457 238
rect 3509 220 3519 238
rect 3699 220 3709 233
rect 3509 186 3709 220
rect 3699 181 3709 186
rect 3761 181 3771 233
rect 2685 164 2747 169
rect 2525 163 2747 164
rect 1895 105 1905 157
rect 1957 105 1967 157
rect 2525 111 2535 163
rect 2587 130 2747 163
rect 2587 111 2597 130
rect 11 63 1088 69
rect 11 29 23 63
rect 489 29 501 63
rect 545 29 557 63
rect 924 29 936 63
rect 1076 29 1088 63
rect 11 23 1088 29
rect 1190 63 2486 69
rect 1190 29 1202 63
rect 2474 29 2486 63
rect 1190 23 2486 29
rect 2599 18 2609 74
rect 2661 70 2671 74
rect 2661 64 3813 70
rect 2661 30 2747 64
rect 3127 30 3139 64
rect 3241 30 3253 64
rect 3668 30 3680 64
rect 3801 30 3813 64
rect 2661 24 3813 30
rect 4089 64 5253 70
rect 4089 30 4101 64
rect 5241 30 5253 64
rect 4089 24 5253 30
rect 2661 18 2671 24
rect 2555 -196 2556 -162
rect 5271 -195 5272 -161
rect -62 -780 -52 -728
rect 0 -780 10 -728
rect 494 -737 633 -731
rect 494 -773 506 -737
rect 621 -773 633 -737
rect 494 -779 633 -773
rect 2549 -778 2731 -730
rect 3219 -736 3342 -730
rect 3219 -772 3231 -736
rect 3330 -772 3342 -736
rect 3219 -778 3342 -772
rect 2819 -1100 2829 -1091
rect 2684 -1134 2829 -1100
rect 2684 -1242 2718 -1134
rect 2819 -1143 2829 -1134
rect 2881 -1143 2891 -1091
rect 3323 -1232 3324 -1201
rect 2411 -1276 2718 -1242
rect 557 -1486 567 -1434
rect 619 -1486 629 -1434
rect 2590 -1466 2600 -1414
rect 2652 -1466 2662 -1414
rect 2599 -1529 2652 -1466
rect 2661 -1529 2671 -1525
rect 2393 -1530 3017 -1529
rect 18 -1535 5302 -1530
rect 18 -1536 2405 -1535
rect 18 -1570 36 -1536
rect 316 -1570 328 -1536
rect 540 -1570 552 -1536
rect 18 -1571 552 -1570
rect 1421 -1570 1433 -1536
rect 2393 -1570 2405 -1536
rect 1421 -1571 2405 -1570
rect 3005 -1536 5302 -1535
rect 3005 -1570 3017 -1536
rect 3256 -1570 3268 -1536
rect 3629 -1570 3641 -1536
rect 3729 -1570 3741 -1536
rect 3901 -1570 3913 -1536
rect 4144 -1570 4156 -1536
rect 5162 -1570 5174 -1536
rect 5290 -1570 5302 -1536
rect 3005 -1571 5302 -1570
rect 18 -1576 5302 -1571
rect 540 -1577 1433 -1576
rect 2393 -1577 3017 -1576
<< via1 >>
rect 2609 1617 2661 1669
rect -52 816 0 868
rect 2684 266 2736 318
rect 2695 169 2747 221
rect 3342 169 3394 221
rect 3457 186 3509 238
rect 3709 181 3761 233
rect 1905 105 1957 157
rect 2535 111 2587 163
rect 2609 18 2661 74
rect -52 -780 0 -728
rect 2829 -1143 2881 -1091
rect 567 -1486 619 -1434
rect 2600 -1466 2652 -1414
<< metal2 >>
rect 2609 1669 2661 1679
rect 2609 1611 2661 1617
rect 2615 1607 2661 1611
rect 33 1207 35 1259
rect -52 868 0 878
rect -52 806 0 816
rect -52 -718 -18 806
rect 382 464 387 516
rect 1905 157 1957 164
rect 2535 163 2587 173
rect 1957 111 2535 129
rect 1957 105 2587 111
rect 1905 101 2587 105
rect 1905 95 2572 101
rect 1905 90 1957 95
rect 2615 84 2649 1607
rect 5179 1298 5180 1350
rect 2684 318 2736 328
rect 2736 266 3509 293
rect 2684 259 3509 266
rect 3457 238 3509 259
rect 2695 221 2747 231
rect 3342 221 3394 231
rect 2747 176 3342 210
rect 2695 159 2747 169
rect 3457 176 3509 186
rect 3342 159 3394 169
rect 3544 131 3579 532
rect 3709 233 3761 243
rect 3761 193 3839 227
rect 5315 204 5349 208
rect 3709 171 3761 181
rect 5146 168 5349 204
rect 2689 97 3579 131
rect 2615 74 2661 84
rect 2600 18 2609 74
rect 2600 8 2661 18
rect 34 -392 35 -340
rect -52 -728 0 -718
rect -52 -790 0 -780
rect 2600 -1404 2634 8
rect 2600 -1414 2652 -1404
rect 567 -1434 619 -1424
rect 2600 -1476 2652 -1466
rect 567 -1496 619 -1486
rect 588 -1514 619 -1496
rect 2689 -1514 2723 97
rect 5180 -301 5181 -249
rect 2829 -1091 2881 -1081
rect 2881 -1143 2949 -1109
rect 2829 -1153 2881 -1143
rect 2915 -1372 2949 -1143
rect 5315 -1325 5349 168
rect 2915 -1406 3895 -1372
rect 5315 -1402 5350 -1325
rect 5138 -1436 5350 -1402
rect 588 -1548 2723 -1514
use bitc  bitc_0
timestamp 1624067212
transform 1 0 1083 0 1 10
box -1084 -8 1577 1677
use bitc  bitc_2
timestamp 1624067212
transform 1 0 1084 0 1 -1589
box -1084 -8 1577 1677
use bitc  bitc_3
timestamp 1624067212
transform 1 0 3800 0 1 -1588
box -1084 -8 1577 1677
use bitc  bitc_1
timestamp 1624067212
transform 1 0 3799 0 1 11
box -1084 -8 1577 1677
<< labels >>
rlabel metal2 384 464 387 516 1 CE
rlabel metal2 33 1207 35 1259 1 Q0
rlabel metal2 34 -392 35 -340 1 Q1
rlabel metal2 5179 1298 5180 1350 1 Q2
rlabel metal2 5180 -301 5181 -249 1 Q3
rlabel metal1 2555 1403 2556 1437 1 Q0n
rlabel metal1 2555 -196 2556 -162 1 Q1n
rlabel metal1 5270 1404 5271 1438 1 Q2n
rlabel metal1 5271 -195 5272 -161 1 Q3n
rlabel metal1 3323 -1232 3324 -1201 1 Sout3
rlabel metal2 2600 -1414 2634 18 1 vss!
rlabel pwell 3741 -1570 3901 -1536 1 vss!
rlabel nwell 603 826 690 860 1 vdd!
rlabel metal1 1106 1288 1183 1359 1 CLK
rlabel metal1 2411 -1276 2718 -1242 1 CLR
<< end >>
