magic
tech sky130A
magscale 1 2
timestamp 1624129585
use sky130_fd_pr__cap_mim_m3_2_2Y8F6P  decap
array 0 4 -6944 0 0 -991
timestamp 1624129585
transform -1 0 3373 0 -1 3102
box -3351 -3261 3373 3261
<< end >>
