magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect 129 919 187 925
rect 129 885 141 919
rect 129 879 187 885
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1042
rect 498 974 556 980
rect 498 940 510 974
rect 668 951 702 969
rect 1090 951 1125 969
rect 498 934 556 940
rect 668 915 738 951
rect 1054 936 1125 951
rect 685 881 756 915
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 881
rect 867 813 925 819
rect 867 779 879 813
rect 867 773 925 779
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1054 477 1124 936
rect 1236 868 1294 874
rect 1236 834 1248 868
rect 1406 845 1440 863
rect 1828 845 1863 863
rect 1236 828 1294 834
rect 1406 809 1476 845
rect 1792 830 1863 845
rect 1423 775 1494 809
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1423 424 1493 775
rect 1605 707 1663 713
rect 1605 673 1617 707
rect 1605 667 1663 673
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1792 371 1862 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 2144 739 2178 757
rect 2566 739 2601 757
rect 1974 722 2032 728
rect 2144 703 2214 739
rect 2530 724 2601 739
rect 2881 724 2916 758
rect 2161 669 2232 703
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2161 318 2231 669
rect 2343 601 2401 607
rect 2343 567 2355 601
rect 2343 561 2401 567
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2161 282 2214 318
rect 2530 265 2600 724
rect 2882 705 2916 724
rect 2712 656 2770 662
rect 2712 622 2724 656
rect 2712 616 2770 622
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
rect 2901 212 2916 705
rect 2935 671 2970 705
rect 2935 212 2969 671
rect 4726 639 4761 673
rect 4727 620 4761 639
rect 3081 603 3139 609
rect 3081 569 3093 603
rect 3251 580 3285 598
rect 3673 580 3708 598
rect 3081 563 3139 569
rect 3251 544 3321 580
rect 3637 565 3708 580
rect 4557 571 4615 577
rect 3268 510 3339 544
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3268 159 3338 510
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3268 123 3321 159
rect 3637 106 3707 565
rect 4557 537 4569 571
rect 4557 531 4615 537
rect 3819 497 3877 503
rect 3819 463 3831 497
rect 3989 474 4023 492
rect 4411 474 4445 492
rect 3819 457 3877 463
rect 3989 438 4059 474
rect 4006 404 4077 438
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3637 70 3690 106
rect 4006 53 4076 404
rect 4188 336 4246 342
rect 4188 302 4200 336
rect 4188 296 4246 302
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4006 17 4059 53
rect 4375 0 4445 474
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4375 -36 4428 0
rect 4746 -53 4761 620
rect 4780 586 4815 620
rect 4780 -53 4814 586
rect 4926 518 4984 524
rect 4926 484 4938 518
rect 4926 478 4984 484
rect 6202 427 6237 461
rect 6203 408 6237 427
rect 6033 359 6091 365
rect 5096 315 5130 333
rect 6033 325 6045 359
rect 6033 319 6091 325
rect 5096 279 5166 315
rect 5113 245 5184 279
rect 5464 245 5499 279
rect 5887 262 5921 280
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5113 -106 5183 245
rect 5465 226 5499 245
rect 5295 177 5353 183
rect 5295 143 5307 177
rect 5295 137 5353 143
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5113 -142 5166 -106
rect 5484 -159 5499 226
rect 5518 192 5553 226
rect 5518 -159 5552 192
rect 5664 124 5722 130
rect 5664 90 5676 124
rect 5664 84 5722 90
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5518 -193 5533 -159
rect 5851 -212 5921 262
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5851 -248 5904 -212
rect 6222 -265 6237 408
rect 6256 374 6291 408
rect 6256 -265 6290 374
rect 6402 306 6460 312
rect 6402 272 6414 306
rect 6402 266 6460 272
rect 6572 103 6606 121
rect 6572 67 6642 103
rect 6589 33 6660 67
rect 6940 33 6975 67
rect 7363 50 7398 68
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6256 -299 6271 -265
rect 6589 -318 6659 33
rect 6941 14 6975 33
rect 7327 35 7398 50
rect 6771 -35 6829 -29
rect 6771 -69 6783 -35
rect 6771 -75 6829 -69
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6589 -354 6642 -318
rect 6960 -371 6975 14
rect 6994 -20 7029 14
rect 6994 -371 7028 -20
rect 7140 -88 7198 -82
rect 7140 -122 7152 -88
rect 7140 -128 7198 -122
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6994 -405 7009 -371
rect 7327 -424 7397 35
rect 7509 -33 7567 -27
rect 7509 -67 7521 -33
rect 7679 -56 7713 -38
rect 8101 -56 8136 -38
rect 7509 -73 7567 -67
rect 7679 -92 7749 -56
rect 8065 -71 8136 -56
rect 7696 -126 7767 -92
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7327 -460 7380 -424
rect 7696 -477 7766 -126
rect 7878 -194 7936 -188
rect 7878 -228 7890 -194
rect 7878 -234 7936 -228
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7696 -513 7749 -477
rect 8065 -530 8135 -71
rect 8247 -139 8305 -133
rect 8247 -173 8259 -139
rect 8417 -162 8451 -144
rect 8247 -179 8305 -173
rect 8417 -198 8487 -162
rect 8434 -232 8505 -198
rect 8247 -447 8305 -441
rect 8247 -481 8259 -447
rect 8247 -487 8305 -481
rect 8065 -566 8118 -530
rect 8434 -583 8504 -232
rect 8616 -300 8674 -294
rect 8616 -334 8628 -300
rect 8616 -340 8674 -334
rect 8616 -500 8674 -494
rect 8616 -534 8628 -500
rect 8616 -540 8674 -534
rect 8434 -619 8487 -583
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__nfet_01v8_HVW3BE  XM6
timestamp 1624053917
transform 1 0 2372 0 1 484
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM7
timestamp 1624053917
transform 1 0 2741 0 1 485
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM8
timestamp 1624053917
transform 1 0 3110 0 1 432
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM10
timestamp 1624053917
transform 1 0 3848 0 1 326
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM15
timestamp 1624053917
transform 1 0 5324 0 1 60
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM14
timestamp 1624053917
transform 1 0 4955 0 1 257
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM13
timestamp 1624053917
transform 1 0 4586 0 1 310
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM11
timestamp 1624053917
transform 1 0 4217 0 1 219
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM19
timestamp 1624053917
transform 1 0 6800 0 1 -152
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM18
timestamp 1624053917
transform 1 0 6431 0 1 45
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM17
timestamp 1624053917
transform 1 0 6062 0 1 98
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM16
timestamp 1624053917
transform 1 0 5693 0 1 7
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM24
timestamp 1624053917
transform 1 0 8645 0 1 -417
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM23
timestamp 1624053917
transform 1 0 8276 0 1 -310
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM22
timestamp 1624053917
transform 1 0 7907 0 1 -311
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM21
timestamp 1624053917
transform 1 0 7538 0 1 -204
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM20
timestamp 1624053917
transform 1 0 7169 0 1 -205
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM1
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM12
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM2
timestamp 1624053917
transform 1 0 896 0 1 696
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM3
timestamp 1624053917
transform 1 0 1265 0 1 697
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1624053917
transform 1 0 1634 0 1 590
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 D
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLK
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLR
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 vss
port 6 nsew
<< end >>
