magic
tech sky130A
timestamp 1616176710
<< pwell >>
rect -1288 -630 1288 630
<< nmos >>
rect -1190 -525 -1000 525
rect -971 -525 -781 525
rect -752 -525 -562 525
rect -533 -525 -343 525
rect -314 -525 -124 525
rect -95 -525 95 525
rect 124 -525 314 525
rect 343 -525 533 525
rect 562 -525 752 525
rect 781 -525 971 525
rect 1000 -525 1190 525
<< ndiff >>
rect -1219 519 -1190 525
rect -1219 -519 -1213 519
rect -1196 -519 -1190 519
rect -1219 -525 -1190 -519
rect -1000 519 -971 525
rect -1000 -519 -994 519
rect -977 -519 -971 519
rect -1000 -525 -971 -519
rect -781 519 -752 525
rect -781 -519 -775 519
rect -758 -519 -752 519
rect -781 -525 -752 -519
rect -562 519 -533 525
rect -562 -519 -556 519
rect -539 -519 -533 519
rect -562 -525 -533 -519
rect -343 519 -314 525
rect -343 -519 -337 519
rect -320 -519 -314 519
rect -343 -525 -314 -519
rect -124 519 -95 525
rect -124 -519 -118 519
rect -101 -519 -95 519
rect -124 -525 -95 -519
rect 95 519 124 525
rect 95 -519 101 519
rect 118 -519 124 519
rect 95 -525 124 -519
rect 314 519 343 525
rect 314 -519 320 519
rect 337 -519 343 519
rect 314 -525 343 -519
rect 533 519 562 525
rect 533 -519 539 519
rect 556 -519 562 519
rect 533 -525 562 -519
rect 752 519 781 525
rect 752 -519 758 519
rect 775 -519 781 519
rect 752 -525 781 -519
rect 971 519 1000 525
rect 971 -519 977 519
rect 994 -519 1000 519
rect 971 -525 1000 -519
rect 1190 519 1219 525
rect 1190 -519 1196 519
rect 1213 -519 1219 519
rect 1190 -525 1219 -519
<< ndiffc >>
rect -1213 -519 -1196 519
rect -994 -519 -977 519
rect -775 -519 -758 519
rect -556 -519 -539 519
rect -337 -519 -320 519
rect -118 -519 -101 519
rect 101 -519 118 519
rect 320 -519 337 519
rect 539 -519 556 519
rect 758 -519 775 519
rect 977 -519 994 519
rect 1196 -519 1213 519
<< psubdiff >>
rect -1270 595 -1222 612
rect 1222 595 1270 612
rect -1270 564 -1253 595
rect 1253 564 1270 595
rect -1270 -595 -1253 -564
rect 1253 -595 1270 -564
rect -1270 -612 -1222 -595
rect 1222 -612 1270 -595
<< psubdiffcont >>
rect -1222 595 1222 612
rect -1270 -564 -1253 564
rect 1253 -564 1270 564
rect -1222 -612 1222 -595
<< poly >>
rect -1190 561 -1000 569
rect -1190 544 -1182 561
rect -1008 544 -1000 561
rect -1190 525 -1000 544
rect -971 561 -781 569
rect -971 544 -963 561
rect -789 544 -781 561
rect -971 525 -781 544
rect -752 561 -562 569
rect -752 544 -744 561
rect -570 544 -562 561
rect -752 525 -562 544
rect -533 561 -343 569
rect -533 544 -525 561
rect -351 544 -343 561
rect -533 525 -343 544
rect -314 561 -124 569
rect -314 544 -306 561
rect -132 544 -124 561
rect -314 525 -124 544
rect -95 561 95 569
rect -95 544 -87 561
rect 87 544 95 561
rect -95 525 95 544
rect 124 561 314 569
rect 124 544 132 561
rect 306 544 314 561
rect 124 525 314 544
rect 343 561 533 569
rect 343 544 351 561
rect 525 544 533 561
rect 343 525 533 544
rect 562 561 752 569
rect 562 544 570 561
rect 744 544 752 561
rect 562 525 752 544
rect 781 561 971 569
rect 781 544 789 561
rect 963 544 971 561
rect 781 525 971 544
rect 1000 561 1190 569
rect 1000 544 1008 561
rect 1182 544 1190 561
rect 1000 525 1190 544
rect -1190 -544 -1000 -525
rect -1190 -561 -1182 -544
rect -1008 -561 -1000 -544
rect -1190 -569 -1000 -561
rect -971 -544 -781 -525
rect -971 -561 -963 -544
rect -789 -561 -781 -544
rect -971 -569 -781 -561
rect -752 -544 -562 -525
rect -752 -561 -744 -544
rect -570 -561 -562 -544
rect -752 -569 -562 -561
rect -533 -544 -343 -525
rect -533 -561 -525 -544
rect -351 -561 -343 -544
rect -533 -569 -343 -561
rect -314 -544 -124 -525
rect -314 -561 -306 -544
rect -132 -561 -124 -544
rect -314 -569 -124 -561
rect -95 -544 95 -525
rect -95 -561 -87 -544
rect 87 -561 95 -544
rect -95 -569 95 -561
rect 124 -544 314 -525
rect 124 -561 132 -544
rect 306 -561 314 -544
rect 124 -569 314 -561
rect 343 -544 533 -525
rect 343 -561 351 -544
rect 525 -561 533 -544
rect 343 -569 533 -561
rect 562 -544 752 -525
rect 562 -561 570 -544
rect 744 -561 752 -544
rect 562 -569 752 -561
rect 781 -544 971 -525
rect 781 -561 789 -544
rect 963 -561 971 -544
rect 781 -569 971 -561
rect 1000 -544 1190 -525
rect 1000 -561 1008 -544
rect 1182 -561 1190 -544
rect 1000 -569 1190 -561
<< polycont >>
rect -1182 544 -1008 561
rect -963 544 -789 561
rect -744 544 -570 561
rect -525 544 -351 561
rect -306 544 -132 561
rect -87 544 87 561
rect 132 544 306 561
rect 351 544 525 561
rect 570 544 744 561
rect 789 544 963 561
rect 1008 544 1182 561
rect -1182 -561 -1008 -544
rect -963 -561 -789 -544
rect -744 -561 -570 -544
rect -525 -561 -351 -544
rect -306 -561 -132 -544
rect -87 -561 87 -544
rect 132 -561 306 -544
rect 351 -561 525 -544
rect 570 -561 744 -544
rect 789 -561 963 -544
rect 1008 -561 1182 -544
<< locali >>
rect -1270 595 -1222 612
rect 1222 595 1270 612
rect -1270 564 -1253 595
rect 1253 564 1270 595
rect -1190 544 -1182 561
rect -1008 544 -1000 561
rect -971 544 -963 561
rect -789 544 -781 561
rect -752 544 -744 561
rect -570 544 -562 561
rect -533 544 -525 561
rect -351 544 -343 561
rect -314 544 -306 561
rect -132 544 -124 561
rect -95 544 -87 561
rect 87 544 95 561
rect 124 544 132 561
rect 306 544 314 561
rect 343 544 351 561
rect 525 544 533 561
rect 562 544 570 561
rect 744 544 752 561
rect 781 544 789 561
rect 963 544 971 561
rect 1000 544 1008 561
rect 1182 544 1190 561
rect -1213 519 -1196 527
rect -1213 -527 -1196 -519
rect -994 519 -977 527
rect -994 -527 -977 -519
rect -775 519 -758 527
rect -775 -527 -758 -519
rect -556 519 -539 527
rect -556 -527 -539 -519
rect -337 519 -320 527
rect -337 -527 -320 -519
rect -118 519 -101 527
rect -118 -527 -101 -519
rect 101 519 118 527
rect 101 -527 118 -519
rect 320 519 337 527
rect 320 -527 337 -519
rect 539 519 556 527
rect 539 -527 556 -519
rect 758 519 775 527
rect 758 -527 775 -519
rect 977 519 994 527
rect 977 -527 994 -519
rect 1196 519 1213 527
rect 1196 -527 1213 -519
rect -1190 -561 -1182 -544
rect -1008 -561 -1000 -544
rect -971 -561 -963 -544
rect -789 -561 -781 -544
rect -752 -561 -744 -544
rect -570 -561 -562 -544
rect -533 -561 -525 -544
rect -351 -561 -343 -544
rect -314 -561 -306 -544
rect -132 -561 -124 -544
rect -95 -561 -87 -544
rect 87 -561 95 -544
rect 124 -561 132 -544
rect 306 -561 314 -544
rect 343 -561 351 -544
rect 525 -561 533 -544
rect 562 -561 570 -544
rect 744 -561 752 -544
rect 781 -561 789 -544
rect 963 -561 971 -544
rect 1000 -561 1008 -544
rect 1182 -561 1190 -544
rect -1270 -595 -1253 -564
rect 1253 -595 1270 -564
rect -1270 -612 -1222 -595
rect 1222 -612 1270 -595
<< viali >>
rect -1182 544 -1008 561
rect -963 544 -789 561
rect -744 544 -570 561
rect -525 544 -351 561
rect -306 544 -132 561
rect -87 544 87 561
rect 132 544 306 561
rect 351 544 525 561
rect 570 544 744 561
rect 789 544 963 561
rect 1008 544 1182 561
rect -1213 -519 -1196 519
rect -994 -519 -977 519
rect -775 -519 -758 519
rect -556 -519 -539 519
rect -337 -519 -320 519
rect -118 -519 -101 519
rect 101 -519 118 519
rect 320 -519 337 519
rect 539 -519 556 519
rect 758 -519 775 519
rect 977 -519 994 519
rect 1196 -519 1213 519
rect -1182 -561 -1008 -544
rect -963 -561 -789 -544
rect -744 -561 -570 -544
rect -525 -561 -351 -544
rect -306 -561 -132 -544
rect -87 -561 87 -544
rect 132 -561 306 -544
rect 351 -561 525 -544
rect 570 -561 744 -544
rect 789 -561 963 -544
rect 1008 -561 1182 -544
<< metal1 >>
rect -1188 561 -1002 564
rect -1188 544 -1182 561
rect -1008 544 -1002 561
rect -1188 541 -1002 544
rect -969 561 -783 564
rect -969 544 -963 561
rect -789 544 -783 561
rect -969 541 -783 544
rect -750 561 -564 564
rect -750 544 -744 561
rect -570 544 -564 561
rect -750 541 -564 544
rect -531 561 -345 564
rect -531 544 -525 561
rect -351 544 -345 561
rect -531 541 -345 544
rect -312 561 -126 564
rect -312 544 -306 561
rect -132 544 -126 561
rect -312 541 -126 544
rect -93 561 93 564
rect -93 544 -87 561
rect 87 544 93 561
rect -93 541 93 544
rect 126 561 312 564
rect 126 544 132 561
rect 306 544 312 561
rect 126 541 312 544
rect 345 561 531 564
rect 345 544 351 561
rect 525 544 531 561
rect 345 541 531 544
rect 564 561 750 564
rect 564 544 570 561
rect 744 544 750 561
rect 564 541 750 544
rect 783 561 969 564
rect 783 544 789 561
rect 963 544 969 561
rect 783 541 969 544
rect 1002 561 1188 564
rect 1002 544 1008 561
rect 1182 544 1188 561
rect 1002 541 1188 544
rect -1216 519 -1193 525
rect -1216 -519 -1213 519
rect -1196 -519 -1193 519
rect -1216 -525 -1193 -519
rect -997 519 -974 525
rect -997 -519 -994 519
rect -977 -519 -974 519
rect -997 -525 -974 -519
rect -778 519 -755 525
rect -778 -519 -775 519
rect -758 -519 -755 519
rect -778 -525 -755 -519
rect -559 519 -536 525
rect -559 -519 -556 519
rect -539 -519 -536 519
rect -559 -525 -536 -519
rect -340 519 -317 525
rect -340 -519 -337 519
rect -320 -519 -317 519
rect -340 -525 -317 -519
rect -121 519 -98 525
rect -121 -519 -118 519
rect -101 -519 -98 519
rect -121 -525 -98 -519
rect 98 519 121 525
rect 98 -519 101 519
rect 118 -519 121 519
rect 98 -525 121 -519
rect 317 519 340 525
rect 317 -519 320 519
rect 337 -519 340 519
rect 317 -525 340 -519
rect 536 519 559 525
rect 536 -519 539 519
rect 556 -519 559 519
rect 536 -525 559 -519
rect 755 519 778 525
rect 755 -519 758 519
rect 775 -519 778 519
rect 755 -525 778 -519
rect 974 519 997 525
rect 974 -519 977 519
rect 994 -519 997 519
rect 974 -525 997 -519
rect 1193 519 1216 525
rect 1193 -519 1196 519
rect 1213 -519 1216 519
rect 1193 -525 1216 -519
rect -1188 -544 -1002 -541
rect -1188 -561 -1182 -544
rect -1008 -561 -1002 -544
rect -1188 -564 -1002 -561
rect -969 -544 -783 -541
rect -969 -561 -963 -544
rect -789 -561 -783 -544
rect -969 -564 -783 -561
rect -750 -544 -564 -541
rect -750 -561 -744 -544
rect -570 -561 -564 -544
rect -750 -564 -564 -561
rect -531 -544 -345 -541
rect -531 -561 -525 -544
rect -351 -561 -345 -544
rect -531 -564 -345 -561
rect -312 -544 -126 -541
rect -312 -561 -306 -544
rect -132 -561 -126 -544
rect -312 -564 -126 -561
rect -93 -544 93 -541
rect -93 -561 -87 -544
rect 87 -561 93 -544
rect -93 -564 93 -561
rect 126 -544 312 -541
rect 126 -561 132 -544
rect 306 -561 312 -544
rect 126 -564 312 -561
rect 345 -544 531 -541
rect 345 -561 351 -544
rect 525 -561 531 -544
rect 345 -564 531 -561
rect 564 -544 750 -541
rect 564 -561 570 -544
rect 744 -561 750 -544
rect 564 -564 750 -561
rect 783 -544 969 -541
rect 783 -561 789 -544
rect 963 -561 969 -544
rect 783 -564 969 -561
rect 1002 -544 1188 -541
rect 1002 -561 1008 -544
rect 1182 -561 1188 -544
rect 1002 -564 1188 -561
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1261 -603 1261 603
string parameters w 10.5 l 1.9 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
