magic
tech sky130A
magscale 1 2
timestamp 1624138001
<< error_p >>
rect 103 650 116 678
rect 150 616 163 650
rect 210 616 231 678
rect 335 650 356 678
rect 599 650 620 678
rect 382 616 403 650
rect 646 616 667 650
rect 670 616 690 650
rect 706 616 727 678
rect 1123 650 1144 678
rect 1188 660 1204 666
rect 1160 650 1214 660
rect 1389 650 1410 678
rect 1454 660 1470 666
rect 1426 650 1480 660
rect 1154 640 1220 650
rect 1154 634 1191 640
rect 1170 616 1191 634
rect 1194 634 1220 640
rect 1420 640 1486 650
rect 1420 634 1457 640
rect 1194 616 1214 634
rect 1436 616 1457 634
rect 1460 634 1486 640
rect 1460 616 1480 634
rect 1496 616 1517 678
rect 1619 650 1642 678
rect 1684 660 1700 666
rect 1656 650 1710 660
rect 1650 640 1716 650
rect 1650 634 1689 640
rect 1666 616 1689 634
rect 1690 634 1716 640
rect 1690 616 1710 634
rect 1728 616 1747 678
rect 1855 650 1874 678
rect 1920 660 1936 666
rect 1892 650 1946 660
rect 1886 640 1952 650
rect 1886 634 1921 640
rect 1902 616 1921 634
rect 1926 634 1952 640
rect 1926 616 1946 634
rect 1960 616 1983 678
rect 219 498 347 519
rect 413 488 414 530
rect 474 498 532 519
rect 1264 498 1322 519
rect 1505 498 1633 519
rect 266 472 268 482
rect 298 472 300 482
rect 266 462 278 472
rect 288 462 300 472
rect 455 472 456 488
rect 1264 482 1280 488
rect 1584 482 1586 488
rect 1236 472 1290 482
rect 1542 472 1554 482
rect 1584 472 1596 482
rect 455 448 465 472
rect 266 438 300 446
rect 455 438 467 448
rect 479 438 499 472
rect 1230 462 1296 472
rect 1230 456 1256 462
rect 1246 438 1256 456
rect 1270 456 1296 462
rect 1536 462 1564 472
rect 1574 462 1602 472
rect 1536 456 1562 462
rect 1270 438 1290 456
rect 1552 448 1562 456
rect 1576 456 1602 462
rect 1576 448 1596 456
rect 1552 438 1596 448
rect 562 404 564 410
rect 520 394 532 404
rect 562 394 574 404
rect 1278 394 1280 436
rect 1570 428 1596 438
rect 1570 422 1586 428
rect 1352 404 1354 410
rect 1570 404 1586 410
rect 1310 394 1322 404
rect 1352 394 1364 404
rect 1542 394 1554 404
rect 1570 396 1596 404
rect 1584 394 1596 396
rect 514 384 542 394
rect 552 384 580 394
rect 514 378 540 384
rect 530 360 540 378
rect 554 378 580 384
rect 1304 384 1332 394
rect 1342 384 1370 394
rect 1304 378 1330 384
rect 554 360 574 378
rect 1320 370 1330 378
rect 1344 378 1370 384
rect 1536 386 1602 394
rect 1536 384 1564 386
rect 1574 384 1602 386
rect 1536 378 1562 384
rect 1344 370 1364 378
rect 1320 360 1364 370
rect 1552 370 1562 378
rect 1576 378 1602 384
rect 1576 370 1596 378
rect 1552 360 1564 370
rect 1574 360 1596 370
rect 530 344 564 354
rect 1338 350 1364 360
rect 1584 350 1596 360
rect 715 318 843 349
rect 1338 344 1354 350
rect 1584 344 1586 350
rect 2057 318 2185 349
rect 794 312 796 318
rect 2136 312 2138 318
rect 752 302 764 312
rect 794 302 806 312
rect 2094 302 2106 312
rect 2136 302 2148 312
rect 746 292 774 302
rect 784 292 812 302
rect 746 286 772 292
rect 762 278 772 286
rect 786 286 812 292
rect 2088 292 2116 302
rect 2126 292 2154 302
rect 2088 286 2114 292
rect 786 278 806 286
rect 762 268 774 278
rect 784 268 806 278
rect 2104 278 2114 286
rect 2128 286 2154 292
rect 2128 278 2148 286
rect 2104 268 2116 278
rect 2126 268 2148 278
rect 794 258 806 268
rect 2136 258 2148 268
rect 794 252 796 258
rect 2136 252 2138 258
rect 1086 244 1088 250
rect 2048 244 2052 250
rect 1044 234 1056 244
rect 1086 234 1098 244
rect 2048 234 2062 244
rect 380 200 390 234
rect 404 200 424 234
rect 1038 224 1066 234
rect 1076 224 1104 234
rect 1038 218 1064 224
rect 1054 210 1064 218
rect 1078 218 1104 224
rect 1078 210 1098 218
rect 1054 200 1066 210
rect 1076 200 1098 210
rect 1436 200 1446 234
rect 1460 200 1480 234
rect 2018 200 2028 234
rect 2038 224 2068 234
rect 2042 218 2068 224
rect 2042 210 2062 218
rect 2038 200 2062 210
rect 1086 190 1098 200
rect 2048 190 2062 200
rect 1086 184 1088 190
rect 2048 184 2052 190
rect 998 176 1014 182
rect 980 166 1024 176
rect 980 156 1030 166
rect 1004 150 1030 156
rect 1004 148 1024 150
rect 980 132 1024 148
rect 1170 148 1180 166
rect 1170 132 1182 148
rect 1194 132 1214 166
rect 998 122 1024 132
rect 998 116 1014 122
rect 112 82 116 110
rect 150 58 160 82
rect 174 58 194 82
rect 150 48 194 58
rect 210 48 222 110
rect 342 82 356 110
rect 608 82 620 110
rect 380 58 394 82
rect 404 58 424 82
rect 380 48 424 58
rect 646 58 658 82
rect 670 58 690 82
rect 646 48 690 58
rect 706 48 718 110
rect 1132 82 1144 110
rect 1398 82 1410 110
rect 1170 58 1182 82
rect 1194 58 1214 82
rect 1170 48 1214 58
rect 1436 58 1448 82
rect 1460 58 1480 82
rect 1436 48 1480 58
rect 1496 48 1508 110
rect 1628 82 1642 110
rect 1666 58 1680 82
rect 1690 58 1710 82
rect 1666 48 1710 58
rect 1728 48 1738 110
rect 1864 82 1874 110
rect 1902 58 1912 82
rect 1926 58 1946 82
rect 1902 48 1946 58
rect 1960 48 1974 110
rect 168 38 194 48
rect 398 38 424 48
rect 664 38 690 48
rect 1188 38 1214 48
rect 1454 38 1480 48
rect 1684 38 1710 48
rect 1920 38 1946 48
rect 168 32 184 38
rect 398 32 414 38
rect 664 32 680 38
rect 1188 32 1204 38
rect 1454 32 1470 38
rect 1684 32 1700 38
rect 1920 32 1936 38
<< nwell >>
rect -66 280 2230 804
<< nmos >>
rect 28 20 58 110
rect 268 20 298 110
rect 532 20 562 110
rect 764 20 794 110
rect 852 20 882 110
rect 1056 20 1086 110
rect 1322 20 1352 110
rect 1554 20 1584 110
rect 1786 20 1816 110
rect 2018 20 2048 110
rect 2106 20 2136 110
<< pmos >>
rect 28 498 58 678
rect 268 498 298 678
rect 532 498 562 678
rect 764 318 794 678
rect 852 318 882 678
rect 1056 498 1086 678
rect 1322 498 1352 678
rect 1554 498 1584 678
rect 1786 498 1816 678
rect 2018 318 2048 678
rect 2106 318 2136 678
<< ndiff >>
rect -30 82 28 110
rect -30 48 -18 82
rect 16 48 28 82
rect -30 20 28 48
rect 58 82 116 110
rect 58 48 70 82
rect 104 48 116 82
rect 210 82 268 110
rect 210 48 222 82
rect 256 48 268 82
rect 58 20 116 48
rect 210 20 268 48
rect 298 82 356 110
rect 298 48 310 82
rect 344 48 356 82
rect 474 82 532 110
rect 474 48 486 82
rect 520 48 532 82
rect 298 20 356 48
rect 474 20 532 48
rect 562 82 620 110
rect 562 48 574 82
rect 608 48 620 82
rect 706 82 764 110
rect 706 48 718 82
rect 752 48 764 82
rect 562 20 620 48
rect 706 20 764 48
rect 794 82 852 110
rect 794 48 806 82
rect 840 48 852 82
rect 794 20 852 48
rect 882 82 940 110
rect 882 48 894 82
rect 928 48 940 82
rect 882 20 940 48
rect 998 82 1056 110
rect 998 48 1010 82
rect 1044 48 1056 82
rect 998 20 1056 48
rect 1086 82 1144 110
rect 1086 48 1098 82
rect 1132 48 1144 82
rect 1264 82 1322 110
rect 1264 48 1276 82
rect 1310 48 1322 82
rect 1086 20 1144 48
rect 1264 20 1322 48
rect 1352 82 1410 110
rect 1352 48 1364 82
rect 1398 48 1410 82
rect 1496 82 1554 110
rect 1496 48 1508 82
rect 1542 48 1554 82
rect 1352 20 1410 48
rect 1496 20 1554 48
rect 1584 82 1642 110
rect 1584 48 1596 82
rect 1630 48 1642 82
rect 1728 82 1786 110
rect 1728 48 1740 82
rect 1774 48 1786 82
rect 1584 20 1642 48
rect 1728 20 1786 48
rect 1816 82 1874 110
rect 1816 48 1828 82
rect 1862 48 1874 82
rect 1960 82 2018 110
rect 1960 48 1972 82
rect 2006 48 2018 82
rect 1816 20 1874 48
rect 1960 20 2018 48
rect 2048 82 2106 110
rect 2048 48 2060 82
rect 2094 48 2106 82
rect 2048 20 2106 48
rect 2136 82 2194 110
rect 2136 48 2148 82
rect 2182 48 2194 82
rect 2136 20 2194 48
<< pdiff >>
rect -30 650 28 678
rect -30 616 -18 650
rect 16 616 28 650
rect -30 498 28 616
rect 58 650 116 678
rect 58 616 70 650
rect 104 616 116 650
rect 58 498 116 616
rect 210 650 268 678
rect 210 616 222 650
rect 256 616 268 650
rect 210 498 268 616
rect 298 650 356 678
rect 298 616 310 650
rect 344 616 356 650
rect 298 498 356 616
rect 474 650 532 678
rect 474 616 486 650
rect 520 616 532 650
rect 474 498 532 616
rect 562 650 620 678
rect 562 616 574 650
rect 608 616 620 650
rect 562 498 620 616
rect 706 650 764 678
rect 706 616 718 650
rect 752 616 764 650
rect 706 318 764 616
rect 794 650 852 678
rect 794 616 806 650
rect 840 616 852 650
rect 794 318 852 616
rect 882 650 940 678
rect 882 616 894 650
rect 928 616 940 650
rect 882 318 940 616
rect 998 650 1056 678
rect 998 616 1010 650
rect 1044 616 1056 650
rect 998 498 1056 616
rect 1086 650 1144 678
rect 1264 650 1322 678
rect 1086 616 1098 650
rect 1132 616 1144 650
rect 1086 498 1144 616
rect 1264 616 1276 650
rect 1310 616 1322 650
rect 1264 498 1322 616
rect 1352 650 1410 678
rect 1496 650 1554 678
rect 1352 616 1364 650
rect 1398 616 1410 650
rect 1352 498 1410 616
rect 1496 616 1508 650
rect 1542 616 1554 650
rect 1496 498 1554 616
rect 1584 650 1642 678
rect 1728 650 1786 678
rect 1584 616 1596 650
rect 1630 616 1642 650
rect 1584 498 1642 616
rect 1728 616 1740 650
rect 1774 616 1786 650
rect 1728 498 1786 616
rect 1816 650 1874 678
rect 1960 650 2018 678
rect 1816 616 1828 650
rect 1862 616 1874 650
rect 1816 498 1874 616
rect 1960 616 1972 650
rect 2006 616 2018 650
rect 1960 318 2018 616
rect 2048 650 2106 678
rect 2048 616 2060 650
rect 2094 616 2106 650
rect 2048 318 2106 616
rect 2136 650 2194 678
rect 2136 616 2148 650
rect 2182 616 2194 650
rect 2136 318 2194 616
<< ndiffc >>
rect -18 48 16 82
rect 70 48 104 82
rect 222 48 256 82
rect 310 48 344 82
rect 486 48 520 82
rect 574 48 608 82
rect 718 48 752 82
rect 806 48 840 82
rect 894 48 928 82
rect 1010 48 1044 82
rect 1098 48 1132 82
rect 1276 48 1310 82
rect 1364 48 1398 82
rect 1508 48 1542 82
rect 1596 48 1630 82
rect 1740 48 1774 82
rect 1828 48 1862 82
rect 1972 48 2006 82
rect 2060 48 2094 82
rect 2148 48 2182 82
<< pdiffc >>
rect -18 616 16 650
rect 70 616 104 650
rect 222 616 256 650
rect 310 616 344 650
rect 486 616 520 650
rect 574 616 608 650
rect 718 616 752 650
rect 806 616 840 650
rect 894 616 928 650
rect 1010 616 1044 650
rect 1098 616 1132 650
rect 1276 616 1310 650
rect 1364 616 1398 650
rect 1508 616 1542 650
rect 1596 616 1630 650
rect 1740 616 1774 650
rect 1828 616 1862 650
rect 1972 616 2006 650
rect 2060 616 2094 650
rect 2148 616 2182 650
<< psubdiff >>
rect 14 -68 58 -34
rect 2106 -68 2154 -34
<< nsubdiff >>
rect 4 732 58 766
rect 2106 732 2154 766
<< psubdiffcont >>
rect 58 -68 2106 -34
<< nsubdiffcont >>
rect 58 732 2106 766
<< poly >>
rect 28 678 58 704
rect 268 678 298 704
rect 532 678 562 704
rect 764 678 794 704
rect 852 678 882 704
rect 1056 678 1086 704
rect 1322 678 1352 704
rect 1554 678 1584 704
rect 1786 678 1816 704
rect 2018 678 2048 704
rect 2106 678 2136 704
rect 140 650 194 666
rect 140 616 150 650
rect 184 616 194 650
rect 140 600 194 616
rect 28 410 58 498
rect 28 394 108 410
rect 28 360 64 394
rect 98 360 108 394
rect 28 344 108 360
rect 28 110 58 344
rect 150 280 184 600
rect 372 650 426 666
rect 372 616 382 650
rect 416 616 426 650
rect 372 606 426 616
rect 380 600 416 606
rect 268 472 298 498
rect 250 438 266 472
rect 300 438 316 472
rect 250 436 316 438
rect 247 384 315 394
rect 247 350 265 384
rect 299 350 315 384
rect 247 333 315 350
rect 140 270 194 280
rect 140 236 150 270
rect 184 236 194 270
rect 140 226 194 236
rect 150 82 184 226
rect 268 110 298 333
rect 380 234 414 600
rect 646 650 680 666
rect 455 472 489 488
rect 457 422 489 438
rect 457 312 487 422
rect 532 394 562 498
rect 530 344 564 360
rect 457 282 562 312
rect 380 82 414 200
rect 532 110 562 282
rect 646 82 680 616
rect 764 302 794 318
rect 764 110 794 268
rect 852 166 882 318
rect 1056 234 1086 498
rect 852 132 980 166
rect 852 110 882 132
rect 1056 110 1086 200
rect 1170 166 1204 616
rect 1246 314 1280 438
rect 1322 394 1352 498
rect 1246 280 1352 314
rect 1170 82 1204 132
rect 1322 110 1352 280
rect 1436 234 1470 616
rect 1554 472 1584 498
rect 1554 394 1584 396
rect 1436 82 1470 200
rect 1554 110 1584 360
rect 1666 82 1700 616
rect 1786 394 1816 498
rect 1902 394 1936 616
rect 1786 360 1936 394
rect 1786 110 1816 360
rect 1902 82 1936 360
rect 2018 234 2048 318
rect 2106 302 2136 318
rect 2018 110 2048 200
rect 2106 110 2136 268
rect 28 -6 58 20
rect 268 -6 298 20
rect 532 -6 562 20
rect 764 -6 794 20
rect 852 -6 882 20
rect 1056 -6 1086 20
rect 1322 -6 1352 20
rect 1554 -6 1584 20
rect 1786 -6 1816 20
rect 2018 -6 2048 20
rect 2106 -6 2136 20
<< polycont >>
rect 150 616 184 650
rect 64 360 98 394
rect 382 616 416 650
rect 266 438 300 472
rect 265 350 299 384
rect 150 236 184 270
rect 646 616 680 650
rect 455 438 489 472
rect 530 360 564 394
rect 380 200 414 234
rect 150 48 184 82
rect 380 48 414 82
rect 1170 616 1204 650
rect 762 268 796 302
rect 1054 200 1088 234
rect 980 132 1014 166
rect 1436 616 1470 650
rect 1246 438 1280 472
rect 1320 360 1354 394
rect 1170 132 1204 166
rect 646 48 680 82
rect 1666 616 1700 650
rect 1552 438 1586 472
rect 1552 360 1586 394
rect 1436 200 1470 234
rect 1170 48 1204 82
rect 1436 48 1470 82
rect 1902 616 1936 650
rect 1666 48 1700 82
rect 2104 268 2138 302
rect 2018 200 2052 234
rect 1902 48 1936 82
<< locali >>
rect 14 732 58 766
rect 2106 732 2182 766
rect -23 650 16 666
rect -23 616 -18 650
rect -23 472 16 616
rect 70 650 104 732
rect 70 600 104 616
rect 150 650 256 666
rect 184 616 222 650
rect 150 600 256 616
rect 310 650 520 666
rect 344 616 382 650
rect 416 616 486 650
rect 310 600 520 616
rect 574 650 752 666
rect 608 616 646 650
rect 680 616 718 650
rect 574 600 752 616
rect 806 650 840 666
rect 806 600 840 616
rect 894 650 928 732
rect 894 600 928 616
rect 1010 650 1044 732
rect 1010 600 1044 616
rect 1098 650 1310 666
rect 1132 616 1170 650
rect 1204 616 1276 650
rect 1098 600 1310 616
rect 1364 650 1542 666
rect 1398 616 1436 650
rect 1470 616 1508 650
rect 1364 600 1542 616
rect 1596 650 1774 666
rect 1630 616 1666 650
rect 1700 616 1740 650
rect 1596 600 1774 616
rect 1828 650 1862 732
rect 1828 600 1862 616
rect 1902 650 2006 666
rect 1936 616 1972 650
rect 1902 600 2006 616
rect 2060 650 2094 666
rect 2060 600 2094 616
rect 2148 650 2182 732
rect 2148 600 2182 616
rect -23 438 266 472
rect 300 438 455 472
rect 489 438 1246 472
rect 1280 438 1552 472
rect 1586 438 1602 472
rect -23 175 14 438
rect 48 360 64 394
rect 98 384 530 394
rect 98 360 265 384
rect 249 350 265 360
rect 299 360 530 384
rect 564 360 1320 394
rect 1354 360 1552 394
rect 1586 360 1602 394
rect 299 350 315 360
rect 249 334 315 350
rect 150 270 184 286
rect 746 268 762 302
rect 796 268 2104 302
rect 2138 268 2154 302
rect 150 220 184 236
rect 364 200 380 234
rect 414 200 1054 234
rect 1088 200 1104 234
rect 1420 200 1436 234
rect 1470 200 2018 234
rect 2052 200 2068 234
rect -23 82 16 175
rect 718 132 928 166
rect 964 132 980 166
rect 1014 132 1170 166
rect 1204 132 1220 166
rect 1972 132 2182 166
rect 718 98 752 132
rect -23 48 -18 82
rect -23 32 16 48
rect 70 82 104 98
rect 70 -34 104 48
rect 150 82 256 98
rect 184 48 222 82
rect 150 32 256 48
rect 310 82 520 98
rect 344 48 380 82
rect 414 48 486 82
rect 310 32 520 48
rect 574 82 752 98
rect 608 48 646 82
rect 680 48 718 82
rect 574 32 752 48
rect 806 82 840 98
rect 806 -34 840 48
rect 894 82 928 132
rect 1972 98 2006 132
rect 894 32 928 48
rect 1010 82 1044 98
rect 1010 -34 1044 48
rect 1098 82 1310 98
rect 1132 48 1170 82
rect 1204 48 1276 82
rect 1098 32 1310 48
rect 1364 82 1542 98
rect 1398 48 1436 82
rect 1470 48 1508 82
rect 1364 32 1542 48
rect 1596 82 1774 98
rect 1630 48 1666 82
rect 1700 48 1740 82
rect 1596 32 1774 48
rect 1828 82 1862 98
rect 1828 -34 1862 48
rect 1902 82 2006 98
rect 1936 48 1972 82
rect 1902 32 2006 48
rect 2060 82 2094 98
rect 2060 -34 2094 48
rect 2148 82 2182 132
rect 2148 32 2182 48
rect 14 -68 58 -34
rect 2106 -68 2138 -34
<< viali >>
rect 58 732 2106 766
rect 64 360 98 394
rect 150 236 184 270
rect 762 268 796 302
rect 1666 48 1700 82
rect 1902 48 1936 82
rect 58 -68 2106 -34
<< metal1 >>
rect -66 766 2230 804
rect -66 732 58 766
rect 2106 732 2230 766
rect -66 694 2230 732
rect 50 394 118 406
rect 50 360 64 394
rect 98 360 118 394
rect 50 348 118 360
rect 750 302 808 314
rect 138 270 196 282
rect 138 236 150 270
rect 184 236 196 270
rect 750 268 762 302
rect 796 268 808 302
rect 750 256 808 268
rect 138 224 196 236
rect 1654 82 1714 94
rect 1654 48 1666 82
rect 1700 48 1714 82
rect 1654 36 1714 48
rect 1890 82 1948 94
rect 1890 48 1902 82
rect 1936 48 1948 82
rect 1890 36 1948 48
rect -66 -34 2230 4
rect -66 -68 58 -34
rect 2106 -68 2230 -34
rect -66 -106 2230 -68
<< labels >>
rlabel metal1 1072 -106 1072 -106 5 VSS
rlabel metal1 1070 804 1070 804 1 VDD
rlabel metal1 88 348 88 348 5 CLK
rlabel metal1 138 252 138 252 7 D
rlabel metal1 780 256 780 256 5 CLR
rlabel metal1 1684 36 1684 36 5 Qb
rlabel metal1 1920 36 1920 36 5 Q
<< end >>
