magic
tech sky130A
magscale 1 2
timestamp 1616184658
<< error_p >>
rect -1445 3131 -1387 3137
rect -1327 3131 -1269 3137
rect -1209 3131 -1151 3137
rect -1091 3131 -1033 3137
rect -973 3131 -915 3137
rect -855 3131 -797 3137
rect -737 3131 -679 3137
rect -619 3131 -561 3137
rect -501 3131 -443 3137
rect -383 3131 -325 3137
rect -265 3131 -207 3137
rect -147 3131 -89 3137
rect -29 3131 29 3137
rect 89 3131 147 3137
rect 207 3131 265 3137
rect 325 3131 383 3137
rect 443 3131 501 3137
rect 561 3131 619 3137
rect 679 3131 737 3137
rect 797 3131 855 3137
rect 915 3131 973 3137
rect 1033 3131 1091 3137
rect 1151 3131 1209 3137
rect 1269 3131 1327 3137
rect 1387 3131 1445 3137
rect -1445 3097 -1433 3131
rect -1327 3097 -1315 3131
rect -1209 3097 -1197 3131
rect -1091 3097 -1079 3131
rect -973 3097 -961 3131
rect -855 3097 -843 3131
rect -737 3097 -725 3131
rect -619 3097 -607 3131
rect -501 3097 -489 3131
rect -383 3097 -371 3131
rect -265 3097 -253 3131
rect -147 3097 -135 3131
rect -29 3097 -17 3131
rect 89 3097 101 3131
rect 207 3097 219 3131
rect 325 3097 337 3131
rect 443 3097 455 3131
rect 561 3097 573 3131
rect 679 3097 691 3131
rect 797 3097 809 3131
rect 915 3097 927 3131
rect 1033 3097 1045 3131
rect 1151 3097 1163 3131
rect 1269 3097 1281 3131
rect 1387 3097 1399 3131
rect -1445 3091 -1387 3097
rect -1327 3091 -1269 3097
rect -1209 3091 -1151 3097
rect -1091 3091 -1033 3097
rect -973 3091 -915 3097
rect -855 3091 -797 3097
rect -737 3091 -679 3097
rect -619 3091 -561 3097
rect -501 3091 -443 3097
rect -383 3091 -325 3097
rect -265 3091 -207 3097
rect -147 3091 -89 3097
rect -29 3091 29 3097
rect 89 3091 147 3097
rect 207 3091 265 3097
rect 325 3091 383 3097
rect 443 3091 501 3097
rect 561 3091 619 3097
rect 679 3091 737 3097
rect 797 3091 855 3097
rect 915 3091 973 3097
rect 1033 3091 1091 3097
rect 1151 3091 1209 3097
rect 1269 3091 1327 3097
rect 1387 3091 1445 3097
rect -1445 2366 -1387 2372
rect -1327 2366 -1269 2372
rect -1209 2366 -1151 2372
rect -1091 2366 -1033 2372
rect -973 2366 -915 2372
rect -855 2366 -797 2372
rect -737 2366 -679 2372
rect -619 2366 -561 2372
rect -501 2366 -443 2372
rect -383 2366 -325 2372
rect -265 2366 -207 2372
rect -147 2366 -89 2372
rect -29 2366 29 2372
rect 89 2366 147 2372
rect 207 2366 265 2372
rect 325 2366 383 2372
rect 443 2366 501 2372
rect 561 2366 619 2372
rect 679 2366 737 2372
rect 797 2366 855 2372
rect 915 2366 973 2372
rect 1033 2366 1091 2372
rect 1151 2366 1209 2372
rect 1269 2366 1327 2372
rect 1387 2366 1445 2372
rect -1445 2332 -1433 2366
rect -1327 2332 -1315 2366
rect -1209 2332 -1197 2366
rect -1091 2332 -1079 2366
rect -973 2332 -961 2366
rect -855 2332 -843 2366
rect -737 2332 -725 2366
rect -619 2332 -607 2366
rect -501 2332 -489 2366
rect -383 2332 -371 2366
rect -265 2332 -253 2366
rect -147 2332 -135 2366
rect -29 2332 -17 2366
rect 89 2332 101 2366
rect 207 2332 219 2366
rect 325 2332 337 2366
rect 443 2332 455 2366
rect 561 2332 573 2366
rect 679 2332 691 2366
rect 797 2332 809 2366
rect 915 2332 927 2366
rect 1033 2332 1045 2366
rect 1151 2332 1163 2366
rect 1269 2332 1281 2366
rect 1387 2332 1399 2366
rect -1445 2326 -1387 2332
rect -1327 2326 -1269 2332
rect -1209 2326 -1151 2332
rect -1091 2326 -1033 2332
rect -973 2326 -915 2332
rect -855 2326 -797 2332
rect -737 2326 -679 2332
rect -619 2326 -561 2332
rect -501 2326 -443 2332
rect -383 2326 -325 2332
rect -265 2326 -207 2332
rect -147 2326 -89 2332
rect -29 2326 29 2332
rect 89 2326 147 2332
rect 207 2326 265 2332
rect 325 2326 383 2332
rect 443 2326 501 2332
rect 561 2326 619 2332
rect 679 2326 737 2332
rect 797 2326 855 2332
rect 915 2326 973 2332
rect 1033 2326 1091 2332
rect 1151 2326 1209 2332
rect 1269 2326 1327 2332
rect 1387 2326 1445 2332
rect -1445 1601 -1387 1607
rect -1327 1601 -1269 1607
rect -1209 1601 -1151 1607
rect -1091 1601 -1033 1607
rect -973 1601 -915 1607
rect -855 1601 -797 1607
rect -737 1601 -679 1607
rect -619 1601 -561 1607
rect -501 1601 -443 1607
rect -383 1601 -325 1607
rect -265 1601 -207 1607
rect -147 1601 -89 1607
rect -29 1601 29 1607
rect 89 1601 147 1607
rect 207 1601 265 1607
rect 325 1601 383 1607
rect 443 1601 501 1607
rect 561 1601 619 1607
rect 679 1601 737 1607
rect 797 1601 855 1607
rect 915 1601 973 1607
rect 1033 1601 1091 1607
rect 1151 1601 1209 1607
rect 1269 1601 1327 1607
rect 1387 1601 1445 1607
rect -1445 1567 -1433 1601
rect -1327 1567 -1315 1601
rect -1209 1567 -1197 1601
rect -1091 1567 -1079 1601
rect -973 1567 -961 1601
rect -855 1567 -843 1601
rect -737 1567 -725 1601
rect -619 1567 -607 1601
rect -501 1567 -489 1601
rect -383 1567 -371 1601
rect -265 1567 -253 1601
rect -147 1567 -135 1601
rect -29 1567 -17 1601
rect 89 1567 101 1601
rect 207 1567 219 1601
rect 325 1567 337 1601
rect 443 1567 455 1601
rect 561 1567 573 1601
rect 679 1567 691 1601
rect 797 1567 809 1601
rect 915 1567 927 1601
rect 1033 1567 1045 1601
rect 1151 1567 1163 1601
rect 1269 1567 1281 1601
rect 1387 1567 1399 1601
rect -1445 1561 -1387 1567
rect -1327 1561 -1269 1567
rect -1209 1561 -1151 1567
rect -1091 1561 -1033 1567
rect -973 1561 -915 1567
rect -855 1561 -797 1567
rect -737 1561 -679 1567
rect -619 1561 -561 1567
rect -501 1561 -443 1567
rect -383 1561 -325 1567
rect -265 1561 -207 1567
rect -147 1561 -89 1567
rect -29 1561 29 1567
rect 89 1561 147 1567
rect 207 1561 265 1567
rect 325 1561 383 1567
rect 443 1561 501 1567
rect 561 1561 619 1567
rect 679 1561 737 1567
rect 797 1561 855 1567
rect 915 1561 973 1567
rect 1033 1561 1091 1567
rect 1151 1561 1209 1567
rect 1269 1561 1327 1567
rect 1387 1561 1445 1567
rect -1445 836 -1387 842
rect -1327 836 -1269 842
rect -1209 836 -1151 842
rect -1091 836 -1033 842
rect -973 836 -915 842
rect -855 836 -797 842
rect -737 836 -679 842
rect -619 836 -561 842
rect -501 836 -443 842
rect -383 836 -325 842
rect -265 836 -207 842
rect -147 836 -89 842
rect -29 836 29 842
rect 89 836 147 842
rect 207 836 265 842
rect 325 836 383 842
rect 443 836 501 842
rect 561 836 619 842
rect 679 836 737 842
rect 797 836 855 842
rect 915 836 973 842
rect 1033 836 1091 842
rect 1151 836 1209 842
rect 1269 836 1327 842
rect 1387 836 1445 842
rect -1445 802 -1433 836
rect -1327 802 -1315 836
rect -1209 802 -1197 836
rect -1091 802 -1079 836
rect -973 802 -961 836
rect -855 802 -843 836
rect -737 802 -725 836
rect -619 802 -607 836
rect -501 802 -489 836
rect -383 802 -371 836
rect -265 802 -253 836
rect -147 802 -135 836
rect -29 802 -17 836
rect 89 802 101 836
rect 207 802 219 836
rect 325 802 337 836
rect 443 802 455 836
rect 561 802 573 836
rect 679 802 691 836
rect 797 802 809 836
rect 915 802 927 836
rect 1033 802 1045 836
rect 1151 802 1163 836
rect 1269 802 1281 836
rect 1387 802 1399 836
rect -1445 796 -1387 802
rect -1327 796 -1269 802
rect -1209 796 -1151 802
rect -1091 796 -1033 802
rect -973 796 -915 802
rect -855 796 -797 802
rect -737 796 -679 802
rect -619 796 -561 802
rect -501 796 -443 802
rect -383 796 -325 802
rect -265 796 -207 802
rect -147 796 -89 802
rect -29 796 29 802
rect 89 796 147 802
rect 207 796 265 802
rect 325 796 383 802
rect 443 796 501 802
rect 561 796 619 802
rect 679 796 737 802
rect 797 796 855 802
rect 915 796 973 802
rect 1033 796 1091 802
rect 1151 796 1209 802
rect 1269 796 1327 802
rect 1387 796 1445 802
rect -1445 71 -1387 77
rect -1327 71 -1269 77
rect -1209 71 -1151 77
rect -1091 71 -1033 77
rect -973 71 -915 77
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect 915 71 973 77
rect 1033 71 1091 77
rect 1151 71 1209 77
rect 1269 71 1327 77
rect 1387 71 1445 77
rect -1445 37 -1433 71
rect -1327 37 -1315 71
rect -1209 37 -1197 71
rect -1091 37 -1079 71
rect -973 37 -961 71
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect 915 37 927 71
rect 1033 37 1045 71
rect 1151 37 1163 71
rect 1269 37 1281 71
rect 1387 37 1399 71
rect -1445 31 -1387 37
rect -1327 31 -1269 37
rect -1209 31 -1151 37
rect -1091 31 -1033 37
rect -973 31 -915 37
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect 915 31 973 37
rect 1033 31 1091 37
rect 1151 31 1209 37
rect 1269 31 1327 37
rect 1387 31 1445 37
rect -1445 -694 -1387 -688
rect -1327 -694 -1269 -688
rect -1209 -694 -1151 -688
rect -1091 -694 -1033 -688
rect -973 -694 -915 -688
rect -855 -694 -797 -688
rect -737 -694 -679 -688
rect -619 -694 -561 -688
rect -501 -694 -443 -688
rect -383 -694 -325 -688
rect -265 -694 -207 -688
rect -147 -694 -89 -688
rect -29 -694 29 -688
rect 89 -694 147 -688
rect 207 -694 265 -688
rect 325 -694 383 -688
rect 443 -694 501 -688
rect 561 -694 619 -688
rect 679 -694 737 -688
rect 797 -694 855 -688
rect 915 -694 973 -688
rect 1033 -694 1091 -688
rect 1151 -694 1209 -688
rect 1269 -694 1327 -688
rect 1387 -694 1445 -688
rect -1445 -728 -1433 -694
rect -1327 -728 -1315 -694
rect -1209 -728 -1197 -694
rect -1091 -728 -1079 -694
rect -973 -728 -961 -694
rect -855 -728 -843 -694
rect -737 -728 -725 -694
rect -619 -728 -607 -694
rect -501 -728 -489 -694
rect -383 -728 -371 -694
rect -265 -728 -253 -694
rect -147 -728 -135 -694
rect -29 -728 -17 -694
rect 89 -728 101 -694
rect 207 -728 219 -694
rect 325 -728 337 -694
rect 443 -728 455 -694
rect 561 -728 573 -694
rect 679 -728 691 -694
rect 797 -728 809 -694
rect 915 -728 927 -694
rect 1033 -728 1045 -694
rect 1151 -728 1163 -694
rect 1269 -728 1281 -694
rect 1387 -728 1399 -694
rect -1445 -734 -1387 -728
rect -1327 -734 -1269 -728
rect -1209 -734 -1151 -728
rect -1091 -734 -1033 -728
rect -973 -734 -915 -728
rect -855 -734 -797 -728
rect -737 -734 -679 -728
rect -619 -734 -561 -728
rect -501 -734 -443 -728
rect -383 -734 -325 -728
rect -265 -734 -207 -728
rect -147 -734 -89 -728
rect -29 -734 29 -728
rect 89 -734 147 -728
rect 207 -734 265 -728
rect 325 -734 383 -728
rect 443 -734 501 -728
rect 561 -734 619 -728
rect 679 -734 737 -728
rect 797 -734 855 -728
rect 915 -734 973 -728
rect 1033 -734 1091 -728
rect 1151 -734 1209 -728
rect 1269 -734 1327 -728
rect 1387 -734 1445 -728
rect -1445 -1459 -1387 -1453
rect -1327 -1459 -1269 -1453
rect -1209 -1459 -1151 -1453
rect -1091 -1459 -1033 -1453
rect -973 -1459 -915 -1453
rect -855 -1459 -797 -1453
rect -737 -1459 -679 -1453
rect -619 -1459 -561 -1453
rect -501 -1459 -443 -1453
rect -383 -1459 -325 -1453
rect -265 -1459 -207 -1453
rect -147 -1459 -89 -1453
rect -29 -1459 29 -1453
rect 89 -1459 147 -1453
rect 207 -1459 265 -1453
rect 325 -1459 383 -1453
rect 443 -1459 501 -1453
rect 561 -1459 619 -1453
rect 679 -1459 737 -1453
rect 797 -1459 855 -1453
rect 915 -1459 973 -1453
rect 1033 -1459 1091 -1453
rect 1151 -1459 1209 -1453
rect 1269 -1459 1327 -1453
rect 1387 -1459 1445 -1453
rect -1445 -1493 -1433 -1459
rect -1327 -1493 -1315 -1459
rect -1209 -1493 -1197 -1459
rect -1091 -1493 -1079 -1459
rect -973 -1493 -961 -1459
rect -855 -1493 -843 -1459
rect -737 -1493 -725 -1459
rect -619 -1493 -607 -1459
rect -501 -1493 -489 -1459
rect -383 -1493 -371 -1459
rect -265 -1493 -253 -1459
rect -147 -1493 -135 -1459
rect -29 -1493 -17 -1459
rect 89 -1493 101 -1459
rect 207 -1493 219 -1459
rect 325 -1493 337 -1459
rect 443 -1493 455 -1459
rect 561 -1493 573 -1459
rect 679 -1493 691 -1459
rect 797 -1493 809 -1459
rect 915 -1493 927 -1459
rect 1033 -1493 1045 -1459
rect 1151 -1493 1163 -1459
rect 1269 -1493 1281 -1459
rect 1387 -1493 1399 -1459
rect -1445 -1499 -1387 -1493
rect -1327 -1499 -1269 -1493
rect -1209 -1499 -1151 -1493
rect -1091 -1499 -1033 -1493
rect -973 -1499 -915 -1493
rect -855 -1499 -797 -1493
rect -737 -1499 -679 -1493
rect -619 -1499 -561 -1493
rect -501 -1499 -443 -1493
rect -383 -1499 -325 -1493
rect -265 -1499 -207 -1493
rect -147 -1499 -89 -1493
rect -29 -1499 29 -1493
rect 89 -1499 147 -1493
rect 207 -1499 265 -1493
rect 325 -1499 383 -1493
rect 443 -1499 501 -1493
rect 561 -1499 619 -1493
rect 679 -1499 737 -1493
rect 797 -1499 855 -1493
rect 915 -1499 973 -1493
rect 1033 -1499 1091 -1493
rect 1151 -1499 1209 -1493
rect 1269 -1499 1327 -1493
rect 1387 -1499 1445 -1493
rect -1445 -2224 -1387 -2218
rect -1327 -2224 -1269 -2218
rect -1209 -2224 -1151 -2218
rect -1091 -2224 -1033 -2218
rect -973 -2224 -915 -2218
rect -855 -2224 -797 -2218
rect -737 -2224 -679 -2218
rect -619 -2224 -561 -2218
rect -501 -2224 -443 -2218
rect -383 -2224 -325 -2218
rect -265 -2224 -207 -2218
rect -147 -2224 -89 -2218
rect -29 -2224 29 -2218
rect 89 -2224 147 -2218
rect 207 -2224 265 -2218
rect 325 -2224 383 -2218
rect 443 -2224 501 -2218
rect 561 -2224 619 -2218
rect 679 -2224 737 -2218
rect 797 -2224 855 -2218
rect 915 -2224 973 -2218
rect 1033 -2224 1091 -2218
rect 1151 -2224 1209 -2218
rect 1269 -2224 1327 -2218
rect 1387 -2224 1445 -2218
rect -1445 -2258 -1433 -2224
rect -1327 -2258 -1315 -2224
rect -1209 -2258 -1197 -2224
rect -1091 -2258 -1079 -2224
rect -973 -2258 -961 -2224
rect -855 -2258 -843 -2224
rect -737 -2258 -725 -2224
rect -619 -2258 -607 -2224
rect -501 -2258 -489 -2224
rect -383 -2258 -371 -2224
rect -265 -2258 -253 -2224
rect -147 -2258 -135 -2224
rect -29 -2258 -17 -2224
rect 89 -2258 101 -2224
rect 207 -2258 219 -2224
rect 325 -2258 337 -2224
rect 443 -2258 455 -2224
rect 561 -2258 573 -2224
rect 679 -2258 691 -2224
rect 797 -2258 809 -2224
rect 915 -2258 927 -2224
rect 1033 -2258 1045 -2224
rect 1151 -2258 1163 -2224
rect 1269 -2258 1281 -2224
rect 1387 -2258 1399 -2224
rect -1445 -2264 -1387 -2258
rect -1327 -2264 -1269 -2258
rect -1209 -2264 -1151 -2258
rect -1091 -2264 -1033 -2258
rect -973 -2264 -915 -2258
rect -855 -2264 -797 -2258
rect -737 -2264 -679 -2258
rect -619 -2264 -561 -2258
rect -501 -2264 -443 -2258
rect -383 -2264 -325 -2258
rect -265 -2264 -207 -2258
rect -147 -2264 -89 -2258
rect -29 -2264 29 -2258
rect 89 -2264 147 -2258
rect 207 -2264 265 -2258
rect 325 -2264 383 -2258
rect 443 -2264 501 -2258
rect 561 -2264 619 -2258
rect 679 -2264 737 -2258
rect 797 -2264 855 -2258
rect 915 -2264 973 -2258
rect 1033 -2264 1091 -2258
rect 1151 -2264 1209 -2258
rect 1269 -2264 1327 -2258
rect 1387 -2264 1445 -2258
rect -1445 -2989 -1387 -2983
rect -1327 -2989 -1269 -2983
rect -1209 -2989 -1151 -2983
rect -1091 -2989 -1033 -2983
rect -973 -2989 -915 -2983
rect -855 -2989 -797 -2983
rect -737 -2989 -679 -2983
rect -619 -2989 -561 -2983
rect -501 -2989 -443 -2983
rect -383 -2989 -325 -2983
rect -265 -2989 -207 -2983
rect -147 -2989 -89 -2983
rect -29 -2989 29 -2983
rect 89 -2989 147 -2983
rect 207 -2989 265 -2983
rect 325 -2989 383 -2983
rect 443 -2989 501 -2983
rect 561 -2989 619 -2983
rect 679 -2989 737 -2983
rect 797 -2989 855 -2983
rect 915 -2989 973 -2983
rect 1033 -2989 1091 -2983
rect 1151 -2989 1209 -2983
rect 1269 -2989 1327 -2983
rect 1387 -2989 1445 -2983
rect -1445 -3023 -1433 -2989
rect -1327 -3023 -1315 -2989
rect -1209 -3023 -1197 -2989
rect -1091 -3023 -1079 -2989
rect -973 -3023 -961 -2989
rect -855 -3023 -843 -2989
rect -737 -3023 -725 -2989
rect -619 -3023 -607 -2989
rect -501 -3023 -489 -2989
rect -383 -3023 -371 -2989
rect -265 -3023 -253 -2989
rect -147 -3023 -135 -2989
rect -29 -3023 -17 -2989
rect 89 -3023 101 -2989
rect 207 -3023 219 -2989
rect 325 -3023 337 -2989
rect 443 -3023 455 -2989
rect 561 -3023 573 -2989
rect 679 -3023 691 -2989
rect 797 -3023 809 -2989
rect 915 -3023 927 -2989
rect 1033 -3023 1045 -2989
rect 1151 -3023 1163 -2989
rect 1269 -3023 1281 -2989
rect 1387 -3023 1399 -2989
rect -1445 -3029 -1387 -3023
rect -1327 -3029 -1269 -3023
rect -1209 -3029 -1151 -3023
rect -1091 -3029 -1033 -3023
rect -973 -3029 -915 -3023
rect -855 -3029 -797 -3023
rect -737 -3029 -679 -3023
rect -619 -3029 -561 -3023
rect -501 -3029 -443 -3023
rect -383 -3029 -325 -3023
rect -265 -3029 -207 -3023
rect -147 -3029 -89 -3023
rect -29 -3029 29 -3023
rect 89 -3029 147 -3023
rect 207 -3029 265 -3023
rect 325 -3029 383 -3023
rect 443 -3029 501 -3023
rect 561 -3029 619 -3023
rect 679 -3029 737 -3023
rect 797 -3029 855 -3023
rect 915 -3029 973 -3023
rect 1033 -3029 1091 -3023
rect 1151 -3029 1209 -3023
rect 1269 -3029 1327 -3023
rect 1387 -3029 1445 -3023
rect -1445 -3754 -1387 -3748
rect -1327 -3754 -1269 -3748
rect -1209 -3754 -1151 -3748
rect -1091 -3754 -1033 -3748
rect -973 -3754 -915 -3748
rect -855 -3754 -797 -3748
rect -737 -3754 -679 -3748
rect -619 -3754 -561 -3748
rect -501 -3754 -443 -3748
rect -383 -3754 -325 -3748
rect -265 -3754 -207 -3748
rect -147 -3754 -89 -3748
rect -29 -3754 29 -3748
rect 89 -3754 147 -3748
rect 207 -3754 265 -3748
rect 325 -3754 383 -3748
rect 443 -3754 501 -3748
rect 561 -3754 619 -3748
rect 679 -3754 737 -3748
rect 797 -3754 855 -3748
rect 915 -3754 973 -3748
rect 1033 -3754 1091 -3748
rect 1151 -3754 1209 -3748
rect 1269 -3754 1327 -3748
rect 1387 -3754 1445 -3748
rect -1445 -3788 -1433 -3754
rect -1327 -3788 -1315 -3754
rect -1209 -3788 -1197 -3754
rect -1091 -3788 -1079 -3754
rect -973 -3788 -961 -3754
rect -855 -3788 -843 -3754
rect -737 -3788 -725 -3754
rect -619 -3788 -607 -3754
rect -501 -3788 -489 -3754
rect -383 -3788 -371 -3754
rect -265 -3788 -253 -3754
rect -147 -3788 -135 -3754
rect -29 -3788 -17 -3754
rect 89 -3788 101 -3754
rect 207 -3788 219 -3754
rect 325 -3788 337 -3754
rect 443 -3788 455 -3754
rect 561 -3788 573 -3754
rect 679 -3788 691 -3754
rect 797 -3788 809 -3754
rect 915 -3788 927 -3754
rect 1033 -3788 1045 -3754
rect 1151 -3788 1163 -3754
rect 1269 -3788 1281 -3754
rect 1387 -3788 1399 -3754
rect -1445 -3794 -1387 -3788
rect -1327 -3794 -1269 -3788
rect -1209 -3794 -1151 -3788
rect -1091 -3794 -1033 -3788
rect -973 -3794 -915 -3788
rect -855 -3794 -797 -3788
rect -737 -3794 -679 -3788
rect -619 -3794 -561 -3788
rect -501 -3794 -443 -3788
rect -383 -3794 -325 -3788
rect -265 -3794 -207 -3788
rect -147 -3794 -89 -3788
rect -29 -3794 29 -3788
rect 89 -3794 147 -3788
rect 207 -3794 265 -3788
rect 325 -3794 383 -3788
rect 443 -3794 501 -3788
rect 561 -3794 619 -3788
rect 679 -3794 737 -3788
rect 797 -3794 855 -3788
rect 915 -3794 973 -3788
rect 1033 -3794 1091 -3788
rect 1151 -3794 1209 -3788
rect 1269 -3794 1327 -3788
rect 1387 -3794 1445 -3788
<< nwell >>
rect -1642 -3926 1642 3926
<< pmos >>
rect -1446 3178 -1386 3778
rect -1328 3178 -1268 3778
rect -1210 3178 -1150 3778
rect -1092 3178 -1032 3778
rect -974 3178 -914 3778
rect -856 3178 -796 3778
rect -738 3178 -678 3778
rect -620 3178 -560 3778
rect -502 3178 -442 3778
rect -384 3178 -324 3778
rect -266 3178 -206 3778
rect -148 3178 -88 3778
rect -30 3178 30 3778
rect 88 3178 148 3778
rect 206 3178 266 3778
rect 324 3178 384 3778
rect 442 3178 502 3778
rect 560 3178 620 3778
rect 678 3178 738 3778
rect 796 3178 856 3778
rect 914 3178 974 3778
rect 1032 3178 1092 3778
rect 1150 3178 1210 3778
rect 1268 3178 1328 3778
rect 1386 3178 1446 3778
rect -1446 2413 -1386 3013
rect -1328 2413 -1268 3013
rect -1210 2413 -1150 3013
rect -1092 2413 -1032 3013
rect -974 2413 -914 3013
rect -856 2413 -796 3013
rect -738 2413 -678 3013
rect -620 2413 -560 3013
rect -502 2413 -442 3013
rect -384 2413 -324 3013
rect -266 2413 -206 3013
rect -148 2413 -88 3013
rect -30 2413 30 3013
rect 88 2413 148 3013
rect 206 2413 266 3013
rect 324 2413 384 3013
rect 442 2413 502 3013
rect 560 2413 620 3013
rect 678 2413 738 3013
rect 796 2413 856 3013
rect 914 2413 974 3013
rect 1032 2413 1092 3013
rect 1150 2413 1210 3013
rect 1268 2413 1328 3013
rect 1386 2413 1446 3013
rect -1446 1648 -1386 2248
rect -1328 1648 -1268 2248
rect -1210 1648 -1150 2248
rect -1092 1648 -1032 2248
rect -974 1648 -914 2248
rect -856 1648 -796 2248
rect -738 1648 -678 2248
rect -620 1648 -560 2248
rect -502 1648 -442 2248
rect -384 1648 -324 2248
rect -266 1648 -206 2248
rect -148 1648 -88 2248
rect -30 1648 30 2248
rect 88 1648 148 2248
rect 206 1648 266 2248
rect 324 1648 384 2248
rect 442 1648 502 2248
rect 560 1648 620 2248
rect 678 1648 738 2248
rect 796 1648 856 2248
rect 914 1648 974 2248
rect 1032 1648 1092 2248
rect 1150 1648 1210 2248
rect 1268 1648 1328 2248
rect 1386 1648 1446 2248
rect -1446 883 -1386 1483
rect -1328 883 -1268 1483
rect -1210 883 -1150 1483
rect -1092 883 -1032 1483
rect -974 883 -914 1483
rect -856 883 -796 1483
rect -738 883 -678 1483
rect -620 883 -560 1483
rect -502 883 -442 1483
rect -384 883 -324 1483
rect -266 883 -206 1483
rect -148 883 -88 1483
rect -30 883 30 1483
rect 88 883 148 1483
rect 206 883 266 1483
rect 324 883 384 1483
rect 442 883 502 1483
rect 560 883 620 1483
rect 678 883 738 1483
rect 796 883 856 1483
rect 914 883 974 1483
rect 1032 883 1092 1483
rect 1150 883 1210 1483
rect 1268 883 1328 1483
rect 1386 883 1446 1483
rect -1446 118 -1386 718
rect -1328 118 -1268 718
rect -1210 118 -1150 718
rect -1092 118 -1032 718
rect -974 118 -914 718
rect -856 118 -796 718
rect -738 118 -678 718
rect -620 118 -560 718
rect -502 118 -442 718
rect -384 118 -324 718
rect -266 118 -206 718
rect -148 118 -88 718
rect -30 118 30 718
rect 88 118 148 718
rect 206 118 266 718
rect 324 118 384 718
rect 442 118 502 718
rect 560 118 620 718
rect 678 118 738 718
rect 796 118 856 718
rect 914 118 974 718
rect 1032 118 1092 718
rect 1150 118 1210 718
rect 1268 118 1328 718
rect 1386 118 1446 718
rect -1446 -647 -1386 -47
rect -1328 -647 -1268 -47
rect -1210 -647 -1150 -47
rect -1092 -647 -1032 -47
rect -974 -647 -914 -47
rect -856 -647 -796 -47
rect -738 -647 -678 -47
rect -620 -647 -560 -47
rect -502 -647 -442 -47
rect -384 -647 -324 -47
rect -266 -647 -206 -47
rect -148 -647 -88 -47
rect -30 -647 30 -47
rect 88 -647 148 -47
rect 206 -647 266 -47
rect 324 -647 384 -47
rect 442 -647 502 -47
rect 560 -647 620 -47
rect 678 -647 738 -47
rect 796 -647 856 -47
rect 914 -647 974 -47
rect 1032 -647 1092 -47
rect 1150 -647 1210 -47
rect 1268 -647 1328 -47
rect 1386 -647 1446 -47
rect -1446 -1412 -1386 -812
rect -1328 -1412 -1268 -812
rect -1210 -1412 -1150 -812
rect -1092 -1412 -1032 -812
rect -974 -1412 -914 -812
rect -856 -1412 -796 -812
rect -738 -1412 -678 -812
rect -620 -1412 -560 -812
rect -502 -1412 -442 -812
rect -384 -1412 -324 -812
rect -266 -1412 -206 -812
rect -148 -1412 -88 -812
rect -30 -1412 30 -812
rect 88 -1412 148 -812
rect 206 -1412 266 -812
rect 324 -1412 384 -812
rect 442 -1412 502 -812
rect 560 -1412 620 -812
rect 678 -1412 738 -812
rect 796 -1412 856 -812
rect 914 -1412 974 -812
rect 1032 -1412 1092 -812
rect 1150 -1412 1210 -812
rect 1268 -1412 1328 -812
rect 1386 -1412 1446 -812
rect -1446 -2177 -1386 -1577
rect -1328 -2177 -1268 -1577
rect -1210 -2177 -1150 -1577
rect -1092 -2177 -1032 -1577
rect -974 -2177 -914 -1577
rect -856 -2177 -796 -1577
rect -738 -2177 -678 -1577
rect -620 -2177 -560 -1577
rect -502 -2177 -442 -1577
rect -384 -2177 -324 -1577
rect -266 -2177 -206 -1577
rect -148 -2177 -88 -1577
rect -30 -2177 30 -1577
rect 88 -2177 148 -1577
rect 206 -2177 266 -1577
rect 324 -2177 384 -1577
rect 442 -2177 502 -1577
rect 560 -2177 620 -1577
rect 678 -2177 738 -1577
rect 796 -2177 856 -1577
rect 914 -2177 974 -1577
rect 1032 -2177 1092 -1577
rect 1150 -2177 1210 -1577
rect 1268 -2177 1328 -1577
rect 1386 -2177 1446 -1577
rect -1446 -2942 -1386 -2342
rect -1328 -2942 -1268 -2342
rect -1210 -2942 -1150 -2342
rect -1092 -2942 -1032 -2342
rect -974 -2942 -914 -2342
rect -856 -2942 -796 -2342
rect -738 -2942 -678 -2342
rect -620 -2942 -560 -2342
rect -502 -2942 -442 -2342
rect -384 -2942 -324 -2342
rect -266 -2942 -206 -2342
rect -148 -2942 -88 -2342
rect -30 -2942 30 -2342
rect 88 -2942 148 -2342
rect 206 -2942 266 -2342
rect 324 -2942 384 -2342
rect 442 -2942 502 -2342
rect 560 -2942 620 -2342
rect 678 -2942 738 -2342
rect 796 -2942 856 -2342
rect 914 -2942 974 -2342
rect 1032 -2942 1092 -2342
rect 1150 -2942 1210 -2342
rect 1268 -2942 1328 -2342
rect 1386 -2942 1446 -2342
rect -1446 -3707 -1386 -3107
rect -1328 -3707 -1268 -3107
rect -1210 -3707 -1150 -3107
rect -1092 -3707 -1032 -3107
rect -974 -3707 -914 -3107
rect -856 -3707 -796 -3107
rect -738 -3707 -678 -3107
rect -620 -3707 -560 -3107
rect -502 -3707 -442 -3107
rect -384 -3707 -324 -3107
rect -266 -3707 -206 -3107
rect -148 -3707 -88 -3107
rect -30 -3707 30 -3107
rect 88 -3707 148 -3107
rect 206 -3707 266 -3107
rect 324 -3707 384 -3107
rect 442 -3707 502 -3107
rect 560 -3707 620 -3107
rect 678 -3707 738 -3107
rect 796 -3707 856 -3107
rect 914 -3707 974 -3107
rect 1032 -3707 1092 -3107
rect 1150 -3707 1210 -3107
rect 1268 -3707 1328 -3107
rect 1386 -3707 1446 -3107
<< pdiff >>
rect -1504 3766 -1446 3778
rect -1504 3190 -1492 3766
rect -1458 3190 -1446 3766
rect -1504 3178 -1446 3190
rect -1386 3766 -1328 3778
rect -1386 3190 -1374 3766
rect -1340 3190 -1328 3766
rect -1386 3178 -1328 3190
rect -1268 3766 -1210 3778
rect -1268 3190 -1256 3766
rect -1222 3190 -1210 3766
rect -1268 3178 -1210 3190
rect -1150 3766 -1092 3778
rect -1150 3190 -1138 3766
rect -1104 3190 -1092 3766
rect -1150 3178 -1092 3190
rect -1032 3766 -974 3778
rect -1032 3190 -1020 3766
rect -986 3190 -974 3766
rect -1032 3178 -974 3190
rect -914 3766 -856 3778
rect -914 3190 -902 3766
rect -868 3190 -856 3766
rect -914 3178 -856 3190
rect -796 3766 -738 3778
rect -796 3190 -784 3766
rect -750 3190 -738 3766
rect -796 3178 -738 3190
rect -678 3766 -620 3778
rect -678 3190 -666 3766
rect -632 3190 -620 3766
rect -678 3178 -620 3190
rect -560 3766 -502 3778
rect -560 3190 -548 3766
rect -514 3190 -502 3766
rect -560 3178 -502 3190
rect -442 3766 -384 3778
rect -442 3190 -430 3766
rect -396 3190 -384 3766
rect -442 3178 -384 3190
rect -324 3766 -266 3778
rect -324 3190 -312 3766
rect -278 3190 -266 3766
rect -324 3178 -266 3190
rect -206 3766 -148 3778
rect -206 3190 -194 3766
rect -160 3190 -148 3766
rect -206 3178 -148 3190
rect -88 3766 -30 3778
rect -88 3190 -76 3766
rect -42 3190 -30 3766
rect -88 3178 -30 3190
rect 30 3766 88 3778
rect 30 3190 42 3766
rect 76 3190 88 3766
rect 30 3178 88 3190
rect 148 3766 206 3778
rect 148 3190 160 3766
rect 194 3190 206 3766
rect 148 3178 206 3190
rect 266 3766 324 3778
rect 266 3190 278 3766
rect 312 3190 324 3766
rect 266 3178 324 3190
rect 384 3766 442 3778
rect 384 3190 396 3766
rect 430 3190 442 3766
rect 384 3178 442 3190
rect 502 3766 560 3778
rect 502 3190 514 3766
rect 548 3190 560 3766
rect 502 3178 560 3190
rect 620 3766 678 3778
rect 620 3190 632 3766
rect 666 3190 678 3766
rect 620 3178 678 3190
rect 738 3766 796 3778
rect 738 3190 750 3766
rect 784 3190 796 3766
rect 738 3178 796 3190
rect 856 3766 914 3778
rect 856 3190 868 3766
rect 902 3190 914 3766
rect 856 3178 914 3190
rect 974 3766 1032 3778
rect 974 3190 986 3766
rect 1020 3190 1032 3766
rect 974 3178 1032 3190
rect 1092 3766 1150 3778
rect 1092 3190 1104 3766
rect 1138 3190 1150 3766
rect 1092 3178 1150 3190
rect 1210 3766 1268 3778
rect 1210 3190 1222 3766
rect 1256 3190 1268 3766
rect 1210 3178 1268 3190
rect 1328 3766 1386 3778
rect 1328 3190 1340 3766
rect 1374 3190 1386 3766
rect 1328 3178 1386 3190
rect 1446 3766 1504 3778
rect 1446 3190 1458 3766
rect 1492 3190 1504 3766
rect 1446 3178 1504 3190
rect -1504 3001 -1446 3013
rect -1504 2425 -1492 3001
rect -1458 2425 -1446 3001
rect -1504 2413 -1446 2425
rect -1386 3001 -1328 3013
rect -1386 2425 -1374 3001
rect -1340 2425 -1328 3001
rect -1386 2413 -1328 2425
rect -1268 3001 -1210 3013
rect -1268 2425 -1256 3001
rect -1222 2425 -1210 3001
rect -1268 2413 -1210 2425
rect -1150 3001 -1092 3013
rect -1150 2425 -1138 3001
rect -1104 2425 -1092 3001
rect -1150 2413 -1092 2425
rect -1032 3001 -974 3013
rect -1032 2425 -1020 3001
rect -986 2425 -974 3001
rect -1032 2413 -974 2425
rect -914 3001 -856 3013
rect -914 2425 -902 3001
rect -868 2425 -856 3001
rect -914 2413 -856 2425
rect -796 3001 -738 3013
rect -796 2425 -784 3001
rect -750 2425 -738 3001
rect -796 2413 -738 2425
rect -678 3001 -620 3013
rect -678 2425 -666 3001
rect -632 2425 -620 3001
rect -678 2413 -620 2425
rect -560 3001 -502 3013
rect -560 2425 -548 3001
rect -514 2425 -502 3001
rect -560 2413 -502 2425
rect -442 3001 -384 3013
rect -442 2425 -430 3001
rect -396 2425 -384 3001
rect -442 2413 -384 2425
rect -324 3001 -266 3013
rect -324 2425 -312 3001
rect -278 2425 -266 3001
rect -324 2413 -266 2425
rect -206 3001 -148 3013
rect -206 2425 -194 3001
rect -160 2425 -148 3001
rect -206 2413 -148 2425
rect -88 3001 -30 3013
rect -88 2425 -76 3001
rect -42 2425 -30 3001
rect -88 2413 -30 2425
rect 30 3001 88 3013
rect 30 2425 42 3001
rect 76 2425 88 3001
rect 30 2413 88 2425
rect 148 3001 206 3013
rect 148 2425 160 3001
rect 194 2425 206 3001
rect 148 2413 206 2425
rect 266 3001 324 3013
rect 266 2425 278 3001
rect 312 2425 324 3001
rect 266 2413 324 2425
rect 384 3001 442 3013
rect 384 2425 396 3001
rect 430 2425 442 3001
rect 384 2413 442 2425
rect 502 3001 560 3013
rect 502 2425 514 3001
rect 548 2425 560 3001
rect 502 2413 560 2425
rect 620 3001 678 3013
rect 620 2425 632 3001
rect 666 2425 678 3001
rect 620 2413 678 2425
rect 738 3001 796 3013
rect 738 2425 750 3001
rect 784 2425 796 3001
rect 738 2413 796 2425
rect 856 3001 914 3013
rect 856 2425 868 3001
rect 902 2425 914 3001
rect 856 2413 914 2425
rect 974 3001 1032 3013
rect 974 2425 986 3001
rect 1020 2425 1032 3001
rect 974 2413 1032 2425
rect 1092 3001 1150 3013
rect 1092 2425 1104 3001
rect 1138 2425 1150 3001
rect 1092 2413 1150 2425
rect 1210 3001 1268 3013
rect 1210 2425 1222 3001
rect 1256 2425 1268 3001
rect 1210 2413 1268 2425
rect 1328 3001 1386 3013
rect 1328 2425 1340 3001
rect 1374 2425 1386 3001
rect 1328 2413 1386 2425
rect 1446 3001 1504 3013
rect 1446 2425 1458 3001
rect 1492 2425 1504 3001
rect 1446 2413 1504 2425
rect -1504 2236 -1446 2248
rect -1504 1660 -1492 2236
rect -1458 1660 -1446 2236
rect -1504 1648 -1446 1660
rect -1386 2236 -1328 2248
rect -1386 1660 -1374 2236
rect -1340 1660 -1328 2236
rect -1386 1648 -1328 1660
rect -1268 2236 -1210 2248
rect -1268 1660 -1256 2236
rect -1222 1660 -1210 2236
rect -1268 1648 -1210 1660
rect -1150 2236 -1092 2248
rect -1150 1660 -1138 2236
rect -1104 1660 -1092 2236
rect -1150 1648 -1092 1660
rect -1032 2236 -974 2248
rect -1032 1660 -1020 2236
rect -986 1660 -974 2236
rect -1032 1648 -974 1660
rect -914 2236 -856 2248
rect -914 1660 -902 2236
rect -868 1660 -856 2236
rect -914 1648 -856 1660
rect -796 2236 -738 2248
rect -796 1660 -784 2236
rect -750 1660 -738 2236
rect -796 1648 -738 1660
rect -678 2236 -620 2248
rect -678 1660 -666 2236
rect -632 1660 -620 2236
rect -678 1648 -620 1660
rect -560 2236 -502 2248
rect -560 1660 -548 2236
rect -514 1660 -502 2236
rect -560 1648 -502 1660
rect -442 2236 -384 2248
rect -442 1660 -430 2236
rect -396 1660 -384 2236
rect -442 1648 -384 1660
rect -324 2236 -266 2248
rect -324 1660 -312 2236
rect -278 1660 -266 2236
rect -324 1648 -266 1660
rect -206 2236 -148 2248
rect -206 1660 -194 2236
rect -160 1660 -148 2236
rect -206 1648 -148 1660
rect -88 2236 -30 2248
rect -88 1660 -76 2236
rect -42 1660 -30 2236
rect -88 1648 -30 1660
rect 30 2236 88 2248
rect 30 1660 42 2236
rect 76 1660 88 2236
rect 30 1648 88 1660
rect 148 2236 206 2248
rect 148 1660 160 2236
rect 194 1660 206 2236
rect 148 1648 206 1660
rect 266 2236 324 2248
rect 266 1660 278 2236
rect 312 1660 324 2236
rect 266 1648 324 1660
rect 384 2236 442 2248
rect 384 1660 396 2236
rect 430 1660 442 2236
rect 384 1648 442 1660
rect 502 2236 560 2248
rect 502 1660 514 2236
rect 548 1660 560 2236
rect 502 1648 560 1660
rect 620 2236 678 2248
rect 620 1660 632 2236
rect 666 1660 678 2236
rect 620 1648 678 1660
rect 738 2236 796 2248
rect 738 1660 750 2236
rect 784 1660 796 2236
rect 738 1648 796 1660
rect 856 2236 914 2248
rect 856 1660 868 2236
rect 902 1660 914 2236
rect 856 1648 914 1660
rect 974 2236 1032 2248
rect 974 1660 986 2236
rect 1020 1660 1032 2236
rect 974 1648 1032 1660
rect 1092 2236 1150 2248
rect 1092 1660 1104 2236
rect 1138 1660 1150 2236
rect 1092 1648 1150 1660
rect 1210 2236 1268 2248
rect 1210 1660 1222 2236
rect 1256 1660 1268 2236
rect 1210 1648 1268 1660
rect 1328 2236 1386 2248
rect 1328 1660 1340 2236
rect 1374 1660 1386 2236
rect 1328 1648 1386 1660
rect 1446 2236 1504 2248
rect 1446 1660 1458 2236
rect 1492 1660 1504 2236
rect 1446 1648 1504 1660
rect -1504 1471 -1446 1483
rect -1504 895 -1492 1471
rect -1458 895 -1446 1471
rect -1504 883 -1446 895
rect -1386 1471 -1328 1483
rect -1386 895 -1374 1471
rect -1340 895 -1328 1471
rect -1386 883 -1328 895
rect -1268 1471 -1210 1483
rect -1268 895 -1256 1471
rect -1222 895 -1210 1471
rect -1268 883 -1210 895
rect -1150 1471 -1092 1483
rect -1150 895 -1138 1471
rect -1104 895 -1092 1471
rect -1150 883 -1092 895
rect -1032 1471 -974 1483
rect -1032 895 -1020 1471
rect -986 895 -974 1471
rect -1032 883 -974 895
rect -914 1471 -856 1483
rect -914 895 -902 1471
rect -868 895 -856 1471
rect -914 883 -856 895
rect -796 1471 -738 1483
rect -796 895 -784 1471
rect -750 895 -738 1471
rect -796 883 -738 895
rect -678 1471 -620 1483
rect -678 895 -666 1471
rect -632 895 -620 1471
rect -678 883 -620 895
rect -560 1471 -502 1483
rect -560 895 -548 1471
rect -514 895 -502 1471
rect -560 883 -502 895
rect -442 1471 -384 1483
rect -442 895 -430 1471
rect -396 895 -384 1471
rect -442 883 -384 895
rect -324 1471 -266 1483
rect -324 895 -312 1471
rect -278 895 -266 1471
rect -324 883 -266 895
rect -206 1471 -148 1483
rect -206 895 -194 1471
rect -160 895 -148 1471
rect -206 883 -148 895
rect -88 1471 -30 1483
rect -88 895 -76 1471
rect -42 895 -30 1471
rect -88 883 -30 895
rect 30 1471 88 1483
rect 30 895 42 1471
rect 76 895 88 1471
rect 30 883 88 895
rect 148 1471 206 1483
rect 148 895 160 1471
rect 194 895 206 1471
rect 148 883 206 895
rect 266 1471 324 1483
rect 266 895 278 1471
rect 312 895 324 1471
rect 266 883 324 895
rect 384 1471 442 1483
rect 384 895 396 1471
rect 430 895 442 1471
rect 384 883 442 895
rect 502 1471 560 1483
rect 502 895 514 1471
rect 548 895 560 1471
rect 502 883 560 895
rect 620 1471 678 1483
rect 620 895 632 1471
rect 666 895 678 1471
rect 620 883 678 895
rect 738 1471 796 1483
rect 738 895 750 1471
rect 784 895 796 1471
rect 738 883 796 895
rect 856 1471 914 1483
rect 856 895 868 1471
rect 902 895 914 1471
rect 856 883 914 895
rect 974 1471 1032 1483
rect 974 895 986 1471
rect 1020 895 1032 1471
rect 974 883 1032 895
rect 1092 1471 1150 1483
rect 1092 895 1104 1471
rect 1138 895 1150 1471
rect 1092 883 1150 895
rect 1210 1471 1268 1483
rect 1210 895 1222 1471
rect 1256 895 1268 1471
rect 1210 883 1268 895
rect 1328 1471 1386 1483
rect 1328 895 1340 1471
rect 1374 895 1386 1471
rect 1328 883 1386 895
rect 1446 1471 1504 1483
rect 1446 895 1458 1471
rect 1492 895 1504 1471
rect 1446 883 1504 895
rect -1504 706 -1446 718
rect -1504 130 -1492 706
rect -1458 130 -1446 706
rect -1504 118 -1446 130
rect -1386 706 -1328 718
rect -1386 130 -1374 706
rect -1340 130 -1328 706
rect -1386 118 -1328 130
rect -1268 706 -1210 718
rect -1268 130 -1256 706
rect -1222 130 -1210 706
rect -1268 118 -1210 130
rect -1150 706 -1092 718
rect -1150 130 -1138 706
rect -1104 130 -1092 706
rect -1150 118 -1092 130
rect -1032 706 -974 718
rect -1032 130 -1020 706
rect -986 130 -974 706
rect -1032 118 -974 130
rect -914 706 -856 718
rect -914 130 -902 706
rect -868 130 -856 706
rect -914 118 -856 130
rect -796 706 -738 718
rect -796 130 -784 706
rect -750 130 -738 706
rect -796 118 -738 130
rect -678 706 -620 718
rect -678 130 -666 706
rect -632 130 -620 706
rect -678 118 -620 130
rect -560 706 -502 718
rect -560 130 -548 706
rect -514 130 -502 706
rect -560 118 -502 130
rect -442 706 -384 718
rect -442 130 -430 706
rect -396 130 -384 706
rect -442 118 -384 130
rect -324 706 -266 718
rect -324 130 -312 706
rect -278 130 -266 706
rect -324 118 -266 130
rect -206 706 -148 718
rect -206 130 -194 706
rect -160 130 -148 706
rect -206 118 -148 130
rect -88 706 -30 718
rect -88 130 -76 706
rect -42 130 -30 706
rect -88 118 -30 130
rect 30 706 88 718
rect 30 130 42 706
rect 76 130 88 706
rect 30 118 88 130
rect 148 706 206 718
rect 148 130 160 706
rect 194 130 206 706
rect 148 118 206 130
rect 266 706 324 718
rect 266 130 278 706
rect 312 130 324 706
rect 266 118 324 130
rect 384 706 442 718
rect 384 130 396 706
rect 430 130 442 706
rect 384 118 442 130
rect 502 706 560 718
rect 502 130 514 706
rect 548 130 560 706
rect 502 118 560 130
rect 620 706 678 718
rect 620 130 632 706
rect 666 130 678 706
rect 620 118 678 130
rect 738 706 796 718
rect 738 130 750 706
rect 784 130 796 706
rect 738 118 796 130
rect 856 706 914 718
rect 856 130 868 706
rect 902 130 914 706
rect 856 118 914 130
rect 974 706 1032 718
rect 974 130 986 706
rect 1020 130 1032 706
rect 974 118 1032 130
rect 1092 706 1150 718
rect 1092 130 1104 706
rect 1138 130 1150 706
rect 1092 118 1150 130
rect 1210 706 1268 718
rect 1210 130 1222 706
rect 1256 130 1268 706
rect 1210 118 1268 130
rect 1328 706 1386 718
rect 1328 130 1340 706
rect 1374 130 1386 706
rect 1328 118 1386 130
rect 1446 706 1504 718
rect 1446 130 1458 706
rect 1492 130 1504 706
rect 1446 118 1504 130
rect -1504 -59 -1446 -47
rect -1504 -635 -1492 -59
rect -1458 -635 -1446 -59
rect -1504 -647 -1446 -635
rect -1386 -59 -1328 -47
rect -1386 -635 -1374 -59
rect -1340 -635 -1328 -59
rect -1386 -647 -1328 -635
rect -1268 -59 -1210 -47
rect -1268 -635 -1256 -59
rect -1222 -635 -1210 -59
rect -1268 -647 -1210 -635
rect -1150 -59 -1092 -47
rect -1150 -635 -1138 -59
rect -1104 -635 -1092 -59
rect -1150 -647 -1092 -635
rect -1032 -59 -974 -47
rect -1032 -635 -1020 -59
rect -986 -635 -974 -59
rect -1032 -647 -974 -635
rect -914 -59 -856 -47
rect -914 -635 -902 -59
rect -868 -635 -856 -59
rect -914 -647 -856 -635
rect -796 -59 -738 -47
rect -796 -635 -784 -59
rect -750 -635 -738 -59
rect -796 -647 -738 -635
rect -678 -59 -620 -47
rect -678 -635 -666 -59
rect -632 -635 -620 -59
rect -678 -647 -620 -635
rect -560 -59 -502 -47
rect -560 -635 -548 -59
rect -514 -635 -502 -59
rect -560 -647 -502 -635
rect -442 -59 -384 -47
rect -442 -635 -430 -59
rect -396 -635 -384 -59
rect -442 -647 -384 -635
rect -324 -59 -266 -47
rect -324 -635 -312 -59
rect -278 -635 -266 -59
rect -324 -647 -266 -635
rect -206 -59 -148 -47
rect -206 -635 -194 -59
rect -160 -635 -148 -59
rect -206 -647 -148 -635
rect -88 -59 -30 -47
rect -88 -635 -76 -59
rect -42 -635 -30 -59
rect -88 -647 -30 -635
rect 30 -59 88 -47
rect 30 -635 42 -59
rect 76 -635 88 -59
rect 30 -647 88 -635
rect 148 -59 206 -47
rect 148 -635 160 -59
rect 194 -635 206 -59
rect 148 -647 206 -635
rect 266 -59 324 -47
rect 266 -635 278 -59
rect 312 -635 324 -59
rect 266 -647 324 -635
rect 384 -59 442 -47
rect 384 -635 396 -59
rect 430 -635 442 -59
rect 384 -647 442 -635
rect 502 -59 560 -47
rect 502 -635 514 -59
rect 548 -635 560 -59
rect 502 -647 560 -635
rect 620 -59 678 -47
rect 620 -635 632 -59
rect 666 -635 678 -59
rect 620 -647 678 -635
rect 738 -59 796 -47
rect 738 -635 750 -59
rect 784 -635 796 -59
rect 738 -647 796 -635
rect 856 -59 914 -47
rect 856 -635 868 -59
rect 902 -635 914 -59
rect 856 -647 914 -635
rect 974 -59 1032 -47
rect 974 -635 986 -59
rect 1020 -635 1032 -59
rect 974 -647 1032 -635
rect 1092 -59 1150 -47
rect 1092 -635 1104 -59
rect 1138 -635 1150 -59
rect 1092 -647 1150 -635
rect 1210 -59 1268 -47
rect 1210 -635 1222 -59
rect 1256 -635 1268 -59
rect 1210 -647 1268 -635
rect 1328 -59 1386 -47
rect 1328 -635 1340 -59
rect 1374 -635 1386 -59
rect 1328 -647 1386 -635
rect 1446 -59 1504 -47
rect 1446 -635 1458 -59
rect 1492 -635 1504 -59
rect 1446 -647 1504 -635
rect -1504 -824 -1446 -812
rect -1504 -1400 -1492 -824
rect -1458 -1400 -1446 -824
rect -1504 -1412 -1446 -1400
rect -1386 -824 -1328 -812
rect -1386 -1400 -1374 -824
rect -1340 -1400 -1328 -824
rect -1386 -1412 -1328 -1400
rect -1268 -824 -1210 -812
rect -1268 -1400 -1256 -824
rect -1222 -1400 -1210 -824
rect -1268 -1412 -1210 -1400
rect -1150 -824 -1092 -812
rect -1150 -1400 -1138 -824
rect -1104 -1400 -1092 -824
rect -1150 -1412 -1092 -1400
rect -1032 -824 -974 -812
rect -1032 -1400 -1020 -824
rect -986 -1400 -974 -824
rect -1032 -1412 -974 -1400
rect -914 -824 -856 -812
rect -914 -1400 -902 -824
rect -868 -1400 -856 -824
rect -914 -1412 -856 -1400
rect -796 -824 -738 -812
rect -796 -1400 -784 -824
rect -750 -1400 -738 -824
rect -796 -1412 -738 -1400
rect -678 -824 -620 -812
rect -678 -1400 -666 -824
rect -632 -1400 -620 -824
rect -678 -1412 -620 -1400
rect -560 -824 -502 -812
rect -560 -1400 -548 -824
rect -514 -1400 -502 -824
rect -560 -1412 -502 -1400
rect -442 -824 -384 -812
rect -442 -1400 -430 -824
rect -396 -1400 -384 -824
rect -442 -1412 -384 -1400
rect -324 -824 -266 -812
rect -324 -1400 -312 -824
rect -278 -1400 -266 -824
rect -324 -1412 -266 -1400
rect -206 -824 -148 -812
rect -206 -1400 -194 -824
rect -160 -1400 -148 -824
rect -206 -1412 -148 -1400
rect -88 -824 -30 -812
rect -88 -1400 -76 -824
rect -42 -1400 -30 -824
rect -88 -1412 -30 -1400
rect 30 -824 88 -812
rect 30 -1400 42 -824
rect 76 -1400 88 -824
rect 30 -1412 88 -1400
rect 148 -824 206 -812
rect 148 -1400 160 -824
rect 194 -1400 206 -824
rect 148 -1412 206 -1400
rect 266 -824 324 -812
rect 266 -1400 278 -824
rect 312 -1400 324 -824
rect 266 -1412 324 -1400
rect 384 -824 442 -812
rect 384 -1400 396 -824
rect 430 -1400 442 -824
rect 384 -1412 442 -1400
rect 502 -824 560 -812
rect 502 -1400 514 -824
rect 548 -1400 560 -824
rect 502 -1412 560 -1400
rect 620 -824 678 -812
rect 620 -1400 632 -824
rect 666 -1400 678 -824
rect 620 -1412 678 -1400
rect 738 -824 796 -812
rect 738 -1400 750 -824
rect 784 -1400 796 -824
rect 738 -1412 796 -1400
rect 856 -824 914 -812
rect 856 -1400 868 -824
rect 902 -1400 914 -824
rect 856 -1412 914 -1400
rect 974 -824 1032 -812
rect 974 -1400 986 -824
rect 1020 -1400 1032 -824
rect 974 -1412 1032 -1400
rect 1092 -824 1150 -812
rect 1092 -1400 1104 -824
rect 1138 -1400 1150 -824
rect 1092 -1412 1150 -1400
rect 1210 -824 1268 -812
rect 1210 -1400 1222 -824
rect 1256 -1400 1268 -824
rect 1210 -1412 1268 -1400
rect 1328 -824 1386 -812
rect 1328 -1400 1340 -824
rect 1374 -1400 1386 -824
rect 1328 -1412 1386 -1400
rect 1446 -824 1504 -812
rect 1446 -1400 1458 -824
rect 1492 -1400 1504 -824
rect 1446 -1412 1504 -1400
rect -1504 -1589 -1446 -1577
rect -1504 -2165 -1492 -1589
rect -1458 -2165 -1446 -1589
rect -1504 -2177 -1446 -2165
rect -1386 -1589 -1328 -1577
rect -1386 -2165 -1374 -1589
rect -1340 -2165 -1328 -1589
rect -1386 -2177 -1328 -2165
rect -1268 -1589 -1210 -1577
rect -1268 -2165 -1256 -1589
rect -1222 -2165 -1210 -1589
rect -1268 -2177 -1210 -2165
rect -1150 -1589 -1092 -1577
rect -1150 -2165 -1138 -1589
rect -1104 -2165 -1092 -1589
rect -1150 -2177 -1092 -2165
rect -1032 -1589 -974 -1577
rect -1032 -2165 -1020 -1589
rect -986 -2165 -974 -1589
rect -1032 -2177 -974 -2165
rect -914 -1589 -856 -1577
rect -914 -2165 -902 -1589
rect -868 -2165 -856 -1589
rect -914 -2177 -856 -2165
rect -796 -1589 -738 -1577
rect -796 -2165 -784 -1589
rect -750 -2165 -738 -1589
rect -796 -2177 -738 -2165
rect -678 -1589 -620 -1577
rect -678 -2165 -666 -1589
rect -632 -2165 -620 -1589
rect -678 -2177 -620 -2165
rect -560 -1589 -502 -1577
rect -560 -2165 -548 -1589
rect -514 -2165 -502 -1589
rect -560 -2177 -502 -2165
rect -442 -1589 -384 -1577
rect -442 -2165 -430 -1589
rect -396 -2165 -384 -1589
rect -442 -2177 -384 -2165
rect -324 -1589 -266 -1577
rect -324 -2165 -312 -1589
rect -278 -2165 -266 -1589
rect -324 -2177 -266 -2165
rect -206 -1589 -148 -1577
rect -206 -2165 -194 -1589
rect -160 -2165 -148 -1589
rect -206 -2177 -148 -2165
rect -88 -1589 -30 -1577
rect -88 -2165 -76 -1589
rect -42 -2165 -30 -1589
rect -88 -2177 -30 -2165
rect 30 -1589 88 -1577
rect 30 -2165 42 -1589
rect 76 -2165 88 -1589
rect 30 -2177 88 -2165
rect 148 -1589 206 -1577
rect 148 -2165 160 -1589
rect 194 -2165 206 -1589
rect 148 -2177 206 -2165
rect 266 -1589 324 -1577
rect 266 -2165 278 -1589
rect 312 -2165 324 -1589
rect 266 -2177 324 -2165
rect 384 -1589 442 -1577
rect 384 -2165 396 -1589
rect 430 -2165 442 -1589
rect 384 -2177 442 -2165
rect 502 -1589 560 -1577
rect 502 -2165 514 -1589
rect 548 -2165 560 -1589
rect 502 -2177 560 -2165
rect 620 -1589 678 -1577
rect 620 -2165 632 -1589
rect 666 -2165 678 -1589
rect 620 -2177 678 -2165
rect 738 -1589 796 -1577
rect 738 -2165 750 -1589
rect 784 -2165 796 -1589
rect 738 -2177 796 -2165
rect 856 -1589 914 -1577
rect 856 -2165 868 -1589
rect 902 -2165 914 -1589
rect 856 -2177 914 -2165
rect 974 -1589 1032 -1577
rect 974 -2165 986 -1589
rect 1020 -2165 1032 -1589
rect 974 -2177 1032 -2165
rect 1092 -1589 1150 -1577
rect 1092 -2165 1104 -1589
rect 1138 -2165 1150 -1589
rect 1092 -2177 1150 -2165
rect 1210 -1589 1268 -1577
rect 1210 -2165 1222 -1589
rect 1256 -2165 1268 -1589
rect 1210 -2177 1268 -2165
rect 1328 -1589 1386 -1577
rect 1328 -2165 1340 -1589
rect 1374 -2165 1386 -1589
rect 1328 -2177 1386 -2165
rect 1446 -1589 1504 -1577
rect 1446 -2165 1458 -1589
rect 1492 -2165 1504 -1589
rect 1446 -2177 1504 -2165
rect -1504 -2354 -1446 -2342
rect -1504 -2930 -1492 -2354
rect -1458 -2930 -1446 -2354
rect -1504 -2942 -1446 -2930
rect -1386 -2354 -1328 -2342
rect -1386 -2930 -1374 -2354
rect -1340 -2930 -1328 -2354
rect -1386 -2942 -1328 -2930
rect -1268 -2354 -1210 -2342
rect -1268 -2930 -1256 -2354
rect -1222 -2930 -1210 -2354
rect -1268 -2942 -1210 -2930
rect -1150 -2354 -1092 -2342
rect -1150 -2930 -1138 -2354
rect -1104 -2930 -1092 -2354
rect -1150 -2942 -1092 -2930
rect -1032 -2354 -974 -2342
rect -1032 -2930 -1020 -2354
rect -986 -2930 -974 -2354
rect -1032 -2942 -974 -2930
rect -914 -2354 -856 -2342
rect -914 -2930 -902 -2354
rect -868 -2930 -856 -2354
rect -914 -2942 -856 -2930
rect -796 -2354 -738 -2342
rect -796 -2930 -784 -2354
rect -750 -2930 -738 -2354
rect -796 -2942 -738 -2930
rect -678 -2354 -620 -2342
rect -678 -2930 -666 -2354
rect -632 -2930 -620 -2354
rect -678 -2942 -620 -2930
rect -560 -2354 -502 -2342
rect -560 -2930 -548 -2354
rect -514 -2930 -502 -2354
rect -560 -2942 -502 -2930
rect -442 -2354 -384 -2342
rect -442 -2930 -430 -2354
rect -396 -2930 -384 -2354
rect -442 -2942 -384 -2930
rect -324 -2354 -266 -2342
rect -324 -2930 -312 -2354
rect -278 -2930 -266 -2354
rect -324 -2942 -266 -2930
rect -206 -2354 -148 -2342
rect -206 -2930 -194 -2354
rect -160 -2930 -148 -2354
rect -206 -2942 -148 -2930
rect -88 -2354 -30 -2342
rect -88 -2930 -76 -2354
rect -42 -2930 -30 -2354
rect -88 -2942 -30 -2930
rect 30 -2354 88 -2342
rect 30 -2930 42 -2354
rect 76 -2930 88 -2354
rect 30 -2942 88 -2930
rect 148 -2354 206 -2342
rect 148 -2930 160 -2354
rect 194 -2930 206 -2354
rect 148 -2942 206 -2930
rect 266 -2354 324 -2342
rect 266 -2930 278 -2354
rect 312 -2930 324 -2354
rect 266 -2942 324 -2930
rect 384 -2354 442 -2342
rect 384 -2930 396 -2354
rect 430 -2930 442 -2354
rect 384 -2942 442 -2930
rect 502 -2354 560 -2342
rect 502 -2930 514 -2354
rect 548 -2930 560 -2354
rect 502 -2942 560 -2930
rect 620 -2354 678 -2342
rect 620 -2930 632 -2354
rect 666 -2930 678 -2354
rect 620 -2942 678 -2930
rect 738 -2354 796 -2342
rect 738 -2930 750 -2354
rect 784 -2930 796 -2354
rect 738 -2942 796 -2930
rect 856 -2354 914 -2342
rect 856 -2930 868 -2354
rect 902 -2930 914 -2354
rect 856 -2942 914 -2930
rect 974 -2354 1032 -2342
rect 974 -2930 986 -2354
rect 1020 -2930 1032 -2354
rect 974 -2942 1032 -2930
rect 1092 -2354 1150 -2342
rect 1092 -2930 1104 -2354
rect 1138 -2930 1150 -2354
rect 1092 -2942 1150 -2930
rect 1210 -2354 1268 -2342
rect 1210 -2930 1222 -2354
rect 1256 -2930 1268 -2354
rect 1210 -2942 1268 -2930
rect 1328 -2354 1386 -2342
rect 1328 -2930 1340 -2354
rect 1374 -2930 1386 -2354
rect 1328 -2942 1386 -2930
rect 1446 -2354 1504 -2342
rect 1446 -2930 1458 -2354
rect 1492 -2930 1504 -2354
rect 1446 -2942 1504 -2930
rect -1504 -3119 -1446 -3107
rect -1504 -3695 -1492 -3119
rect -1458 -3695 -1446 -3119
rect -1504 -3707 -1446 -3695
rect -1386 -3119 -1328 -3107
rect -1386 -3695 -1374 -3119
rect -1340 -3695 -1328 -3119
rect -1386 -3707 -1328 -3695
rect -1268 -3119 -1210 -3107
rect -1268 -3695 -1256 -3119
rect -1222 -3695 -1210 -3119
rect -1268 -3707 -1210 -3695
rect -1150 -3119 -1092 -3107
rect -1150 -3695 -1138 -3119
rect -1104 -3695 -1092 -3119
rect -1150 -3707 -1092 -3695
rect -1032 -3119 -974 -3107
rect -1032 -3695 -1020 -3119
rect -986 -3695 -974 -3119
rect -1032 -3707 -974 -3695
rect -914 -3119 -856 -3107
rect -914 -3695 -902 -3119
rect -868 -3695 -856 -3119
rect -914 -3707 -856 -3695
rect -796 -3119 -738 -3107
rect -796 -3695 -784 -3119
rect -750 -3695 -738 -3119
rect -796 -3707 -738 -3695
rect -678 -3119 -620 -3107
rect -678 -3695 -666 -3119
rect -632 -3695 -620 -3119
rect -678 -3707 -620 -3695
rect -560 -3119 -502 -3107
rect -560 -3695 -548 -3119
rect -514 -3695 -502 -3119
rect -560 -3707 -502 -3695
rect -442 -3119 -384 -3107
rect -442 -3695 -430 -3119
rect -396 -3695 -384 -3119
rect -442 -3707 -384 -3695
rect -324 -3119 -266 -3107
rect -324 -3695 -312 -3119
rect -278 -3695 -266 -3119
rect -324 -3707 -266 -3695
rect -206 -3119 -148 -3107
rect -206 -3695 -194 -3119
rect -160 -3695 -148 -3119
rect -206 -3707 -148 -3695
rect -88 -3119 -30 -3107
rect -88 -3695 -76 -3119
rect -42 -3695 -30 -3119
rect -88 -3707 -30 -3695
rect 30 -3119 88 -3107
rect 30 -3695 42 -3119
rect 76 -3695 88 -3119
rect 30 -3707 88 -3695
rect 148 -3119 206 -3107
rect 148 -3695 160 -3119
rect 194 -3695 206 -3119
rect 148 -3707 206 -3695
rect 266 -3119 324 -3107
rect 266 -3695 278 -3119
rect 312 -3695 324 -3119
rect 266 -3707 324 -3695
rect 384 -3119 442 -3107
rect 384 -3695 396 -3119
rect 430 -3695 442 -3119
rect 384 -3707 442 -3695
rect 502 -3119 560 -3107
rect 502 -3695 514 -3119
rect 548 -3695 560 -3119
rect 502 -3707 560 -3695
rect 620 -3119 678 -3107
rect 620 -3695 632 -3119
rect 666 -3695 678 -3119
rect 620 -3707 678 -3695
rect 738 -3119 796 -3107
rect 738 -3695 750 -3119
rect 784 -3695 796 -3119
rect 738 -3707 796 -3695
rect 856 -3119 914 -3107
rect 856 -3695 868 -3119
rect 902 -3695 914 -3119
rect 856 -3707 914 -3695
rect 974 -3119 1032 -3107
rect 974 -3695 986 -3119
rect 1020 -3695 1032 -3119
rect 974 -3707 1032 -3695
rect 1092 -3119 1150 -3107
rect 1092 -3695 1104 -3119
rect 1138 -3695 1150 -3119
rect 1092 -3707 1150 -3695
rect 1210 -3119 1268 -3107
rect 1210 -3695 1222 -3119
rect 1256 -3695 1268 -3119
rect 1210 -3707 1268 -3695
rect 1328 -3119 1386 -3107
rect 1328 -3695 1340 -3119
rect 1374 -3695 1386 -3119
rect 1328 -3707 1386 -3695
rect 1446 -3119 1504 -3107
rect 1446 -3695 1458 -3119
rect 1492 -3695 1504 -3119
rect 1446 -3707 1504 -3695
<< pdiffc >>
rect -1492 3190 -1458 3766
rect -1374 3190 -1340 3766
rect -1256 3190 -1222 3766
rect -1138 3190 -1104 3766
rect -1020 3190 -986 3766
rect -902 3190 -868 3766
rect -784 3190 -750 3766
rect -666 3190 -632 3766
rect -548 3190 -514 3766
rect -430 3190 -396 3766
rect -312 3190 -278 3766
rect -194 3190 -160 3766
rect -76 3190 -42 3766
rect 42 3190 76 3766
rect 160 3190 194 3766
rect 278 3190 312 3766
rect 396 3190 430 3766
rect 514 3190 548 3766
rect 632 3190 666 3766
rect 750 3190 784 3766
rect 868 3190 902 3766
rect 986 3190 1020 3766
rect 1104 3190 1138 3766
rect 1222 3190 1256 3766
rect 1340 3190 1374 3766
rect 1458 3190 1492 3766
rect -1492 2425 -1458 3001
rect -1374 2425 -1340 3001
rect -1256 2425 -1222 3001
rect -1138 2425 -1104 3001
rect -1020 2425 -986 3001
rect -902 2425 -868 3001
rect -784 2425 -750 3001
rect -666 2425 -632 3001
rect -548 2425 -514 3001
rect -430 2425 -396 3001
rect -312 2425 -278 3001
rect -194 2425 -160 3001
rect -76 2425 -42 3001
rect 42 2425 76 3001
rect 160 2425 194 3001
rect 278 2425 312 3001
rect 396 2425 430 3001
rect 514 2425 548 3001
rect 632 2425 666 3001
rect 750 2425 784 3001
rect 868 2425 902 3001
rect 986 2425 1020 3001
rect 1104 2425 1138 3001
rect 1222 2425 1256 3001
rect 1340 2425 1374 3001
rect 1458 2425 1492 3001
rect -1492 1660 -1458 2236
rect -1374 1660 -1340 2236
rect -1256 1660 -1222 2236
rect -1138 1660 -1104 2236
rect -1020 1660 -986 2236
rect -902 1660 -868 2236
rect -784 1660 -750 2236
rect -666 1660 -632 2236
rect -548 1660 -514 2236
rect -430 1660 -396 2236
rect -312 1660 -278 2236
rect -194 1660 -160 2236
rect -76 1660 -42 2236
rect 42 1660 76 2236
rect 160 1660 194 2236
rect 278 1660 312 2236
rect 396 1660 430 2236
rect 514 1660 548 2236
rect 632 1660 666 2236
rect 750 1660 784 2236
rect 868 1660 902 2236
rect 986 1660 1020 2236
rect 1104 1660 1138 2236
rect 1222 1660 1256 2236
rect 1340 1660 1374 2236
rect 1458 1660 1492 2236
rect -1492 895 -1458 1471
rect -1374 895 -1340 1471
rect -1256 895 -1222 1471
rect -1138 895 -1104 1471
rect -1020 895 -986 1471
rect -902 895 -868 1471
rect -784 895 -750 1471
rect -666 895 -632 1471
rect -548 895 -514 1471
rect -430 895 -396 1471
rect -312 895 -278 1471
rect -194 895 -160 1471
rect -76 895 -42 1471
rect 42 895 76 1471
rect 160 895 194 1471
rect 278 895 312 1471
rect 396 895 430 1471
rect 514 895 548 1471
rect 632 895 666 1471
rect 750 895 784 1471
rect 868 895 902 1471
rect 986 895 1020 1471
rect 1104 895 1138 1471
rect 1222 895 1256 1471
rect 1340 895 1374 1471
rect 1458 895 1492 1471
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect -1492 -635 -1458 -59
rect -1374 -635 -1340 -59
rect -1256 -635 -1222 -59
rect -1138 -635 -1104 -59
rect -1020 -635 -986 -59
rect -902 -635 -868 -59
rect -784 -635 -750 -59
rect -666 -635 -632 -59
rect -548 -635 -514 -59
rect -430 -635 -396 -59
rect -312 -635 -278 -59
rect -194 -635 -160 -59
rect -76 -635 -42 -59
rect 42 -635 76 -59
rect 160 -635 194 -59
rect 278 -635 312 -59
rect 396 -635 430 -59
rect 514 -635 548 -59
rect 632 -635 666 -59
rect 750 -635 784 -59
rect 868 -635 902 -59
rect 986 -635 1020 -59
rect 1104 -635 1138 -59
rect 1222 -635 1256 -59
rect 1340 -635 1374 -59
rect 1458 -635 1492 -59
rect -1492 -1400 -1458 -824
rect -1374 -1400 -1340 -824
rect -1256 -1400 -1222 -824
rect -1138 -1400 -1104 -824
rect -1020 -1400 -986 -824
rect -902 -1400 -868 -824
rect -784 -1400 -750 -824
rect -666 -1400 -632 -824
rect -548 -1400 -514 -824
rect -430 -1400 -396 -824
rect -312 -1400 -278 -824
rect -194 -1400 -160 -824
rect -76 -1400 -42 -824
rect 42 -1400 76 -824
rect 160 -1400 194 -824
rect 278 -1400 312 -824
rect 396 -1400 430 -824
rect 514 -1400 548 -824
rect 632 -1400 666 -824
rect 750 -1400 784 -824
rect 868 -1400 902 -824
rect 986 -1400 1020 -824
rect 1104 -1400 1138 -824
rect 1222 -1400 1256 -824
rect 1340 -1400 1374 -824
rect 1458 -1400 1492 -824
rect -1492 -2165 -1458 -1589
rect -1374 -2165 -1340 -1589
rect -1256 -2165 -1222 -1589
rect -1138 -2165 -1104 -1589
rect -1020 -2165 -986 -1589
rect -902 -2165 -868 -1589
rect -784 -2165 -750 -1589
rect -666 -2165 -632 -1589
rect -548 -2165 -514 -1589
rect -430 -2165 -396 -1589
rect -312 -2165 -278 -1589
rect -194 -2165 -160 -1589
rect -76 -2165 -42 -1589
rect 42 -2165 76 -1589
rect 160 -2165 194 -1589
rect 278 -2165 312 -1589
rect 396 -2165 430 -1589
rect 514 -2165 548 -1589
rect 632 -2165 666 -1589
rect 750 -2165 784 -1589
rect 868 -2165 902 -1589
rect 986 -2165 1020 -1589
rect 1104 -2165 1138 -1589
rect 1222 -2165 1256 -1589
rect 1340 -2165 1374 -1589
rect 1458 -2165 1492 -1589
rect -1492 -2930 -1458 -2354
rect -1374 -2930 -1340 -2354
rect -1256 -2930 -1222 -2354
rect -1138 -2930 -1104 -2354
rect -1020 -2930 -986 -2354
rect -902 -2930 -868 -2354
rect -784 -2930 -750 -2354
rect -666 -2930 -632 -2354
rect -548 -2930 -514 -2354
rect -430 -2930 -396 -2354
rect -312 -2930 -278 -2354
rect -194 -2930 -160 -2354
rect -76 -2930 -42 -2354
rect 42 -2930 76 -2354
rect 160 -2930 194 -2354
rect 278 -2930 312 -2354
rect 396 -2930 430 -2354
rect 514 -2930 548 -2354
rect 632 -2930 666 -2354
rect 750 -2930 784 -2354
rect 868 -2930 902 -2354
rect 986 -2930 1020 -2354
rect 1104 -2930 1138 -2354
rect 1222 -2930 1256 -2354
rect 1340 -2930 1374 -2354
rect 1458 -2930 1492 -2354
rect -1492 -3695 -1458 -3119
rect -1374 -3695 -1340 -3119
rect -1256 -3695 -1222 -3119
rect -1138 -3695 -1104 -3119
rect -1020 -3695 -986 -3119
rect -902 -3695 -868 -3119
rect -784 -3695 -750 -3119
rect -666 -3695 -632 -3119
rect -548 -3695 -514 -3119
rect -430 -3695 -396 -3119
rect -312 -3695 -278 -3119
rect -194 -3695 -160 -3119
rect -76 -3695 -42 -3119
rect 42 -3695 76 -3119
rect 160 -3695 194 -3119
rect 278 -3695 312 -3119
rect 396 -3695 430 -3119
rect 514 -3695 548 -3119
rect 632 -3695 666 -3119
rect 750 -3695 784 -3119
rect 868 -3695 902 -3119
rect 986 -3695 1020 -3119
rect 1104 -3695 1138 -3119
rect 1222 -3695 1256 -3119
rect 1340 -3695 1374 -3119
rect 1458 -3695 1492 -3119
<< nsubdiff >>
rect -1606 3856 -1510 3890
rect 1510 3856 1606 3890
rect -1606 3794 -1572 3856
rect 1572 3794 1606 3856
rect -1606 -3856 -1572 -3794
rect 1572 -3856 1606 -3794
rect -1606 -3890 -1510 -3856
rect 1510 -3890 1606 -3856
<< nsubdiffcont >>
rect -1510 3856 1510 3890
rect -1606 -3794 -1572 3794
rect 1572 -3794 1606 3794
rect -1510 -3890 1510 -3856
<< poly >>
rect -1446 3778 -1386 3804
rect -1328 3778 -1268 3804
rect -1210 3778 -1150 3804
rect -1092 3778 -1032 3804
rect -974 3778 -914 3804
rect -856 3778 -796 3804
rect -738 3778 -678 3804
rect -620 3778 -560 3804
rect -502 3778 -442 3804
rect -384 3778 -324 3804
rect -266 3778 -206 3804
rect -148 3778 -88 3804
rect -30 3778 30 3804
rect 88 3778 148 3804
rect 206 3778 266 3804
rect 324 3778 384 3804
rect 442 3778 502 3804
rect 560 3778 620 3804
rect 678 3778 738 3804
rect 796 3778 856 3804
rect 914 3778 974 3804
rect 1032 3778 1092 3804
rect 1150 3778 1210 3804
rect 1268 3778 1328 3804
rect 1386 3778 1446 3804
rect -1446 3147 -1386 3178
rect -1328 3147 -1268 3178
rect -1210 3147 -1150 3178
rect -1092 3147 -1032 3178
rect -974 3147 -914 3178
rect -856 3147 -796 3178
rect -738 3147 -678 3178
rect -620 3147 -560 3178
rect -502 3147 -442 3178
rect -384 3147 -324 3178
rect -266 3147 -206 3178
rect -148 3147 -88 3178
rect -30 3147 30 3178
rect 88 3147 148 3178
rect 206 3147 266 3178
rect 324 3147 384 3178
rect 442 3147 502 3178
rect 560 3147 620 3178
rect 678 3147 738 3178
rect 796 3147 856 3178
rect 914 3147 974 3178
rect 1032 3147 1092 3178
rect 1150 3147 1210 3178
rect 1268 3147 1328 3178
rect 1386 3147 1446 3178
rect -1449 3131 -1383 3147
rect -1449 3097 -1433 3131
rect -1399 3097 -1383 3131
rect -1449 3081 -1383 3097
rect -1331 3131 -1265 3147
rect -1331 3097 -1315 3131
rect -1281 3097 -1265 3131
rect -1331 3081 -1265 3097
rect -1213 3131 -1147 3147
rect -1213 3097 -1197 3131
rect -1163 3097 -1147 3131
rect -1213 3081 -1147 3097
rect -1095 3131 -1029 3147
rect -1095 3097 -1079 3131
rect -1045 3097 -1029 3131
rect -1095 3081 -1029 3097
rect -977 3131 -911 3147
rect -977 3097 -961 3131
rect -927 3097 -911 3131
rect -977 3081 -911 3097
rect -859 3131 -793 3147
rect -859 3097 -843 3131
rect -809 3097 -793 3131
rect -859 3081 -793 3097
rect -741 3131 -675 3147
rect -741 3097 -725 3131
rect -691 3097 -675 3131
rect -741 3081 -675 3097
rect -623 3131 -557 3147
rect -623 3097 -607 3131
rect -573 3097 -557 3131
rect -623 3081 -557 3097
rect -505 3131 -439 3147
rect -505 3097 -489 3131
rect -455 3097 -439 3131
rect -505 3081 -439 3097
rect -387 3131 -321 3147
rect -387 3097 -371 3131
rect -337 3097 -321 3131
rect -387 3081 -321 3097
rect -269 3131 -203 3147
rect -269 3097 -253 3131
rect -219 3097 -203 3131
rect -269 3081 -203 3097
rect -151 3131 -85 3147
rect -151 3097 -135 3131
rect -101 3097 -85 3131
rect -151 3081 -85 3097
rect -33 3131 33 3147
rect -33 3097 -17 3131
rect 17 3097 33 3131
rect -33 3081 33 3097
rect 85 3131 151 3147
rect 85 3097 101 3131
rect 135 3097 151 3131
rect 85 3081 151 3097
rect 203 3131 269 3147
rect 203 3097 219 3131
rect 253 3097 269 3131
rect 203 3081 269 3097
rect 321 3131 387 3147
rect 321 3097 337 3131
rect 371 3097 387 3131
rect 321 3081 387 3097
rect 439 3131 505 3147
rect 439 3097 455 3131
rect 489 3097 505 3131
rect 439 3081 505 3097
rect 557 3131 623 3147
rect 557 3097 573 3131
rect 607 3097 623 3131
rect 557 3081 623 3097
rect 675 3131 741 3147
rect 675 3097 691 3131
rect 725 3097 741 3131
rect 675 3081 741 3097
rect 793 3131 859 3147
rect 793 3097 809 3131
rect 843 3097 859 3131
rect 793 3081 859 3097
rect 911 3131 977 3147
rect 911 3097 927 3131
rect 961 3097 977 3131
rect 911 3081 977 3097
rect 1029 3131 1095 3147
rect 1029 3097 1045 3131
rect 1079 3097 1095 3131
rect 1029 3081 1095 3097
rect 1147 3131 1213 3147
rect 1147 3097 1163 3131
rect 1197 3097 1213 3131
rect 1147 3081 1213 3097
rect 1265 3131 1331 3147
rect 1265 3097 1281 3131
rect 1315 3097 1331 3131
rect 1265 3081 1331 3097
rect 1383 3131 1449 3147
rect 1383 3097 1399 3131
rect 1433 3097 1449 3131
rect 1383 3081 1449 3097
rect -1446 3013 -1386 3039
rect -1328 3013 -1268 3039
rect -1210 3013 -1150 3039
rect -1092 3013 -1032 3039
rect -974 3013 -914 3039
rect -856 3013 -796 3039
rect -738 3013 -678 3039
rect -620 3013 -560 3039
rect -502 3013 -442 3039
rect -384 3013 -324 3039
rect -266 3013 -206 3039
rect -148 3013 -88 3039
rect -30 3013 30 3039
rect 88 3013 148 3039
rect 206 3013 266 3039
rect 324 3013 384 3039
rect 442 3013 502 3039
rect 560 3013 620 3039
rect 678 3013 738 3039
rect 796 3013 856 3039
rect 914 3013 974 3039
rect 1032 3013 1092 3039
rect 1150 3013 1210 3039
rect 1268 3013 1328 3039
rect 1386 3013 1446 3039
rect -1446 2382 -1386 2413
rect -1328 2382 -1268 2413
rect -1210 2382 -1150 2413
rect -1092 2382 -1032 2413
rect -974 2382 -914 2413
rect -856 2382 -796 2413
rect -738 2382 -678 2413
rect -620 2382 -560 2413
rect -502 2382 -442 2413
rect -384 2382 -324 2413
rect -266 2382 -206 2413
rect -148 2382 -88 2413
rect -30 2382 30 2413
rect 88 2382 148 2413
rect 206 2382 266 2413
rect 324 2382 384 2413
rect 442 2382 502 2413
rect 560 2382 620 2413
rect 678 2382 738 2413
rect 796 2382 856 2413
rect 914 2382 974 2413
rect 1032 2382 1092 2413
rect 1150 2382 1210 2413
rect 1268 2382 1328 2413
rect 1386 2382 1446 2413
rect -1449 2366 -1383 2382
rect -1449 2332 -1433 2366
rect -1399 2332 -1383 2366
rect -1449 2316 -1383 2332
rect -1331 2366 -1265 2382
rect -1331 2332 -1315 2366
rect -1281 2332 -1265 2366
rect -1331 2316 -1265 2332
rect -1213 2366 -1147 2382
rect -1213 2332 -1197 2366
rect -1163 2332 -1147 2366
rect -1213 2316 -1147 2332
rect -1095 2366 -1029 2382
rect -1095 2332 -1079 2366
rect -1045 2332 -1029 2366
rect -1095 2316 -1029 2332
rect -977 2366 -911 2382
rect -977 2332 -961 2366
rect -927 2332 -911 2366
rect -977 2316 -911 2332
rect -859 2366 -793 2382
rect -859 2332 -843 2366
rect -809 2332 -793 2366
rect -859 2316 -793 2332
rect -741 2366 -675 2382
rect -741 2332 -725 2366
rect -691 2332 -675 2366
rect -741 2316 -675 2332
rect -623 2366 -557 2382
rect -623 2332 -607 2366
rect -573 2332 -557 2366
rect -623 2316 -557 2332
rect -505 2366 -439 2382
rect -505 2332 -489 2366
rect -455 2332 -439 2366
rect -505 2316 -439 2332
rect -387 2366 -321 2382
rect -387 2332 -371 2366
rect -337 2332 -321 2366
rect -387 2316 -321 2332
rect -269 2366 -203 2382
rect -269 2332 -253 2366
rect -219 2332 -203 2366
rect -269 2316 -203 2332
rect -151 2366 -85 2382
rect -151 2332 -135 2366
rect -101 2332 -85 2366
rect -151 2316 -85 2332
rect -33 2366 33 2382
rect -33 2332 -17 2366
rect 17 2332 33 2366
rect -33 2316 33 2332
rect 85 2366 151 2382
rect 85 2332 101 2366
rect 135 2332 151 2366
rect 85 2316 151 2332
rect 203 2366 269 2382
rect 203 2332 219 2366
rect 253 2332 269 2366
rect 203 2316 269 2332
rect 321 2366 387 2382
rect 321 2332 337 2366
rect 371 2332 387 2366
rect 321 2316 387 2332
rect 439 2366 505 2382
rect 439 2332 455 2366
rect 489 2332 505 2366
rect 439 2316 505 2332
rect 557 2366 623 2382
rect 557 2332 573 2366
rect 607 2332 623 2366
rect 557 2316 623 2332
rect 675 2366 741 2382
rect 675 2332 691 2366
rect 725 2332 741 2366
rect 675 2316 741 2332
rect 793 2366 859 2382
rect 793 2332 809 2366
rect 843 2332 859 2366
rect 793 2316 859 2332
rect 911 2366 977 2382
rect 911 2332 927 2366
rect 961 2332 977 2366
rect 911 2316 977 2332
rect 1029 2366 1095 2382
rect 1029 2332 1045 2366
rect 1079 2332 1095 2366
rect 1029 2316 1095 2332
rect 1147 2366 1213 2382
rect 1147 2332 1163 2366
rect 1197 2332 1213 2366
rect 1147 2316 1213 2332
rect 1265 2366 1331 2382
rect 1265 2332 1281 2366
rect 1315 2332 1331 2366
rect 1265 2316 1331 2332
rect 1383 2366 1449 2382
rect 1383 2332 1399 2366
rect 1433 2332 1449 2366
rect 1383 2316 1449 2332
rect -1446 2248 -1386 2274
rect -1328 2248 -1268 2274
rect -1210 2248 -1150 2274
rect -1092 2248 -1032 2274
rect -974 2248 -914 2274
rect -856 2248 -796 2274
rect -738 2248 -678 2274
rect -620 2248 -560 2274
rect -502 2248 -442 2274
rect -384 2248 -324 2274
rect -266 2248 -206 2274
rect -148 2248 -88 2274
rect -30 2248 30 2274
rect 88 2248 148 2274
rect 206 2248 266 2274
rect 324 2248 384 2274
rect 442 2248 502 2274
rect 560 2248 620 2274
rect 678 2248 738 2274
rect 796 2248 856 2274
rect 914 2248 974 2274
rect 1032 2248 1092 2274
rect 1150 2248 1210 2274
rect 1268 2248 1328 2274
rect 1386 2248 1446 2274
rect -1446 1617 -1386 1648
rect -1328 1617 -1268 1648
rect -1210 1617 -1150 1648
rect -1092 1617 -1032 1648
rect -974 1617 -914 1648
rect -856 1617 -796 1648
rect -738 1617 -678 1648
rect -620 1617 -560 1648
rect -502 1617 -442 1648
rect -384 1617 -324 1648
rect -266 1617 -206 1648
rect -148 1617 -88 1648
rect -30 1617 30 1648
rect 88 1617 148 1648
rect 206 1617 266 1648
rect 324 1617 384 1648
rect 442 1617 502 1648
rect 560 1617 620 1648
rect 678 1617 738 1648
rect 796 1617 856 1648
rect 914 1617 974 1648
rect 1032 1617 1092 1648
rect 1150 1617 1210 1648
rect 1268 1617 1328 1648
rect 1386 1617 1446 1648
rect -1449 1601 -1383 1617
rect -1449 1567 -1433 1601
rect -1399 1567 -1383 1601
rect -1449 1551 -1383 1567
rect -1331 1601 -1265 1617
rect -1331 1567 -1315 1601
rect -1281 1567 -1265 1601
rect -1331 1551 -1265 1567
rect -1213 1601 -1147 1617
rect -1213 1567 -1197 1601
rect -1163 1567 -1147 1601
rect -1213 1551 -1147 1567
rect -1095 1601 -1029 1617
rect -1095 1567 -1079 1601
rect -1045 1567 -1029 1601
rect -1095 1551 -1029 1567
rect -977 1601 -911 1617
rect -977 1567 -961 1601
rect -927 1567 -911 1601
rect -977 1551 -911 1567
rect -859 1601 -793 1617
rect -859 1567 -843 1601
rect -809 1567 -793 1601
rect -859 1551 -793 1567
rect -741 1601 -675 1617
rect -741 1567 -725 1601
rect -691 1567 -675 1601
rect -741 1551 -675 1567
rect -623 1601 -557 1617
rect -623 1567 -607 1601
rect -573 1567 -557 1601
rect -623 1551 -557 1567
rect -505 1601 -439 1617
rect -505 1567 -489 1601
rect -455 1567 -439 1601
rect -505 1551 -439 1567
rect -387 1601 -321 1617
rect -387 1567 -371 1601
rect -337 1567 -321 1601
rect -387 1551 -321 1567
rect -269 1601 -203 1617
rect -269 1567 -253 1601
rect -219 1567 -203 1601
rect -269 1551 -203 1567
rect -151 1601 -85 1617
rect -151 1567 -135 1601
rect -101 1567 -85 1601
rect -151 1551 -85 1567
rect -33 1601 33 1617
rect -33 1567 -17 1601
rect 17 1567 33 1601
rect -33 1551 33 1567
rect 85 1601 151 1617
rect 85 1567 101 1601
rect 135 1567 151 1601
rect 85 1551 151 1567
rect 203 1601 269 1617
rect 203 1567 219 1601
rect 253 1567 269 1601
rect 203 1551 269 1567
rect 321 1601 387 1617
rect 321 1567 337 1601
rect 371 1567 387 1601
rect 321 1551 387 1567
rect 439 1601 505 1617
rect 439 1567 455 1601
rect 489 1567 505 1601
rect 439 1551 505 1567
rect 557 1601 623 1617
rect 557 1567 573 1601
rect 607 1567 623 1601
rect 557 1551 623 1567
rect 675 1601 741 1617
rect 675 1567 691 1601
rect 725 1567 741 1601
rect 675 1551 741 1567
rect 793 1601 859 1617
rect 793 1567 809 1601
rect 843 1567 859 1601
rect 793 1551 859 1567
rect 911 1601 977 1617
rect 911 1567 927 1601
rect 961 1567 977 1601
rect 911 1551 977 1567
rect 1029 1601 1095 1617
rect 1029 1567 1045 1601
rect 1079 1567 1095 1601
rect 1029 1551 1095 1567
rect 1147 1601 1213 1617
rect 1147 1567 1163 1601
rect 1197 1567 1213 1601
rect 1147 1551 1213 1567
rect 1265 1601 1331 1617
rect 1265 1567 1281 1601
rect 1315 1567 1331 1601
rect 1265 1551 1331 1567
rect 1383 1601 1449 1617
rect 1383 1567 1399 1601
rect 1433 1567 1449 1601
rect 1383 1551 1449 1567
rect -1446 1483 -1386 1509
rect -1328 1483 -1268 1509
rect -1210 1483 -1150 1509
rect -1092 1483 -1032 1509
rect -974 1483 -914 1509
rect -856 1483 -796 1509
rect -738 1483 -678 1509
rect -620 1483 -560 1509
rect -502 1483 -442 1509
rect -384 1483 -324 1509
rect -266 1483 -206 1509
rect -148 1483 -88 1509
rect -30 1483 30 1509
rect 88 1483 148 1509
rect 206 1483 266 1509
rect 324 1483 384 1509
rect 442 1483 502 1509
rect 560 1483 620 1509
rect 678 1483 738 1509
rect 796 1483 856 1509
rect 914 1483 974 1509
rect 1032 1483 1092 1509
rect 1150 1483 1210 1509
rect 1268 1483 1328 1509
rect 1386 1483 1446 1509
rect -1446 852 -1386 883
rect -1328 852 -1268 883
rect -1210 852 -1150 883
rect -1092 852 -1032 883
rect -974 852 -914 883
rect -856 852 -796 883
rect -738 852 -678 883
rect -620 852 -560 883
rect -502 852 -442 883
rect -384 852 -324 883
rect -266 852 -206 883
rect -148 852 -88 883
rect -30 852 30 883
rect 88 852 148 883
rect 206 852 266 883
rect 324 852 384 883
rect 442 852 502 883
rect 560 852 620 883
rect 678 852 738 883
rect 796 852 856 883
rect 914 852 974 883
rect 1032 852 1092 883
rect 1150 852 1210 883
rect 1268 852 1328 883
rect 1386 852 1446 883
rect -1449 836 -1383 852
rect -1449 802 -1433 836
rect -1399 802 -1383 836
rect -1449 786 -1383 802
rect -1331 836 -1265 852
rect -1331 802 -1315 836
rect -1281 802 -1265 836
rect -1331 786 -1265 802
rect -1213 836 -1147 852
rect -1213 802 -1197 836
rect -1163 802 -1147 836
rect -1213 786 -1147 802
rect -1095 836 -1029 852
rect -1095 802 -1079 836
rect -1045 802 -1029 836
rect -1095 786 -1029 802
rect -977 836 -911 852
rect -977 802 -961 836
rect -927 802 -911 836
rect -977 786 -911 802
rect -859 836 -793 852
rect -859 802 -843 836
rect -809 802 -793 836
rect -859 786 -793 802
rect -741 836 -675 852
rect -741 802 -725 836
rect -691 802 -675 836
rect -741 786 -675 802
rect -623 836 -557 852
rect -623 802 -607 836
rect -573 802 -557 836
rect -623 786 -557 802
rect -505 836 -439 852
rect -505 802 -489 836
rect -455 802 -439 836
rect -505 786 -439 802
rect -387 836 -321 852
rect -387 802 -371 836
rect -337 802 -321 836
rect -387 786 -321 802
rect -269 836 -203 852
rect -269 802 -253 836
rect -219 802 -203 836
rect -269 786 -203 802
rect -151 836 -85 852
rect -151 802 -135 836
rect -101 802 -85 836
rect -151 786 -85 802
rect -33 836 33 852
rect -33 802 -17 836
rect 17 802 33 836
rect -33 786 33 802
rect 85 836 151 852
rect 85 802 101 836
rect 135 802 151 836
rect 85 786 151 802
rect 203 836 269 852
rect 203 802 219 836
rect 253 802 269 836
rect 203 786 269 802
rect 321 836 387 852
rect 321 802 337 836
rect 371 802 387 836
rect 321 786 387 802
rect 439 836 505 852
rect 439 802 455 836
rect 489 802 505 836
rect 439 786 505 802
rect 557 836 623 852
rect 557 802 573 836
rect 607 802 623 836
rect 557 786 623 802
rect 675 836 741 852
rect 675 802 691 836
rect 725 802 741 836
rect 675 786 741 802
rect 793 836 859 852
rect 793 802 809 836
rect 843 802 859 836
rect 793 786 859 802
rect 911 836 977 852
rect 911 802 927 836
rect 961 802 977 836
rect 911 786 977 802
rect 1029 836 1095 852
rect 1029 802 1045 836
rect 1079 802 1095 836
rect 1029 786 1095 802
rect 1147 836 1213 852
rect 1147 802 1163 836
rect 1197 802 1213 836
rect 1147 786 1213 802
rect 1265 836 1331 852
rect 1265 802 1281 836
rect 1315 802 1331 836
rect 1265 786 1331 802
rect 1383 836 1449 852
rect 1383 802 1399 836
rect 1433 802 1449 836
rect 1383 786 1449 802
rect -1446 718 -1386 744
rect -1328 718 -1268 744
rect -1210 718 -1150 744
rect -1092 718 -1032 744
rect -974 718 -914 744
rect -856 718 -796 744
rect -738 718 -678 744
rect -620 718 -560 744
rect -502 718 -442 744
rect -384 718 -324 744
rect -266 718 -206 744
rect -148 718 -88 744
rect -30 718 30 744
rect 88 718 148 744
rect 206 718 266 744
rect 324 718 384 744
rect 442 718 502 744
rect 560 718 620 744
rect 678 718 738 744
rect 796 718 856 744
rect 914 718 974 744
rect 1032 718 1092 744
rect 1150 718 1210 744
rect 1268 718 1328 744
rect 1386 718 1446 744
rect -1446 87 -1386 118
rect -1328 87 -1268 118
rect -1210 87 -1150 118
rect -1092 87 -1032 118
rect -974 87 -914 118
rect -856 87 -796 118
rect -738 87 -678 118
rect -620 87 -560 118
rect -502 87 -442 118
rect -384 87 -324 118
rect -266 87 -206 118
rect -148 87 -88 118
rect -30 87 30 118
rect 88 87 148 118
rect 206 87 266 118
rect 324 87 384 118
rect 442 87 502 118
rect 560 87 620 118
rect 678 87 738 118
rect 796 87 856 118
rect 914 87 974 118
rect 1032 87 1092 118
rect 1150 87 1210 118
rect 1268 87 1328 118
rect 1386 87 1446 118
rect -1449 71 -1383 87
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1449 21 -1383 37
rect -1331 71 -1265 87
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1331 21 -1265 37
rect -1213 71 -1147 87
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1213 21 -1147 37
rect -1095 71 -1029 87
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -1095 21 -1029 37
rect -977 71 -911 87
rect -977 37 -961 71
rect -927 37 -911 71
rect -977 21 -911 37
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect 911 71 977 87
rect 911 37 927 71
rect 961 37 977 71
rect 911 21 977 37
rect 1029 71 1095 87
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1029 21 1095 37
rect 1147 71 1213 87
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1147 21 1213 37
rect 1265 71 1331 87
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1265 21 1331 37
rect 1383 71 1449 87
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1383 21 1449 37
rect -1446 -47 -1386 -21
rect -1328 -47 -1268 -21
rect -1210 -47 -1150 -21
rect -1092 -47 -1032 -21
rect -974 -47 -914 -21
rect -856 -47 -796 -21
rect -738 -47 -678 -21
rect -620 -47 -560 -21
rect -502 -47 -442 -21
rect -384 -47 -324 -21
rect -266 -47 -206 -21
rect -148 -47 -88 -21
rect -30 -47 30 -21
rect 88 -47 148 -21
rect 206 -47 266 -21
rect 324 -47 384 -21
rect 442 -47 502 -21
rect 560 -47 620 -21
rect 678 -47 738 -21
rect 796 -47 856 -21
rect 914 -47 974 -21
rect 1032 -47 1092 -21
rect 1150 -47 1210 -21
rect 1268 -47 1328 -21
rect 1386 -47 1446 -21
rect -1446 -678 -1386 -647
rect -1328 -678 -1268 -647
rect -1210 -678 -1150 -647
rect -1092 -678 -1032 -647
rect -974 -678 -914 -647
rect -856 -678 -796 -647
rect -738 -678 -678 -647
rect -620 -678 -560 -647
rect -502 -678 -442 -647
rect -384 -678 -324 -647
rect -266 -678 -206 -647
rect -148 -678 -88 -647
rect -30 -678 30 -647
rect 88 -678 148 -647
rect 206 -678 266 -647
rect 324 -678 384 -647
rect 442 -678 502 -647
rect 560 -678 620 -647
rect 678 -678 738 -647
rect 796 -678 856 -647
rect 914 -678 974 -647
rect 1032 -678 1092 -647
rect 1150 -678 1210 -647
rect 1268 -678 1328 -647
rect 1386 -678 1446 -647
rect -1449 -694 -1383 -678
rect -1449 -728 -1433 -694
rect -1399 -728 -1383 -694
rect -1449 -744 -1383 -728
rect -1331 -694 -1265 -678
rect -1331 -728 -1315 -694
rect -1281 -728 -1265 -694
rect -1331 -744 -1265 -728
rect -1213 -694 -1147 -678
rect -1213 -728 -1197 -694
rect -1163 -728 -1147 -694
rect -1213 -744 -1147 -728
rect -1095 -694 -1029 -678
rect -1095 -728 -1079 -694
rect -1045 -728 -1029 -694
rect -1095 -744 -1029 -728
rect -977 -694 -911 -678
rect -977 -728 -961 -694
rect -927 -728 -911 -694
rect -977 -744 -911 -728
rect -859 -694 -793 -678
rect -859 -728 -843 -694
rect -809 -728 -793 -694
rect -859 -744 -793 -728
rect -741 -694 -675 -678
rect -741 -728 -725 -694
rect -691 -728 -675 -694
rect -741 -744 -675 -728
rect -623 -694 -557 -678
rect -623 -728 -607 -694
rect -573 -728 -557 -694
rect -623 -744 -557 -728
rect -505 -694 -439 -678
rect -505 -728 -489 -694
rect -455 -728 -439 -694
rect -505 -744 -439 -728
rect -387 -694 -321 -678
rect -387 -728 -371 -694
rect -337 -728 -321 -694
rect -387 -744 -321 -728
rect -269 -694 -203 -678
rect -269 -728 -253 -694
rect -219 -728 -203 -694
rect -269 -744 -203 -728
rect -151 -694 -85 -678
rect -151 -728 -135 -694
rect -101 -728 -85 -694
rect -151 -744 -85 -728
rect -33 -694 33 -678
rect -33 -728 -17 -694
rect 17 -728 33 -694
rect -33 -744 33 -728
rect 85 -694 151 -678
rect 85 -728 101 -694
rect 135 -728 151 -694
rect 85 -744 151 -728
rect 203 -694 269 -678
rect 203 -728 219 -694
rect 253 -728 269 -694
rect 203 -744 269 -728
rect 321 -694 387 -678
rect 321 -728 337 -694
rect 371 -728 387 -694
rect 321 -744 387 -728
rect 439 -694 505 -678
rect 439 -728 455 -694
rect 489 -728 505 -694
rect 439 -744 505 -728
rect 557 -694 623 -678
rect 557 -728 573 -694
rect 607 -728 623 -694
rect 557 -744 623 -728
rect 675 -694 741 -678
rect 675 -728 691 -694
rect 725 -728 741 -694
rect 675 -744 741 -728
rect 793 -694 859 -678
rect 793 -728 809 -694
rect 843 -728 859 -694
rect 793 -744 859 -728
rect 911 -694 977 -678
rect 911 -728 927 -694
rect 961 -728 977 -694
rect 911 -744 977 -728
rect 1029 -694 1095 -678
rect 1029 -728 1045 -694
rect 1079 -728 1095 -694
rect 1029 -744 1095 -728
rect 1147 -694 1213 -678
rect 1147 -728 1163 -694
rect 1197 -728 1213 -694
rect 1147 -744 1213 -728
rect 1265 -694 1331 -678
rect 1265 -728 1281 -694
rect 1315 -728 1331 -694
rect 1265 -744 1331 -728
rect 1383 -694 1449 -678
rect 1383 -728 1399 -694
rect 1433 -728 1449 -694
rect 1383 -744 1449 -728
rect -1446 -812 -1386 -786
rect -1328 -812 -1268 -786
rect -1210 -812 -1150 -786
rect -1092 -812 -1032 -786
rect -974 -812 -914 -786
rect -856 -812 -796 -786
rect -738 -812 -678 -786
rect -620 -812 -560 -786
rect -502 -812 -442 -786
rect -384 -812 -324 -786
rect -266 -812 -206 -786
rect -148 -812 -88 -786
rect -30 -812 30 -786
rect 88 -812 148 -786
rect 206 -812 266 -786
rect 324 -812 384 -786
rect 442 -812 502 -786
rect 560 -812 620 -786
rect 678 -812 738 -786
rect 796 -812 856 -786
rect 914 -812 974 -786
rect 1032 -812 1092 -786
rect 1150 -812 1210 -786
rect 1268 -812 1328 -786
rect 1386 -812 1446 -786
rect -1446 -1443 -1386 -1412
rect -1328 -1443 -1268 -1412
rect -1210 -1443 -1150 -1412
rect -1092 -1443 -1032 -1412
rect -974 -1443 -914 -1412
rect -856 -1443 -796 -1412
rect -738 -1443 -678 -1412
rect -620 -1443 -560 -1412
rect -502 -1443 -442 -1412
rect -384 -1443 -324 -1412
rect -266 -1443 -206 -1412
rect -148 -1443 -88 -1412
rect -30 -1443 30 -1412
rect 88 -1443 148 -1412
rect 206 -1443 266 -1412
rect 324 -1443 384 -1412
rect 442 -1443 502 -1412
rect 560 -1443 620 -1412
rect 678 -1443 738 -1412
rect 796 -1443 856 -1412
rect 914 -1443 974 -1412
rect 1032 -1443 1092 -1412
rect 1150 -1443 1210 -1412
rect 1268 -1443 1328 -1412
rect 1386 -1443 1446 -1412
rect -1449 -1459 -1383 -1443
rect -1449 -1493 -1433 -1459
rect -1399 -1493 -1383 -1459
rect -1449 -1509 -1383 -1493
rect -1331 -1459 -1265 -1443
rect -1331 -1493 -1315 -1459
rect -1281 -1493 -1265 -1459
rect -1331 -1509 -1265 -1493
rect -1213 -1459 -1147 -1443
rect -1213 -1493 -1197 -1459
rect -1163 -1493 -1147 -1459
rect -1213 -1509 -1147 -1493
rect -1095 -1459 -1029 -1443
rect -1095 -1493 -1079 -1459
rect -1045 -1493 -1029 -1459
rect -1095 -1509 -1029 -1493
rect -977 -1459 -911 -1443
rect -977 -1493 -961 -1459
rect -927 -1493 -911 -1459
rect -977 -1509 -911 -1493
rect -859 -1459 -793 -1443
rect -859 -1493 -843 -1459
rect -809 -1493 -793 -1459
rect -859 -1509 -793 -1493
rect -741 -1459 -675 -1443
rect -741 -1493 -725 -1459
rect -691 -1493 -675 -1459
rect -741 -1509 -675 -1493
rect -623 -1459 -557 -1443
rect -623 -1493 -607 -1459
rect -573 -1493 -557 -1459
rect -623 -1509 -557 -1493
rect -505 -1459 -439 -1443
rect -505 -1493 -489 -1459
rect -455 -1493 -439 -1459
rect -505 -1509 -439 -1493
rect -387 -1459 -321 -1443
rect -387 -1493 -371 -1459
rect -337 -1493 -321 -1459
rect -387 -1509 -321 -1493
rect -269 -1459 -203 -1443
rect -269 -1493 -253 -1459
rect -219 -1493 -203 -1459
rect -269 -1509 -203 -1493
rect -151 -1459 -85 -1443
rect -151 -1493 -135 -1459
rect -101 -1493 -85 -1459
rect -151 -1509 -85 -1493
rect -33 -1459 33 -1443
rect -33 -1493 -17 -1459
rect 17 -1493 33 -1459
rect -33 -1509 33 -1493
rect 85 -1459 151 -1443
rect 85 -1493 101 -1459
rect 135 -1493 151 -1459
rect 85 -1509 151 -1493
rect 203 -1459 269 -1443
rect 203 -1493 219 -1459
rect 253 -1493 269 -1459
rect 203 -1509 269 -1493
rect 321 -1459 387 -1443
rect 321 -1493 337 -1459
rect 371 -1493 387 -1459
rect 321 -1509 387 -1493
rect 439 -1459 505 -1443
rect 439 -1493 455 -1459
rect 489 -1493 505 -1459
rect 439 -1509 505 -1493
rect 557 -1459 623 -1443
rect 557 -1493 573 -1459
rect 607 -1493 623 -1459
rect 557 -1509 623 -1493
rect 675 -1459 741 -1443
rect 675 -1493 691 -1459
rect 725 -1493 741 -1459
rect 675 -1509 741 -1493
rect 793 -1459 859 -1443
rect 793 -1493 809 -1459
rect 843 -1493 859 -1459
rect 793 -1509 859 -1493
rect 911 -1459 977 -1443
rect 911 -1493 927 -1459
rect 961 -1493 977 -1459
rect 911 -1509 977 -1493
rect 1029 -1459 1095 -1443
rect 1029 -1493 1045 -1459
rect 1079 -1493 1095 -1459
rect 1029 -1509 1095 -1493
rect 1147 -1459 1213 -1443
rect 1147 -1493 1163 -1459
rect 1197 -1493 1213 -1459
rect 1147 -1509 1213 -1493
rect 1265 -1459 1331 -1443
rect 1265 -1493 1281 -1459
rect 1315 -1493 1331 -1459
rect 1265 -1509 1331 -1493
rect 1383 -1459 1449 -1443
rect 1383 -1493 1399 -1459
rect 1433 -1493 1449 -1459
rect 1383 -1509 1449 -1493
rect -1446 -1577 -1386 -1551
rect -1328 -1577 -1268 -1551
rect -1210 -1577 -1150 -1551
rect -1092 -1577 -1032 -1551
rect -974 -1577 -914 -1551
rect -856 -1577 -796 -1551
rect -738 -1577 -678 -1551
rect -620 -1577 -560 -1551
rect -502 -1577 -442 -1551
rect -384 -1577 -324 -1551
rect -266 -1577 -206 -1551
rect -148 -1577 -88 -1551
rect -30 -1577 30 -1551
rect 88 -1577 148 -1551
rect 206 -1577 266 -1551
rect 324 -1577 384 -1551
rect 442 -1577 502 -1551
rect 560 -1577 620 -1551
rect 678 -1577 738 -1551
rect 796 -1577 856 -1551
rect 914 -1577 974 -1551
rect 1032 -1577 1092 -1551
rect 1150 -1577 1210 -1551
rect 1268 -1577 1328 -1551
rect 1386 -1577 1446 -1551
rect -1446 -2208 -1386 -2177
rect -1328 -2208 -1268 -2177
rect -1210 -2208 -1150 -2177
rect -1092 -2208 -1032 -2177
rect -974 -2208 -914 -2177
rect -856 -2208 -796 -2177
rect -738 -2208 -678 -2177
rect -620 -2208 -560 -2177
rect -502 -2208 -442 -2177
rect -384 -2208 -324 -2177
rect -266 -2208 -206 -2177
rect -148 -2208 -88 -2177
rect -30 -2208 30 -2177
rect 88 -2208 148 -2177
rect 206 -2208 266 -2177
rect 324 -2208 384 -2177
rect 442 -2208 502 -2177
rect 560 -2208 620 -2177
rect 678 -2208 738 -2177
rect 796 -2208 856 -2177
rect 914 -2208 974 -2177
rect 1032 -2208 1092 -2177
rect 1150 -2208 1210 -2177
rect 1268 -2208 1328 -2177
rect 1386 -2208 1446 -2177
rect -1449 -2224 -1383 -2208
rect -1449 -2258 -1433 -2224
rect -1399 -2258 -1383 -2224
rect -1449 -2274 -1383 -2258
rect -1331 -2224 -1265 -2208
rect -1331 -2258 -1315 -2224
rect -1281 -2258 -1265 -2224
rect -1331 -2274 -1265 -2258
rect -1213 -2224 -1147 -2208
rect -1213 -2258 -1197 -2224
rect -1163 -2258 -1147 -2224
rect -1213 -2274 -1147 -2258
rect -1095 -2224 -1029 -2208
rect -1095 -2258 -1079 -2224
rect -1045 -2258 -1029 -2224
rect -1095 -2274 -1029 -2258
rect -977 -2224 -911 -2208
rect -977 -2258 -961 -2224
rect -927 -2258 -911 -2224
rect -977 -2274 -911 -2258
rect -859 -2224 -793 -2208
rect -859 -2258 -843 -2224
rect -809 -2258 -793 -2224
rect -859 -2274 -793 -2258
rect -741 -2224 -675 -2208
rect -741 -2258 -725 -2224
rect -691 -2258 -675 -2224
rect -741 -2274 -675 -2258
rect -623 -2224 -557 -2208
rect -623 -2258 -607 -2224
rect -573 -2258 -557 -2224
rect -623 -2274 -557 -2258
rect -505 -2224 -439 -2208
rect -505 -2258 -489 -2224
rect -455 -2258 -439 -2224
rect -505 -2274 -439 -2258
rect -387 -2224 -321 -2208
rect -387 -2258 -371 -2224
rect -337 -2258 -321 -2224
rect -387 -2274 -321 -2258
rect -269 -2224 -203 -2208
rect -269 -2258 -253 -2224
rect -219 -2258 -203 -2224
rect -269 -2274 -203 -2258
rect -151 -2224 -85 -2208
rect -151 -2258 -135 -2224
rect -101 -2258 -85 -2224
rect -151 -2274 -85 -2258
rect -33 -2224 33 -2208
rect -33 -2258 -17 -2224
rect 17 -2258 33 -2224
rect -33 -2274 33 -2258
rect 85 -2224 151 -2208
rect 85 -2258 101 -2224
rect 135 -2258 151 -2224
rect 85 -2274 151 -2258
rect 203 -2224 269 -2208
rect 203 -2258 219 -2224
rect 253 -2258 269 -2224
rect 203 -2274 269 -2258
rect 321 -2224 387 -2208
rect 321 -2258 337 -2224
rect 371 -2258 387 -2224
rect 321 -2274 387 -2258
rect 439 -2224 505 -2208
rect 439 -2258 455 -2224
rect 489 -2258 505 -2224
rect 439 -2274 505 -2258
rect 557 -2224 623 -2208
rect 557 -2258 573 -2224
rect 607 -2258 623 -2224
rect 557 -2274 623 -2258
rect 675 -2224 741 -2208
rect 675 -2258 691 -2224
rect 725 -2258 741 -2224
rect 675 -2274 741 -2258
rect 793 -2224 859 -2208
rect 793 -2258 809 -2224
rect 843 -2258 859 -2224
rect 793 -2274 859 -2258
rect 911 -2224 977 -2208
rect 911 -2258 927 -2224
rect 961 -2258 977 -2224
rect 911 -2274 977 -2258
rect 1029 -2224 1095 -2208
rect 1029 -2258 1045 -2224
rect 1079 -2258 1095 -2224
rect 1029 -2274 1095 -2258
rect 1147 -2224 1213 -2208
rect 1147 -2258 1163 -2224
rect 1197 -2258 1213 -2224
rect 1147 -2274 1213 -2258
rect 1265 -2224 1331 -2208
rect 1265 -2258 1281 -2224
rect 1315 -2258 1331 -2224
rect 1265 -2274 1331 -2258
rect 1383 -2224 1449 -2208
rect 1383 -2258 1399 -2224
rect 1433 -2258 1449 -2224
rect 1383 -2274 1449 -2258
rect -1446 -2342 -1386 -2316
rect -1328 -2342 -1268 -2316
rect -1210 -2342 -1150 -2316
rect -1092 -2342 -1032 -2316
rect -974 -2342 -914 -2316
rect -856 -2342 -796 -2316
rect -738 -2342 -678 -2316
rect -620 -2342 -560 -2316
rect -502 -2342 -442 -2316
rect -384 -2342 -324 -2316
rect -266 -2342 -206 -2316
rect -148 -2342 -88 -2316
rect -30 -2342 30 -2316
rect 88 -2342 148 -2316
rect 206 -2342 266 -2316
rect 324 -2342 384 -2316
rect 442 -2342 502 -2316
rect 560 -2342 620 -2316
rect 678 -2342 738 -2316
rect 796 -2342 856 -2316
rect 914 -2342 974 -2316
rect 1032 -2342 1092 -2316
rect 1150 -2342 1210 -2316
rect 1268 -2342 1328 -2316
rect 1386 -2342 1446 -2316
rect -1446 -2973 -1386 -2942
rect -1328 -2973 -1268 -2942
rect -1210 -2973 -1150 -2942
rect -1092 -2973 -1032 -2942
rect -974 -2973 -914 -2942
rect -856 -2973 -796 -2942
rect -738 -2973 -678 -2942
rect -620 -2973 -560 -2942
rect -502 -2973 -442 -2942
rect -384 -2973 -324 -2942
rect -266 -2973 -206 -2942
rect -148 -2973 -88 -2942
rect -30 -2973 30 -2942
rect 88 -2973 148 -2942
rect 206 -2973 266 -2942
rect 324 -2973 384 -2942
rect 442 -2973 502 -2942
rect 560 -2973 620 -2942
rect 678 -2973 738 -2942
rect 796 -2973 856 -2942
rect 914 -2973 974 -2942
rect 1032 -2973 1092 -2942
rect 1150 -2973 1210 -2942
rect 1268 -2973 1328 -2942
rect 1386 -2973 1446 -2942
rect -1449 -2989 -1383 -2973
rect -1449 -3023 -1433 -2989
rect -1399 -3023 -1383 -2989
rect -1449 -3039 -1383 -3023
rect -1331 -2989 -1265 -2973
rect -1331 -3023 -1315 -2989
rect -1281 -3023 -1265 -2989
rect -1331 -3039 -1265 -3023
rect -1213 -2989 -1147 -2973
rect -1213 -3023 -1197 -2989
rect -1163 -3023 -1147 -2989
rect -1213 -3039 -1147 -3023
rect -1095 -2989 -1029 -2973
rect -1095 -3023 -1079 -2989
rect -1045 -3023 -1029 -2989
rect -1095 -3039 -1029 -3023
rect -977 -2989 -911 -2973
rect -977 -3023 -961 -2989
rect -927 -3023 -911 -2989
rect -977 -3039 -911 -3023
rect -859 -2989 -793 -2973
rect -859 -3023 -843 -2989
rect -809 -3023 -793 -2989
rect -859 -3039 -793 -3023
rect -741 -2989 -675 -2973
rect -741 -3023 -725 -2989
rect -691 -3023 -675 -2989
rect -741 -3039 -675 -3023
rect -623 -2989 -557 -2973
rect -623 -3023 -607 -2989
rect -573 -3023 -557 -2989
rect -623 -3039 -557 -3023
rect -505 -2989 -439 -2973
rect -505 -3023 -489 -2989
rect -455 -3023 -439 -2989
rect -505 -3039 -439 -3023
rect -387 -2989 -321 -2973
rect -387 -3023 -371 -2989
rect -337 -3023 -321 -2989
rect -387 -3039 -321 -3023
rect -269 -2989 -203 -2973
rect -269 -3023 -253 -2989
rect -219 -3023 -203 -2989
rect -269 -3039 -203 -3023
rect -151 -2989 -85 -2973
rect -151 -3023 -135 -2989
rect -101 -3023 -85 -2989
rect -151 -3039 -85 -3023
rect -33 -2989 33 -2973
rect -33 -3023 -17 -2989
rect 17 -3023 33 -2989
rect -33 -3039 33 -3023
rect 85 -2989 151 -2973
rect 85 -3023 101 -2989
rect 135 -3023 151 -2989
rect 85 -3039 151 -3023
rect 203 -2989 269 -2973
rect 203 -3023 219 -2989
rect 253 -3023 269 -2989
rect 203 -3039 269 -3023
rect 321 -2989 387 -2973
rect 321 -3023 337 -2989
rect 371 -3023 387 -2989
rect 321 -3039 387 -3023
rect 439 -2989 505 -2973
rect 439 -3023 455 -2989
rect 489 -3023 505 -2989
rect 439 -3039 505 -3023
rect 557 -2989 623 -2973
rect 557 -3023 573 -2989
rect 607 -3023 623 -2989
rect 557 -3039 623 -3023
rect 675 -2989 741 -2973
rect 675 -3023 691 -2989
rect 725 -3023 741 -2989
rect 675 -3039 741 -3023
rect 793 -2989 859 -2973
rect 793 -3023 809 -2989
rect 843 -3023 859 -2989
rect 793 -3039 859 -3023
rect 911 -2989 977 -2973
rect 911 -3023 927 -2989
rect 961 -3023 977 -2989
rect 911 -3039 977 -3023
rect 1029 -2989 1095 -2973
rect 1029 -3023 1045 -2989
rect 1079 -3023 1095 -2989
rect 1029 -3039 1095 -3023
rect 1147 -2989 1213 -2973
rect 1147 -3023 1163 -2989
rect 1197 -3023 1213 -2989
rect 1147 -3039 1213 -3023
rect 1265 -2989 1331 -2973
rect 1265 -3023 1281 -2989
rect 1315 -3023 1331 -2989
rect 1265 -3039 1331 -3023
rect 1383 -2989 1449 -2973
rect 1383 -3023 1399 -2989
rect 1433 -3023 1449 -2989
rect 1383 -3039 1449 -3023
rect -1446 -3107 -1386 -3081
rect -1328 -3107 -1268 -3081
rect -1210 -3107 -1150 -3081
rect -1092 -3107 -1032 -3081
rect -974 -3107 -914 -3081
rect -856 -3107 -796 -3081
rect -738 -3107 -678 -3081
rect -620 -3107 -560 -3081
rect -502 -3107 -442 -3081
rect -384 -3107 -324 -3081
rect -266 -3107 -206 -3081
rect -148 -3107 -88 -3081
rect -30 -3107 30 -3081
rect 88 -3107 148 -3081
rect 206 -3107 266 -3081
rect 324 -3107 384 -3081
rect 442 -3107 502 -3081
rect 560 -3107 620 -3081
rect 678 -3107 738 -3081
rect 796 -3107 856 -3081
rect 914 -3107 974 -3081
rect 1032 -3107 1092 -3081
rect 1150 -3107 1210 -3081
rect 1268 -3107 1328 -3081
rect 1386 -3107 1446 -3081
rect -1446 -3738 -1386 -3707
rect -1328 -3738 -1268 -3707
rect -1210 -3738 -1150 -3707
rect -1092 -3738 -1032 -3707
rect -974 -3738 -914 -3707
rect -856 -3738 -796 -3707
rect -738 -3738 -678 -3707
rect -620 -3738 -560 -3707
rect -502 -3738 -442 -3707
rect -384 -3738 -324 -3707
rect -266 -3738 -206 -3707
rect -148 -3738 -88 -3707
rect -30 -3738 30 -3707
rect 88 -3738 148 -3707
rect 206 -3738 266 -3707
rect 324 -3738 384 -3707
rect 442 -3738 502 -3707
rect 560 -3738 620 -3707
rect 678 -3738 738 -3707
rect 796 -3738 856 -3707
rect 914 -3738 974 -3707
rect 1032 -3738 1092 -3707
rect 1150 -3738 1210 -3707
rect 1268 -3738 1328 -3707
rect 1386 -3738 1446 -3707
rect -1449 -3754 -1383 -3738
rect -1449 -3788 -1433 -3754
rect -1399 -3788 -1383 -3754
rect -1449 -3804 -1383 -3788
rect -1331 -3754 -1265 -3738
rect -1331 -3788 -1315 -3754
rect -1281 -3788 -1265 -3754
rect -1331 -3804 -1265 -3788
rect -1213 -3754 -1147 -3738
rect -1213 -3788 -1197 -3754
rect -1163 -3788 -1147 -3754
rect -1213 -3804 -1147 -3788
rect -1095 -3754 -1029 -3738
rect -1095 -3788 -1079 -3754
rect -1045 -3788 -1029 -3754
rect -1095 -3804 -1029 -3788
rect -977 -3754 -911 -3738
rect -977 -3788 -961 -3754
rect -927 -3788 -911 -3754
rect -977 -3804 -911 -3788
rect -859 -3754 -793 -3738
rect -859 -3788 -843 -3754
rect -809 -3788 -793 -3754
rect -859 -3804 -793 -3788
rect -741 -3754 -675 -3738
rect -741 -3788 -725 -3754
rect -691 -3788 -675 -3754
rect -741 -3804 -675 -3788
rect -623 -3754 -557 -3738
rect -623 -3788 -607 -3754
rect -573 -3788 -557 -3754
rect -623 -3804 -557 -3788
rect -505 -3754 -439 -3738
rect -505 -3788 -489 -3754
rect -455 -3788 -439 -3754
rect -505 -3804 -439 -3788
rect -387 -3754 -321 -3738
rect -387 -3788 -371 -3754
rect -337 -3788 -321 -3754
rect -387 -3804 -321 -3788
rect -269 -3754 -203 -3738
rect -269 -3788 -253 -3754
rect -219 -3788 -203 -3754
rect -269 -3804 -203 -3788
rect -151 -3754 -85 -3738
rect -151 -3788 -135 -3754
rect -101 -3788 -85 -3754
rect -151 -3804 -85 -3788
rect -33 -3754 33 -3738
rect -33 -3788 -17 -3754
rect 17 -3788 33 -3754
rect -33 -3804 33 -3788
rect 85 -3754 151 -3738
rect 85 -3788 101 -3754
rect 135 -3788 151 -3754
rect 85 -3804 151 -3788
rect 203 -3754 269 -3738
rect 203 -3788 219 -3754
rect 253 -3788 269 -3754
rect 203 -3804 269 -3788
rect 321 -3754 387 -3738
rect 321 -3788 337 -3754
rect 371 -3788 387 -3754
rect 321 -3804 387 -3788
rect 439 -3754 505 -3738
rect 439 -3788 455 -3754
rect 489 -3788 505 -3754
rect 439 -3804 505 -3788
rect 557 -3754 623 -3738
rect 557 -3788 573 -3754
rect 607 -3788 623 -3754
rect 557 -3804 623 -3788
rect 675 -3754 741 -3738
rect 675 -3788 691 -3754
rect 725 -3788 741 -3754
rect 675 -3804 741 -3788
rect 793 -3754 859 -3738
rect 793 -3788 809 -3754
rect 843 -3788 859 -3754
rect 793 -3804 859 -3788
rect 911 -3754 977 -3738
rect 911 -3788 927 -3754
rect 961 -3788 977 -3754
rect 911 -3804 977 -3788
rect 1029 -3754 1095 -3738
rect 1029 -3788 1045 -3754
rect 1079 -3788 1095 -3754
rect 1029 -3804 1095 -3788
rect 1147 -3754 1213 -3738
rect 1147 -3788 1163 -3754
rect 1197 -3788 1213 -3754
rect 1147 -3804 1213 -3788
rect 1265 -3754 1331 -3738
rect 1265 -3788 1281 -3754
rect 1315 -3788 1331 -3754
rect 1265 -3804 1331 -3788
rect 1383 -3754 1449 -3738
rect 1383 -3788 1399 -3754
rect 1433 -3788 1449 -3754
rect 1383 -3804 1449 -3788
<< polycont >>
rect -1433 3097 -1399 3131
rect -1315 3097 -1281 3131
rect -1197 3097 -1163 3131
rect -1079 3097 -1045 3131
rect -961 3097 -927 3131
rect -843 3097 -809 3131
rect -725 3097 -691 3131
rect -607 3097 -573 3131
rect -489 3097 -455 3131
rect -371 3097 -337 3131
rect -253 3097 -219 3131
rect -135 3097 -101 3131
rect -17 3097 17 3131
rect 101 3097 135 3131
rect 219 3097 253 3131
rect 337 3097 371 3131
rect 455 3097 489 3131
rect 573 3097 607 3131
rect 691 3097 725 3131
rect 809 3097 843 3131
rect 927 3097 961 3131
rect 1045 3097 1079 3131
rect 1163 3097 1197 3131
rect 1281 3097 1315 3131
rect 1399 3097 1433 3131
rect -1433 2332 -1399 2366
rect -1315 2332 -1281 2366
rect -1197 2332 -1163 2366
rect -1079 2332 -1045 2366
rect -961 2332 -927 2366
rect -843 2332 -809 2366
rect -725 2332 -691 2366
rect -607 2332 -573 2366
rect -489 2332 -455 2366
rect -371 2332 -337 2366
rect -253 2332 -219 2366
rect -135 2332 -101 2366
rect -17 2332 17 2366
rect 101 2332 135 2366
rect 219 2332 253 2366
rect 337 2332 371 2366
rect 455 2332 489 2366
rect 573 2332 607 2366
rect 691 2332 725 2366
rect 809 2332 843 2366
rect 927 2332 961 2366
rect 1045 2332 1079 2366
rect 1163 2332 1197 2366
rect 1281 2332 1315 2366
rect 1399 2332 1433 2366
rect -1433 1567 -1399 1601
rect -1315 1567 -1281 1601
rect -1197 1567 -1163 1601
rect -1079 1567 -1045 1601
rect -961 1567 -927 1601
rect -843 1567 -809 1601
rect -725 1567 -691 1601
rect -607 1567 -573 1601
rect -489 1567 -455 1601
rect -371 1567 -337 1601
rect -253 1567 -219 1601
rect -135 1567 -101 1601
rect -17 1567 17 1601
rect 101 1567 135 1601
rect 219 1567 253 1601
rect 337 1567 371 1601
rect 455 1567 489 1601
rect 573 1567 607 1601
rect 691 1567 725 1601
rect 809 1567 843 1601
rect 927 1567 961 1601
rect 1045 1567 1079 1601
rect 1163 1567 1197 1601
rect 1281 1567 1315 1601
rect 1399 1567 1433 1601
rect -1433 802 -1399 836
rect -1315 802 -1281 836
rect -1197 802 -1163 836
rect -1079 802 -1045 836
rect -961 802 -927 836
rect -843 802 -809 836
rect -725 802 -691 836
rect -607 802 -573 836
rect -489 802 -455 836
rect -371 802 -337 836
rect -253 802 -219 836
rect -135 802 -101 836
rect -17 802 17 836
rect 101 802 135 836
rect 219 802 253 836
rect 337 802 371 836
rect 455 802 489 836
rect 573 802 607 836
rect 691 802 725 836
rect 809 802 843 836
rect 927 802 961 836
rect 1045 802 1079 836
rect 1163 802 1197 836
rect 1281 802 1315 836
rect 1399 802 1433 836
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1433 -728 -1399 -694
rect -1315 -728 -1281 -694
rect -1197 -728 -1163 -694
rect -1079 -728 -1045 -694
rect -961 -728 -927 -694
rect -843 -728 -809 -694
rect -725 -728 -691 -694
rect -607 -728 -573 -694
rect -489 -728 -455 -694
rect -371 -728 -337 -694
rect -253 -728 -219 -694
rect -135 -728 -101 -694
rect -17 -728 17 -694
rect 101 -728 135 -694
rect 219 -728 253 -694
rect 337 -728 371 -694
rect 455 -728 489 -694
rect 573 -728 607 -694
rect 691 -728 725 -694
rect 809 -728 843 -694
rect 927 -728 961 -694
rect 1045 -728 1079 -694
rect 1163 -728 1197 -694
rect 1281 -728 1315 -694
rect 1399 -728 1433 -694
rect -1433 -1493 -1399 -1459
rect -1315 -1493 -1281 -1459
rect -1197 -1493 -1163 -1459
rect -1079 -1493 -1045 -1459
rect -961 -1493 -927 -1459
rect -843 -1493 -809 -1459
rect -725 -1493 -691 -1459
rect -607 -1493 -573 -1459
rect -489 -1493 -455 -1459
rect -371 -1493 -337 -1459
rect -253 -1493 -219 -1459
rect -135 -1493 -101 -1459
rect -17 -1493 17 -1459
rect 101 -1493 135 -1459
rect 219 -1493 253 -1459
rect 337 -1493 371 -1459
rect 455 -1493 489 -1459
rect 573 -1493 607 -1459
rect 691 -1493 725 -1459
rect 809 -1493 843 -1459
rect 927 -1493 961 -1459
rect 1045 -1493 1079 -1459
rect 1163 -1493 1197 -1459
rect 1281 -1493 1315 -1459
rect 1399 -1493 1433 -1459
rect -1433 -2258 -1399 -2224
rect -1315 -2258 -1281 -2224
rect -1197 -2258 -1163 -2224
rect -1079 -2258 -1045 -2224
rect -961 -2258 -927 -2224
rect -843 -2258 -809 -2224
rect -725 -2258 -691 -2224
rect -607 -2258 -573 -2224
rect -489 -2258 -455 -2224
rect -371 -2258 -337 -2224
rect -253 -2258 -219 -2224
rect -135 -2258 -101 -2224
rect -17 -2258 17 -2224
rect 101 -2258 135 -2224
rect 219 -2258 253 -2224
rect 337 -2258 371 -2224
rect 455 -2258 489 -2224
rect 573 -2258 607 -2224
rect 691 -2258 725 -2224
rect 809 -2258 843 -2224
rect 927 -2258 961 -2224
rect 1045 -2258 1079 -2224
rect 1163 -2258 1197 -2224
rect 1281 -2258 1315 -2224
rect 1399 -2258 1433 -2224
rect -1433 -3023 -1399 -2989
rect -1315 -3023 -1281 -2989
rect -1197 -3023 -1163 -2989
rect -1079 -3023 -1045 -2989
rect -961 -3023 -927 -2989
rect -843 -3023 -809 -2989
rect -725 -3023 -691 -2989
rect -607 -3023 -573 -2989
rect -489 -3023 -455 -2989
rect -371 -3023 -337 -2989
rect -253 -3023 -219 -2989
rect -135 -3023 -101 -2989
rect -17 -3023 17 -2989
rect 101 -3023 135 -2989
rect 219 -3023 253 -2989
rect 337 -3023 371 -2989
rect 455 -3023 489 -2989
rect 573 -3023 607 -2989
rect 691 -3023 725 -2989
rect 809 -3023 843 -2989
rect 927 -3023 961 -2989
rect 1045 -3023 1079 -2989
rect 1163 -3023 1197 -2989
rect 1281 -3023 1315 -2989
rect 1399 -3023 1433 -2989
rect -1433 -3788 -1399 -3754
rect -1315 -3788 -1281 -3754
rect -1197 -3788 -1163 -3754
rect -1079 -3788 -1045 -3754
rect -961 -3788 -927 -3754
rect -843 -3788 -809 -3754
rect -725 -3788 -691 -3754
rect -607 -3788 -573 -3754
rect -489 -3788 -455 -3754
rect -371 -3788 -337 -3754
rect -253 -3788 -219 -3754
rect -135 -3788 -101 -3754
rect -17 -3788 17 -3754
rect 101 -3788 135 -3754
rect 219 -3788 253 -3754
rect 337 -3788 371 -3754
rect 455 -3788 489 -3754
rect 573 -3788 607 -3754
rect 691 -3788 725 -3754
rect 809 -3788 843 -3754
rect 927 -3788 961 -3754
rect 1045 -3788 1079 -3754
rect 1163 -3788 1197 -3754
rect 1281 -3788 1315 -3754
rect 1399 -3788 1433 -3754
<< locali >>
rect -1606 3856 -1510 3890
rect 1510 3856 1606 3890
rect -1606 3794 -1572 3856
rect 1572 3794 1606 3856
rect -1492 3766 -1458 3782
rect -1492 3174 -1458 3190
rect -1374 3766 -1340 3782
rect -1374 3174 -1340 3190
rect -1256 3766 -1222 3782
rect -1256 3174 -1222 3190
rect -1138 3766 -1104 3782
rect -1138 3174 -1104 3190
rect -1020 3766 -986 3782
rect -1020 3174 -986 3190
rect -902 3766 -868 3782
rect -902 3174 -868 3190
rect -784 3766 -750 3782
rect -784 3174 -750 3190
rect -666 3766 -632 3782
rect -666 3174 -632 3190
rect -548 3766 -514 3782
rect -548 3174 -514 3190
rect -430 3766 -396 3782
rect -430 3174 -396 3190
rect -312 3766 -278 3782
rect -312 3174 -278 3190
rect -194 3766 -160 3782
rect -194 3174 -160 3190
rect -76 3766 -42 3782
rect -76 3174 -42 3190
rect 42 3766 76 3782
rect 42 3174 76 3190
rect 160 3766 194 3782
rect 160 3174 194 3190
rect 278 3766 312 3782
rect 278 3174 312 3190
rect 396 3766 430 3782
rect 396 3174 430 3190
rect 514 3766 548 3782
rect 514 3174 548 3190
rect 632 3766 666 3782
rect 632 3174 666 3190
rect 750 3766 784 3782
rect 750 3174 784 3190
rect 868 3766 902 3782
rect 868 3174 902 3190
rect 986 3766 1020 3782
rect 986 3174 1020 3190
rect 1104 3766 1138 3782
rect 1104 3174 1138 3190
rect 1222 3766 1256 3782
rect 1222 3174 1256 3190
rect 1340 3766 1374 3782
rect 1340 3174 1374 3190
rect 1458 3766 1492 3782
rect 1458 3174 1492 3190
rect -1449 3097 -1433 3131
rect -1399 3097 -1383 3131
rect -1331 3097 -1315 3131
rect -1281 3097 -1265 3131
rect -1213 3097 -1197 3131
rect -1163 3097 -1147 3131
rect -1095 3097 -1079 3131
rect -1045 3097 -1029 3131
rect -977 3097 -961 3131
rect -927 3097 -911 3131
rect -859 3097 -843 3131
rect -809 3097 -793 3131
rect -741 3097 -725 3131
rect -691 3097 -675 3131
rect -623 3097 -607 3131
rect -573 3097 -557 3131
rect -505 3097 -489 3131
rect -455 3097 -439 3131
rect -387 3097 -371 3131
rect -337 3097 -321 3131
rect -269 3097 -253 3131
rect -219 3097 -203 3131
rect -151 3097 -135 3131
rect -101 3097 -85 3131
rect -33 3097 -17 3131
rect 17 3097 33 3131
rect 85 3097 101 3131
rect 135 3097 151 3131
rect 203 3097 219 3131
rect 253 3097 269 3131
rect 321 3097 337 3131
rect 371 3097 387 3131
rect 439 3097 455 3131
rect 489 3097 505 3131
rect 557 3097 573 3131
rect 607 3097 623 3131
rect 675 3097 691 3131
rect 725 3097 741 3131
rect 793 3097 809 3131
rect 843 3097 859 3131
rect 911 3097 927 3131
rect 961 3097 977 3131
rect 1029 3097 1045 3131
rect 1079 3097 1095 3131
rect 1147 3097 1163 3131
rect 1197 3097 1213 3131
rect 1265 3097 1281 3131
rect 1315 3097 1331 3131
rect 1383 3097 1399 3131
rect 1433 3097 1449 3131
rect -1492 3001 -1458 3017
rect -1492 2409 -1458 2425
rect -1374 3001 -1340 3017
rect -1374 2409 -1340 2425
rect -1256 3001 -1222 3017
rect -1256 2409 -1222 2425
rect -1138 3001 -1104 3017
rect -1138 2409 -1104 2425
rect -1020 3001 -986 3017
rect -1020 2409 -986 2425
rect -902 3001 -868 3017
rect -902 2409 -868 2425
rect -784 3001 -750 3017
rect -784 2409 -750 2425
rect -666 3001 -632 3017
rect -666 2409 -632 2425
rect -548 3001 -514 3017
rect -548 2409 -514 2425
rect -430 3001 -396 3017
rect -430 2409 -396 2425
rect -312 3001 -278 3017
rect -312 2409 -278 2425
rect -194 3001 -160 3017
rect -194 2409 -160 2425
rect -76 3001 -42 3017
rect -76 2409 -42 2425
rect 42 3001 76 3017
rect 42 2409 76 2425
rect 160 3001 194 3017
rect 160 2409 194 2425
rect 278 3001 312 3017
rect 278 2409 312 2425
rect 396 3001 430 3017
rect 396 2409 430 2425
rect 514 3001 548 3017
rect 514 2409 548 2425
rect 632 3001 666 3017
rect 632 2409 666 2425
rect 750 3001 784 3017
rect 750 2409 784 2425
rect 868 3001 902 3017
rect 868 2409 902 2425
rect 986 3001 1020 3017
rect 986 2409 1020 2425
rect 1104 3001 1138 3017
rect 1104 2409 1138 2425
rect 1222 3001 1256 3017
rect 1222 2409 1256 2425
rect 1340 3001 1374 3017
rect 1340 2409 1374 2425
rect 1458 3001 1492 3017
rect 1458 2409 1492 2425
rect -1449 2332 -1433 2366
rect -1399 2332 -1383 2366
rect -1331 2332 -1315 2366
rect -1281 2332 -1265 2366
rect -1213 2332 -1197 2366
rect -1163 2332 -1147 2366
rect -1095 2332 -1079 2366
rect -1045 2332 -1029 2366
rect -977 2332 -961 2366
rect -927 2332 -911 2366
rect -859 2332 -843 2366
rect -809 2332 -793 2366
rect -741 2332 -725 2366
rect -691 2332 -675 2366
rect -623 2332 -607 2366
rect -573 2332 -557 2366
rect -505 2332 -489 2366
rect -455 2332 -439 2366
rect -387 2332 -371 2366
rect -337 2332 -321 2366
rect -269 2332 -253 2366
rect -219 2332 -203 2366
rect -151 2332 -135 2366
rect -101 2332 -85 2366
rect -33 2332 -17 2366
rect 17 2332 33 2366
rect 85 2332 101 2366
rect 135 2332 151 2366
rect 203 2332 219 2366
rect 253 2332 269 2366
rect 321 2332 337 2366
rect 371 2332 387 2366
rect 439 2332 455 2366
rect 489 2332 505 2366
rect 557 2332 573 2366
rect 607 2332 623 2366
rect 675 2332 691 2366
rect 725 2332 741 2366
rect 793 2332 809 2366
rect 843 2332 859 2366
rect 911 2332 927 2366
rect 961 2332 977 2366
rect 1029 2332 1045 2366
rect 1079 2332 1095 2366
rect 1147 2332 1163 2366
rect 1197 2332 1213 2366
rect 1265 2332 1281 2366
rect 1315 2332 1331 2366
rect 1383 2332 1399 2366
rect 1433 2332 1449 2366
rect -1492 2236 -1458 2252
rect -1492 1644 -1458 1660
rect -1374 2236 -1340 2252
rect -1374 1644 -1340 1660
rect -1256 2236 -1222 2252
rect -1256 1644 -1222 1660
rect -1138 2236 -1104 2252
rect -1138 1644 -1104 1660
rect -1020 2236 -986 2252
rect -1020 1644 -986 1660
rect -902 2236 -868 2252
rect -902 1644 -868 1660
rect -784 2236 -750 2252
rect -784 1644 -750 1660
rect -666 2236 -632 2252
rect -666 1644 -632 1660
rect -548 2236 -514 2252
rect -548 1644 -514 1660
rect -430 2236 -396 2252
rect -430 1644 -396 1660
rect -312 2236 -278 2252
rect -312 1644 -278 1660
rect -194 2236 -160 2252
rect -194 1644 -160 1660
rect -76 2236 -42 2252
rect -76 1644 -42 1660
rect 42 2236 76 2252
rect 42 1644 76 1660
rect 160 2236 194 2252
rect 160 1644 194 1660
rect 278 2236 312 2252
rect 278 1644 312 1660
rect 396 2236 430 2252
rect 396 1644 430 1660
rect 514 2236 548 2252
rect 514 1644 548 1660
rect 632 2236 666 2252
rect 632 1644 666 1660
rect 750 2236 784 2252
rect 750 1644 784 1660
rect 868 2236 902 2252
rect 868 1644 902 1660
rect 986 2236 1020 2252
rect 986 1644 1020 1660
rect 1104 2236 1138 2252
rect 1104 1644 1138 1660
rect 1222 2236 1256 2252
rect 1222 1644 1256 1660
rect 1340 2236 1374 2252
rect 1340 1644 1374 1660
rect 1458 2236 1492 2252
rect 1458 1644 1492 1660
rect -1449 1567 -1433 1601
rect -1399 1567 -1383 1601
rect -1331 1567 -1315 1601
rect -1281 1567 -1265 1601
rect -1213 1567 -1197 1601
rect -1163 1567 -1147 1601
rect -1095 1567 -1079 1601
rect -1045 1567 -1029 1601
rect -977 1567 -961 1601
rect -927 1567 -911 1601
rect -859 1567 -843 1601
rect -809 1567 -793 1601
rect -741 1567 -725 1601
rect -691 1567 -675 1601
rect -623 1567 -607 1601
rect -573 1567 -557 1601
rect -505 1567 -489 1601
rect -455 1567 -439 1601
rect -387 1567 -371 1601
rect -337 1567 -321 1601
rect -269 1567 -253 1601
rect -219 1567 -203 1601
rect -151 1567 -135 1601
rect -101 1567 -85 1601
rect -33 1567 -17 1601
rect 17 1567 33 1601
rect 85 1567 101 1601
rect 135 1567 151 1601
rect 203 1567 219 1601
rect 253 1567 269 1601
rect 321 1567 337 1601
rect 371 1567 387 1601
rect 439 1567 455 1601
rect 489 1567 505 1601
rect 557 1567 573 1601
rect 607 1567 623 1601
rect 675 1567 691 1601
rect 725 1567 741 1601
rect 793 1567 809 1601
rect 843 1567 859 1601
rect 911 1567 927 1601
rect 961 1567 977 1601
rect 1029 1567 1045 1601
rect 1079 1567 1095 1601
rect 1147 1567 1163 1601
rect 1197 1567 1213 1601
rect 1265 1567 1281 1601
rect 1315 1567 1331 1601
rect 1383 1567 1399 1601
rect 1433 1567 1449 1601
rect -1492 1471 -1458 1487
rect -1492 879 -1458 895
rect -1374 1471 -1340 1487
rect -1374 879 -1340 895
rect -1256 1471 -1222 1487
rect -1256 879 -1222 895
rect -1138 1471 -1104 1487
rect -1138 879 -1104 895
rect -1020 1471 -986 1487
rect -1020 879 -986 895
rect -902 1471 -868 1487
rect -902 879 -868 895
rect -784 1471 -750 1487
rect -784 879 -750 895
rect -666 1471 -632 1487
rect -666 879 -632 895
rect -548 1471 -514 1487
rect -548 879 -514 895
rect -430 1471 -396 1487
rect -430 879 -396 895
rect -312 1471 -278 1487
rect -312 879 -278 895
rect -194 1471 -160 1487
rect -194 879 -160 895
rect -76 1471 -42 1487
rect -76 879 -42 895
rect 42 1471 76 1487
rect 42 879 76 895
rect 160 1471 194 1487
rect 160 879 194 895
rect 278 1471 312 1487
rect 278 879 312 895
rect 396 1471 430 1487
rect 396 879 430 895
rect 514 1471 548 1487
rect 514 879 548 895
rect 632 1471 666 1487
rect 632 879 666 895
rect 750 1471 784 1487
rect 750 879 784 895
rect 868 1471 902 1487
rect 868 879 902 895
rect 986 1471 1020 1487
rect 986 879 1020 895
rect 1104 1471 1138 1487
rect 1104 879 1138 895
rect 1222 1471 1256 1487
rect 1222 879 1256 895
rect 1340 1471 1374 1487
rect 1340 879 1374 895
rect 1458 1471 1492 1487
rect 1458 879 1492 895
rect -1449 802 -1433 836
rect -1399 802 -1383 836
rect -1331 802 -1315 836
rect -1281 802 -1265 836
rect -1213 802 -1197 836
rect -1163 802 -1147 836
rect -1095 802 -1079 836
rect -1045 802 -1029 836
rect -977 802 -961 836
rect -927 802 -911 836
rect -859 802 -843 836
rect -809 802 -793 836
rect -741 802 -725 836
rect -691 802 -675 836
rect -623 802 -607 836
rect -573 802 -557 836
rect -505 802 -489 836
rect -455 802 -439 836
rect -387 802 -371 836
rect -337 802 -321 836
rect -269 802 -253 836
rect -219 802 -203 836
rect -151 802 -135 836
rect -101 802 -85 836
rect -33 802 -17 836
rect 17 802 33 836
rect 85 802 101 836
rect 135 802 151 836
rect 203 802 219 836
rect 253 802 269 836
rect 321 802 337 836
rect 371 802 387 836
rect 439 802 455 836
rect 489 802 505 836
rect 557 802 573 836
rect 607 802 623 836
rect 675 802 691 836
rect 725 802 741 836
rect 793 802 809 836
rect 843 802 859 836
rect 911 802 927 836
rect 961 802 977 836
rect 1029 802 1045 836
rect 1079 802 1095 836
rect 1147 802 1163 836
rect 1197 802 1213 836
rect 1265 802 1281 836
rect 1315 802 1331 836
rect 1383 802 1399 836
rect 1433 802 1449 836
rect -1492 706 -1458 722
rect -1492 114 -1458 130
rect -1374 706 -1340 722
rect -1374 114 -1340 130
rect -1256 706 -1222 722
rect -1256 114 -1222 130
rect -1138 706 -1104 722
rect -1138 114 -1104 130
rect -1020 706 -986 722
rect -1020 114 -986 130
rect -902 706 -868 722
rect -902 114 -868 130
rect -784 706 -750 722
rect -784 114 -750 130
rect -666 706 -632 722
rect -666 114 -632 130
rect -548 706 -514 722
rect -548 114 -514 130
rect -430 706 -396 722
rect -430 114 -396 130
rect -312 706 -278 722
rect -312 114 -278 130
rect -194 706 -160 722
rect -194 114 -160 130
rect -76 706 -42 722
rect -76 114 -42 130
rect 42 706 76 722
rect 42 114 76 130
rect 160 706 194 722
rect 160 114 194 130
rect 278 706 312 722
rect 278 114 312 130
rect 396 706 430 722
rect 396 114 430 130
rect 514 706 548 722
rect 514 114 548 130
rect 632 706 666 722
rect 632 114 666 130
rect 750 706 784 722
rect 750 114 784 130
rect 868 706 902 722
rect 868 114 902 130
rect 986 706 1020 722
rect 986 114 1020 130
rect 1104 706 1138 722
rect 1104 114 1138 130
rect 1222 706 1256 722
rect 1222 114 1256 130
rect 1340 706 1374 722
rect 1340 114 1374 130
rect 1458 706 1492 722
rect 1458 114 1492 130
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -977 37 -961 71
rect -927 37 -911 71
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect 911 37 927 71
rect 961 37 977 71
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1383 37 1399 71
rect 1433 37 1449 71
rect -1492 -59 -1458 -43
rect -1492 -651 -1458 -635
rect -1374 -59 -1340 -43
rect -1374 -651 -1340 -635
rect -1256 -59 -1222 -43
rect -1256 -651 -1222 -635
rect -1138 -59 -1104 -43
rect -1138 -651 -1104 -635
rect -1020 -59 -986 -43
rect -1020 -651 -986 -635
rect -902 -59 -868 -43
rect -902 -651 -868 -635
rect -784 -59 -750 -43
rect -784 -651 -750 -635
rect -666 -59 -632 -43
rect -666 -651 -632 -635
rect -548 -59 -514 -43
rect -548 -651 -514 -635
rect -430 -59 -396 -43
rect -430 -651 -396 -635
rect -312 -59 -278 -43
rect -312 -651 -278 -635
rect -194 -59 -160 -43
rect -194 -651 -160 -635
rect -76 -59 -42 -43
rect -76 -651 -42 -635
rect 42 -59 76 -43
rect 42 -651 76 -635
rect 160 -59 194 -43
rect 160 -651 194 -635
rect 278 -59 312 -43
rect 278 -651 312 -635
rect 396 -59 430 -43
rect 396 -651 430 -635
rect 514 -59 548 -43
rect 514 -651 548 -635
rect 632 -59 666 -43
rect 632 -651 666 -635
rect 750 -59 784 -43
rect 750 -651 784 -635
rect 868 -59 902 -43
rect 868 -651 902 -635
rect 986 -59 1020 -43
rect 986 -651 1020 -635
rect 1104 -59 1138 -43
rect 1104 -651 1138 -635
rect 1222 -59 1256 -43
rect 1222 -651 1256 -635
rect 1340 -59 1374 -43
rect 1340 -651 1374 -635
rect 1458 -59 1492 -43
rect 1458 -651 1492 -635
rect -1449 -728 -1433 -694
rect -1399 -728 -1383 -694
rect -1331 -728 -1315 -694
rect -1281 -728 -1265 -694
rect -1213 -728 -1197 -694
rect -1163 -728 -1147 -694
rect -1095 -728 -1079 -694
rect -1045 -728 -1029 -694
rect -977 -728 -961 -694
rect -927 -728 -911 -694
rect -859 -728 -843 -694
rect -809 -728 -793 -694
rect -741 -728 -725 -694
rect -691 -728 -675 -694
rect -623 -728 -607 -694
rect -573 -728 -557 -694
rect -505 -728 -489 -694
rect -455 -728 -439 -694
rect -387 -728 -371 -694
rect -337 -728 -321 -694
rect -269 -728 -253 -694
rect -219 -728 -203 -694
rect -151 -728 -135 -694
rect -101 -728 -85 -694
rect -33 -728 -17 -694
rect 17 -728 33 -694
rect 85 -728 101 -694
rect 135 -728 151 -694
rect 203 -728 219 -694
rect 253 -728 269 -694
rect 321 -728 337 -694
rect 371 -728 387 -694
rect 439 -728 455 -694
rect 489 -728 505 -694
rect 557 -728 573 -694
rect 607 -728 623 -694
rect 675 -728 691 -694
rect 725 -728 741 -694
rect 793 -728 809 -694
rect 843 -728 859 -694
rect 911 -728 927 -694
rect 961 -728 977 -694
rect 1029 -728 1045 -694
rect 1079 -728 1095 -694
rect 1147 -728 1163 -694
rect 1197 -728 1213 -694
rect 1265 -728 1281 -694
rect 1315 -728 1331 -694
rect 1383 -728 1399 -694
rect 1433 -728 1449 -694
rect -1492 -824 -1458 -808
rect -1492 -1416 -1458 -1400
rect -1374 -824 -1340 -808
rect -1374 -1416 -1340 -1400
rect -1256 -824 -1222 -808
rect -1256 -1416 -1222 -1400
rect -1138 -824 -1104 -808
rect -1138 -1416 -1104 -1400
rect -1020 -824 -986 -808
rect -1020 -1416 -986 -1400
rect -902 -824 -868 -808
rect -902 -1416 -868 -1400
rect -784 -824 -750 -808
rect -784 -1416 -750 -1400
rect -666 -824 -632 -808
rect -666 -1416 -632 -1400
rect -548 -824 -514 -808
rect -548 -1416 -514 -1400
rect -430 -824 -396 -808
rect -430 -1416 -396 -1400
rect -312 -824 -278 -808
rect -312 -1416 -278 -1400
rect -194 -824 -160 -808
rect -194 -1416 -160 -1400
rect -76 -824 -42 -808
rect -76 -1416 -42 -1400
rect 42 -824 76 -808
rect 42 -1416 76 -1400
rect 160 -824 194 -808
rect 160 -1416 194 -1400
rect 278 -824 312 -808
rect 278 -1416 312 -1400
rect 396 -824 430 -808
rect 396 -1416 430 -1400
rect 514 -824 548 -808
rect 514 -1416 548 -1400
rect 632 -824 666 -808
rect 632 -1416 666 -1400
rect 750 -824 784 -808
rect 750 -1416 784 -1400
rect 868 -824 902 -808
rect 868 -1416 902 -1400
rect 986 -824 1020 -808
rect 986 -1416 1020 -1400
rect 1104 -824 1138 -808
rect 1104 -1416 1138 -1400
rect 1222 -824 1256 -808
rect 1222 -1416 1256 -1400
rect 1340 -824 1374 -808
rect 1340 -1416 1374 -1400
rect 1458 -824 1492 -808
rect 1458 -1416 1492 -1400
rect -1449 -1493 -1433 -1459
rect -1399 -1493 -1383 -1459
rect -1331 -1493 -1315 -1459
rect -1281 -1493 -1265 -1459
rect -1213 -1493 -1197 -1459
rect -1163 -1493 -1147 -1459
rect -1095 -1493 -1079 -1459
rect -1045 -1493 -1029 -1459
rect -977 -1493 -961 -1459
rect -927 -1493 -911 -1459
rect -859 -1493 -843 -1459
rect -809 -1493 -793 -1459
rect -741 -1493 -725 -1459
rect -691 -1493 -675 -1459
rect -623 -1493 -607 -1459
rect -573 -1493 -557 -1459
rect -505 -1493 -489 -1459
rect -455 -1493 -439 -1459
rect -387 -1493 -371 -1459
rect -337 -1493 -321 -1459
rect -269 -1493 -253 -1459
rect -219 -1493 -203 -1459
rect -151 -1493 -135 -1459
rect -101 -1493 -85 -1459
rect -33 -1493 -17 -1459
rect 17 -1493 33 -1459
rect 85 -1493 101 -1459
rect 135 -1493 151 -1459
rect 203 -1493 219 -1459
rect 253 -1493 269 -1459
rect 321 -1493 337 -1459
rect 371 -1493 387 -1459
rect 439 -1493 455 -1459
rect 489 -1493 505 -1459
rect 557 -1493 573 -1459
rect 607 -1493 623 -1459
rect 675 -1493 691 -1459
rect 725 -1493 741 -1459
rect 793 -1493 809 -1459
rect 843 -1493 859 -1459
rect 911 -1493 927 -1459
rect 961 -1493 977 -1459
rect 1029 -1493 1045 -1459
rect 1079 -1493 1095 -1459
rect 1147 -1493 1163 -1459
rect 1197 -1493 1213 -1459
rect 1265 -1493 1281 -1459
rect 1315 -1493 1331 -1459
rect 1383 -1493 1399 -1459
rect 1433 -1493 1449 -1459
rect -1492 -1589 -1458 -1573
rect -1492 -2181 -1458 -2165
rect -1374 -1589 -1340 -1573
rect -1374 -2181 -1340 -2165
rect -1256 -1589 -1222 -1573
rect -1256 -2181 -1222 -2165
rect -1138 -1589 -1104 -1573
rect -1138 -2181 -1104 -2165
rect -1020 -1589 -986 -1573
rect -1020 -2181 -986 -2165
rect -902 -1589 -868 -1573
rect -902 -2181 -868 -2165
rect -784 -1589 -750 -1573
rect -784 -2181 -750 -2165
rect -666 -1589 -632 -1573
rect -666 -2181 -632 -2165
rect -548 -1589 -514 -1573
rect -548 -2181 -514 -2165
rect -430 -1589 -396 -1573
rect -430 -2181 -396 -2165
rect -312 -1589 -278 -1573
rect -312 -2181 -278 -2165
rect -194 -1589 -160 -1573
rect -194 -2181 -160 -2165
rect -76 -1589 -42 -1573
rect -76 -2181 -42 -2165
rect 42 -1589 76 -1573
rect 42 -2181 76 -2165
rect 160 -1589 194 -1573
rect 160 -2181 194 -2165
rect 278 -1589 312 -1573
rect 278 -2181 312 -2165
rect 396 -1589 430 -1573
rect 396 -2181 430 -2165
rect 514 -1589 548 -1573
rect 514 -2181 548 -2165
rect 632 -1589 666 -1573
rect 632 -2181 666 -2165
rect 750 -1589 784 -1573
rect 750 -2181 784 -2165
rect 868 -1589 902 -1573
rect 868 -2181 902 -2165
rect 986 -1589 1020 -1573
rect 986 -2181 1020 -2165
rect 1104 -1589 1138 -1573
rect 1104 -2181 1138 -2165
rect 1222 -1589 1256 -1573
rect 1222 -2181 1256 -2165
rect 1340 -1589 1374 -1573
rect 1340 -2181 1374 -2165
rect 1458 -1589 1492 -1573
rect 1458 -2181 1492 -2165
rect -1449 -2258 -1433 -2224
rect -1399 -2258 -1383 -2224
rect -1331 -2258 -1315 -2224
rect -1281 -2258 -1265 -2224
rect -1213 -2258 -1197 -2224
rect -1163 -2258 -1147 -2224
rect -1095 -2258 -1079 -2224
rect -1045 -2258 -1029 -2224
rect -977 -2258 -961 -2224
rect -927 -2258 -911 -2224
rect -859 -2258 -843 -2224
rect -809 -2258 -793 -2224
rect -741 -2258 -725 -2224
rect -691 -2258 -675 -2224
rect -623 -2258 -607 -2224
rect -573 -2258 -557 -2224
rect -505 -2258 -489 -2224
rect -455 -2258 -439 -2224
rect -387 -2258 -371 -2224
rect -337 -2258 -321 -2224
rect -269 -2258 -253 -2224
rect -219 -2258 -203 -2224
rect -151 -2258 -135 -2224
rect -101 -2258 -85 -2224
rect -33 -2258 -17 -2224
rect 17 -2258 33 -2224
rect 85 -2258 101 -2224
rect 135 -2258 151 -2224
rect 203 -2258 219 -2224
rect 253 -2258 269 -2224
rect 321 -2258 337 -2224
rect 371 -2258 387 -2224
rect 439 -2258 455 -2224
rect 489 -2258 505 -2224
rect 557 -2258 573 -2224
rect 607 -2258 623 -2224
rect 675 -2258 691 -2224
rect 725 -2258 741 -2224
rect 793 -2258 809 -2224
rect 843 -2258 859 -2224
rect 911 -2258 927 -2224
rect 961 -2258 977 -2224
rect 1029 -2258 1045 -2224
rect 1079 -2258 1095 -2224
rect 1147 -2258 1163 -2224
rect 1197 -2258 1213 -2224
rect 1265 -2258 1281 -2224
rect 1315 -2258 1331 -2224
rect 1383 -2258 1399 -2224
rect 1433 -2258 1449 -2224
rect -1492 -2354 -1458 -2338
rect -1492 -2946 -1458 -2930
rect -1374 -2354 -1340 -2338
rect -1374 -2946 -1340 -2930
rect -1256 -2354 -1222 -2338
rect -1256 -2946 -1222 -2930
rect -1138 -2354 -1104 -2338
rect -1138 -2946 -1104 -2930
rect -1020 -2354 -986 -2338
rect -1020 -2946 -986 -2930
rect -902 -2354 -868 -2338
rect -902 -2946 -868 -2930
rect -784 -2354 -750 -2338
rect -784 -2946 -750 -2930
rect -666 -2354 -632 -2338
rect -666 -2946 -632 -2930
rect -548 -2354 -514 -2338
rect -548 -2946 -514 -2930
rect -430 -2354 -396 -2338
rect -430 -2946 -396 -2930
rect -312 -2354 -278 -2338
rect -312 -2946 -278 -2930
rect -194 -2354 -160 -2338
rect -194 -2946 -160 -2930
rect -76 -2354 -42 -2338
rect -76 -2946 -42 -2930
rect 42 -2354 76 -2338
rect 42 -2946 76 -2930
rect 160 -2354 194 -2338
rect 160 -2946 194 -2930
rect 278 -2354 312 -2338
rect 278 -2946 312 -2930
rect 396 -2354 430 -2338
rect 396 -2946 430 -2930
rect 514 -2354 548 -2338
rect 514 -2946 548 -2930
rect 632 -2354 666 -2338
rect 632 -2946 666 -2930
rect 750 -2354 784 -2338
rect 750 -2946 784 -2930
rect 868 -2354 902 -2338
rect 868 -2946 902 -2930
rect 986 -2354 1020 -2338
rect 986 -2946 1020 -2930
rect 1104 -2354 1138 -2338
rect 1104 -2946 1138 -2930
rect 1222 -2354 1256 -2338
rect 1222 -2946 1256 -2930
rect 1340 -2354 1374 -2338
rect 1340 -2946 1374 -2930
rect 1458 -2354 1492 -2338
rect 1458 -2946 1492 -2930
rect -1449 -3023 -1433 -2989
rect -1399 -3023 -1383 -2989
rect -1331 -3023 -1315 -2989
rect -1281 -3023 -1265 -2989
rect -1213 -3023 -1197 -2989
rect -1163 -3023 -1147 -2989
rect -1095 -3023 -1079 -2989
rect -1045 -3023 -1029 -2989
rect -977 -3023 -961 -2989
rect -927 -3023 -911 -2989
rect -859 -3023 -843 -2989
rect -809 -3023 -793 -2989
rect -741 -3023 -725 -2989
rect -691 -3023 -675 -2989
rect -623 -3023 -607 -2989
rect -573 -3023 -557 -2989
rect -505 -3023 -489 -2989
rect -455 -3023 -439 -2989
rect -387 -3023 -371 -2989
rect -337 -3023 -321 -2989
rect -269 -3023 -253 -2989
rect -219 -3023 -203 -2989
rect -151 -3023 -135 -2989
rect -101 -3023 -85 -2989
rect -33 -3023 -17 -2989
rect 17 -3023 33 -2989
rect 85 -3023 101 -2989
rect 135 -3023 151 -2989
rect 203 -3023 219 -2989
rect 253 -3023 269 -2989
rect 321 -3023 337 -2989
rect 371 -3023 387 -2989
rect 439 -3023 455 -2989
rect 489 -3023 505 -2989
rect 557 -3023 573 -2989
rect 607 -3023 623 -2989
rect 675 -3023 691 -2989
rect 725 -3023 741 -2989
rect 793 -3023 809 -2989
rect 843 -3023 859 -2989
rect 911 -3023 927 -2989
rect 961 -3023 977 -2989
rect 1029 -3023 1045 -2989
rect 1079 -3023 1095 -2989
rect 1147 -3023 1163 -2989
rect 1197 -3023 1213 -2989
rect 1265 -3023 1281 -2989
rect 1315 -3023 1331 -2989
rect 1383 -3023 1399 -2989
rect 1433 -3023 1449 -2989
rect -1492 -3119 -1458 -3103
rect -1492 -3711 -1458 -3695
rect -1374 -3119 -1340 -3103
rect -1374 -3711 -1340 -3695
rect -1256 -3119 -1222 -3103
rect -1256 -3711 -1222 -3695
rect -1138 -3119 -1104 -3103
rect -1138 -3711 -1104 -3695
rect -1020 -3119 -986 -3103
rect -1020 -3711 -986 -3695
rect -902 -3119 -868 -3103
rect -902 -3711 -868 -3695
rect -784 -3119 -750 -3103
rect -784 -3711 -750 -3695
rect -666 -3119 -632 -3103
rect -666 -3711 -632 -3695
rect -548 -3119 -514 -3103
rect -548 -3711 -514 -3695
rect -430 -3119 -396 -3103
rect -430 -3711 -396 -3695
rect -312 -3119 -278 -3103
rect -312 -3711 -278 -3695
rect -194 -3119 -160 -3103
rect -194 -3711 -160 -3695
rect -76 -3119 -42 -3103
rect -76 -3711 -42 -3695
rect 42 -3119 76 -3103
rect 42 -3711 76 -3695
rect 160 -3119 194 -3103
rect 160 -3711 194 -3695
rect 278 -3119 312 -3103
rect 278 -3711 312 -3695
rect 396 -3119 430 -3103
rect 396 -3711 430 -3695
rect 514 -3119 548 -3103
rect 514 -3711 548 -3695
rect 632 -3119 666 -3103
rect 632 -3711 666 -3695
rect 750 -3119 784 -3103
rect 750 -3711 784 -3695
rect 868 -3119 902 -3103
rect 868 -3711 902 -3695
rect 986 -3119 1020 -3103
rect 986 -3711 1020 -3695
rect 1104 -3119 1138 -3103
rect 1104 -3711 1138 -3695
rect 1222 -3119 1256 -3103
rect 1222 -3711 1256 -3695
rect 1340 -3119 1374 -3103
rect 1340 -3711 1374 -3695
rect 1458 -3119 1492 -3103
rect 1458 -3711 1492 -3695
rect -1449 -3788 -1433 -3754
rect -1399 -3788 -1383 -3754
rect -1331 -3788 -1315 -3754
rect -1281 -3788 -1265 -3754
rect -1213 -3788 -1197 -3754
rect -1163 -3788 -1147 -3754
rect -1095 -3788 -1079 -3754
rect -1045 -3788 -1029 -3754
rect -977 -3788 -961 -3754
rect -927 -3788 -911 -3754
rect -859 -3788 -843 -3754
rect -809 -3788 -793 -3754
rect -741 -3788 -725 -3754
rect -691 -3788 -675 -3754
rect -623 -3788 -607 -3754
rect -573 -3788 -557 -3754
rect -505 -3788 -489 -3754
rect -455 -3788 -439 -3754
rect -387 -3788 -371 -3754
rect -337 -3788 -321 -3754
rect -269 -3788 -253 -3754
rect -219 -3788 -203 -3754
rect -151 -3788 -135 -3754
rect -101 -3788 -85 -3754
rect -33 -3788 -17 -3754
rect 17 -3788 33 -3754
rect 85 -3788 101 -3754
rect 135 -3788 151 -3754
rect 203 -3788 219 -3754
rect 253 -3788 269 -3754
rect 321 -3788 337 -3754
rect 371 -3788 387 -3754
rect 439 -3788 455 -3754
rect 489 -3788 505 -3754
rect 557 -3788 573 -3754
rect 607 -3788 623 -3754
rect 675 -3788 691 -3754
rect 725 -3788 741 -3754
rect 793 -3788 809 -3754
rect 843 -3788 859 -3754
rect 911 -3788 927 -3754
rect 961 -3788 977 -3754
rect 1029 -3788 1045 -3754
rect 1079 -3788 1095 -3754
rect 1147 -3788 1163 -3754
rect 1197 -3788 1213 -3754
rect 1265 -3788 1281 -3754
rect 1315 -3788 1331 -3754
rect 1383 -3788 1399 -3754
rect 1433 -3788 1449 -3754
rect -1606 -3856 -1572 -3794
rect 1572 -3856 1606 -3794
rect -1606 -3890 -1510 -3856
rect 1510 -3890 1606 -3856
<< viali >>
rect -1492 3190 -1458 3766
rect -1374 3190 -1340 3766
rect -1256 3190 -1222 3766
rect -1138 3190 -1104 3766
rect -1020 3190 -986 3766
rect -902 3190 -868 3766
rect -784 3190 -750 3766
rect -666 3190 -632 3766
rect -548 3190 -514 3766
rect -430 3190 -396 3766
rect -312 3190 -278 3766
rect -194 3190 -160 3766
rect -76 3190 -42 3766
rect 42 3190 76 3766
rect 160 3190 194 3766
rect 278 3190 312 3766
rect 396 3190 430 3766
rect 514 3190 548 3766
rect 632 3190 666 3766
rect 750 3190 784 3766
rect 868 3190 902 3766
rect 986 3190 1020 3766
rect 1104 3190 1138 3766
rect 1222 3190 1256 3766
rect 1340 3190 1374 3766
rect 1458 3190 1492 3766
rect -1433 3097 -1399 3131
rect -1315 3097 -1281 3131
rect -1197 3097 -1163 3131
rect -1079 3097 -1045 3131
rect -961 3097 -927 3131
rect -843 3097 -809 3131
rect -725 3097 -691 3131
rect -607 3097 -573 3131
rect -489 3097 -455 3131
rect -371 3097 -337 3131
rect -253 3097 -219 3131
rect -135 3097 -101 3131
rect -17 3097 17 3131
rect 101 3097 135 3131
rect 219 3097 253 3131
rect 337 3097 371 3131
rect 455 3097 489 3131
rect 573 3097 607 3131
rect 691 3097 725 3131
rect 809 3097 843 3131
rect 927 3097 961 3131
rect 1045 3097 1079 3131
rect 1163 3097 1197 3131
rect 1281 3097 1315 3131
rect 1399 3097 1433 3131
rect -1492 2425 -1458 3001
rect -1374 2425 -1340 3001
rect -1256 2425 -1222 3001
rect -1138 2425 -1104 3001
rect -1020 2425 -986 3001
rect -902 2425 -868 3001
rect -784 2425 -750 3001
rect -666 2425 -632 3001
rect -548 2425 -514 3001
rect -430 2425 -396 3001
rect -312 2425 -278 3001
rect -194 2425 -160 3001
rect -76 2425 -42 3001
rect 42 2425 76 3001
rect 160 2425 194 3001
rect 278 2425 312 3001
rect 396 2425 430 3001
rect 514 2425 548 3001
rect 632 2425 666 3001
rect 750 2425 784 3001
rect 868 2425 902 3001
rect 986 2425 1020 3001
rect 1104 2425 1138 3001
rect 1222 2425 1256 3001
rect 1340 2425 1374 3001
rect 1458 2425 1492 3001
rect -1433 2332 -1399 2366
rect -1315 2332 -1281 2366
rect -1197 2332 -1163 2366
rect -1079 2332 -1045 2366
rect -961 2332 -927 2366
rect -843 2332 -809 2366
rect -725 2332 -691 2366
rect -607 2332 -573 2366
rect -489 2332 -455 2366
rect -371 2332 -337 2366
rect -253 2332 -219 2366
rect -135 2332 -101 2366
rect -17 2332 17 2366
rect 101 2332 135 2366
rect 219 2332 253 2366
rect 337 2332 371 2366
rect 455 2332 489 2366
rect 573 2332 607 2366
rect 691 2332 725 2366
rect 809 2332 843 2366
rect 927 2332 961 2366
rect 1045 2332 1079 2366
rect 1163 2332 1197 2366
rect 1281 2332 1315 2366
rect 1399 2332 1433 2366
rect -1492 1660 -1458 2236
rect -1374 1660 -1340 2236
rect -1256 1660 -1222 2236
rect -1138 1660 -1104 2236
rect -1020 1660 -986 2236
rect -902 1660 -868 2236
rect -784 1660 -750 2236
rect -666 1660 -632 2236
rect -548 1660 -514 2236
rect -430 1660 -396 2236
rect -312 1660 -278 2236
rect -194 1660 -160 2236
rect -76 1660 -42 2236
rect 42 1660 76 2236
rect 160 1660 194 2236
rect 278 1660 312 2236
rect 396 1660 430 2236
rect 514 1660 548 2236
rect 632 1660 666 2236
rect 750 1660 784 2236
rect 868 1660 902 2236
rect 986 1660 1020 2236
rect 1104 1660 1138 2236
rect 1222 1660 1256 2236
rect 1340 1660 1374 2236
rect 1458 1660 1492 2236
rect -1433 1567 -1399 1601
rect -1315 1567 -1281 1601
rect -1197 1567 -1163 1601
rect -1079 1567 -1045 1601
rect -961 1567 -927 1601
rect -843 1567 -809 1601
rect -725 1567 -691 1601
rect -607 1567 -573 1601
rect -489 1567 -455 1601
rect -371 1567 -337 1601
rect -253 1567 -219 1601
rect -135 1567 -101 1601
rect -17 1567 17 1601
rect 101 1567 135 1601
rect 219 1567 253 1601
rect 337 1567 371 1601
rect 455 1567 489 1601
rect 573 1567 607 1601
rect 691 1567 725 1601
rect 809 1567 843 1601
rect 927 1567 961 1601
rect 1045 1567 1079 1601
rect 1163 1567 1197 1601
rect 1281 1567 1315 1601
rect 1399 1567 1433 1601
rect -1492 895 -1458 1471
rect -1374 895 -1340 1471
rect -1256 895 -1222 1471
rect -1138 895 -1104 1471
rect -1020 895 -986 1471
rect -902 895 -868 1471
rect -784 895 -750 1471
rect -666 895 -632 1471
rect -548 895 -514 1471
rect -430 895 -396 1471
rect -312 895 -278 1471
rect -194 895 -160 1471
rect -76 895 -42 1471
rect 42 895 76 1471
rect 160 895 194 1471
rect 278 895 312 1471
rect 396 895 430 1471
rect 514 895 548 1471
rect 632 895 666 1471
rect 750 895 784 1471
rect 868 895 902 1471
rect 986 895 1020 1471
rect 1104 895 1138 1471
rect 1222 895 1256 1471
rect 1340 895 1374 1471
rect 1458 895 1492 1471
rect -1433 802 -1399 836
rect -1315 802 -1281 836
rect -1197 802 -1163 836
rect -1079 802 -1045 836
rect -961 802 -927 836
rect -843 802 -809 836
rect -725 802 -691 836
rect -607 802 -573 836
rect -489 802 -455 836
rect -371 802 -337 836
rect -253 802 -219 836
rect -135 802 -101 836
rect -17 802 17 836
rect 101 802 135 836
rect 219 802 253 836
rect 337 802 371 836
rect 455 802 489 836
rect 573 802 607 836
rect 691 802 725 836
rect 809 802 843 836
rect 927 802 961 836
rect 1045 802 1079 836
rect 1163 802 1197 836
rect 1281 802 1315 836
rect 1399 802 1433 836
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1492 -635 -1458 -59
rect -1374 -635 -1340 -59
rect -1256 -635 -1222 -59
rect -1138 -635 -1104 -59
rect -1020 -635 -986 -59
rect -902 -635 -868 -59
rect -784 -635 -750 -59
rect -666 -635 -632 -59
rect -548 -635 -514 -59
rect -430 -635 -396 -59
rect -312 -635 -278 -59
rect -194 -635 -160 -59
rect -76 -635 -42 -59
rect 42 -635 76 -59
rect 160 -635 194 -59
rect 278 -635 312 -59
rect 396 -635 430 -59
rect 514 -635 548 -59
rect 632 -635 666 -59
rect 750 -635 784 -59
rect 868 -635 902 -59
rect 986 -635 1020 -59
rect 1104 -635 1138 -59
rect 1222 -635 1256 -59
rect 1340 -635 1374 -59
rect 1458 -635 1492 -59
rect -1433 -728 -1399 -694
rect -1315 -728 -1281 -694
rect -1197 -728 -1163 -694
rect -1079 -728 -1045 -694
rect -961 -728 -927 -694
rect -843 -728 -809 -694
rect -725 -728 -691 -694
rect -607 -728 -573 -694
rect -489 -728 -455 -694
rect -371 -728 -337 -694
rect -253 -728 -219 -694
rect -135 -728 -101 -694
rect -17 -728 17 -694
rect 101 -728 135 -694
rect 219 -728 253 -694
rect 337 -728 371 -694
rect 455 -728 489 -694
rect 573 -728 607 -694
rect 691 -728 725 -694
rect 809 -728 843 -694
rect 927 -728 961 -694
rect 1045 -728 1079 -694
rect 1163 -728 1197 -694
rect 1281 -728 1315 -694
rect 1399 -728 1433 -694
rect -1492 -1400 -1458 -824
rect -1374 -1400 -1340 -824
rect -1256 -1400 -1222 -824
rect -1138 -1400 -1104 -824
rect -1020 -1400 -986 -824
rect -902 -1400 -868 -824
rect -784 -1400 -750 -824
rect -666 -1400 -632 -824
rect -548 -1400 -514 -824
rect -430 -1400 -396 -824
rect -312 -1400 -278 -824
rect -194 -1400 -160 -824
rect -76 -1400 -42 -824
rect 42 -1400 76 -824
rect 160 -1400 194 -824
rect 278 -1400 312 -824
rect 396 -1400 430 -824
rect 514 -1400 548 -824
rect 632 -1400 666 -824
rect 750 -1400 784 -824
rect 868 -1400 902 -824
rect 986 -1400 1020 -824
rect 1104 -1400 1138 -824
rect 1222 -1400 1256 -824
rect 1340 -1400 1374 -824
rect 1458 -1400 1492 -824
rect -1433 -1493 -1399 -1459
rect -1315 -1493 -1281 -1459
rect -1197 -1493 -1163 -1459
rect -1079 -1493 -1045 -1459
rect -961 -1493 -927 -1459
rect -843 -1493 -809 -1459
rect -725 -1493 -691 -1459
rect -607 -1493 -573 -1459
rect -489 -1493 -455 -1459
rect -371 -1493 -337 -1459
rect -253 -1493 -219 -1459
rect -135 -1493 -101 -1459
rect -17 -1493 17 -1459
rect 101 -1493 135 -1459
rect 219 -1493 253 -1459
rect 337 -1493 371 -1459
rect 455 -1493 489 -1459
rect 573 -1493 607 -1459
rect 691 -1493 725 -1459
rect 809 -1493 843 -1459
rect 927 -1493 961 -1459
rect 1045 -1493 1079 -1459
rect 1163 -1493 1197 -1459
rect 1281 -1493 1315 -1459
rect 1399 -1493 1433 -1459
rect -1492 -2165 -1458 -1589
rect -1374 -2165 -1340 -1589
rect -1256 -2165 -1222 -1589
rect -1138 -2165 -1104 -1589
rect -1020 -2165 -986 -1589
rect -902 -2165 -868 -1589
rect -784 -2165 -750 -1589
rect -666 -2165 -632 -1589
rect -548 -2165 -514 -1589
rect -430 -2165 -396 -1589
rect -312 -2165 -278 -1589
rect -194 -2165 -160 -1589
rect -76 -2165 -42 -1589
rect 42 -2165 76 -1589
rect 160 -2165 194 -1589
rect 278 -2165 312 -1589
rect 396 -2165 430 -1589
rect 514 -2165 548 -1589
rect 632 -2165 666 -1589
rect 750 -2165 784 -1589
rect 868 -2165 902 -1589
rect 986 -2165 1020 -1589
rect 1104 -2165 1138 -1589
rect 1222 -2165 1256 -1589
rect 1340 -2165 1374 -1589
rect 1458 -2165 1492 -1589
rect -1433 -2258 -1399 -2224
rect -1315 -2258 -1281 -2224
rect -1197 -2258 -1163 -2224
rect -1079 -2258 -1045 -2224
rect -961 -2258 -927 -2224
rect -843 -2258 -809 -2224
rect -725 -2258 -691 -2224
rect -607 -2258 -573 -2224
rect -489 -2258 -455 -2224
rect -371 -2258 -337 -2224
rect -253 -2258 -219 -2224
rect -135 -2258 -101 -2224
rect -17 -2258 17 -2224
rect 101 -2258 135 -2224
rect 219 -2258 253 -2224
rect 337 -2258 371 -2224
rect 455 -2258 489 -2224
rect 573 -2258 607 -2224
rect 691 -2258 725 -2224
rect 809 -2258 843 -2224
rect 927 -2258 961 -2224
rect 1045 -2258 1079 -2224
rect 1163 -2258 1197 -2224
rect 1281 -2258 1315 -2224
rect 1399 -2258 1433 -2224
rect -1492 -2930 -1458 -2354
rect -1374 -2930 -1340 -2354
rect -1256 -2930 -1222 -2354
rect -1138 -2930 -1104 -2354
rect -1020 -2930 -986 -2354
rect -902 -2930 -868 -2354
rect -784 -2930 -750 -2354
rect -666 -2930 -632 -2354
rect -548 -2930 -514 -2354
rect -430 -2930 -396 -2354
rect -312 -2930 -278 -2354
rect -194 -2930 -160 -2354
rect -76 -2930 -42 -2354
rect 42 -2930 76 -2354
rect 160 -2930 194 -2354
rect 278 -2930 312 -2354
rect 396 -2930 430 -2354
rect 514 -2930 548 -2354
rect 632 -2930 666 -2354
rect 750 -2930 784 -2354
rect 868 -2930 902 -2354
rect 986 -2930 1020 -2354
rect 1104 -2930 1138 -2354
rect 1222 -2930 1256 -2354
rect 1340 -2930 1374 -2354
rect 1458 -2930 1492 -2354
rect -1433 -3023 -1399 -2989
rect -1315 -3023 -1281 -2989
rect -1197 -3023 -1163 -2989
rect -1079 -3023 -1045 -2989
rect -961 -3023 -927 -2989
rect -843 -3023 -809 -2989
rect -725 -3023 -691 -2989
rect -607 -3023 -573 -2989
rect -489 -3023 -455 -2989
rect -371 -3023 -337 -2989
rect -253 -3023 -219 -2989
rect -135 -3023 -101 -2989
rect -17 -3023 17 -2989
rect 101 -3023 135 -2989
rect 219 -3023 253 -2989
rect 337 -3023 371 -2989
rect 455 -3023 489 -2989
rect 573 -3023 607 -2989
rect 691 -3023 725 -2989
rect 809 -3023 843 -2989
rect 927 -3023 961 -2989
rect 1045 -3023 1079 -2989
rect 1163 -3023 1197 -2989
rect 1281 -3023 1315 -2989
rect 1399 -3023 1433 -2989
rect -1492 -3695 -1458 -3119
rect -1374 -3695 -1340 -3119
rect -1256 -3695 -1222 -3119
rect -1138 -3695 -1104 -3119
rect -1020 -3695 -986 -3119
rect -902 -3695 -868 -3119
rect -784 -3695 -750 -3119
rect -666 -3695 -632 -3119
rect -548 -3695 -514 -3119
rect -430 -3695 -396 -3119
rect -312 -3695 -278 -3119
rect -194 -3695 -160 -3119
rect -76 -3695 -42 -3119
rect 42 -3695 76 -3119
rect 160 -3695 194 -3119
rect 278 -3695 312 -3119
rect 396 -3695 430 -3119
rect 514 -3695 548 -3119
rect 632 -3695 666 -3119
rect 750 -3695 784 -3119
rect 868 -3695 902 -3119
rect 986 -3695 1020 -3119
rect 1104 -3695 1138 -3119
rect 1222 -3695 1256 -3119
rect 1340 -3695 1374 -3119
rect 1458 -3695 1492 -3119
rect -1433 -3788 -1399 -3754
rect -1315 -3788 -1281 -3754
rect -1197 -3788 -1163 -3754
rect -1079 -3788 -1045 -3754
rect -961 -3788 -927 -3754
rect -843 -3788 -809 -3754
rect -725 -3788 -691 -3754
rect -607 -3788 -573 -3754
rect -489 -3788 -455 -3754
rect -371 -3788 -337 -3754
rect -253 -3788 -219 -3754
rect -135 -3788 -101 -3754
rect -17 -3788 17 -3754
rect 101 -3788 135 -3754
rect 219 -3788 253 -3754
rect 337 -3788 371 -3754
rect 455 -3788 489 -3754
rect 573 -3788 607 -3754
rect 691 -3788 725 -3754
rect 809 -3788 843 -3754
rect 927 -3788 961 -3754
rect 1045 -3788 1079 -3754
rect 1163 -3788 1197 -3754
rect 1281 -3788 1315 -3754
rect 1399 -3788 1433 -3754
<< metal1 >>
rect -1498 3766 -1452 3778
rect -1498 3190 -1492 3766
rect -1458 3190 -1452 3766
rect -1498 3178 -1452 3190
rect -1380 3766 -1334 3778
rect -1380 3190 -1374 3766
rect -1340 3190 -1334 3766
rect -1380 3178 -1334 3190
rect -1262 3766 -1216 3778
rect -1262 3190 -1256 3766
rect -1222 3190 -1216 3766
rect -1262 3178 -1216 3190
rect -1144 3766 -1098 3778
rect -1144 3190 -1138 3766
rect -1104 3190 -1098 3766
rect -1144 3178 -1098 3190
rect -1026 3766 -980 3778
rect -1026 3190 -1020 3766
rect -986 3190 -980 3766
rect -1026 3178 -980 3190
rect -908 3766 -862 3778
rect -908 3190 -902 3766
rect -868 3190 -862 3766
rect -908 3178 -862 3190
rect -790 3766 -744 3778
rect -790 3190 -784 3766
rect -750 3190 -744 3766
rect -790 3178 -744 3190
rect -672 3766 -626 3778
rect -672 3190 -666 3766
rect -632 3190 -626 3766
rect -672 3178 -626 3190
rect -554 3766 -508 3778
rect -554 3190 -548 3766
rect -514 3190 -508 3766
rect -554 3178 -508 3190
rect -436 3766 -390 3778
rect -436 3190 -430 3766
rect -396 3190 -390 3766
rect -436 3178 -390 3190
rect -318 3766 -272 3778
rect -318 3190 -312 3766
rect -278 3190 -272 3766
rect -318 3178 -272 3190
rect -200 3766 -154 3778
rect -200 3190 -194 3766
rect -160 3190 -154 3766
rect -200 3178 -154 3190
rect -82 3766 -36 3778
rect -82 3190 -76 3766
rect -42 3190 -36 3766
rect -82 3178 -36 3190
rect 36 3766 82 3778
rect 36 3190 42 3766
rect 76 3190 82 3766
rect 36 3178 82 3190
rect 154 3766 200 3778
rect 154 3190 160 3766
rect 194 3190 200 3766
rect 154 3178 200 3190
rect 272 3766 318 3778
rect 272 3190 278 3766
rect 312 3190 318 3766
rect 272 3178 318 3190
rect 390 3766 436 3778
rect 390 3190 396 3766
rect 430 3190 436 3766
rect 390 3178 436 3190
rect 508 3766 554 3778
rect 508 3190 514 3766
rect 548 3190 554 3766
rect 508 3178 554 3190
rect 626 3766 672 3778
rect 626 3190 632 3766
rect 666 3190 672 3766
rect 626 3178 672 3190
rect 744 3766 790 3778
rect 744 3190 750 3766
rect 784 3190 790 3766
rect 744 3178 790 3190
rect 862 3766 908 3778
rect 862 3190 868 3766
rect 902 3190 908 3766
rect 862 3178 908 3190
rect 980 3766 1026 3778
rect 980 3190 986 3766
rect 1020 3190 1026 3766
rect 980 3178 1026 3190
rect 1098 3766 1144 3778
rect 1098 3190 1104 3766
rect 1138 3190 1144 3766
rect 1098 3178 1144 3190
rect 1216 3766 1262 3778
rect 1216 3190 1222 3766
rect 1256 3190 1262 3766
rect 1216 3178 1262 3190
rect 1334 3766 1380 3778
rect 1334 3190 1340 3766
rect 1374 3190 1380 3766
rect 1334 3178 1380 3190
rect 1452 3766 1498 3778
rect 1452 3190 1458 3766
rect 1492 3190 1498 3766
rect 1452 3178 1498 3190
rect -1445 3131 -1387 3137
rect -1445 3097 -1433 3131
rect -1399 3097 -1387 3131
rect -1445 3091 -1387 3097
rect -1327 3131 -1269 3137
rect -1327 3097 -1315 3131
rect -1281 3097 -1269 3131
rect -1327 3091 -1269 3097
rect -1209 3131 -1151 3137
rect -1209 3097 -1197 3131
rect -1163 3097 -1151 3131
rect -1209 3091 -1151 3097
rect -1091 3131 -1033 3137
rect -1091 3097 -1079 3131
rect -1045 3097 -1033 3131
rect -1091 3091 -1033 3097
rect -973 3131 -915 3137
rect -973 3097 -961 3131
rect -927 3097 -915 3131
rect -973 3091 -915 3097
rect -855 3131 -797 3137
rect -855 3097 -843 3131
rect -809 3097 -797 3131
rect -855 3091 -797 3097
rect -737 3131 -679 3137
rect -737 3097 -725 3131
rect -691 3097 -679 3131
rect -737 3091 -679 3097
rect -619 3131 -561 3137
rect -619 3097 -607 3131
rect -573 3097 -561 3131
rect -619 3091 -561 3097
rect -501 3131 -443 3137
rect -501 3097 -489 3131
rect -455 3097 -443 3131
rect -501 3091 -443 3097
rect -383 3131 -325 3137
rect -383 3097 -371 3131
rect -337 3097 -325 3131
rect -383 3091 -325 3097
rect -265 3131 -207 3137
rect -265 3097 -253 3131
rect -219 3097 -207 3131
rect -265 3091 -207 3097
rect -147 3131 -89 3137
rect -147 3097 -135 3131
rect -101 3097 -89 3131
rect -147 3091 -89 3097
rect -29 3131 29 3137
rect -29 3097 -17 3131
rect 17 3097 29 3131
rect -29 3091 29 3097
rect 89 3131 147 3137
rect 89 3097 101 3131
rect 135 3097 147 3131
rect 89 3091 147 3097
rect 207 3131 265 3137
rect 207 3097 219 3131
rect 253 3097 265 3131
rect 207 3091 265 3097
rect 325 3131 383 3137
rect 325 3097 337 3131
rect 371 3097 383 3131
rect 325 3091 383 3097
rect 443 3131 501 3137
rect 443 3097 455 3131
rect 489 3097 501 3131
rect 443 3091 501 3097
rect 561 3131 619 3137
rect 561 3097 573 3131
rect 607 3097 619 3131
rect 561 3091 619 3097
rect 679 3131 737 3137
rect 679 3097 691 3131
rect 725 3097 737 3131
rect 679 3091 737 3097
rect 797 3131 855 3137
rect 797 3097 809 3131
rect 843 3097 855 3131
rect 797 3091 855 3097
rect 915 3131 973 3137
rect 915 3097 927 3131
rect 961 3097 973 3131
rect 915 3091 973 3097
rect 1033 3131 1091 3137
rect 1033 3097 1045 3131
rect 1079 3097 1091 3131
rect 1033 3091 1091 3097
rect 1151 3131 1209 3137
rect 1151 3097 1163 3131
rect 1197 3097 1209 3131
rect 1151 3091 1209 3097
rect 1269 3131 1327 3137
rect 1269 3097 1281 3131
rect 1315 3097 1327 3131
rect 1269 3091 1327 3097
rect 1387 3131 1445 3137
rect 1387 3097 1399 3131
rect 1433 3097 1445 3131
rect 1387 3091 1445 3097
rect -1498 3001 -1452 3013
rect -1498 2425 -1492 3001
rect -1458 2425 -1452 3001
rect -1498 2413 -1452 2425
rect -1380 3001 -1334 3013
rect -1380 2425 -1374 3001
rect -1340 2425 -1334 3001
rect -1380 2413 -1334 2425
rect -1262 3001 -1216 3013
rect -1262 2425 -1256 3001
rect -1222 2425 -1216 3001
rect -1262 2413 -1216 2425
rect -1144 3001 -1098 3013
rect -1144 2425 -1138 3001
rect -1104 2425 -1098 3001
rect -1144 2413 -1098 2425
rect -1026 3001 -980 3013
rect -1026 2425 -1020 3001
rect -986 2425 -980 3001
rect -1026 2413 -980 2425
rect -908 3001 -862 3013
rect -908 2425 -902 3001
rect -868 2425 -862 3001
rect -908 2413 -862 2425
rect -790 3001 -744 3013
rect -790 2425 -784 3001
rect -750 2425 -744 3001
rect -790 2413 -744 2425
rect -672 3001 -626 3013
rect -672 2425 -666 3001
rect -632 2425 -626 3001
rect -672 2413 -626 2425
rect -554 3001 -508 3013
rect -554 2425 -548 3001
rect -514 2425 -508 3001
rect -554 2413 -508 2425
rect -436 3001 -390 3013
rect -436 2425 -430 3001
rect -396 2425 -390 3001
rect -436 2413 -390 2425
rect -318 3001 -272 3013
rect -318 2425 -312 3001
rect -278 2425 -272 3001
rect -318 2413 -272 2425
rect -200 3001 -154 3013
rect -200 2425 -194 3001
rect -160 2425 -154 3001
rect -200 2413 -154 2425
rect -82 3001 -36 3013
rect -82 2425 -76 3001
rect -42 2425 -36 3001
rect -82 2413 -36 2425
rect 36 3001 82 3013
rect 36 2425 42 3001
rect 76 2425 82 3001
rect 36 2413 82 2425
rect 154 3001 200 3013
rect 154 2425 160 3001
rect 194 2425 200 3001
rect 154 2413 200 2425
rect 272 3001 318 3013
rect 272 2425 278 3001
rect 312 2425 318 3001
rect 272 2413 318 2425
rect 390 3001 436 3013
rect 390 2425 396 3001
rect 430 2425 436 3001
rect 390 2413 436 2425
rect 508 3001 554 3013
rect 508 2425 514 3001
rect 548 2425 554 3001
rect 508 2413 554 2425
rect 626 3001 672 3013
rect 626 2425 632 3001
rect 666 2425 672 3001
rect 626 2413 672 2425
rect 744 3001 790 3013
rect 744 2425 750 3001
rect 784 2425 790 3001
rect 744 2413 790 2425
rect 862 3001 908 3013
rect 862 2425 868 3001
rect 902 2425 908 3001
rect 862 2413 908 2425
rect 980 3001 1026 3013
rect 980 2425 986 3001
rect 1020 2425 1026 3001
rect 980 2413 1026 2425
rect 1098 3001 1144 3013
rect 1098 2425 1104 3001
rect 1138 2425 1144 3001
rect 1098 2413 1144 2425
rect 1216 3001 1262 3013
rect 1216 2425 1222 3001
rect 1256 2425 1262 3001
rect 1216 2413 1262 2425
rect 1334 3001 1380 3013
rect 1334 2425 1340 3001
rect 1374 2425 1380 3001
rect 1334 2413 1380 2425
rect 1452 3001 1498 3013
rect 1452 2425 1458 3001
rect 1492 2425 1498 3001
rect 1452 2413 1498 2425
rect -1445 2366 -1387 2372
rect -1445 2332 -1433 2366
rect -1399 2332 -1387 2366
rect -1445 2326 -1387 2332
rect -1327 2366 -1269 2372
rect -1327 2332 -1315 2366
rect -1281 2332 -1269 2366
rect -1327 2326 -1269 2332
rect -1209 2366 -1151 2372
rect -1209 2332 -1197 2366
rect -1163 2332 -1151 2366
rect -1209 2326 -1151 2332
rect -1091 2366 -1033 2372
rect -1091 2332 -1079 2366
rect -1045 2332 -1033 2366
rect -1091 2326 -1033 2332
rect -973 2366 -915 2372
rect -973 2332 -961 2366
rect -927 2332 -915 2366
rect -973 2326 -915 2332
rect -855 2366 -797 2372
rect -855 2332 -843 2366
rect -809 2332 -797 2366
rect -855 2326 -797 2332
rect -737 2366 -679 2372
rect -737 2332 -725 2366
rect -691 2332 -679 2366
rect -737 2326 -679 2332
rect -619 2366 -561 2372
rect -619 2332 -607 2366
rect -573 2332 -561 2366
rect -619 2326 -561 2332
rect -501 2366 -443 2372
rect -501 2332 -489 2366
rect -455 2332 -443 2366
rect -501 2326 -443 2332
rect -383 2366 -325 2372
rect -383 2332 -371 2366
rect -337 2332 -325 2366
rect -383 2326 -325 2332
rect -265 2366 -207 2372
rect -265 2332 -253 2366
rect -219 2332 -207 2366
rect -265 2326 -207 2332
rect -147 2366 -89 2372
rect -147 2332 -135 2366
rect -101 2332 -89 2366
rect -147 2326 -89 2332
rect -29 2366 29 2372
rect -29 2332 -17 2366
rect 17 2332 29 2366
rect -29 2326 29 2332
rect 89 2366 147 2372
rect 89 2332 101 2366
rect 135 2332 147 2366
rect 89 2326 147 2332
rect 207 2366 265 2372
rect 207 2332 219 2366
rect 253 2332 265 2366
rect 207 2326 265 2332
rect 325 2366 383 2372
rect 325 2332 337 2366
rect 371 2332 383 2366
rect 325 2326 383 2332
rect 443 2366 501 2372
rect 443 2332 455 2366
rect 489 2332 501 2366
rect 443 2326 501 2332
rect 561 2366 619 2372
rect 561 2332 573 2366
rect 607 2332 619 2366
rect 561 2326 619 2332
rect 679 2366 737 2372
rect 679 2332 691 2366
rect 725 2332 737 2366
rect 679 2326 737 2332
rect 797 2366 855 2372
rect 797 2332 809 2366
rect 843 2332 855 2366
rect 797 2326 855 2332
rect 915 2366 973 2372
rect 915 2332 927 2366
rect 961 2332 973 2366
rect 915 2326 973 2332
rect 1033 2366 1091 2372
rect 1033 2332 1045 2366
rect 1079 2332 1091 2366
rect 1033 2326 1091 2332
rect 1151 2366 1209 2372
rect 1151 2332 1163 2366
rect 1197 2332 1209 2366
rect 1151 2326 1209 2332
rect 1269 2366 1327 2372
rect 1269 2332 1281 2366
rect 1315 2332 1327 2366
rect 1269 2326 1327 2332
rect 1387 2366 1445 2372
rect 1387 2332 1399 2366
rect 1433 2332 1445 2366
rect 1387 2326 1445 2332
rect -1498 2236 -1452 2248
rect -1498 1660 -1492 2236
rect -1458 1660 -1452 2236
rect -1498 1648 -1452 1660
rect -1380 2236 -1334 2248
rect -1380 1660 -1374 2236
rect -1340 1660 -1334 2236
rect -1380 1648 -1334 1660
rect -1262 2236 -1216 2248
rect -1262 1660 -1256 2236
rect -1222 1660 -1216 2236
rect -1262 1648 -1216 1660
rect -1144 2236 -1098 2248
rect -1144 1660 -1138 2236
rect -1104 1660 -1098 2236
rect -1144 1648 -1098 1660
rect -1026 2236 -980 2248
rect -1026 1660 -1020 2236
rect -986 1660 -980 2236
rect -1026 1648 -980 1660
rect -908 2236 -862 2248
rect -908 1660 -902 2236
rect -868 1660 -862 2236
rect -908 1648 -862 1660
rect -790 2236 -744 2248
rect -790 1660 -784 2236
rect -750 1660 -744 2236
rect -790 1648 -744 1660
rect -672 2236 -626 2248
rect -672 1660 -666 2236
rect -632 1660 -626 2236
rect -672 1648 -626 1660
rect -554 2236 -508 2248
rect -554 1660 -548 2236
rect -514 1660 -508 2236
rect -554 1648 -508 1660
rect -436 2236 -390 2248
rect -436 1660 -430 2236
rect -396 1660 -390 2236
rect -436 1648 -390 1660
rect -318 2236 -272 2248
rect -318 1660 -312 2236
rect -278 1660 -272 2236
rect -318 1648 -272 1660
rect -200 2236 -154 2248
rect -200 1660 -194 2236
rect -160 1660 -154 2236
rect -200 1648 -154 1660
rect -82 2236 -36 2248
rect -82 1660 -76 2236
rect -42 1660 -36 2236
rect -82 1648 -36 1660
rect 36 2236 82 2248
rect 36 1660 42 2236
rect 76 1660 82 2236
rect 36 1648 82 1660
rect 154 2236 200 2248
rect 154 1660 160 2236
rect 194 1660 200 2236
rect 154 1648 200 1660
rect 272 2236 318 2248
rect 272 1660 278 2236
rect 312 1660 318 2236
rect 272 1648 318 1660
rect 390 2236 436 2248
rect 390 1660 396 2236
rect 430 1660 436 2236
rect 390 1648 436 1660
rect 508 2236 554 2248
rect 508 1660 514 2236
rect 548 1660 554 2236
rect 508 1648 554 1660
rect 626 2236 672 2248
rect 626 1660 632 2236
rect 666 1660 672 2236
rect 626 1648 672 1660
rect 744 2236 790 2248
rect 744 1660 750 2236
rect 784 1660 790 2236
rect 744 1648 790 1660
rect 862 2236 908 2248
rect 862 1660 868 2236
rect 902 1660 908 2236
rect 862 1648 908 1660
rect 980 2236 1026 2248
rect 980 1660 986 2236
rect 1020 1660 1026 2236
rect 980 1648 1026 1660
rect 1098 2236 1144 2248
rect 1098 1660 1104 2236
rect 1138 1660 1144 2236
rect 1098 1648 1144 1660
rect 1216 2236 1262 2248
rect 1216 1660 1222 2236
rect 1256 1660 1262 2236
rect 1216 1648 1262 1660
rect 1334 2236 1380 2248
rect 1334 1660 1340 2236
rect 1374 1660 1380 2236
rect 1334 1648 1380 1660
rect 1452 2236 1498 2248
rect 1452 1660 1458 2236
rect 1492 1660 1498 2236
rect 1452 1648 1498 1660
rect -1445 1601 -1387 1607
rect -1445 1567 -1433 1601
rect -1399 1567 -1387 1601
rect -1445 1561 -1387 1567
rect -1327 1601 -1269 1607
rect -1327 1567 -1315 1601
rect -1281 1567 -1269 1601
rect -1327 1561 -1269 1567
rect -1209 1601 -1151 1607
rect -1209 1567 -1197 1601
rect -1163 1567 -1151 1601
rect -1209 1561 -1151 1567
rect -1091 1601 -1033 1607
rect -1091 1567 -1079 1601
rect -1045 1567 -1033 1601
rect -1091 1561 -1033 1567
rect -973 1601 -915 1607
rect -973 1567 -961 1601
rect -927 1567 -915 1601
rect -973 1561 -915 1567
rect -855 1601 -797 1607
rect -855 1567 -843 1601
rect -809 1567 -797 1601
rect -855 1561 -797 1567
rect -737 1601 -679 1607
rect -737 1567 -725 1601
rect -691 1567 -679 1601
rect -737 1561 -679 1567
rect -619 1601 -561 1607
rect -619 1567 -607 1601
rect -573 1567 -561 1601
rect -619 1561 -561 1567
rect -501 1601 -443 1607
rect -501 1567 -489 1601
rect -455 1567 -443 1601
rect -501 1561 -443 1567
rect -383 1601 -325 1607
rect -383 1567 -371 1601
rect -337 1567 -325 1601
rect -383 1561 -325 1567
rect -265 1601 -207 1607
rect -265 1567 -253 1601
rect -219 1567 -207 1601
rect -265 1561 -207 1567
rect -147 1601 -89 1607
rect -147 1567 -135 1601
rect -101 1567 -89 1601
rect -147 1561 -89 1567
rect -29 1601 29 1607
rect -29 1567 -17 1601
rect 17 1567 29 1601
rect -29 1561 29 1567
rect 89 1601 147 1607
rect 89 1567 101 1601
rect 135 1567 147 1601
rect 89 1561 147 1567
rect 207 1601 265 1607
rect 207 1567 219 1601
rect 253 1567 265 1601
rect 207 1561 265 1567
rect 325 1601 383 1607
rect 325 1567 337 1601
rect 371 1567 383 1601
rect 325 1561 383 1567
rect 443 1601 501 1607
rect 443 1567 455 1601
rect 489 1567 501 1601
rect 443 1561 501 1567
rect 561 1601 619 1607
rect 561 1567 573 1601
rect 607 1567 619 1601
rect 561 1561 619 1567
rect 679 1601 737 1607
rect 679 1567 691 1601
rect 725 1567 737 1601
rect 679 1561 737 1567
rect 797 1601 855 1607
rect 797 1567 809 1601
rect 843 1567 855 1601
rect 797 1561 855 1567
rect 915 1601 973 1607
rect 915 1567 927 1601
rect 961 1567 973 1601
rect 915 1561 973 1567
rect 1033 1601 1091 1607
rect 1033 1567 1045 1601
rect 1079 1567 1091 1601
rect 1033 1561 1091 1567
rect 1151 1601 1209 1607
rect 1151 1567 1163 1601
rect 1197 1567 1209 1601
rect 1151 1561 1209 1567
rect 1269 1601 1327 1607
rect 1269 1567 1281 1601
rect 1315 1567 1327 1601
rect 1269 1561 1327 1567
rect 1387 1601 1445 1607
rect 1387 1567 1399 1601
rect 1433 1567 1445 1601
rect 1387 1561 1445 1567
rect -1498 1471 -1452 1483
rect -1498 895 -1492 1471
rect -1458 895 -1452 1471
rect -1498 883 -1452 895
rect -1380 1471 -1334 1483
rect -1380 895 -1374 1471
rect -1340 895 -1334 1471
rect -1380 883 -1334 895
rect -1262 1471 -1216 1483
rect -1262 895 -1256 1471
rect -1222 895 -1216 1471
rect -1262 883 -1216 895
rect -1144 1471 -1098 1483
rect -1144 895 -1138 1471
rect -1104 895 -1098 1471
rect -1144 883 -1098 895
rect -1026 1471 -980 1483
rect -1026 895 -1020 1471
rect -986 895 -980 1471
rect -1026 883 -980 895
rect -908 1471 -862 1483
rect -908 895 -902 1471
rect -868 895 -862 1471
rect -908 883 -862 895
rect -790 1471 -744 1483
rect -790 895 -784 1471
rect -750 895 -744 1471
rect -790 883 -744 895
rect -672 1471 -626 1483
rect -672 895 -666 1471
rect -632 895 -626 1471
rect -672 883 -626 895
rect -554 1471 -508 1483
rect -554 895 -548 1471
rect -514 895 -508 1471
rect -554 883 -508 895
rect -436 1471 -390 1483
rect -436 895 -430 1471
rect -396 895 -390 1471
rect -436 883 -390 895
rect -318 1471 -272 1483
rect -318 895 -312 1471
rect -278 895 -272 1471
rect -318 883 -272 895
rect -200 1471 -154 1483
rect -200 895 -194 1471
rect -160 895 -154 1471
rect -200 883 -154 895
rect -82 1471 -36 1483
rect -82 895 -76 1471
rect -42 895 -36 1471
rect -82 883 -36 895
rect 36 1471 82 1483
rect 36 895 42 1471
rect 76 895 82 1471
rect 36 883 82 895
rect 154 1471 200 1483
rect 154 895 160 1471
rect 194 895 200 1471
rect 154 883 200 895
rect 272 1471 318 1483
rect 272 895 278 1471
rect 312 895 318 1471
rect 272 883 318 895
rect 390 1471 436 1483
rect 390 895 396 1471
rect 430 895 436 1471
rect 390 883 436 895
rect 508 1471 554 1483
rect 508 895 514 1471
rect 548 895 554 1471
rect 508 883 554 895
rect 626 1471 672 1483
rect 626 895 632 1471
rect 666 895 672 1471
rect 626 883 672 895
rect 744 1471 790 1483
rect 744 895 750 1471
rect 784 895 790 1471
rect 744 883 790 895
rect 862 1471 908 1483
rect 862 895 868 1471
rect 902 895 908 1471
rect 862 883 908 895
rect 980 1471 1026 1483
rect 980 895 986 1471
rect 1020 895 1026 1471
rect 980 883 1026 895
rect 1098 1471 1144 1483
rect 1098 895 1104 1471
rect 1138 895 1144 1471
rect 1098 883 1144 895
rect 1216 1471 1262 1483
rect 1216 895 1222 1471
rect 1256 895 1262 1471
rect 1216 883 1262 895
rect 1334 1471 1380 1483
rect 1334 895 1340 1471
rect 1374 895 1380 1471
rect 1334 883 1380 895
rect 1452 1471 1498 1483
rect 1452 895 1458 1471
rect 1492 895 1498 1471
rect 1452 883 1498 895
rect -1445 836 -1387 842
rect -1445 802 -1433 836
rect -1399 802 -1387 836
rect -1445 796 -1387 802
rect -1327 836 -1269 842
rect -1327 802 -1315 836
rect -1281 802 -1269 836
rect -1327 796 -1269 802
rect -1209 836 -1151 842
rect -1209 802 -1197 836
rect -1163 802 -1151 836
rect -1209 796 -1151 802
rect -1091 836 -1033 842
rect -1091 802 -1079 836
rect -1045 802 -1033 836
rect -1091 796 -1033 802
rect -973 836 -915 842
rect -973 802 -961 836
rect -927 802 -915 836
rect -973 796 -915 802
rect -855 836 -797 842
rect -855 802 -843 836
rect -809 802 -797 836
rect -855 796 -797 802
rect -737 836 -679 842
rect -737 802 -725 836
rect -691 802 -679 836
rect -737 796 -679 802
rect -619 836 -561 842
rect -619 802 -607 836
rect -573 802 -561 836
rect -619 796 -561 802
rect -501 836 -443 842
rect -501 802 -489 836
rect -455 802 -443 836
rect -501 796 -443 802
rect -383 836 -325 842
rect -383 802 -371 836
rect -337 802 -325 836
rect -383 796 -325 802
rect -265 836 -207 842
rect -265 802 -253 836
rect -219 802 -207 836
rect -265 796 -207 802
rect -147 836 -89 842
rect -147 802 -135 836
rect -101 802 -89 836
rect -147 796 -89 802
rect -29 836 29 842
rect -29 802 -17 836
rect 17 802 29 836
rect -29 796 29 802
rect 89 836 147 842
rect 89 802 101 836
rect 135 802 147 836
rect 89 796 147 802
rect 207 836 265 842
rect 207 802 219 836
rect 253 802 265 836
rect 207 796 265 802
rect 325 836 383 842
rect 325 802 337 836
rect 371 802 383 836
rect 325 796 383 802
rect 443 836 501 842
rect 443 802 455 836
rect 489 802 501 836
rect 443 796 501 802
rect 561 836 619 842
rect 561 802 573 836
rect 607 802 619 836
rect 561 796 619 802
rect 679 836 737 842
rect 679 802 691 836
rect 725 802 737 836
rect 679 796 737 802
rect 797 836 855 842
rect 797 802 809 836
rect 843 802 855 836
rect 797 796 855 802
rect 915 836 973 842
rect 915 802 927 836
rect 961 802 973 836
rect 915 796 973 802
rect 1033 836 1091 842
rect 1033 802 1045 836
rect 1079 802 1091 836
rect 1033 796 1091 802
rect 1151 836 1209 842
rect 1151 802 1163 836
rect 1197 802 1209 836
rect 1151 796 1209 802
rect 1269 836 1327 842
rect 1269 802 1281 836
rect 1315 802 1327 836
rect 1269 796 1327 802
rect 1387 836 1445 842
rect 1387 802 1399 836
rect 1433 802 1445 836
rect 1387 796 1445 802
rect -1498 706 -1452 718
rect -1498 130 -1492 706
rect -1458 130 -1452 706
rect -1498 118 -1452 130
rect -1380 706 -1334 718
rect -1380 130 -1374 706
rect -1340 130 -1334 706
rect -1380 118 -1334 130
rect -1262 706 -1216 718
rect -1262 130 -1256 706
rect -1222 130 -1216 706
rect -1262 118 -1216 130
rect -1144 706 -1098 718
rect -1144 130 -1138 706
rect -1104 130 -1098 706
rect -1144 118 -1098 130
rect -1026 706 -980 718
rect -1026 130 -1020 706
rect -986 130 -980 706
rect -1026 118 -980 130
rect -908 706 -862 718
rect -908 130 -902 706
rect -868 130 -862 706
rect -908 118 -862 130
rect -790 706 -744 718
rect -790 130 -784 706
rect -750 130 -744 706
rect -790 118 -744 130
rect -672 706 -626 718
rect -672 130 -666 706
rect -632 130 -626 706
rect -672 118 -626 130
rect -554 706 -508 718
rect -554 130 -548 706
rect -514 130 -508 706
rect -554 118 -508 130
rect -436 706 -390 718
rect -436 130 -430 706
rect -396 130 -390 706
rect -436 118 -390 130
rect -318 706 -272 718
rect -318 130 -312 706
rect -278 130 -272 706
rect -318 118 -272 130
rect -200 706 -154 718
rect -200 130 -194 706
rect -160 130 -154 706
rect -200 118 -154 130
rect -82 706 -36 718
rect -82 130 -76 706
rect -42 130 -36 706
rect -82 118 -36 130
rect 36 706 82 718
rect 36 130 42 706
rect 76 130 82 706
rect 36 118 82 130
rect 154 706 200 718
rect 154 130 160 706
rect 194 130 200 706
rect 154 118 200 130
rect 272 706 318 718
rect 272 130 278 706
rect 312 130 318 706
rect 272 118 318 130
rect 390 706 436 718
rect 390 130 396 706
rect 430 130 436 706
rect 390 118 436 130
rect 508 706 554 718
rect 508 130 514 706
rect 548 130 554 706
rect 508 118 554 130
rect 626 706 672 718
rect 626 130 632 706
rect 666 130 672 706
rect 626 118 672 130
rect 744 706 790 718
rect 744 130 750 706
rect 784 130 790 706
rect 744 118 790 130
rect 862 706 908 718
rect 862 130 868 706
rect 902 130 908 706
rect 862 118 908 130
rect 980 706 1026 718
rect 980 130 986 706
rect 1020 130 1026 706
rect 980 118 1026 130
rect 1098 706 1144 718
rect 1098 130 1104 706
rect 1138 130 1144 706
rect 1098 118 1144 130
rect 1216 706 1262 718
rect 1216 130 1222 706
rect 1256 130 1262 706
rect 1216 118 1262 130
rect 1334 706 1380 718
rect 1334 130 1340 706
rect 1374 130 1380 706
rect 1334 118 1380 130
rect 1452 706 1498 718
rect 1452 130 1458 706
rect 1492 130 1498 706
rect 1452 118 1498 130
rect -1445 71 -1387 77
rect -1445 37 -1433 71
rect -1399 37 -1387 71
rect -1445 31 -1387 37
rect -1327 71 -1269 77
rect -1327 37 -1315 71
rect -1281 37 -1269 71
rect -1327 31 -1269 37
rect -1209 71 -1151 77
rect -1209 37 -1197 71
rect -1163 37 -1151 71
rect -1209 31 -1151 37
rect -1091 71 -1033 77
rect -1091 37 -1079 71
rect -1045 37 -1033 71
rect -1091 31 -1033 37
rect -973 71 -915 77
rect -973 37 -961 71
rect -927 37 -915 71
rect -973 31 -915 37
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect 915 71 973 77
rect 915 37 927 71
rect 961 37 973 71
rect 915 31 973 37
rect 1033 71 1091 77
rect 1033 37 1045 71
rect 1079 37 1091 71
rect 1033 31 1091 37
rect 1151 71 1209 77
rect 1151 37 1163 71
rect 1197 37 1209 71
rect 1151 31 1209 37
rect 1269 71 1327 77
rect 1269 37 1281 71
rect 1315 37 1327 71
rect 1269 31 1327 37
rect 1387 71 1445 77
rect 1387 37 1399 71
rect 1433 37 1445 71
rect 1387 31 1445 37
rect -1498 -59 -1452 -47
rect -1498 -635 -1492 -59
rect -1458 -635 -1452 -59
rect -1498 -647 -1452 -635
rect -1380 -59 -1334 -47
rect -1380 -635 -1374 -59
rect -1340 -635 -1334 -59
rect -1380 -647 -1334 -635
rect -1262 -59 -1216 -47
rect -1262 -635 -1256 -59
rect -1222 -635 -1216 -59
rect -1262 -647 -1216 -635
rect -1144 -59 -1098 -47
rect -1144 -635 -1138 -59
rect -1104 -635 -1098 -59
rect -1144 -647 -1098 -635
rect -1026 -59 -980 -47
rect -1026 -635 -1020 -59
rect -986 -635 -980 -59
rect -1026 -647 -980 -635
rect -908 -59 -862 -47
rect -908 -635 -902 -59
rect -868 -635 -862 -59
rect -908 -647 -862 -635
rect -790 -59 -744 -47
rect -790 -635 -784 -59
rect -750 -635 -744 -59
rect -790 -647 -744 -635
rect -672 -59 -626 -47
rect -672 -635 -666 -59
rect -632 -635 -626 -59
rect -672 -647 -626 -635
rect -554 -59 -508 -47
rect -554 -635 -548 -59
rect -514 -635 -508 -59
rect -554 -647 -508 -635
rect -436 -59 -390 -47
rect -436 -635 -430 -59
rect -396 -635 -390 -59
rect -436 -647 -390 -635
rect -318 -59 -272 -47
rect -318 -635 -312 -59
rect -278 -635 -272 -59
rect -318 -647 -272 -635
rect -200 -59 -154 -47
rect -200 -635 -194 -59
rect -160 -635 -154 -59
rect -200 -647 -154 -635
rect -82 -59 -36 -47
rect -82 -635 -76 -59
rect -42 -635 -36 -59
rect -82 -647 -36 -635
rect 36 -59 82 -47
rect 36 -635 42 -59
rect 76 -635 82 -59
rect 36 -647 82 -635
rect 154 -59 200 -47
rect 154 -635 160 -59
rect 194 -635 200 -59
rect 154 -647 200 -635
rect 272 -59 318 -47
rect 272 -635 278 -59
rect 312 -635 318 -59
rect 272 -647 318 -635
rect 390 -59 436 -47
rect 390 -635 396 -59
rect 430 -635 436 -59
rect 390 -647 436 -635
rect 508 -59 554 -47
rect 508 -635 514 -59
rect 548 -635 554 -59
rect 508 -647 554 -635
rect 626 -59 672 -47
rect 626 -635 632 -59
rect 666 -635 672 -59
rect 626 -647 672 -635
rect 744 -59 790 -47
rect 744 -635 750 -59
rect 784 -635 790 -59
rect 744 -647 790 -635
rect 862 -59 908 -47
rect 862 -635 868 -59
rect 902 -635 908 -59
rect 862 -647 908 -635
rect 980 -59 1026 -47
rect 980 -635 986 -59
rect 1020 -635 1026 -59
rect 980 -647 1026 -635
rect 1098 -59 1144 -47
rect 1098 -635 1104 -59
rect 1138 -635 1144 -59
rect 1098 -647 1144 -635
rect 1216 -59 1262 -47
rect 1216 -635 1222 -59
rect 1256 -635 1262 -59
rect 1216 -647 1262 -635
rect 1334 -59 1380 -47
rect 1334 -635 1340 -59
rect 1374 -635 1380 -59
rect 1334 -647 1380 -635
rect 1452 -59 1498 -47
rect 1452 -635 1458 -59
rect 1492 -635 1498 -59
rect 1452 -647 1498 -635
rect -1445 -694 -1387 -688
rect -1445 -728 -1433 -694
rect -1399 -728 -1387 -694
rect -1445 -734 -1387 -728
rect -1327 -694 -1269 -688
rect -1327 -728 -1315 -694
rect -1281 -728 -1269 -694
rect -1327 -734 -1269 -728
rect -1209 -694 -1151 -688
rect -1209 -728 -1197 -694
rect -1163 -728 -1151 -694
rect -1209 -734 -1151 -728
rect -1091 -694 -1033 -688
rect -1091 -728 -1079 -694
rect -1045 -728 -1033 -694
rect -1091 -734 -1033 -728
rect -973 -694 -915 -688
rect -973 -728 -961 -694
rect -927 -728 -915 -694
rect -973 -734 -915 -728
rect -855 -694 -797 -688
rect -855 -728 -843 -694
rect -809 -728 -797 -694
rect -855 -734 -797 -728
rect -737 -694 -679 -688
rect -737 -728 -725 -694
rect -691 -728 -679 -694
rect -737 -734 -679 -728
rect -619 -694 -561 -688
rect -619 -728 -607 -694
rect -573 -728 -561 -694
rect -619 -734 -561 -728
rect -501 -694 -443 -688
rect -501 -728 -489 -694
rect -455 -728 -443 -694
rect -501 -734 -443 -728
rect -383 -694 -325 -688
rect -383 -728 -371 -694
rect -337 -728 -325 -694
rect -383 -734 -325 -728
rect -265 -694 -207 -688
rect -265 -728 -253 -694
rect -219 -728 -207 -694
rect -265 -734 -207 -728
rect -147 -694 -89 -688
rect -147 -728 -135 -694
rect -101 -728 -89 -694
rect -147 -734 -89 -728
rect -29 -694 29 -688
rect -29 -728 -17 -694
rect 17 -728 29 -694
rect -29 -734 29 -728
rect 89 -694 147 -688
rect 89 -728 101 -694
rect 135 -728 147 -694
rect 89 -734 147 -728
rect 207 -694 265 -688
rect 207 -728 219 -694
rect 253 -728 265 -694
rect 207 -734 265 -728
rect 325 -694 383 -688
rect 325 -728 337 -694
rect 371 -728 383 -694
rect 325 -734 383 -728
rect 443 -694 501 -688
rect 443 -728 455 -694
rect 489 -728 501 -694
rect 443 -734 501 -728
rect 561 -694 619 -688
rect 561 -728 573 -694
rect 607 -728 619 -694
rect 561 -734 619 -728
rect 679 -694 737 -688
rect 679 -728 691 -694
rect 725 -728 737 -694
rect 679 -734 737 -728
rect 797 -694 855 -688
rect 797 -728 809 -694
rect 843 -728 855 -694
rect 797 -734 855 -728
rect 915 -694 973 -688
rect 915 -728 927 -694
rect 961 -728 973 -694
rect 915 -734 973 -728
rect 1033 -694 1091 -688
rect 1033 -728 1045 -694
rect 1079 -728 1091 -694
rect 1033 -734 1091 -728
rect 1151 -694 1209 -688
rect 1151 -728 1163 -694
rect 1197 -728 1209 -694
rect 1151 -734 1209 -728
rect 1269 -694 1327 -688
rect 1269 -728 1281 -694
rect 1315 -728 1327 -694
rect 1269 -734 1327 -728
rect 1387 -694 1445 -688
rect 1387 -728 1399 -694
rect 1433 -728 1445 -694
rect 1387 -734 1445 -728
rect -1498 -824 -1452 -812
rect -1498 -1400 -1492 -824
rect -1458 -1400 -1452 -824
rect -1498 -1412 -1452 -1400
rect -1380 -824 -1334 -812
rect -1380 -1400 -1374 -824
rect -1340 -1400 -1334 -824
rect -1380 -1412 -1334 -1400
rect -1262 -824 -1216 -812
rect -1262 -1400 -1256 -824
rect -1222 -1400 -1216 -824
rect -1262 -1412 -1216 -1400
rect -1144 -824 -1098 -812
rect -1144 -1400 -1138 -824
rect -1104 -1400 -1098 -824
rect -1144 -1412 -1098 -1400
rect -1026 -824 -980 -812
rect -1026 -1400 -1020 -824
rect -986 -1400 -980 -824
rect -1026 -1412 -980 -1400
rect -908 -824 -862 -812
rect -908 -1400 -902 -824
rect -868 -1400 -862 -824
rect -908 -1412 -862 -1400
rect -790 -824 -744 -812
rect -790 -1400 -784 -824
rect -750 -1400 -744 -824
rect -790 -1412 -744 -1400
rect -672 -824 -626 -812
rect -672 -1400 -666 -824
rect -632 -1400 -626 -824
rect -672 -1412 -626 -1400
rect -554 -824 -508 -812
rect -554 -1400 -548 -824
rect -514 -1400 -508 -824
rect -554 -1412 -508 -1400
rect -436 -824 -390 -812
rect -436 -1400 -430 -824
rect -396 -1400 -390 -824
rect -436 -1412 -390 -1400
rect -318 -824 -272 -812
rect -318 -1400 -312 -824
rect -278 -1400 -272 -824
rect -318 -1412 -272 -1400
rect -200 -824 -154 -812
rect -200 -1400 -194 -824
rect -160 -1400 -154 -824
rect -200 -1412 -154 -1400
rect -82 -824 -36 -812
rect -82 -1400 -76 -824
rect -42 -1400 -36 -824
rect -82 -1412 -36 -1400
rect 36 -824 82 -812
rect 36 -1400 42 -824
rect 76 -1400 82 -824
rect 36 -1412 82 -1400
rect 154 -824 200 -812
rect 154 -1400 160 -824
rect 194 -1400 200 -824
rect 154 -1412 200 -1400
rect 272 -824 318 -812
rect 272 -1400 278 -824
rect 312 -1400 318 -824
rect 272 -1412 318 -1400
rect 390 -824 436 -812
rect 390 -1400 396 -824
rect 430 -1400 436 -824
rect 390 -1412 436 -1400
rect 508 -824 554 -812
rect 508 -1400 514 -824
rect 548 -1400 554 -824
rect 508 -1412 554 -1400
rect 626 -824 672 -812
rect 626 -1400 632 -824
rect 666 -1400 672 -824
rect 626 -1412 672 -1400
rect 744 -824 790 -812
rect 744 -1400 750 -824
rect 784 -1400 790 -824
rect 744 -1412 790 -1400
rect 862 -824 908 -812
rect 862 -1400 868 -824
rect 902 -1400 908 -824
rect 862 -1412 908 -1400
rect 980 -824 1026 -812
rect 980 -1400 986 -824
rect 1020 -1400 1026 -824
rect 980 -1412 1026 -1400
rect 1098 -824 1144 -812
rect 1098 -1400 1104 -824
rect 1138 -1400 1144 -824
rect 1098 -1412 1144 -1400
rect 1216 -824 1262 -812
rect 1216 -1400 1222 -824
rect 1256 -1400 1262 -824
rect 1216 -1412 1262 -1400
rect 1334 -824 1380 -812
rect 1334 -1400 1340 -824
rect 1374 -1400 1380 -824
rect 1334 -1412 1380 -1400
rect 1452 -824 1498 -812
rect 1452 -1400 1458 -824
rect 1492 -1400 1498 -824
rect 1452 -1412 1498 -1400
rect -1445 -1459 -1387 -1453
rect -1445 -1493 -1433 -1459
rect -1399 -1493 -1387 -1459
rect -1445 -1499 -1387 -1493
rect -1327 -1459 -1269 -1453
rect -1327 -1493 -1315 -1459
rect -1281 -1493 -1269 -1459
rect -1327 -1499 -1269 -1493
rect -1209 -1459 -1151 -1453
rect -1209 -1493 -1197 -1459
rect -1163 -1493 -1151 -1459
rect -1209 -1499 -1151 -1493
rect -1091 -1459 -1033 -1453
rect -1091 -1493 -1079 -1459
rect -1045 -1493 -1033 -1459
rect -1091 -1499 -1033 -1493
rect -973 -1459 -915 -1453
rect -973 -1493 -961 -1459
rect -927 -1493 -915 -1459
rect -973 -1499 -915 -1493
rect -855 -1459 -797 -1453
rect -855 -1493 -843 -1459
rect -809 -1493 -797 -1459
rect -855 -1499 -797 -1493
rect -737 -1459 -679 -1453
rect -737 -1493 -725 -1459
rect -691 -1493 -679 -1459
rect -737 -1499 -679 -1493
rect -619 -1459 -561 -1453
rect -619 -1493 -607 -1459
rect -573 -1493 -561 -1459
rect -619 -1499 -561 -1493
rect -501 -1459 -443 -1453
rect -501 -1493 -489 -1459
rect -455 -1493 -443 -1459
rect -501 -1499 -443 -1493
rect -383 -1459 -325 -1453
rect -383 -1493 -371 -1459
rect -337 -1493 -325 -1459
rect -383 -1499 -325 -1493
rect -265 -1459 -207 -1453
rect -265 -1493 -253 -1459
rect -219 -1493 -207 -1459
rect -265 -1499 -207 -1493
rect -147 -1459 -89 -1453
rect -147 -1493 -135 -1459
rect -101 -1493 -89 -1459
rect -147 -1499 -89 -1493
rect -29 -1459 29 -1453
rect -29 -1493 -17 -1459
rect 17 -1493 29 -1459
rect -29 -1499 29 -1493
rect 89 -1459 147 -1453
rect 89 -1493 101 -1459
rect 135 -1493 147 -1459
rect 89 -1499 147 -1493
rect 207 -1459 265 -1453
rect 207 -1493 219 -1459
rect 253 -1493 265 -1459
rect 207 -1499 265 -1493
rect 325 -1459 383 -1453
rect 325 -1493 337 -1459
rect 371 -1493 383 -1459
rect 325 -1499 383 -1493
rect 443 -1459 501 -1453
rect 443 -1493 455 -1459
rect 489 -1493 501 -1459
rect 443 -1499 501 -1493
rect 561 -1459 619 -1453
rect 561 -1493 573 -1459
rect 607 -1493 619 -1459
rect 561 -1499 619 -1493
rect 679 -1459 737 -1453
rect 679 -1493 691 -1459
rect 725 -1493 737 -1459
rect 679 -1499 737 -1493
rect 797 -1459 855 -1453
rect 797 -1493 809 -1459
rect 843 -1493 855 -1459
rect 797 -1499 855 -1493
rect 915 -1459 973 -1453
rect 915 -1493 927 -1459
rect 961 -1493 973 -1459
rect 915 -1499 973 -1493
rect 1033 -1459 1091 -1453
rect 1033 -1493 1045 -1459
rect 1079 -1493 1091 -1459
rect 1033 -1499 1091 -1493
rect 1151 -1459 1209 -1453
rect 1151 -1493 1163 -1459
rect 1197 -1493 1209 -1459
rect 1151 -1499 1209 -1493
rect 1269 -1459 1327 -1453
rect 1269 -1493 1281 -1459
rect 1315 -1493 1327 -1459
rect 1269 -1499 1327 -1493
rect 1387 -1459 1445 -1453
rect 1387 -1493 1399 -1459
rect 1433 -1493 1445 -1459
rect 1387 -1499 1445 -1493
rect -1498 -1589 -1452 -1577
rect -1498 -2165 -1492 -1589
rect -1458 -2165 -1452 -1589
rect -1498 -2177 -1452 -2165
rect -1380 -1589 -1334 -1577
rect -1380 -2165 -1374 -1589
rect -1340 -2165 -1334 -1589
rect -1380 -2177 -1334 -2165
rect -1262 -1589 -1216 -1577
rect -1262 -2165 -1256 -1589
rect -1222 -2165 -1216 -1589
rect -1262 -2177 -1216 -2165
rect -1144 -1589 -1098 -1577
rect -1144 -2165 -1138 -1589
rect -1104 -2165 -1098 -1589
rect -1144 -2177 -1098 -2165
rect -1026 -1589 -980 -1577
rect -1026 -2165 -1020 -1589
rect -986 -2165 -980 -1589
rect -1026 -2177 -980 -2165
rect -908 -1589 -862 -1577
rect -908 -2165 -902 -1589
rect -868 -2165 -862 -1589
rect -908 -2177 -862 -2165
rect -790 -1589 -744 -1577
rect -790 -2165 -784 -1589
rect -750 -2165 -744 -1589
rect -790 -2177 -744 -2165
rect -672 -1589 -626 -1577
rect -672 -2165 -666 -1589
rect -632 -2165 -626 -1589
rect -672 -2177 -626 -2165
rect -554 -1589 -508 -1577
rect -554 -2165 -548 -1589
rect -514 -2165 -508 -1589
rect -554 -2177 -508 -2165
rect -436 -1589 -390 -1577
rect -436 -2165 -430 -1589
rect -396 -2165 -390 -1589
rect -436 -2177 -390 -2165
rect -318 -1589 -272 -1577
rect -318 -2165 -312 -1589
rect -278 -2165 -272 -1589
rect -318 -2177 -272 -2165
rect -200 -1589 -154 -1577
rect -200 -2165 -194 -1589
rect -160 -2165 -154 -1589
rect -200 -2177 -154 -2165
rect -82 -1589 -36 -1577
rect -82 -2165 -76 -1589
rect -42 -2165 -36 -1589
rect -82 -2177 -36 -2165
rect 36 -1589 82 -1577
rect 36 -2165 42 -1589
rect 76 -2165 82 -1589
rect 36 -2177 82 -2165
rect 154 -1589 200 -1577
rect 154 -2165 160 -1589
rect 194 -2165 200 -1589
rect 154 -2177 200 -2165
rect 272 -1589 318 -1577
rect 272 -2165 278 -1589
rect 312 -2165 318 -1589
rect 272 -2177 318 -2165
rect 390 -1589 436 -1577
rect 390 -2165 396 -1589
rect 430 -2165 436 -1589
rect 390 -2177 436 -2165
rect 508 -1589 554 -1577
rect 508 -2165 514 -1589
rect 548 -2165 554 -1589
rect 508 -2177 554 -2165
rect 626 -1589 672 -1577
rect 626 -2165 632 -1589
rect 666 -2165 672 -1589
rect 626 -2177 672 -2165
rect 744 -1589 790 -1577
rect 744 -2165 750 -1589
rect 784 -2165 790 -1589
rect 744 -2177 790 -2165
rect 862 -1589 908 -1577
rect 862 -2165 868 -1589
rect 902 -2165 908 -1589
rect 862 -2177 908 -2165
rect 980 -1589 1026 -1577
rect 980 -2165 986 -1589
rect 1020 -2165 1026 -1589
rect 980 -2177 1026 -2165
rect 1098 -1589 1144 -1577
rect 1098 -2165 1104 -1589
rect 1138 -2165 1144 -1589
rect 1098 -2177 1144 -2165
rect 1216 -1589 1262 -1577
rect 1216 -2165 1222 -1589
rect 1256 -2165 1262 -1589
rect 1216 -2177 1262 -2165
rect 1334 -1589 1380 -1577
rect 1334 -2165 1340 -1589
rect 1374 -2165 1380 -1589
rect 1334 -2177 1380 -2165
rect 1452 -1589 1498 -1577
rect 1452 -2165 1458 -1589
rect 1492 -2165 1498 -1589
rect 1452 -2177 1498 -2165
rect -1445 -2224 -1387 -2218
rect -1445 -2258 -1433 -2224
rect -1399 -2258 -1387 -2224
rect -1445 -2264 -1387 -2258
rect -1327 -2224 -1269 -2218
rect -1327 -2258 -1315 -2224
rect -1281 -2258 -1269 -2224
rect -1327 -2264 -1269 -2258
rect -1209 -2224 -1151 -2218
rect -1209 -2258 -1197 -2224
rect -1163 -2258 -1151 -2224
rect -1209 -2264 -1151 -2258
rect -1091 -2224 -1033 -2218
rect -1091 -2258 -1079 -2224
rect -1045 -2258 -1033 -2224
rect -1091 -2264 -1033 -2258
rect -973 -2224 -915 -2218
rect -973 -2258 -961 -2224
rect -927 -2258 -915 -2224
rect -973 -2264 -915 -2258
rect -855 -2224 -797 -2218
rect -855 -2258 -843 -2224
rect -809 -2258 -797 -2224
rect -855 -2264 -797 -2258
rect -737 -2224 -679 -2218
rect -737 -2258 -725 -2224
rect -691 -2258 -679 -2224
rect -737 -2264 -679 -2258
rect -619 -2224 -561 -2218
rect -619 -2258 -607 -2224
rect -573 -2258 -561 -2224
rect -619 -2264 -561 -2258
rect -501 -2224 -443 -2218
rect -501 -2258 -489 -2224
rect -455 -2258 -443 -2224
rect -501 -2264 -443 -2258
rect -383 -2224 -325 -2218
rect -383 -2258 -371 -2224
rect -337 -2258 -325 -2224
rect -383 -2264 -325 -2258
rect -265 -2224 -207 -2218
rect -265 -2258 -253 -2224
rect -219 -2258 -207 -2224
rect -265 -2264 -207 -2258
rect -147 -2224 -89 -2218
rect -147 -2258 -135 -2224
rect -101 -2258 -89 -2224
rect -147 -2264 -89 -2258
rect -29 -2224 29 -2218
rect -29 -2258 -17 -2224
rect 17 -2258 29 -2224
rect -29 -2264 29 -2258
rect 89 -2224 147 -2218
rect 89 -2258 101 -2224
rect 135 -2258 147 -2224
rect 89 -2264 147 -2258
rect 207 -2224 265 -2218
rect 207 -2258 219 -2224
rect 253 -2258 265 -2224
rect 207 -2264 265 -2258
rect 325 -2224 383 -2218
rect 325 -2258 337 -2224
rect 371 -2258 383 -2224
rect 325 -2264 383 -2258
rect 443 -2224 501 -2218
rect 443 -2258 455 -2224
rect 489 -2258 501 -2224
rect 443 -2264 501 -2258
rect 561 -2224 619 -2218
rect 561 -2258 573 -2224
rect 607 -2258 619 -2224
rect 561 -2264 619 -2258
rect 679 -2224 737 -2218
rect 679 -2258 691 -2224
rect 725 -2258 737 -2224
rect 679 -2264 737 -2258
rect 797 -2224 855 -2218
rect 797 -2258 809 -2224
rect 843 -2258 855 -2224
rect 797 -2264 855 -2258
rect 915 -2224 973 -2218
rect 915 -2258 927 -2224
rect 961 -2258 973 -2224
rect 915 -2264 973 -2258
rect 1033 -2224 1091 -2218
rect 1033 -2258 1045 -2224
rect 1079 -2258 1091 -2224
rect 1033 -2264 1091 -2258
rect 1151 -2224 1209 -2218
rect 1151 -2258 1163 -2224
rect 1197 -2258 1209 -2224
rect 1151 -2264 1209 -2258
rect 1269 -2224 1327 -2218
rect 1269 -2258 1281 -2224
rect 1315 -2258 1327 -2224
rect 1269 -2264 1327 -2258
rect 1387 -2224 1445 -2218
rect 1387 -2258 1399 -2224
rect 1433 -2258 1445 -2224
rect 1387 -2264 1445 -2258
rect -1498 -2354 -1452 -2342
rect -1498 -2930 -1492 -2354
rect -1458 -2930 -1452 -2354
rect -1498 -2942 -1452 -2930
rect -1380 -2354 -1334 -2342
rect -1380 -2930 -1374 -2354
rect -1340 -2930 -1334 -2354
rect -1380 -2942 -1334 -2930
rect -1262 -2354 -1216 -2342
rect -1262 -2930 -1256 -2354
rect -1222 -2930 -1216 -2354
rect -1262 -2942 -1216 -2930
rect -1144 -2354 -1098 -2342
rect -1144 -2930 -1138 -2354
rect -1104 -2930 -1098 -2354
rect -1144 -2942 -1098 -2930
rect -1026 -2354 -980 -2342
rect -1026 -2930 -1020 -2354
rect -986 -2930 -980 -2354
rect -1026 -2942 -980 -2930
rect -908 -2354 -862 -2342
rect -908 -2930 -902 -2354
rect -868 -2930 -862 -2354
rect -908 -2942 -862 -2930
rect -790 -2354 -744 -2342
rect -790 -2930 -784 -2354
rect -750 -2930 -744 -2354
rect -790 -2942 -744 -2930
rect -672 -2354 -626 -2342
rect -672 -2930 -666 -2354
rect -632 -2930 -626 -2354
rect -672 -2942 -626 -2930
rect -554 -2354 -508 -2342
rect -554 -2930 -548 -2354
rect -514 -2930 -508 -2354
rect -554 -2942 -508 -2930
rect -436 -2354 -390 -2342
rect -436 -2930 -430 -2354
rect -396 -2930 -390 -2354
rect -436 -2942 -390 -2930
rect -318 -2354 -272 -2342
rect -318 -2930 -312 -2354
rect -278 -2930 -272 -2354
rect -318 -2942 -272 -2930
rect -200 -2354 -154 -2342
rect -200 -2930 -194 -2354
rect -160 -2930 -154 -2354
rect -200 -2942 -154 -2930
rect -82 -2354 -36 -2342
rect -82 -2930 -76 -2354
rect -42 -2930 -36 -2354
rect -82 -2942 -36 -2930
rect 36 -2354 82 -2342
rect 36 -2930 42 -2354
rect 76 -2930 82 -2354
rect 36 -2942 82 -2930
rect 154 -2354 200 -2342
rect 154 -2930 160 -2354
rect 194 -2930 200 -2354
rect 154 -2942 200 -2930
rect 272 -2354 318 -2342
rect 272 -2930 278 -2354
rect 312 -2930 318 -2354
rect 272 -2942 318 -2930
rect 390 -2354 436 -2342
rect 390 -2930 396 -2354
rect 430 -2930 436 -2354
rect 390 -2942 436 -2930
rect 508 -2354 554 -2342
rect 508 -2930 514 -2354
rect 548 -2930 554 -2354
rect 508 -2942 554 -2930
rect 626 -2354 672 -2342
rect 626 -2930 632 -2354
rect 666 -2930 672 -2354
rect 626 -2942 672 -2930
rect 744 -2354 790 -2342
rect 744 -2930 750 -2354
rect 784 -2930 790 -2354
rect 744 -2942 790 -2930
rect 862 -2354 908 -2342
rect 862 -2930 868 -2354
rect 902 -2930 908 -2354
rect 862 -2942 908 -2930
rect 980 -2354 1026 -2342
rect 980 -2930 986 -2354
rect 1020 -2930 1026 -2354
rect 980 -2942 1026 -2930
rect 1098 -2354 1144 -2342
rect 1098 -2930 1104 -2354
rect 1138 -2930 1144 -2354
rect 1098 -2942 1144 -2930
rect 1216 -2354 1262 -2342
rect 1216 -2930 1222 -2354
rect 1256 -2930 1262 -2354
rect 1216 -2942 1262 -2930
rect 1334 -2354 1380 -2342
rect 1334 -2930 1340 -2354
rect 1374 -2930 1380 -2354
rect 1334 -2942 1380 -2930
rect 1452 -2354 1498 -2342
rect 1452 -2930 1458 -2354
rect 1492 -2930 1498 -2354
rect 1452 -2942 1498 -2930
rect -1445 -2989 -1387 -2983
rect -1445 -3023 -1433 -2989
rect -1399 -3023 -1387 -2989
rect -1445 -3029 -1387 -3023
rect -1327 -2989 -1269 -2983
rect -1327 -3023 -1315 -2989
rect -1281 -3023 -1269 -2989
rect -1327 -3029 -1269 -3023
rect -1209 -2989 -1151 -2983
rect -1209 -3023 -1197 -2989
rect -1163 -3023 -1151 -2989
rect -1209 -3029 -1151 -3023
rect -1091 -2989 -1033 -2983
rect -1091 -3023 -1079 -2989
rect -1045 -3023 -1033 -2989
rect -1091 -3029 -1033 -3023
rect -973 -2989 -915 -2983
rect -973 -3023 -961 -2989
rect -927 -3023 -915 -2989
rect -973 -3029 -915 -3023
rect -855 -2989 -797 -2983
rect -855 -3023 -843 -2989
rect -809 -3023 -797 -2989
rect -855 -3029 -797 -3023
rect -737 -2989 -679 -2983
rect -737 -3023 -725 -2989
rect -691 -3023 -679 -2989
rect -737 -3029 -679 -3023
rect -619 -2989 -561 -2983
rect -619 -3023 -607 -2989
rect -573 -3023 -561 -2989
rect -619 -3029 -561 -3023
rect -501 -2989 -443 -2983
rect -501 -3023 -489 -2989
rect -455 -3023 -443 -2989
rect -501 -3029 -443 -3023
rect -383 -2989 -325 -2983
rect -383 -3023 -371 -2989
rect -337 -3023 -325 -2989
rect -383 -3029 -325 -3023
rect -265 -2989 -207 -2983
rect -265 -3023 -253 -2989
rect -219 -3023 -207 -2989
rect -265 -3029 -207 -3023
rect -147 -2989 -89 -2983
rect -147 -3023 -135 -2989
rect -101 -3023 -89 -2989
rect -147 -3029 -89 -3023
rect -29 -2989 29 -2983
rect -29 -3023 -17 -2989
rect 17 -3023 29 -2989
rect -29 -3029 29 -3023
rect 89 -2989 147 -2983
rect 89 -3023 101 -2989
rect 135 -3023 147 -2989
rect 89 -3029 147 -3023
rect 207 -2989 265 -2983
rect 207 -3023 219 -2989
rect 253 -3023 265 -2989
rect 207 -3029 265 -3023
rect 325 -2989 383 -2983
rect 325 -3023 337 -2989
rect 371 -3023 383 -2989
rect 325 -3029 383 -3023
rect 443 -2989 501 -2983
rect 443 -3023 455 -2989
rect 489 -3023 501 -2989
rect 443 -3029 501 -3023
rect 561 -2989 619 -2983
rect 561 -3023 573 -2989
rect 607 -3023 619 -2989
rect 561 -3029 619 -3023
rect 679 -2989 737 -2983
rect 679 -3023 691 -2989
rect 725 -3023 737 -2989
rect 679 -3029 737 -3023
rect 797 -2989 855 -2983
rect 797 -3023 809 -2989
rect 843 -3023 855 -2989
rect 797 -3029 855 -3023
rect 915 -2989 973 -2983
rect 915 -3023 927 -2989
rect 961 -3023 973 -2989
rect 915 -3029 973 -3023
rect 1033 -2989 1091 -2983
rect 1033 -3023 1045 -2989
rect 1079 -3023 1091 -2989
rect 1033 -3029 1091 -3023
rect 1151 -2989 1209 -2983
rect 1151 -3023 1163 -2989
rect 1197 -3023 1209 -2989
rect 1151 -3029 1209 -3023
rect 1269 -2989 1327 -2983
rect 1269 -3023 1281 -2989
rect 1315 -3023 1327 -2989
rect 1269 -3029 1327 -3023
rect 1387 -2989 1445 -2983
rect 1387 -3023 1399 -2989
rect 1433 -3023 1445 -2989
rect 1387 -3029 1445 -3023
rect -1498 -3119 -1452 -3107
rect -1498 -3695 -1492 -3119
rect -1458 -3695 -1452 -3119
rect -1498 -3707 -1452 -3695
rect -1380 -3119 -1334 -3107
rect -1380 -3695 -1374 -3119
rect -1340 -3695 -1334 -3119
rect -1380 -3707 -1334 -3695
rect -1262 -3119 -1216 -3107
rect -1262 -3695 -1256 -3119
rect -1222 -3695 -1216 -3119
rect -1262 -3707 -1216 -3695
rect -1144 -3119 -1098 -3107
rect -1144 -3695 -1138 -3119
rect -1104 -3695 -1098 -3119
rect -1144 -3707 -1098 -3695
rect -1026 -3119 -980 -3107
rect -1026 -3695 -1020 -3119
rect -986 -3695 -980 -3119
rect -1026 -3707 -980 -3695
rect -908 -3119 -862 -3107
rect -908 -3695 -902 -3119
rect -868 -3695 -862 -3119
rect -908 -3707 -862 -3695
rect -790 -3119 -744 -3107
rect -790 -3695 -784 -3119
rect -750 -3695 -744 -3119
rect -790 -3707 -744 -3695
rect -672 -3119 -626 -3107
rect -672 -3695 -666 -3119
rect -632 -3695 -626 -3119
rect -672 -3707 -626 -3695
rect -554 -3119 -508 -3107
rect -554 -3695 -548 -3119
rect -514 -3695 -508 -3119
rect -554 -3707 -508 -3695
rect -436 -3119 -390 -3107
rect -436 -3695 -430 -3119
rect -396 -3695 -390 -3119
rect -436 -3707 -390 -3695
rect -318 -3119 -272 -3107
rect -318 -3695 -312 -3119
rect -278 -3695 -272 -3119
rect -318 -3707 -272 -3695
rect -200 -3119 -154 -3107
rect -200 -3695 -194 -3119
rect -160 -3695 -154 -3119
rect -200 -3707 -154 -3695
rect -82 -3119 -36 -3107
rect -82 -3695 -76 -3119
rect -42 -3695 -36 -3119
rect -82 -3707 -36 -3695
rect 36 -3119 82 -3107
rect 36 -3695 42 -3119
rect 76 -3695 82 -3119
rect 36 -3707 82 -3695
rect 154 -3119 200 -3107
rect 154 -3695 160 -3119
rect 194 -3695 200 -3119
rect 154 -3707 200 -3695
rect 272 -3119 318 -3107
rect 272 -3695 278 -3119
rect 312 -3695 318 -3119
rect 272 -3707 318 -3695
rect 390 -3119 436 -3107
rect 390 -3695 396 -3119
rect 430 -3695 436 -3119
rect 390 -3707 436 -3695
rect 508 -3119 554 -3107
rect 508 -3695 514 -3119
rect 548 -3695 554 -3119
rect 508 -3707 554 -3695
rect 626 -3119 672 -3107
rect 626 -3695 632 -3119
rect 666 -3695 672 -3119
rect 626 -3707 672 -3695
rect 744 -3119 790 -3107
rect 744 -3695 750 -3119
rect 784 -3695 790 -3119
rect 744 -3707 790 -3695
rect 862 -3119 908 -3107
rect 862 -3695 868 -3119
rect 902 -3695 908 -3119
rect 862 -3707 908 -3695
rect 980 -3119 1026 -3107
rect 980 -3695 986 -3119
rect 1020 -3695 1026 -3119
rect 980 -3707 1026 -3695
rect 1098 -3119 1144 -3107
rect 1098 -3695 1104 -3119
rect 1138 -3695 1144 -3119
rect 1098 -3707 1144 -3695
rect 1216 -3119 1262 -3107
rect 1216 -3695 1222 -3119
rect 1256 -3695 1262 -3119
rect 1216 -3707 1262 -3695
rect 1334 -3119 1380 -3107
rect 1334 -3695 1340 -3119
rect 1374 -3695 1380 -3119
rect 1334 -3707 1380 -3695
rect 1452 -3119 1498 -3107
rect 1452 -3695 1458 -3119
rect 1492 -3695 1498 -3119
rect 1452 -3707 1498 -3695
rect -1445 -3754 -1387 -3748
rect -1445 -3788 -1433 -3754
rect -1399 -3788 -1387 -3754
rect -1445 -3794 -1387 -3788
rect -1327 -3754 -1269 -3748
rect -1327 -3788 -1315 -3754
rect -1281 -3788 -1269 -3754
rect -1327 -3794 -1269 -3788
rect -1209 -3754 -1151 -3748
rect -1209 -3788 -1197 -3754
rect -1163 -3788 -1151 -3754
rect -1209 -3794 -1151 -3788
rect -1091 -3754 -1033 -3748
rect -1091 -3788 -1079 -3754
rect -1045 -3788 -1033 -3754
rect -1091 -3794 -1033 -3788
rect -973 -3754 -915 -3748
rect -973 -3788 -961 -3754
rect -927 -3788 -915 -3754
rect -973 -3794 -915 -3788
rect -855 -3754 -797 -3748
rect -855 -3788 -843 -3754
rect -809 -3788 -797 -3754
rect -855 -3794 -797 -3788
rect -737 -3754 -679 -3748
rect -737 -3788 -725 -3754
rect -691 -3788 -679 -3754
rect -737 -3794 -679 -3788
rect -619 -3754 -561 -3748
rect -619 -3788 -607 -3754
rect -573 -3788 -561 -3754
rect -619 -3794 -561 -3788
rect -501 -3754 -443 -3748
rect -501 -3788 -489 -3754
rect -455 -3788 -443 -3754
rect -501 -3794 -443 -3788
rect -383 -3754 -325 -3748
rect -383 -3788 -371 -3754
rect -337 -3788 -325 -3754
rect -383 -3794 -325 -3788
rect -265 -3754 -207 -3748
rect -265 -3788 -253 -3754
rect -219 -3788 -207 -3754
rect -265 -3794 -207 -3788
rect -147 -3754 -89 -3748
rect -147 -3788 -135 -3754
rect -101 -3788 -89 -3754
rect -147 -3794 -89 -3788
rect -29 -3754 29 -3748
rect -29 -3788 -17 -3754
rect 17 -3788 29 -3754
rect -29 -3794 29 -3788
rect 89 -3754 147 -3748
rect 89 -3788 101 -3754
rect 135 -3788 147 -3754
rect 89 -3794 147 -3788
rect 207 -3754 265 -3748
rect 207 -3788 219 -3754
rect 253 -3788 265 -3754
rect 207 -3794 265 -3788
rect 325 -3754 383 -3748
rect 325 -3788 337 -3754
rect 371 -3788 383 -3754
rect 325 -3794 383 -3788
rect 443 -3754 501 -3748
rect 443 -3788 455 -3754
rect 489 -3788 501 -3754
rect 443 -3794 501 -3788
rect 561 -3754 619 -3748
rect 561 -3788 573 -3754
rect 607 -3788 619 -3754
rect 561 -3794 619 -3788
rect 679 -3754 737 -3748
rect 679 -3788 691 -3754
rect 725 -3788 737 -3754
rect 679 -3794 737 -3788
rect 797 -3754 855 -3748
rect 797 -3788 809 -3754
rect 843 -3788 855 -3754
rect 797 -3794 855 -3788
rect 915 -3754 973 -3748
rect 915 -3788 927 -3754
rect 961 -3788 973 -3754
rect 915 -3794 973 -3788
rect 1033 -3754 1091 -3748
rect 1033 -3788 1045 -3754
rect 1079 -3788 1091 -3754
rect 1033 -3794 1091 -3788
rect 1151 -3754 1209 -3748
rect 1151 -3788 1163 -3754
rect 1197 -3788 1209 -3754
rect 1151 -3794 1209 -3788
rect 1269 -3754 1327 -3748
rect 1269 -3788 1281 -3754
rect 1315 -3788 1327 -3754
rect 1269 -3794 1327 -3788
rect 1387 -3754 1445 -3748
rect 1387 -3788 1399 -3754
rect 1433 -3788 1445 -3754
rect 1387 -3794 1445 -3788
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1589 -3873 1589 3873
string parameters w 3 l 0.3 m 10 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
