magic
tech sky130A
magscale 1 2
timestamp 1624067212
<< nwell >>
rect -67 720 2436 852
rect -67 696 1642 720
rect 1650 696 2436 720
rect -67 672 2436 696
rect -67 669 1973 672
rect -67 658 1575 669
rect -67 655 1514 658
rect -67 513 485 655
rect 648 573 1514 655
rect 1775 599 1973 669
rect 2015 669 2436 672
rect -67 486 427 513
rect 648 504 1496 573
rect 648 488 1492 504
rect 1493 488 1496 504
rect 1526 492 1852 542
rect 648 486 1505 488
rect 209 380 427 486
rect 681 484 711 486
rect 716 456 1505 486
rect 1533 456 1852 492
rect 716 436 1852 456
rect 716 424 1534 436
rect 716 422 937 424
rect 967 422 1534 424
rect 716 419 1534 422
rect 716 414 1276 419
rect 209 361 479 380
rect 716 364 1017 414
rect 2015 412 2073 669
rect 2353 400 2436 669
<< psubdiff >>
rect -67 -17 82 17
rect 2265 -17 2436 17
<< nsubdiff >>
rect -31 782 129 816
rect 354 782 1299 816
rect 1529 782 2051 816
rect 2233 782 2400 816
<< psubdiffcont >>
rect 82 -17 2265 17
<< nsubdiffcont >>
rect 129 782 354 816
rect 1299 782 1529 816
rect 2051 782 2233 816
<< poly >>
rect 138 742 1419 756
rect 138 740 1369 742
rect 138 706 155 740
rect 189 726 1369 740
rect 189 706 205 726
rect 138 696 205 706
rect 1352 708 1369 726
rect 1403 708 1419 742
rect 1783 742 2259 752
rect 1352 698 1419 708
rect 1496 684 1629 714
rect 1783 708 1800 742
rect 1834 722 2259 742
rect 1834 708 1850 722
rect 1783 698 1850 708
rect 250 659 759 682
rect 250 652 710 659
rect 250 648 280 652
rect 85 618 280 648
rect 693 625 710 652
rect 744 625 761 659
rect 1149 645 1203 647
rect 1132 630 1203 645
rect 1132 626 1159 630
rect 85 600 115 618
rect 693 615 759 625
rect 1035 596 1159 626
rect 1193 596 1203 630
rect 1149 580 1203 596
rect 197 543 269 573
rect 85 188 115 400
rect 197 331 227 543
rect 1035 508 1168 538
rect 1138 488 1168 508
rect 1245 488 1277 603
rect 1496 573 1526 684
rect 2229 654 2259 722
rect 171 314 227 331
rect 171 280 181 314
rect 215 280 227 314
rect 171 264 227 280
rect 197 248 227 264
rect 681 248 711 485
rect 1138 458 1328 488
rect 1184 356 1251 366
rect 1184 342 1201 356
rect 197 218 415 248
rect 385 188 415 218
rect 473 218 711 248
rect 849 322 1201 342
rect 1235 322 1251 356
rect 849 312 1251 322
rect 1298 342 1328 458
rect 1416 428 1484 438
rect 1416 394 1433 428
rect 1467 414 1484 428
rect 1687 414 1717 457
rect 1467 394 1717 414
rect 1416 384 1717 394
rect 1891 418 1921 456
rect 1989 420 2043 437
rect 1989 418 1999 420
rect 1891 388 1999 418
rect 1298 312 1717 342
rect 849 242 879 312
rect 1298 270 1328 312
rect 937 244 1328 270
rect 1438 269 1629 270
rect 937 240 1121 244
rect 1094 220 1121 240
rect 473 188 503 218
rect 1104 210 1121 220
rect 1155 240 1328 244
rect 1155 210 1171 240
rect 1104 200 1171 210
rect 1298 189 1328 240
rect 1431 259 1629 269
rect 1431 225 1447 259
rect 1481 240 1629 259
rect 1687 240 1717 312
rect 1481 225 1499 240
rect 1431 211 1499 225
rect 1891 208 1921 388
rect 1989 386 1999 388
rect 2033 386 2043 420
rect 1989 370 2043 386
rect 2141 189 2171 279
rect 2229 164 2259 295
rect 654 104 721 108
rect 643 98 721 104
rect 473 58 503 76
rect 643 64 671 98
rect 705 64 722 98
rect 641 58 735 64
rect 473 28 2171 58
<< polycont >>
rect 155 706 189 740
rect 1369 708 1403 742
rect 1800 708 1834 742
rect 710 625 744 659
rect 1159 596 1193 630
rect 181 280 215 314
rect 1201 322 1235 356
rect 1433 394 1467 428
rect 1121 210 1155 244
rect 1447 225 1481 259
rect 1999 386 2033 420
rect 671 64 705 98
<< locali >>
rect -31 782 129 816
rect 354 782 1299 816
rect 1529 782 2051 816
rect 2233 782 2400 816
rect 138 706 155 740
rect 189 706 205 740
rect 1352 708 1369 742
rect 1403 708 1419 742
rect 1783 708 1800 742
rect 1834 708 1850 742
rect 693 625 710 659
rect 744 625 761 659
rect 1159 630 1193 647
rect 1159 580 1193 596
rect 1416 394 1433 428
rect 1467 394 1483 428
rect 1999 420 2033 437
rect 1999 370 2033 386
rect 181 314 215 331
rect 1184 322 1201 356
rect 1235 322 1251 356
rect 181 264 215 280
rect 1104 210 1121 244
rect 1155 210 1171 244
rect 1431 225 1447 259
rect 1481 225 1498 259
rect 654 64 671 98
rect 705 64 721 98
rect -59 -17 82 17
rect 2265 -17 2428 17
<< viali >>
rect 129 782 354 816
rect 1299 782 1529 816
rect 2051 782 2233 816
rect 155 706 189 740
rect 1369 708 1403 742
rect 1800 708 1834 742
rect 710 625 744 659
rect 1159 596 1193 630
rect 1433 394 1467 428
rect 1999 386 2033 420
rect 1201 322 1235 356
rect 181 280 215 314
rect 1121 210 1155 244
rect 1447 225 1481 259
rect 671 64 705 98
rect 82 -17 2265 17
<< metal1 >>
rect -31 816 2400 822
rect -31 782 129 816
rect 354 782 1299 816
rect 1529 782 2051 816
rect 2233 782 2400 816
rect -31 776 2400 782
rect 33 574 61 776
rect 138 740 206 748
rect 138 726 155 740
rect 127 706 155 726
rect 189 706 206 740
rect 127 698 206 706
rect 127 574 155 698
rect 295 622 323 776
rect 723 667 759 684
rect 692 659 759 667
rect 692 625 710 659
rect 744 632 759 659
rect 832 638 842 690
rect 894 638 904 690
rect 1009 632 1123 660
rect 1292 647 1320 776
rect 1352 742 1554 748
rect 1352 708 1369 742
rect 1403 720 1554 742
rect 1403 708 1419 720
rect 1352 700 1419 708
rect 744 625 761 632
rect 692 615 761 625
rect 733 578 761 615
rect 825 578 841 584
rect 733 550 841 578
rect 825 547 841 550
rect 1009 544 1067 572
rect 803 439 831 492
rect 655 411 831 439
rect 1039 428 1067 544
rect 139 331 167 394
rect 139 314 223 331
rect 139 280 181 314
rect 215 280 223 314
rect 431 290 459 406
rect 139 263 223 280
rect 139 162 167 263
rect 339 262 549 290
rect 339 157 373 262
rect 515 156 549 262
rect 803 215 831 411
rect 894 400 1067 428
rect 894 216 922 400
rect 1095 372 1123 632
rect 1151 630 1201 647
rect 1526 630 1554 720
rect 1635 742 1851 748
rect 1635 720 1800 742
rect 1151 596 1159 630
rect 1193 617 1201 630
rect 1635 629 1663 720
rect 1783 708 1800 720
rect 1834 708 1851 742
rect 1783 696 1851 708
rect 1927 654 1955 776
rect 2089 654 2119 776
rect 1193 596 1212 617
rect 1151 579 1212 596
rect 982 344 1123 372
rect 1184 364 1212 579
rect 1334 423 1362 521
rect 1769 484 1839 512
rect 1416 428 1484 436
rect 1416 423 1433 428
rect 1334 395 1433 423
rect 1184 356 1252 364
rect 982 216 1010 344
rect 1184 322 1201 356
rect 1235 351 1252 356
rect 1334 351 1362 395
rect 1416 394 1433 395
rect 1467 394 1484 428
rect 1416 386 1484 394
rect 1235 323 1362 351
rect 1235 322 1252 323
rect 1184 314 1252 322
rect 1094 211 1104 265
rect 1172 211 1182 265
rect 1334 245 1362 323
rect 1431 259 1498 267
rect 1431 245 1447 259
rect 1334 225 1447 245
rect 1481 225 1498 259
rect 1334 217 1498 225
rect 1334 216 1431 217
rect 1556 216 1584 482
rect 1644 216 1672 482
rect 1848 216 1876 482
rect 1991 431 2041 437
rect 1979 376 1989 431
rect 2041 376 2051 431
rect 1989 368 2048 376
rect 2020 219 2048 368
rect 2269 219 2297 300
rect 1104 210 1121 211
rect 1155 210 1172 211
rect 1104 202 1172 210
rect 1334 163 1362 216
rect 2020 191 2297 219
rect 1769 160 1839 188
rect 2098 163 2126 191
rect 2269 163 2297 191
rect 39 23 67 72
rect 430 23 458 103
rect 644 65 654 119
rect 722 65 732 119
rect 654 64 671 65
rect 705 64 722 65
rect 654 56 722 64
rect 1253 23 1281 126
rect 1927 24 1955 126
rect 2186 24 2214 73
rect 1870 23 2277 24
rect -67 17 2436 23
rect -67 -17 82 17
rect 2265 -17 2436 17
rect -67 -23 2436 -17
<< via1 >>
rect 842 638 894 690
rect 1104 244 1172 265
rect 1104 211 1121 244
rect 1121 211 1155 244
rect 1155 211 1172 244
rect 1989 420 2041 431
rect 1989 386 1999 420
rect 1999 386 2033 420
rect 2033 386 2041 420
rect 1989 376 2041 386
rect 654 98 722 119
rect 654 65 671 98
rect 671 65 705 98
rect 705 65 722 98
<< metal2 >>
rect 842 690 894 700
rect 842 628 894 638
rect 1989 431 2041 441
rect 1989 366 2041 376
rect 1104 265 1172 275
rect 1104 201 1172 211
rect 654 119 722 129
rect 654 55 722 65
<< comment >>
rect 0 799 464 800
rect 1275 799 1529 800
rect 1866 799 2395 800
rect 0 1 1 799
rect 2394 1 2395 799
rect 0 0 2395 1
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_1
timestamp 1615600491
transform 1 0 400 0 1 147
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_2
timestamp 1615600491
transform 1 0 488 0 1 147
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615600491
transform 1 0 100 0 1 117
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_1
timestamp 1615600491
transform 0 1 475 -1 0 558
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_0
timestamp 1615600491
transform 0 1 475 -1 0 470
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_0
timestamp 1615851015
transform 1 0 100 0 1 484
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_3
timestamp 1615600491
transform 1 0 864 0 1 171
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_4
timestamp 1615600491
transform 1 0 952 0 1 171
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_1
timestamp 1615851015
transform 0 1 919 -1 0 611
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_3
timestamp 1615851015
transform 0 1 919 -1 0 523
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_5
timestamp 1615600491
transform 1 0 1313 0 1 171
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_2
timestamp 1615851015
transform 0 1 1382 -1 0 588
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_7
timestamp 1615600491
transform 1 0 1702 0 1 171
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_6
timestamp 1615600491
transform 1 0 1614 0 1 171
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_8
timestamp 1615600491
transform 1 0 1906 0 1 171
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_5
timestamp 1615851015
transform 1 0 1906 0 1 564
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_4
timestamp 1615851015
transform 1 0 1614 0 1 572
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_6
timestamp 1615851015
transform 1 0 1702 0 1 572
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_9
timestamp 1615600491
transform 1 0 2244 0 1 118
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_10
timestamp 1615600491
transform 1 0 2156 0 1 118
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_3
timestamp 1615600491
transform 1 0 2244 0 1 474
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_2
timestamp 1615600491
transform 1 0 2156 0 1 474
box -109 -242 109 242
<< labels >>
rlabel metal2 1104 211 1172 265 1 CLK
rlabel via1 842 638 894 690 1 D
rlabel metal2 654 65 722 119 1 CLR
rlabel metal1 1857 325 1860 329 1 Qb
rlabel metal1 660 -13 690 14 1 vss
rlabel metal1 640 791 674 813 1 vdd
rlabel metal2 1989 376 2041 431 1 Q
<< end >>
