magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 8885 3173 8920 3190
rect 8849 3156 8920 3173
rect 8516 3120 8551 3137
rect 8480 3103 8551 3120
rect 8147 3067 8182 3084
rect 8111 3050 8182 3067
rect 7778 3014 7813 3031
rect 7742 2997 7813 3014
rect 7409 2961 7444 2978
rect 7373 2944 7444 2961
rect 7040 2891 7075 2925
rect 6671 2838 6706 2872
rect 6302 2802 6337 2819
rect 6266 2785 6337 2802
rect 5933 2732 5968 2766
rect 449 2680 467 2732
rect 477 2680 495 2732
rect 5564 2679 5599 2713
rect 449 2644 467 2650
rect 477 2644 495 2650
rect 1335 2606 1353 2644
rect 501 2560 510 2603
rect 348 2492 456 2549
rect 501 2526 647 2560
rect 398 2459 524 2492
rect 709 2486 906 2560
rect 721 2482 838 2486
rect 1329 2484 1353 2606
rect 1363 2578 1381 2644
rect 5195 2643 5230 2660
rect 5159 2626 5230 2643
rect 1357 2488 1381 2578
rect 4826 2573 4861 2607
rect 4457 2520 4492 2554
rect 4122 2492 4385 2501
rect 418 2455 444 2459
rect 731 2456 838 2482
rect 1153 2460 1353 2484
rect 4052 2467 4385 2492
rect 452 2455 478 2456
rect 452 2437 487 2455
rect 652 2448 838 2456
rect 652 2445 704 2448
rect 533 2440 643 2444
rect 49 2370 68 2435
rect 416 2422 487 2437
rect 521 2433 655 2440
rect 663 2433 693 2445
rect 521 2422 704 2433
rect 83 2374 256 2401
rect 357 2390 409 2401
rect 368 2378 398 2390
rect 83 2306 110 2374
rect 157 2367 209 2374
rect 357 2367 409 2378
rect 183 2332 198 2357
rect 209 2356 286 2360
rect 181 2328 258 2332
rect 183 2315 198 2328
rect 225 2306 240 2315
rect 244 2306 258 2328
rect 272 2306 286 2356
rect 399 2306 409 2367
rect 416 2306 486 2422
rect 731 2418 838 2448
rect 1001 2418 1092 2436
rect 1125 2432 1381 2456
rect 1559 2420 1644 2454
rect 1750 2420 1969 2452
rect 3981 2448 4016 2455
rect 3753 2437 4016 2448
rect 3683 2431 4016 2437
rect 555 2388 621 2406
rect 663 2388 693 2412
rect 560 2372 693 2388
rect 621 2368 693 2372
rect 621 2360 626 2368
rect 621 2354 656 2360
rect 594 2340 656 2354
rect 594 2338 655 2340
rect 598 2334 643 2338
rect 47 2250 486 2306
rect 570 2286 587 2328
rect 598 2314 615 2334
rect 663 2314 693 2368
rect 768 2331 802 2349
rect 985 2331 1092 2418
rect 3576 2414 4016 2431
rect 4052 2414 4367 2467
rect 1564 2384 1576 2386
rect 1156 2331 1171 2378
rect 1252 2350 1259 2362
rect 1190 2331 1271 2350
rect 768 2295 838 2331
rect 985 2316 1271 2331
rect 1286 2339 1380 2350
rect 1414 2349 1466 2350
rect 1414 2339 1499 2349
rect 1818 2346 1830 2384
rect 3350 2378 3385 2395
rect 3314 2361 3385 2378
rect 1286 2316 1293 2339
rect 1303 2332 1369 2339
rect 1425 2331 1499 2339
rect 1870 2338 2030 2348
rect 1870 2337 1911 2338
rect 1529 2331 1540 2337
rect 1881 2331 1911 2337
rect 1953 2337 2030 2338
rect 2092 2337 2144 2348
rect 2180 2347 2204 2348
rect 1425 2327 1871 2331
rect 1414 2316 1871 2327
rect 985 2295 1224 2316
rect 785 2294 928 2295
rect 948 2294 1224 2295
rect 566 2273 600 2284
rect 612 2273 642 2284
rect 654 2273 688 2284
rect 564 2261 612 2273
rect 642 2269 700 2273
rect 651 2263 700 2269
rect 642 2261 700 2263
rect 566 2258 612 2261
rect 566 2250 609 2258
rect 654 2250 700 2261
rect 47 2243 755 2250
rect 47 2225 768 2243
rect 785 2242 1224 2294
rect 1225 2242 1258 2316
rect 1308 2270 1422 2282
rect 1348 2260 1404 2270
rect 1332 2242 1404 2260
rect 1449 2263 1871 2316
rect 1881 2314 1943 2331
rect 1953 2324 2019 2337
rect 2103 2325 2133 2337
rect 2092 2316 2133 2325
rect 2193 2316 2204 2327
rect 2322 2325 2499 2346
rect 2981 2325 3016 2342
rect 2092 2314 2204 2316
rect 1881 2297 1888 2314
rect 1881 2263 1909 2297
rect 785 2225 1271 2242
rect 1276 2240 1420 2242
rect 1276 2236 1447 2240
rect 1449 2236 1909 2263
rect 1996 2244 2023 2262
rect 2103 2244 2104 2282
rect 2170 2271 2204 2314
rect 2576 2272 2787 2325
rect 2945 2308 3016 2325
rect 2175 2266 2204 2271
rect 2170 2244 2204 2252
rect 1276 2231 1909 2236
rect 47 2216 1271 2225
rect 1287 2221 1317 2231
rect 1325 2222 1909 2231
rect 1325 2221 1889 2222
rect 1287 2219 1889 2221
rect 47 2160 486 2216
rect 579 2170 609 2216
rect 654 2208 1271 2216
rect 1276 2208 1889 2219
rect 654 2192 1224 2208
rect 667 2178 700 2192
rect 46 2154 486 2160
rect 47 2136 486 2154
rect 566 2142 609 2170
rect 642 2148 700 2178
rect 642 2142 670 2148
rect 685 2142 700 2148
rect 566 2136 629 2142
rect 642 2136 700 2142
rect 711 2136 1224 2192
rect 47 2119 1224 2136
rect -14 2113 1224 2119
rect 1225 2187 1258 2208
rect 1332 2202 1359 2208
rect 1332 2198 1426 2202
rect 1225 2113 1271 2187
rect 1350 2182 1426 2198
rect 1432 2201 1889 2208
rect 1894 2201 1909 2222
rect 1350 2174 1430 2182
rect 1304 2171 1342 2174
rect 1304 2168 1338 2171
rect 1304 2167 1342 2168
rect 1350 2167 1372 2174
rect 1375 2168 1430 2174
rect 1292 2140 1351 2167
rect 1274 2113 1351 2140
rect 1359 2113 1372 2167
rect 1380 2167 1430 2168
rect 1432 2167 1909 2201
rect 1928 2237 2204 2244
rect 2207 2237 2533 2272
rect 1928 2236 2533 2237
rect 2576 2255 2647 2272
rect 1928 2227 2559 2236
rect 2576 2227 2646 2255
rect 1928 2210 2646 2227
rect 1928 2183 1962 2210
rect 1996 2196 2023 2210
rect 2103 2196 2104 2210
rect 2014 2187 2023 2196
rect 1970 2183 2124 2187
rect 2170 2183 2204 2210
rect 2207 2183 2646 2210
rect 1380 2152 1909 2167
rect 1392 2150 1909 2152
rect 1934 2150 1939 2183
rect 1951 2174 2646 2183
rect 2758 2187 2816 2193
rect 1951 2156 2647 2174
rect 2758 2167 2770 2187
rect 2758 2156 2772 2167
rect 2802 2156 2804 2167
rect 2945 2156 3015 2308
rect 3127 2240 3185 2246
rect 3127 2206 3139 2240
rect 3127 2200 3185 2206
rect 1951 2150 3015 2156
rect 1392 2149 3015 2150
rect 1392 2130 1909 2149
rect 1398 2113 1909 2130
rect -14 2102 1909 2113
rect -14 1952 486 2102
rect 519 2100 629 2102
rect 553 2093 629 2100
rect 553 2089 628 2093
rect 553 2088 587 2089
rect 594 2088 628 2089
rect 641 2089 1909 2102
rect 641 2088 675 2089
rect 682 2088 1909 2089
rect 506 2072 540 2076
rect 541 2073 628 2088
rect 547 2072 628 2073
rect 629 2072 1909 2088
rect 506 2050 546 2072
rect 547 2052 1909 2072
rect 547 2050 628 2052
rect 506 2046 628 2050
rect 629 2046 640 2052
rect 641 2046 1909 2052
rect 506 2012 1909 2046
rect 506 2006 628 2012
rect 629 2006 640 2012
rect 641 2006 675 2012
rect 506 2000 675 2006
rect 506 1957 587 2000
rect 492 1954 587 1957
rect 594 1996 675 2000
rect 594 1954 634 1996
rect 492 1953 634 1954
rect 492 1952 546 1953
rect -14 1944 546 1952
rect 547 1944 634 1953
rect 635 1944 675 1996
rect 682 1944 1909 2012
rect -14 1927 1909 1944
rect -14 1920 412 1927
rect 418 1920 446 1927
rect 452 1920 1909 1927
rect -14 1910 1909 1920
rect -14 1892 464 1910
rect 492 1906 546 1910
rect 547 1908 574 1910
rect 486 1894 546 1906
rect 553 1904 574 1908
rect 580 1908 1909 1910
rect 580 1894 640 1908
rect 480 1892 546 1894
rect 568 1892 640 1894
rect 641 1892 1909 1908
rect -14 1878 412 1892
rect 418 1888 452 1892
rect 480 1880 540 1892
rect 568 1888 628 1892
rect 480 1878 526 1880
rect 568 1878 626 1888
rect 640 1878 675 1892
rect 682 1888 1909 1892
rect 694 1878 1909 1888
rect -14 1866 467 1878
rect 477 1866 526 1878
rect 540 1867 1909 1878
rect 540 1866 614 1867
rect 620 1866 1909 1867
rect -14 1864 1909 1866
rect -14 1847 412 1864
rect 438 1847 1909 1864
rect -14 1842 1909 1847
rect -14 1837 1871 1842
rect 1874 1837 1909 1842
rect 1928 2138 2002 2149
rect 2014 2138 2033 2149
rect 1928 2097 2033 2138
rect 2050 2128 2065 2149
rect 2070 2142 2102 2149
rect 2070 2128 2136 2142
rect 2050 2115 2136 2128
rect 2170 2120 3015 2149
rect 2050 2097 2102 2115
rect 2120 2108 2124 2115
rect 1928 2083 2039 2097
rect 2044 2083 2102 2097
rect 1928 2061 2102 2083
rect 2136 2061 2164 2065
rect 1928 2049 2103 2061
rect 1928 2047 2090 2049
rect 1928 2041 2039 2047
rect 2042 2041 2090 2047
rect 1928 2034 2090 2041
rect 1928 2031 2039 2034
rect 1928 2000 2027 2031
rect 2033 2013 2039 2031
rect 2034 2000 2039 2013
rect 2042 2004 2090 2034
rect 2118 2046 2164 2061
rect 2118 2038 2133 2046
rect 2136 2038 2164 2046
rect 2042 2000 2110 2004
rect 2118 2003 2164 2038
rect 2170 2003 3016 2120
rect 3083 2078 3141 2121
rect 3171 2078 3229 2121
rect 3314 2103 3384 2361
rect 3496 2293 3554 2299
rect 3496 2259 3508 2293
rect 3496 2253 3554 2259
rect 3576 2250 4015 2414
rect 4035 2295 4367 2414
rect 4423 2329 4438 2501
rect 4412 2304 4438 2329
rect 4404 2295 4438 2304
rect 4457 2295 4491 2520
rect 4603 2452 4661 2458
rect 4603 2418 4615 2452
rect 4603 2412 4661 2418
rect 4792 2386 4807 2554
rect 4826 2386 4860 2573
rect 4972 2505 5030 2511
rect 4972 2471 4984 2505
rect 4972 2465 5030 2471
rect 4683 2380 5105 2386
rect 4665 2350 5105 2380
rect 4683 2333 5105 2350
rect 5159 2333 5229 2626
rect 5341 2558 5399 2564
rect 5341 2524 5353 2558
rect 5341 2518 5399 2524
rect 4571 2302 4605 2329
rect 4683 2297 5229 2333
rect 5309 2309 5343 2331
rect 5297 2297 5354 2309
rect 5438 2297 5443 2322
rect 4683 2295 5342 2297
rect 4035 2288 5342 2295
rect 5355 2288 5385 2297
rect 5403 2288 5438 2297
rect 4035 2263 5438 2288
rect 5530 2278 5545 2660
rect 4035 2261 5229 2263
rect 4035 2250 4493 2261
rect 4603 2252 4661 2258
rect 3576 2216 4493 2250
rect 3576 2212 4015 2216
rect 3573 2134 4015 2212
rect 3314 2101 3421 2103
rect 3095 2074 3129 2078
rect 3183 2074 3217 2078
rect 2118 2000 3016 2003
rect 1928 1985 2033 2000
rect 2036 1997 3016 2000
rect 2036 1990 2076 1997
rect 2088 1990 3016 1997
rect 1928 1837 1962 1985
rect 1968 1981 2034 1985
rect 1988 1972 2034 1981
rect 1978 1970 2034 1972
rect 1976 1944 2034 1970
rect 2036 1944 3016 1990
rect 1976 1942 3016 1944
rect 1976 1938 2034 1942
rect 2042 1938 3016 1942
rect 3035 2040 3251 2067
rect 3297 2050 3421 2101
rect 3576 2050 4015 2134
rect 3035 2033 3070 2040
rect 3112 2033 3200 2040
rect 3297 2033 4015 2050
rect 3035 1938 3069 2033
rect 3127 2023 3139 2033
rect 3127 2000 3189 2023
rect 3135 1990 3189 2000
rect 3314 1997 4015 2033
rect 4035 2193 4493 2216
rect 4599 2227 4665 2252
rect 4599 2202 4600 2227
rect 4603 2218 4615 2227
rect 4632 2218 4665 2227
rect 4603 2212 4661 2218
rect 4496 2193 4554 2199
rect 4035 2184 4538 2193
rect 4035 2159 4558 2184
rect 4666 2172 5229 2261
rect 5342 2256 5355 2263
rect 5385 2256 5438 2263
rect 5341 2250 5438 2256
rect 5337 2239 5438 2250
rect 5519 2244 5545 2278
rect 5564 2244 5598 2679
rect 5710 2611 5768 2617
rect 5710 2577 5722 2611
rect 5710 2571 5768 2577
rect 5337 2229 5403 2239
rect 5234 2195 5292 2201
rect 5337 2200 5338 2229
rect 5341 2216 5353 2229
rect 5370 2216 5403 2229
rect 5341 2210 5399 2216
rect 5230 2182 5267 2195
rect 5230 2172 5296 2182
rect 4666 2161 5296 2172
rect 4035 2150 4493 2159
rect 4496 2153 4554 2159
rect 4666 2155 5292 2161
rect 4666 2150 5248 2155
rect 4035 2148 5248 2150
rect 5278 2148 5291 2155
rect 5404 2148 5438 2239
rect 5457 2210 5492 2244
rect 5553 2210 5812 2244
rect 5899 2225 5914 2713
rect 5457 2148 5491 2210
rect 5511 2148 5545 2210
rect 4035 2133 5449 2148
rect 4035 2125 4861 2133
rect 4035 2121 4493 2125
rect 4510 2121 4540 2125
rect 4553 2121 4861 2125
rect 4035 2116 4861 2121
rect 4035 2027 4493 2116
rect 4035 1997 4069 2027
rect 4123 2012 4223 2027
rect 4123 1997 4169 2012
rect 4177 2006 4185 2012
rect 3314 1996 4169 1997
rect 3193 1971 3227 1972
rect 3181 1965 3239 1971
rect 3181 1938 3193 1965
rect 3314 1947 4159 1996
rect 4205 1978 4223 2012
rect 4297 1962 4493 2027
rect 4666 2080 4843 2116
rect 4666 2034 4753 2080
rect 4666 2008 4818 2034
rect 4496 1993 4554 1999
rect 4496 1964 4508 1993
rect 4496 1962 4530 1964
rect 3297 1944 4159 1947
rect 4204 1944 4245 1960
rect 4297 1959 4530 1962
rect 4297 1953 4554 1959
rect 4666 1953 4846 2008
rect 4297 1944 4528 1953
rect 3297 1938 4257 1944
rect 1976 1906 3016 1938
rect 1976 1898 2116 1906
rect 1976 1888 2034 1898
rect 2036 1893 2116 1898
rect 2036 1890 2070 1893
rect 2076 1890 2116 1893
rect 1976 1878 2028 1888
rect 2036 1881 2116 1890
rect 2122 1881 3016 1906
rect 3017 1926 4257 1938
rect 3017 1910 4272 1926
rect 3017 1904 4275 1910
rect 2042 1878 2118 1881
rect 2130 1878 2164 1881
rect 2170 1878 3016 1881
rect 1976 1877 3016 1878
rect 1976 1856 2070 1877
rect 2076 1856 3016 1877
rect 1976 1837 3016 1856
rect -14 1790 3016 1837
rect -14 1785 526 1790
rect -14 1779 520 1785
rect -14 1773 538 1779
rect 549 1773 690 1790
rect -14 1754 486 1773
rect 492 1769 520 1773
rect 9 1734 43 1754
rect 9 1566 30 1734
rect 32 1723 43 1734
rect 35 1589 43 1723
rect 69 1734 486 1754
rect 580 1762 690 1773
rect 580 1754 648 1762
rect 694 1754 1539 1790
rect 580 1735 660 1754
rect 69 1696 117 1734
rect 123 1729 151 1734
rect 169 1729 257 1734
rect 119 1725 206 1729
rect 211 1725 245 1729
rect 119 1714 169 1725
rect 211 1709 248 1725
rect 325 1721 520 1734
rect 580 1732 644 1735
rect 646 1732 660 1735
rect 556 1730 660 1732
rect 556 1726 582 1730
rect 584 1728 660 1730
rect 694 1746 964 1754
rect 1063 1750 1539 1754
rect 1559 1788 2136 1790
rect 2190 1788 3016 1790
rect 1559 1784 3016 1788
rect 1559 1782 2106 1784
rect 2110 1782 3016 1784
rect 1559 1779 2026 1782
rect 1559 1773 2078 1779
rect 1559 1751 2082 1773
rect 2190 1762 3016 1782
rect 2190 1760 2224 1762
rect 694 1729 838 1746
rect 1063 1734 1540 1750
rect 865 1729 884 1734
rect 584 1726 656 1728
rect 546 1721 656 1726
rect 325 1720 660 1721
rect 325 1714 656 1720
rect 694 1718 868 1729
rect 1063 1723 1074 1734
rect 325 1712 586 1714
rect 594 1712 628 1714
rect 325 1710 628 1712
rect 183 1699 277 1709
rect 183 1696 275 1699
rect 325 1696 486 1710
rect 58 1664 486 1696
rect 520 1704 628 1710
rect 694 1705 840 1718
rect 694 1704 1061 1705
rect 1080 1704 1540 1734
rect 1587 1739 2082 1751
rect 2138 1754 2224 1760
rect 2138 1752 2184 1754
rect 1587 1734 2078 1739
rect 2138 1734 2150 1752
rect 2190 1734 2224 1754
rect 1587 1732 2082 1734
rect 2134 1732 2152 1734
rect 2182 1732 2224 1734
rect 2244 1732 2278 1762
rect 1587 1723 2255 1732
rect 1587 1720 2222 1723
rect 1587 1707 2200 1720
rect 520 1694 684 1704
rect 694 1694 1540 1704
rect 520 1692 1540 1694
rect 540 1683 546 1692
rect 548 1686 1540 1692
rect 548 1683 600 1686
rect 540 1670 600 1683
rect 606 1683 634 1686
rect 640 1683 1540 1686
rect 606 1670 1540 1683
rect 518 1668 600 1670
rect 628 1668 1540 1670
rect 540 1664 600 1668
rect 606 1664 1540 1668
rect 58 1650 1540 1664
rect 1545 1704 2200 1707
rect 2224 1708 2262 1711
rect 2263 1708 2278 1732
rect 1545 1703 2193 1704
rect 2224 1703 2278 1708
rect 1545 1698 2201 1703
rect 1545 1671 2026 1698
rect 2072 1688 2128 1695
rect 2190 1692 2201 1698
rect 2213 1698 2278 1703
rect 2213 1692 2224 1698
rect 2072 1673 2140 1688
rect 2190 1684 2224 1692
rect 2190 1673 2228 1684
rect 2297 1679 2342 1762
rect 2361 1679 2395 1762
rect 2455 1759 2477 1762
rect 2455 1752 2611 1759
rect 2461 1734 2611 1752
rect 2612 1743 3016 1762
rect 2439 1731 2505 1734
rect 2613 1707 3016 1743
rect 2507 1701 2565 1707
rect 2507 1688 2519 1701
rect 2507 1686 2553 1688
rect 2613 1686 2747 1707
rect 2812 1694 2824 1707
rect 2812 1688 2870 1694
rect 2982 1688 3016 1707
rect 2982 1686 2996 1688
rect 3001 1686 3016 1688
rect 3035 1733 3069 1904
rect 3167 1897 3305 1904
rect 3149 1893 3305 1897
rect 3137 1885 3305 1893
rect 3314 1892 4275 1904
rect 4311 1894 4528 1944
rect 3314 1885 4176 1892
rect 4211 1888 4245 1890
rect 3071 1870 4176 1885
rect 3071 1851 3123 1870
rect 3137 1851 3283 1870
rect 3314 1856 4176 1870
rect 4314 1856 4528 1894
rect 3314 1854 4528 1856
rect 3071 1733 3105 1851
rect 3137 1765 3159 1851
rect 3314 1830 4235 1854
rect 3314 1822 4253 1830
rect 4262 1824 4528 1854
rect 4264 1822 4528 1824
rect 3237 1817 3275 1821
rect 3179 1765 3183 1817
rect 3237 1799 3297 1817
rect 3137 1733 3195 1765
rect 3213 1749 3217 1783
rect 3225 1749 3297 1799
rect 3314 1815 4176 1822
rect 4297 1821 4528 1822
rect 3314 1796 4195 1815
rect 3314 1762 4219 1796
rect 4297 1765 4331 1821
rect 4332 1774 4350 1806
rect 3225 1733 3283 1749
rect 3314 1744 4207 1762
rect 4274 1752 4412 1765
rect 4274 1747 4431 1752
rect 4263 1744 4431 1747
rect 4458 1744 4492 1821
rect 4683 1750 4846 1953
rect 4865 1940 4923 1946
rect 4865 1906 4877 1940
rect 4865 1900 4923 1906
rect 5054 1804 5069 2133
rect 5088 1837 5122 2133
rect 5196 2127 5449 2133
rect 5248 2114 5278 2127
rect 5291 2114 5449 2127
rect 5457 2114 5483 2148
rect 5530 2114 5545 2148
rect 5190 2089 5195 2114
rect 5234 1887 5292 1893
rect 5234 1853 5246 1887
rect 5234 1847 5292 1853
rect 5404 1847 5438 2114
rect 5423 1837 5438 1847
rect 5457 1837 5491 2114
rect 5564 2021 5598 2210
rect 5772 2191 5812 2210
rect 5888 2191 5914 2225
rect 5933 2191 5967 2732
rect 6079 2664 6137 2670
rect 6079 2630 6091 2664
rect 6079 2624 6137 2630
rect 6266 2415 6336 2785
rect 6448 2717 6506 2723
rect 6448 2683 6460 2717
rect 6448 2677 6506 2683
rect 6448 2517 6506 2523
rect 6448 2483 6460 2517
rect 6448 2477 6506 2483
rect 6266 2381 6337 2415
rect 6637 2400 6652 2819
rect 6671 2468 6705 2838
rect 6817 2770 6875 2776
rect 6817 2736 6829 2770
rect 6817 2730 6875 2736
rect 6817 2570 6875 2576
rect 6817 2536 6829 2570
rect 6817 2530 6875 2536
rect 6671 2434 6706 2468
rect 7006 2453 7021 2872
rect 7040 2521 7074 2891
rect 7186 2823 7244 2829
rect 7186 2789 7198 2823
rect 7186 2783 7244 2789
rect 7186 2623 7244 2629
rect 7186 2589 7198 2623
rect 7186 2583 7244 2589
rect 7040 2487 7075 2521
rect 7373 2487 7443 2944
rect 7555 2876 7613 2882
rect 7555 2842 7567 2876
rect 7555 2836 7613 2842
rect 7742 2627 7812 2997
rect 7924 2929 7982 2935
rect 7924 2895 7936 2929
rect 7924 2889 7982 2895
rect 7924 2729 7982 2735
rect 7924 2695 7936 2729
rect 7924 2689 7982 2695
rect 7742 2593 7813 2627
rect 8111 2593 8181 3050
rect 8293 2982 8351 2988
rect 8293 2948 8305 2982
rect 8293 2942 8351 2948
rect 8480 2733 8550 3103
rect 8662 3035 8720 3041
rect 8662 3001 8674 3035
rect 8662 2995 8720 3001
rect 8662 2835 8720 2841
rect 8662 2801 8674 2835
rect 8662 2795 8720 2801
rect 8480 2699 8551 2733
rect 8849 2699 8919 3156
rect 9031 3088 9089 3094
rect 9031 3054 9043 3088
rect 9031 3048 9089 3054
rect 9031 2780 9089 2786
rect 9031 2746 9043 2780
rect 9031 2740 9089 2746
rect 8293 2674 8351 2680
rect 8293 2640 8305 2674
rect 8480 2663 8533 2699
rect 8849 2663 8902 2699
rect 8293 2634 8351 2640
rect 7555 2568 7613 2574
rect 7555 2534 7567 2568
rect 7742 2557 7795 2593
rect 8111 2557 8164 2593
rect 7555 2528 7613 2534
rect 7373 2451 7426 2487
rect 6266 2345 6319 2381
rect 6035 2225 6075 2245
rect 6141 2225 6181 2245
rect 6035 2223 6081 2225
rect 6047 2219 6081 2223
rect 6135 2223 6181 2225
rect 6135 2219 6169 2223
rect 5666 2182 5678 2189
rect 5666 2176 5696 2182
rect 5666 2170 5699 2176
rect 5773 2170 5812 2191
rect 5826 2170 5866 2191
rect 5922 2185 6176 2191
rect 5922 2174 6163 2185
rect 5678 2166 5699 2170
rect 5792 2161 5807 2170
rect 5603 2142 5661 2148
rect 5664 2142 5665 2158
rect 5599 2108 5636 2142
rect 5649 2132 5665 2142
rect 5603 2102 5661 2108
rect 5706 2099 5707 2139
rect 5710 2123 5768 2129
rect 5710 2108 5722 2123
rect 5739 2108 5772 2123
rect 5710 2099 5772 2108
rect 5706 2089 5772 2099
rect 5710 2083 5768 2089
rect 5672 2061 5693 2065
rect 5672 2058 5705 2061
rect 5672 2055 5699 2058
rect 5626 2049 5693 2055
rect 5626 2021 5659 2049
rect 5773 2021 5807 2161
rect 5826 2157 5861 2170
rect 5922 2157 6176 2174
rect 5564 1987 5818 2021
rect 5559 1881 5617 1910
rect 5647 1881 5705 1910
rect 5571 1877 5605 1881
rect 5659 1877 5693 1881
rect 5617 1856 5683 1868
rect 5773 1856 5807 1987
rect 5521 1843 5807 1856
rect 5521 1837 5556 1843
rect 5088 1822 5556 1837
rect 5577 1834 5807 1843
rect 5599 1833 5807 1834
rect 5588 1822 5807 1833
rect 5088 1801 5555 1822
rect 5603 1806 5615 1822
rect 5621 1806 5665 1812
rect 5088 1764 5103 1801
rect 5116 1764 5555 1801
rect 5599 1784 5665 1806
rect 5773 1794 5807 1822
rect 5088 1751 5555 1764
rect 5773 1764 5784 1775
rect 5792 1764 5807 1794
rect 3314 1734 4528 1744
rect 3314 1733 4432 1734
rect 3035 1731 4432 1733
rect 4458 1731 4492 1734
rect 4517 1731 4528 1734
rect 4683 1734 5069 1750
rect 4683 1731 4846 1734
rect 3035 1728 4592 1731
rect 3035 1720 4207 1728
rect 3035 1704 4199 1720
rect 4244 1704 4592 1728
rect 3035 1692 4213 1704
rect 4240 1695 4592 1704
rect 4683 1716 4754 1731
rect 5034 1716 5069 1734
rect 4240 1692 4666 1695
rect 4683 1692 4753 1716
rect 3035 1686 4753 1692
rect 2507 1679 2565 1686
rect 2613 1679 4753 1686
rect 5035 1697 5069 1716
rect 5116 1732 5555 1751
rect 5667 1754 5725 1760
rect 5667 1734 5679 1754
rect 5773 1734 5807 1764
rect 5663 1732 5681 1734
rect 5711 1732 5729 1734
rect 5773 1732 5784 1734
rect 5116 1723 5784 1732
rect 5116 1720 5751 1723
rect 5116 1712 5729 1720
rect 5116 1711 5761 1712
rect 5116 1704 5791 1711
rect 5792 1704 5807 1734
rect 5116 1698 5807 1704
rect 5826 1856 5860 2157
rect 5880 2021 5914 2157
rect 5933 2074 5967 2157
rect 6079 2142 6091 2157
rect 6108 2142 6141 2157
rect 6142 2156 6176 2157
rect 6079 2136 6137 2142
rect 6142 2108 6319 2156
rect 6159 2095 6319 2108
rect 5972 2089 6030 2095
rect 5968 2074 6005 2089
rect 6142 2074 6319 2095
rect 6510 2086 6545 2120
rect 5933 2040 6319 2074
rect 6511 2067 6545 2086
rect 5874 2008 5914 2021
rect 5940 2008 5974 2012
rect 5899 2006 5914 2008
rect 5903 1987 5914 2006
rect 5928 2006 5974 2008
rect 6028 2006 6062 2012
rect 5928 1987 5968 2006
rect 6142 2004 6319 2040
rect 6341 2018 6399 2024
rect 5940 1953 5948 1987
rect 5116 1697 5555 1698
rect 5035 1692 5046 1697
rect 5054 1692 5069 1697
rect 2072 1671 2152 1673
rect 2182 1671 2240 1673
rect 1545 1654 2240 1671
rect 2297 1670 4753 1679
rect 2297 1662 4240 1670
rect 2297 1655 2342 1662
rect 2361 1658 2569 1662
rect 2630 1658 4240 1662
rect 4244 1658 4753 1670
rect 2361 1655 2593 1658
rect 2630 1655 4753 1658
rect 1545 1650 2264 1654
rect 2297 1650 2593 1655
rect 2609 1650 4753 1655
rect 4843 1650 4945 1682
rect 5035 1662 5069 1692
rect 5035 1654 5046 1662
rect 5054 1654 5069 1662
rect 5035 1650 5069 1654
rect 5088 1650 5555 1697
rect 5631 1673 5681 1698
rect 5623 1662 5681 1673
rect 5711 1673 5761 1698
rect 5826 1679 5871 1856
rect 5928 1828 5986 1857
rect 6016 1828 6074 1857
rect 6142 1839 6229 2004
rect 6341 1984 6353 2018
rect 6341 1978 6399 1984
rect 5940 1824 5974 1828
rect 6028 1824 6062 1828
rect 5986 1803 6052 1815
rect 6142 1803 6276 1839
rect 5890 1790 6276 1803
rect 5890 1775 5925 1790
rect 5946 1781 6276 1790
rect 5968 1780 6276 1781
rect 5957 1775 6276 1780
rect 5890 1769 6276 1775
rect 5890 1679 5924 1769
rect 5972 1747 5984 1769
rect 5990 1747 6140 1759
rect 5972 1741 6140 1747
rect 5990 1734 6140 1741
rect 5968 1731 6034 1734
rect 6036 1701 6094 1707
rect 6036 1688 6048 1701
rect 6036 1686 6082 1688
rect 6142 1686 6276 1769
rect 6297 1766 6355 1779
rect 6385 1766 6443 1779
rect 6511 1764 6522 1775
rect 6530 1764 6545 2067
rect 6511 1734 6545 1764
rect 6341 1728 6399 1734
rect 6341 1694 6353 1728
rect 6511 1723 6522 1734
rect 6341 1688 6399 1694
rect 6511 1692 6522 1703
rect 6511 1686 6525 1692
rect 6530 1686 6545 1734
rect 6564 2033 6599 2067
rect 6879 2033 6914 2067
rect 6564 1733 6598 2033
rect 6880 2014 6914 2033
rect 6710 1965 6768 1971
rect 6710 1931 6722 1965
rect 6710 1925 6768 1931
rect 6696 1885 6834 1915
rect 6600 1851 6652 1885
rect 6666 1851 6812 1885
rect 6880 1851 6888 1919
rect 6899 1885 6914 2014
rect 6933 1980 6968 2014
rect 7248 1980 7283 2014
rect 6933 1886 6967 1980
rect 7249 1961 7283 1980
rect 7635 1961 7688 1962
rect 7079 1912 7137 1918
rect 7079 1888 7091 1912
rect 7079 1886 7093 1888
rect 7123 1886 7125 1888
rect 7268 1886 7283 1961
rect 7302 1927 7337 1961
rect 7617 1927 7688 1961
rect 7302 1886 7336 1927
rect 7618 1926 7688 1927
rect 7635 1892 7706 1926
rect 6933 1885 7355 1886
rect 6915 1851 7355 1885
rect 6600 1733 6634 1851
rect 6666 1765 6688 1851
rect 6766 1817 6804 1821
rect 6708 1765 6712 1817
rect 6766 1799 6826 1817
rect 6666 1733 6724 1765
rect 6742 1749 6746 1783
rect 6754 1749 6826 1799
rect 6882 1765 6914 1851
rect 6754 1733 6812 1749
rect 6880 1733 6914 1765
rect 6916 1807 7355 1851
rect 7448 1859 7506 1865
rect 7448 1825 7460 1859
rect 7448 1819 7506 1825
rect 7635 1815 7705 1892
rect 7817 1824 7875 1830
rect 7434 1807 7572 1809
rect 7618 1807 7626 1813
rect 7635 1807 7724 1815
rect 6916 1733 7724 1807
rect 7817 1790 7829 1824
rect 7817 1784 7875 1790
rect 7803 1744 7941 1765
rect 7803 1743 7872 1744
rect 6564 1686 7724 1733
rect 6036 1679 6094 1686
rect 6142 1679 7724 1686
rect 7773 1718 7961 1743
rect 7987 1718 8021 1830
rect 7773 1684 8021 1718
rect 5711 1662 5769 1673
rect 5623 1650 5669 1662
rect 5723 1650 5769 1662
rect 5826 1662 7724 1679
rect 5826 1651 5871 1662
rect 5837 1650 5871 1651
rect 5890 1658 6098 1662
rect 5890 1650 6122 1658
rect 6159 1650 7724 1662
rect 58 1648 7724 1650
rect 58 1622 7741 1648
rect 7748 1622 7769 1684
rect 58 1616 7769 1622
rect 58 1590 728 1616
rect 754 1603 1540 1616
rect 754 1590 1224 1603
rect 58 1572 486 1590
rect 506 1588 1224 1590
rect 9 1555 41 1566
rect 58 1562 500 1572
rect 58 1544 486 1562
rect 506 1548 728 1588
rect 754 1548 1224 1588
rect 1286 1577 1336 1603
rect 1492 1598 1540 1603
rect 1545 1601 1579 1611
rect 1587 1610 2278 1616
rect 1587 1601 2026 1610
rect 1545 1598 2026 1601
rect 1492 1584 2026 1598
rect 2094 1598 2109 1610
rect 2196 1598 2228 1610
rect 2229 1601 2278 1610
rect 2308 1601 2342 1616
rect 2361 1601 2395 1616
rect 2475 1601 2509 1616
rect 2630 1610 5769 1616
rect 5792 1610 5807 1616
rect 2563 1601 2597 1608
rect 2630 1604 5555 1610
rect 2630 1601 4950 1604
rect 2230 1598 2278 1601
rect 2094 1586 2152 1598
rect 1378 1580 1412 1581
rect 1278 1568 1336 1577
rect 1366 1568 1424 1577
rect 1278 1565 1293 1568
rect 1294 1565 1324 1568
rect 1366 1567 1380 1568
rect 1278 1555 1324 1565
rect 1336 1555 1338 1566
rect 1367 1565 1380 1567
rect 1409 1567 1424 1568
rect 1409 1565 1438 1567
rect 1278 1553 1338 1555
rect 58 1534 500 1544
rect 58 1510 486 1534
rect 506 1533 1224 1548
rect 58 1500 500 1510
rect 506 1505 722 1533
rect 58 1482 486 1500
rect 506 1499 716 1505
rect 506 1486 552 1499
rect 554 1493 716 1499
rect 566 1489 716 1493
rect 594 1486 668 1489
rect 682 1486 716 1489
rect 492 1482 552 1486
rect 580 1482 716 1486
rect 58 1474 716 1482
rect 58 1472 714 1474
rect 728 1472 1224 1533
rect 1290 1474 1338 1553
rect 1378 1553 1438 1565
rect 1378 1541 1426 1553
rect 1378 1498 1438 1541
rect 1344 1474 1370 1498
rect 58 1462 728 1472
rect 58 1354 486 1462
rect 492 1460 526 1462
rect 532 1460 540 1462
rect 492 1382 540 1460
rect 576 1456 628 1462
rect 630 1460 702 1462
rect 630 1456 716 1460
rect 576 1446 716 1456
rect 580 1412 716 1446
rect 580 1382 628 1412
rect 634 1406 656 1412
rect 662 1409 716 1412
rect 662 1396 728 1409
rect 634 1382 728 1396
rect 492 1354 728 1382
rect 754 1354 1224 1472
rect 1248 1470 1282 1474
rect 58 1353 765 1354
rect 58 1348 728 1353
rect 768 1348 1224 1354
rect 58 1327 1224 1348
rect 142 1314 1224 1327
rect 282 1274 286 1308
rect 310 1302 314 1308
rect 330 1304 364 1314
rect 384 1310 732 1314
rect 384 1304 452 1310
rect 494 1304 540 1310
rect 347 1302 362 1304
rect 384 1302 450 1304
rect 494 1302 538 1304
rect 347 1301 376 1302
rect 318 1292 376 1301
rect 384 1292 464 1302
rect 494 1300 552 1302
rect 582 1300 640 1310
rect 670 1300 728 1310
rect 768 1304 1224 1314
rect 492 1298 552 1300
rect 580 1298 640 1300
rect 668 1298 728 1300
rect 494 1292 552 1298
rect 582 1292 640 1298
rect 670 1292 728 1298
rect 418 1288 452 1292
rect 506 1288 540 1292
rect 594 1288 628 1292
rect 640 1266 670 1290
rect 682 1288 716 1292
rect 771 1266 1224 1304
rect 1236 1397 1282 1470
rect 1290 1399 1370 1474
rect 1372 1481 1438 1498
rect 1372 1470 1426 1481
rect 1290 1397 1324 1399
rect 1336 1397 1370 1399
rect 1378 1458 1426 1470
rect 1378 1399 1458 1458
rect 1236 1359 1288 1397
rect 1290 1393 1316 1397
rect 1298 1387 1316 1393
rect 1336 1387 1376 1397
rect 1378 1393 1412 1399
rect 1382 1387 1412 1393
rect 1424 1387 1458 1399
rect 1304 1384 1316 1387
rect 1323 1384 1458 1387
rect 1304 1383 1458 1384
rect 1323 1374 1458 1383
rect 1236 1349 1282 1359
rect 1236 1302 1278 1349
rect 1314 1340 1458 1374
rect 1324 1306 1458 1340
rect 1236 1290 1294 1302
rect 1324 1290 1382 1306
rect 1390 1300 1394 1306
rect 1418 1290 1422 1306
rect 1424 1302 1458 1306
rect 1248 1286 1258 1290
rect 1424 1286 1432 1302
rect 1467 1290 1470 1470
rect 1492 1290 1540 1584
rect 16 1212 30 1254
rect 224 1247 406 1256
rect 438 1254 1224 1266
rect 438 1247 494 1254
rect 58 1243 494 1247
rect 538 1243 582 1254
rect 732 1248 1224 1254
rect 588 1243 692 1244
rect 732 1243 1242 1248
rect 58 1232 505 1243
rect 527 1240 692 1243
rect 527 1232 710 1240
rect 721 1232 1242 1243
rect 58 1174 472 1232
rect 754 1231 1242 1232
rect 538 1206 610 1222
rect 538 1198 676 1206
rect 754 1202 776 1231
rect 785 1221 1242 1231
rect 1176 1216 1242 1221
rect 1154 1214 1242 1216
rect 1272 1244 1487 1248
rect 1272 1238 1430 1244
rect 1272 1215 1444 1238
rect 1446 1237 1487 1244
rect 1446 1215 1476 1237
rect 1272 1214 1487 1215
rect 1154 1204 1231 1214
rect 1283 1204 1487 1214
rect 1524 1204 1540 1290
rect 1545 1344 2026 1584
rect 2032 1576 2152 1586
rect 2032 1568 2154 1576
rect 2182 1568 2278 1598
rect 2032 1562 2122 1568
rect 2094 1558 2122 1562
rect 2060 1552 2136 1558
rect 2056 1542 2136 1552
rect 2140 1542 2154 1568
rect 2056 1524 2154 1542
rect 2196 1524 2228 1568
rect 2230 1524 2278 1568
rect 2056 1518 2278 1524
rect 2060 1512 2278 1518
rect 2070 1508 2278 1512
rect 2074 1502 2278 1508
rect 2028 1498 2062 1502
rect 2028 1471 2074 1498
rect 2094 1493 2278 1502
rect 2106 1489 2140 1493
rect 2152 1492 2178 1493
rect 2152 1480 2162 1492
rect 2194 1489 2228 1493
rect 2116 1471 2164 1480
rect 2230 1474 2278 1493
rect 2028 1449 2062 1471
rect 2104 1461 2164 1471
rect 2216 1470 2278 1474
rect 2074 1449 2076 1460
rect 2028 1344 2076 1449
rect 2104 1381 2176 1461
rect 2178 1412 2200 1446
rect 2182 1406 2196 1412
rect 2104 1344 2164 1381
rect 2204 1344 2278 1470
rect 2283 1576 4950 1601
rect 5035 1594 5069 1604
rect 5088 1594 5555 1604
rect 5623 1598 5638 1610
rect 5739 1598 5769 1610
rect 2283 1559 4984 1576
rect 5035 1570 5555 1594
rect 5034 1562 5555 1570
rect 5557 1576 5619 1598
rect 5623 1589 5681 1598
rect 5623 1576 5682 1589
rect 5557 1568 5683 1576
rect 5711 1568 5769 1598
rect 5575 1562 5683 1568
rect 2283 1557 4274 1559
rect 2283 1344 2342 1557
rect 1545 1327 2176 1344
rect 2204 1336 2342 1344
rect 1545 1247 1593 1327
rect 1624 1247 1658 1327
rect 1670 1287 1771 1327
rect 1774 1287 1804 1327
rect 1687 1263 1692 1287
rect 1663 1247 1664 1260
rect 1691 1257 1692 1260
rect 1700 1253 1804 1287
rect 1818 1260 1826 1327
rect 1846 1306 1854 1327
rect 1861 1306 1909 1327
rect 1828 1272 1909 1306
rect 1914 1314 1974 1327
rect 1992 1320 2176 1327
rect 2196 1320 2342 1336
rect 1700 1247 1758 1253
rect 1774 1247 1804 1253
rect 1846 1247 1854 1272
rect 1861 1247 1912 1272
rect 1914 1247 1962 1314
rect 1992 1310 2342 1320
rect 2361 1499 2395 1557
rect 2463 1515 2478 1530
rect 2463 1505 2491 1515
rect 2509 1505 2523 1523
rect 2548 1518 2563 1552
rect 2565 1539 2597 1557
rect 2598 1548 4274 1557
rect 4280 1548 4984 1559
rect 2598 1539 4984 1548
rect 2463 1499 2523 1505
rect 2361 1470 2438 1499
rect 2361 1458 2395 1470
rect 2410 1465 2438 1470
rect 2441 1469 2523 1499
rect 2565 1474 4984 1539
rect 2565 1472 4240 1474
rect 4257 1472 4984 1474
rect 2441 1465 2525 1469
rect 2405 1458 2438 1465
rect 2361 1449 2438 1458
rect 2439 1455 2525 1465
rect 2443 1449 2460 1455
rect 2361 1421 2432 1449
rect 2468 1440 2514 1455
rect 2521 1440 2525 1455
rect 2565 1462 4257 1472
rect 4284 1470 4984 1472
rect 5035 1542 5069 1562
rect 5088 1542 5555 1562
rect 5623 1548 5683 1562
rect 5035 1534 5555 1542
rect 5603 1536 5683 1548
rect 4284 1466 4999 1470
rect 4297 1462 4999 1466
rect 2565 1460 4240 1462
rect 2468 1427 2526 1440
rect 2565 1436 4274 1460
rect 2590 1427 4274 1436
rect 2361 1406 2426 1421
rect 2468 1418 2533 1427
rect 2438 1407 2443 1418
rect 2473 1408 2533 1418
rect 2539 1414 4274 1427
rect 4280 1455 4999 1462
rect 5035 1455 5069 1534
rect 2539 1408 4257 1414
rect 2361 1396 2431 1406
rect 2438 1396 2445 1407
rect 2016 1291 2076 1310
rect 2104 1291 2176 1310
rect 2028 1287 2176 1291
rect 2204 1290 2278 1310
rect 2030 1281 2176 1287
rect 2216 1286 2278 1290
rect 2042 1278 2076 1281
rect 2130 1278 2164 1281
rect 2042 1277 2164 1278
rect 2074 1268 2140 1277
rect 2074 1266 2154 1268
rect 2230 1266 2278 1286
rect 2283 1286 2338 1310
rect 2361 1302 2445 1396
rect 2361 1291 2395 1302
rect 2397 1291 2445 1302
rect 2446 1291 2451 1408
rect 2474 1291 2479 1408
rect 2480 1406 4257 1408
rect 2480 1399 2545 1406
rect 2590 1402 4257 1406
rect 4280 1402 4987 1455
rect 2480 1393 2565 1399
rect 2480 1378 2569 1393
rect 2480 1328 2545 1378
rect 2553 1359 2569 1378
rect 2590 1380 4987 1402
rect 2590 1374 4274 1380
rect 4292 1377 4987 1380
rect 4297 1374 4987 1377
rect 2590 1360 4987 1374
rect 5018 1414 5069 1455
rect 5088 1426 5555 1534
rect 5599 1524 5683 1536
rect 5739 1524 5769 1568
rect 5599 1508 5769 1524
rect 5603 1502 5680 1508
rect 5084 1425 5555 1426
rect 5076 1414 5555 1425
rect 5018 1360 5555 1414
rect 2590 1344 5555 1360
rect 5557 1498 5591 1502
rect 5557 1477 5603 1498
rect 5623 1493 5680 1502
rect 5681 1493 5769 1508
rect 5557 1474 5597 1477
rect 5557 1449 5591 1474
rect 5602 1461 5603 1477
rect 5621 1489 5669 1493
rect 5681 1492 5707 1493
rect 5621 1480 5649 1489
rect 5681 1480 5691 1492
rect 5723 1489 5757 1493
rect 5621 1462 5693 1480
rect 5773 1474 5807 1610
rect 5837 1591 5871 1616
rect 5890 1591 5924 1616
rect 6004 1591 6038 1608
rect 6092 1591 6126 1608
rect 6159 1591 7769 1616
rect 5745 1470 5807 1474
rect 5645 1461 5693 1462
rect 5557 1344 5605 1449
rect 5645 1446 5705 1461
rect 5733 1455 5807 1470
rect 5647 1344 5649 1446
rect 5663 1396 5705 1446
rect 5707 1412 5729 1446
rect 5711 1406 5725 1412
rect 5690 1381 5705 1396
rect 5733 1378 5763 1455
rect 5659 1344 5693 1378
rect 5733 1344 5759 1378
rect 5773 1344 5807 1455
rect 5826 1582 7769 1591
rect 5826 1557 6138 1582
rect 6159 1574 7769 1582
rect 6141 1557 7769 1574
rect 7773 1615 7823 1684
rect 7873 1676 7919 1684
rect 7860 1658 7861 1663
rect 7873 1658 7933 1676
rect 7773 1565 7831 1615
rect 7849 1608 7853 1642
rect 7860 1616 7933 1658
rect 7861 1599 7919 1616
rect 7927 1608 7941 1616
rect 7925 1599 7941 1608
rect 7861 1582 7943 1599
rect 7861 1576 7939 1582
rect 7861 1565 7919 1576
rect 7773 1563 7855 1565
rect 7861 1563 7943 1565
rect 7785 1561 7819 1563
rect 7821 1561 7855 1563
rect 7867 1561 7907 1563
rect 7909 1561 7943 1563
rect 7785 1559 7867 1561
rect 7873 1559 7955 1561
rect 5826 1344 5871 1557
rect 2590 1343 5727 1344
rect 2480 1302 2533 1328
rect 2485 1291 2533 1302
rect 2599 1327 5727 1343
rect 2599 1307 5333 1327
rect 5404 1307 5438 1327
rect 5457 1314 5503 1327
rect 5457 1307 5491 1314
rect 5521 1310 5727 1327
rect 5733 1326 5871 1344
rect 5890 1458 5924 1557
rect 6004 1523 6051 1536
rect 5944 1520 5998 1523
rect 6004 1520 6052 1523
rect 5944 1500 6052 1520
rect 6077 1518 6092 1552
rect 6108 1534 6138 1557
rect 5992 1495 6052 1500
rect 5972 1489 6052 1495
rect 5934 1470 5955 1474
rect 5934 1458 5961 1470
rect 5890 1421 5961 1458
rect 5968 1469 6052 1489
rect 6095 1487 6138 1534
rect 6142 1487 7769 1557
rect 7809 1550 7867 1559
rect 7897 1551 7955 1559
rect 7897 1550 7949 1551
rect 7795 1548 7949 1550
rect 7795 1535 7943 1548
rect 7795 1516 7897 1535
rect 6095 1484 7769 1487
rect 5968 1455 6054 1469
rect 6095 1468 6138 1484
rect 5972 1449 5989 1455
rect 5997 1440 6043 1455
rect 6050 1453 6054 1455
rect 6108 1453 6138 1468
rect 6142 1453 7769 1484
rect 6050 1440 7769 1453
rect 5997 1431 6080 1440
rect 6119 1431 7769 1440
rect 5890 1396 5955 1421
rect 5997 1419 7769 1431
rect 5997 1408 6140 1419
rect 5967 1396 5974 1407
rect 5890 1326 5974 1396
rect 5975 1326 5980 1408
rect 6003 1326 6008 1408
rect 6009 1406 6140 1408
rect 6009 1399 6085 1406
rect 6009 1393 6094 1399
rect 6009 1385 6098 1393
rect 6009 1359 6096 1385
rect 6009 1357 6085 1359
rect 6009 1326 6096 1357
rect 6119 1343 6140 1406
rect 6142 1414 7769 1419
rect 7809 1482 7897 1516
rect 7903 1523 7943 1535
rect 7953 1535 7971 1539
rect 7953 1523 7983 1535
rect 7809 1414 7889 1482
rect 7903 1414 7983 1523
rect 7987 1414 8021 1684
rect 6142 1380 7983 1414
rect 7989 1380 8021 1414
rect 8023 1622 8075 1684
rect 8023 1619 8085 1622
rect 8445 1619 8480 1637
rect 5559 1307 5617 1310
rect 5647 1307 5717 1310
rect 2599 1292 5717 1307
rect 5733 1292 6096 1326
rect 2599 1291 4199 1292
rect 2283 1266 2331 1286
rect 1978 1247 2331 1266
rect 2361 1266 4199 1291
rect 2361 1257 4195 1266
rect 2397 1250 2445 1257
rect 2485 1250 2545 1257
rect 2411 1247 2445 1250
rect 2487 1247 2545 1250
rect 1545 1243 2331 1247
rect 1545 1232 2027 1243
rect 2045 1232 2331 1243
rect 2397 1238 2445 1247
rect 2485 1238 2545 1247
rect 2397 1234 2545 1238
rect 538 1192 624 1198
rect 552 1182 624 1192
rect 56 1144 472 1174
rect 568 1164 580 1174
rect 610 1172 624 1182
rect 626 1172 674 1198
rect 690 1178 898 1202
rect 1154 1198 1220 1204
rect 1545 1194 2012 1232
rect 2056 1216 2058 1232
rect 2072 1222 2120 1232
rect 2072 1216 2136 1222
rect 2230 1216 2278 1232
rect 2056 1204 2218 1216
rect 2230 1204 2280 1216
rect 1536 1189 2012 1194
rect 754 1174 776 1178
rect 777 1174 788 1178
rect 612 1164 624 1172
rect 16 1102 30 1144
rect 56 1110 538 1144
rect 568 1140 630 1164
rect 640 1162 674 1172
rect 690 1150 926 1174
rect 1126 1170 1248 1174
rect 1524 1160 2012 1189
rect 2046 1194 2218 1204
rect 2244 1200 2280 1204
rect 2244 1194 2278 1200
rect 2046 1174 2062 1194
rect 2070 1186 2218 1194
rect 2070 1184 2136 1186
rect 2188 1174 2218 1186
rect 2230 1174 2241 1185
rect 2249 1174 2278 1194
rect 2046 1166 2160 1174
rect 580 1138 630 1140
rect 582 1134 630 1138
rect 582 1122 598 1134
rect 602 1130 630 1134
rect 754 1141 788 1150
rect 870 1144 926 1150
rect 1176 1144 2012 1160
rect 1176 1141 1180 1144
rect 548 1114 598 1122
rect 56 1074 472 1110
rect 548 1102 624 1114
rect 754 1102 1193 1141
rect 1374 1137 1404 1144
rect 1446 1137 1476 1144
rect 1363 1126 1415 1137
rect 1435 1126 1487 1137
rect 1502 1126 1526 1144
rect 1492 1114 1526 1126
rect 1536 1114 1560 1144
rect 1199 1102 1210 1113
rect 480 1074 536 1102
rect 548 1083 598 1102
rect 640 1083 674 1094
rect 540 1074 598 1083
rect 628 1074 686 1083
rect 56 1060 686 1074
rect 754 1072 1210 1102
rect 1492 1107 1560 1114
rect 1573 1142 2012 1144
rect 2188 1142 2218 1144
rect 2230 1142 2278 1174
rect 1573 1133 2241 1142
rect 1573 1131 2229 1133
rect 1573 1122 2186 1131
rect 2188 1122 2218 1131
rect 1573 1121 2218 1122
rect 1573 1114 2248 1121
rect 2249 1114 2278 1142
rect 1573 1108 2278 1114
rect 1573 1107 2012 1108
rect 1492 1102 2012 1107
rect 2024 1102 2278 1108
rect 1492 1098 2278 1102
rect 754 1064 1193 1072
rect 1199 1064 1210 1072
rect 754 1060 1210 1064
rect 1300 1060 1402 1092
rect 1492 1088 2012 1098
rect 1492 1083 2080 1088
rect 2088 1083 2138 1098
rect 1492 1072 2138 1083
rect 2168 1083 2218 1098
rect 2283 1089 2331 1232
rect 2399 1228 2545 1234
rect 2599 1234 4195 1257
rect 4206 1234 4240 1292
rect 4314 1287 5716 1292
rect 5733 1290 5770 1292
rect 4308 1250 5716 1287
rect 5745 1286 5750 1290
rect 2599 1232 4240 1234
rect 4270 1232 4274 1234
rect 4308 1232 5699 1250
rect 2411 1225 2445 1228
rect 2499 1225 2533 1228
rect 2401 1224 2533 1225
rect 2401 1216 2426 1224
rect 2398 1213 2426 1216
rect 2443 1215 2509 1224
rect 2443 1213 2523 1215
rect 2544 1213 2567 1216
rect 2599 1213 4241 1232
rect 4259 1230 5699 1232
rect 4259 1221 5716 1230
rect 2347 1208 4241 1213
rect 4262 1209 4492 1221
rect 4259 1208 4492 1209
rect 4511 1208 5716 1221
rect 2347 1198 5716 1208
rect 2347 1196 4187 1198
rect 4206 1196 4240 1198
rect 2347 1181 4240 1196
rect 4284 1190 4300 1191
rect 4308 1190 4368 1198
rect 4308 1181 4366 1190
rect 4396 1181 4492 1198
rect 2347 1179 4492 1181
rect 2347 1089 2381 1179
rect 2401 1174 2489 1179
rect 2599 1178 4492 1179
rect 2599 1174 4240 1178
rect 4308 1175 4366 1178
rect 4396 1175 4492 1178
rect 2441 1169 2489 1174
rect 2580 1169 4240 1174
rect 2441 1162 4240 1169
rect 2441 1158 4187 1162
rect 2398 1154 4187 1158
rect 4206 1154 4240 1162
rect 4260 1165 4398 1175
rect 4408 1171 4442 1175
rect 4260 1162 4412 1165
rect 4260 1157 4432 1162
rect 4242 1154 4432 1157
rect 4444 1154 4492 1175
rect 4511 1154 5716 1198
rect 5773 1194 5807 1292
rect 5826 1286 5867 1292
rect 5890 1291 5924 1292
rect 5940 1291 5974 1292
rect 5975 1291 5980 1292
rect 5998 1291 6096 1292
rect 6142 1326 7769 1380
rect 7831 1350 7849 1368
rect 7867 1360 7895 1380
rect 7865 1350 7895 1360
rect 7831 1334 7895 1350
rect 7899 1334 7971 1380
rect 7849 1326 7971 1334
rect 6142 1294 7983 1326
rect 6142 1291 7724 1294
rect 5890 1290 7724 1291
rect 5826 1240 5860 1286
rect 5890 1282 5914 1290
rect 5879 1262 5914 1282
rect 5928 1268 7724 1290
rect 5928 1262 7058 1268
rect 5890 1257 7058 1262
rect 5940 1240 5986 1257
rect 5826 1224 5890 1240
rect 5952 1233 5986 1240
rect 5928 1228 5986 1233
rect 5998 1240 6096 1257
rect 6142 1244 7058 1257
rect 7097 1262 7141 1268
rect 7157 1262 7183 1268
rect 7097 1250 7123 1262
rect 7155 1250 7203 1262
rect 7139 1244 7203 1250
rect 6142 1240 7065 1244
rect 7135 1240 7203 1244
rect 5998 1228 6032 1240
rect 6045 1228 6085 1240
rect 5964 1224 5974 1228
rect 5790 1156 5807 1194
rect 5824 1218 5890 1224
rect 5998 1219 6016 1228
rect 6017 1219 6032 1224
rect 5824 1190 5860 1218
rect 2398 1144 2597 1154
rect 2425 1141 2505 1144
rect 2439 1131 2505 1141
rect 2456 1100 2490 1123
rect 2467 1098 2490 1100
rect 2456 1089 2490 1098
rect 2505 1098 2528 1111
rect 2590 1102 2597 1144
rect 2599 1153 4240 1154
rect 4260 1153 5716 1154
rect 2599 1146 5716 1153
rect 5792 1147 5807 1156
rect 2599 1145 4823 1146
rect 2599 1137 4609 1145
rect 2599 1128 4435 1137
rect 4444 1128 4609 1137
rect 2505 1089 2539 1098
rect 2599 1089 4199 1128
rect 2283 1088 4199 1089
rect 4206 1094 4492 1128
rect 4511 1109 4609 1128
rect 4677 1125 4723 1145
rect 4880 1132 5716 1146
rect 5798 1143 5807 1147
rect 5826 1171 5860 1190
rect 5897 1188 5932 1218
rect 5998 1215 6032 1219
rect 6051 1216 6085 1228
rect 6051 1215 6096 1216
rect 5897 1174 5927 1188
rect 5897 1171 5914 1174
rect 5944 1171 5955 1215
rect 5998 1200 6096 1215
rect 5826 1143 5864 1171
rect 5885 1166 5955 1171
rect 5884 1143 5894 1147
rect 5897 1143 5914 1166
rect 5968 1158 5969 1188
rect 5998 1187 6085 1200
rect 5972 1181 6085 1187
rect 5972 1158 5984 1181
rect 5998 1158 6085 1181
rect 5968 1147 6085 1158
rect 4677 1113 4724 1125
rect 4880 1121 5758 1132
rect 5784 1128 5864 1143
rect 5882 1131 5930 1143
rect 5968 1134 6034 1147
rect 6051 1134 6085 1147
rect 5968 1131 6085 1134
rect 4206 1088 4240 1094
rect 2226 1083 2230 1088
rect 2168 1072 2230 1083
rect 1492 1066 2134 1072
rect 1492 1060 1526 1066
rect 1536 1062 2134 1066
rect 1545 1060 2134 1062
rect 2180 1060 2230 1072
rect 2264 1072 4199 1088
rect 2264 1061 2555 1072
rect 2590 1064 4199 1072
rect 4208 1064 4240 1088
rect 2264 1060 2551 1061
rect 2590 1060 4240 1064
rect 56 1052 708 1060
rect 56 1042 714 1052
rect 721 1049 4240 1060
rect 732 1046 4240 1049
rect 732 1042 4226 1046
rect 4230 1042 4240 1046
rect 4242 1086 4290 1094
rect 4242 1070 4324 1086
rect 4330 1084 4413 1094
rect 4444 1084 4492 1094
rect 4522 1092 4526 1109
rect 4539 1102 4609 1109
rect 4537 1092 4609 1102
rect 4522 1088 4609 1092
rect 4679 1109 4723 1113
rect 4679 1091 4709 1109
rect 4735 1091 4751 1113
rect 4537 1084 4609 1088
rect 4242 1042 4296 1070
rect 4330 1068 4442 1084
rect 4318 1058 4442 1068
rect 4310 1054 4442 1058
rect 4444 1054 4609 1084
rect 4310 1052 4390 1054
rect 56 1037 728 1042
rect 732 1037 4296 1042
rect 56 1026 4296 1037
rect 4306 1026 4390 1052
rect 4444 1032 4514 1054
rect 4537 1040 4609 1054
rect 4621 1040 4643 1068
rect 4537 1035 4643 1040
rect 4537 1034 4621 1035
rect 4537 1032 4609 1034
rect 4444 1026 4609 1032
rect 56 972 486 1026
rect 58 888 486 972
rect 492 1003 716 1026
rect 717 1022 1210 1026
rect 1492 1022 1526 1026
rect 717 1003 1278 1022
rect 492 988 1278 1003
rect 492 958 728 988
rect 754 977 1278 988
rect 1424 982 1526 1022
rect 1330 977 1364 982
rect 1418 977 1526 982
rect 754 976 1364 977
rect 1366 976 1526 977
rect 754 972 1526 976
rect 754 963 1336 972
rect 1350 963 1526 972
rect 754 962 1324 963
rect 1350 962 1419 963
rect 754 958 1310 962
rect 492 954 1310 958
rect 1350 954 1412 962
rect 1424 954 1526 963
rect 1545 1020 2452 1026
rect 1545 956 2012 1020
rect 2046 1008 2061 1020
rect 2080 1008 2226 1020
rect 2230 1008 2268 1020
rect 2288 1008 2390 1020
rect 2046 986 2280 1008
rect 2294 1001 2390 1008
rect 2410 1001 2444 1020
rect 2449 1001 2456 1020
rect 2461 1018 2478 1026
rect 2461 1001 2495 1018
rect 2549 1001 2583 1018
rect 2590 1016 2595 1026
rect 2590 1001 2599 1016
rect 2616 1001 4609 1026
rect 4717 1025 4751 1091
rect 4880 1109 5716 1121
rect 5717 1109 5747 1121
rect 4880 1098 5758 1109
rect 5784 1098 5807 1128
rect 4880 1088 5716 1098
rect 4880 1084 5784 1088
rect 4866 1074 5784 1084
rect 5809 1079 5864 1128
rect 5884 1128 5930 1131
rect 5884 1079 5894 1128
rect 5897 1117 5927 1128
rect 5897 1088 5930 1117
rect 5998 1116 6085 1131
rect 5969 1113 6085 1116
rect 5998 1088 6085 1113
rect 5897 1079 6085 1088
rect 6142 1132 7085 1240
rect 7117 1234 7203 1240
rect 7124 1225 7181 1234
rect 7139 1184 7181 1225
rect 7189 1200 7203 1234
rect 7166 1169 7181 1184
rect 7135 1132 7169 1166
rect 7249 1132 7283 1268
rect 6142 1124 7283 1132
rect 6142 1079 6149 1124
rect 4866 1062 5805 1074
rect 4866 1042 5561 1062
rect 492 943 1210 954
rect 1242 944 1248 954
rect 1262 951 1424 954
rect 1430 951 1526 954
rect 492 903 716 943
rect 492 888 540 903
rect 552 899 574 903
rect 580 890 628 903
rect 640 899 662 903
rect 668 894 716 903
rect 58 882 540 888
rect 562 882 628 890
rect 630 882 716 894
rect 58 874 716 882
rect 728 942 1210 943
rect 1262 942 1526 951
rect 728 894 1244 942
rect 1278 936 1526 942
rect 1278 906 1446 936
rect 1492 914 1526 936
rect 1532 914 2012 956
rect 2038 978 2280 986
rect 2283 993 4609 1001
rect 4866 1022 5507 1042
rect 4866 1008 5347 1022
rect 4866 993 5397 1008
rect 5415 1007 5470 1015
rect 5473 1014 5497 1022
rect 2283 992 4592 993
rect 2038 952 2226 978
rect 2230 972 2268 978
rect 2283 975 4312 992
rect 4324 982 4400 992
rect 4444 988 4592 992
rect 2046 934 2226 952
rect 2228 934 2274 972
rect 2283 969 4260 975
rect 4290 973 4312 975
rect 4288 971 4312 973
rect 4323 973 4424 982
rect 4440 973 4592 988
rect 2283 967 4279 969
rect 2283 957 2390 967
rect 2283 948 2398 957
rect 2280 942 2398 948
rect 2280 934 2381 942
rect 2382 934 2398 942
rect 2410 937 2415 967
rect 2423 946 2482 967
rect 2549 963 4279 967
rect 4288 963 4318 971
rect 4323 968 4592 973
rect 4629 980 4787 993
rect 4857 984 5397 993
rect 5431 984 5467 1003
rect 5473 985 5501 1014
rect 5509 1007 5561 1042
rect 5595 1020 5621 1024
rect 5575 1007 5621 1020
rect 4857 980 5294 984
rect 5313 980 5347 984
rect 4629 976 4813 980
rect 4629 968 4829 976
rect 4857 973 5369 980
rect 5481 979 5501 985
rect 4323 963 4829 968
rect 2549 956 4829 963
rect 2549 952 4400 956
rect 2544 948 4400 952
rect 4406 954 4829 956
rect 4866 956 5369 973
rect 5459 969 5467 975
rect 5529 974 5559 1007
rect 5581 979 5583 1007
rect 5471 969 5559 974
rect 4866 954 5294 956
rect 4406 948 5294 954
rect 2423 944 2508 946
rect 2423 942 2444 944
rect 2427 937 2444 942
rect 2449 937 2456 944
rect 2403 934 2456 937
rect 2046 930 2456 934
rect 2461 933 2508 944
rect 2532 942 4400 948
rect 4410 945 4428 948
rect 4440 945 5294 948
rect 4406 942 5294 945
rect 2532 939 5294 942
rect 2461 930 2509 933
rect 1492 908 2012 914
rect 2056 918 2226 930
rect 2014 908 2048 912
rect 2056 908 2137 918
rect 1492 906 2137 908
rect 728 884 1268 894
rect 728 880 1244 884
rect 1248 880 1268 884
rect 1278 880 1526 906
rect 728 876 1456 880
rect 58 863 714 874
rect 728 865 1210 876
rect 1222 868 1430 876
rect 1431 868 1456 876
rect 1222 865 1456 868
rect 728 864 1444 865
rect 728 863 1210 864
rect 58 862 1210 863
rect 58 758 472 862
rect 480 836 526 862
rect 562 858 628 862
rect 562 856 626 858
rect 630 856 702 862
rect 568 836 702 856
rect 480 804 506 836
rect 580 822 680 836
rect 580 816 642 822
rect 580 806 626 816
rect 662 806 680 822
rect 620 804 680 806
rect 699 804 714 819
rect 480 788 538 804
rect 568 788 714 804
rect 480 784 714 788
rect 754 784 1210 862
rect 480 774 1210 784
rect 1222 796 1280 864
rect 1284 809 1362 864
rect 1366 838 1368 864
rect 1372 838 1444 864
rect 1284 797 1316 809
rect 1322 797 1362 809
rect 1368 809 1444 838
rect 1368 797 1404 809
rect 1290 796 1302 797
rect 1322 796 1366 797
rect 1368 796 1398 797
rect 1222 790 1316 796
rect 1322 790 1404 796
rect 1410 790 1444 809
rect 1446 790 1456 865
rect 1492 836 1526 880
rect 1536 903 2137 906
rect 2138 903 2226 918
rect 2230 926 2268 930
rect 1536 899 2126 903
rect 2138 902 2164 903
rect 1536 890 2106 899
rect 2138 890 2148 902
rect 2180 899 2214 903
rect 1536 887 2150 890
rect 1536 871 2054 887
rect 2058 872 2150 887
rect 2230 884 2264 926
rect 2202 880 2264 884
rect 2280 882 2328 930
rect 2058 871 2092 872
rect 1536 862 2048 871
rect 2082 868 2092 871
rect 2102 871 2150 872
rect 1536 836 2074 862
rect 2102 856 2162 871
rect 2190 865 2264 880
rect 2278 865 2328 882
rect 2190 862 2220 865
rect 2230 862 2264 865
rect 2280 862 2328 865
rect 1492 832 2074 836
rect 1492 824 2012 832
rect 1222 774 1456 790
rect 1510 798 2012 824
rect 1510 782 1526 798
rect 1492 774 1526 782
rect 480 769 1526 774
rect 480 764 1280 769
rect 492 760 1280 764
rect 492 758 1268 760
rect 58 748 1268 758
rect 1300 750 1526 769
rect 1318 748 1526 750
rect 1545 790 2012 798
rect 2014 790 2062 832
rect 2082 796 2092 834
rect 2104 832 2162 856
rect 2164 832 2186 856
rect 2104 790 2106 832
rect 2110 806 2186 832
rect 2190 832 2264 862
rect 2278 832 2328 862
rect 2110 796 2120 806
rect 2147 796 2162 806
rect 2190 796 2220 832
rect 2147 790 2220 796
rect 2230 790 2264 832
rect 2283 790 2328 832
rect 2347 868 2381 930
rect 2382 906 2398 930
rect 2410 926 2509 930
rect 2425 910 2440 915
rect 2444 910 2509 926
rect 2425 906 2444 910
rect 2424 905 2444 906
rect 2449 905 2509 910
rect 2424 904 2440 905
rect 2444 899 2509 905
rect 2391 868 2412 884
rect 2347 806 2412 868
rect 2425 879 2509 899
rect 2532 920 4578 939
rect 2532 908 4440 920
rect 4444 908 4578 920
rect 2532 897 4578 908
rect 4617 914 4651 918
rect 4617 905 4663 914
rect 2425 865 2511 879
rect 2427 822 2444 859
rect 2424 806 2431 817
rect 1545 782 2074 790
rect 2104 788 2264 790
rect 2104 782 2162 788
rect 2190 782 2264 788
rect 1545 760 2264 782
rect 2278 760 2336 790
rect 1545 754 2012 760
rect 2014 754 2062 760
rect 2074 754 2216 760
rect 2230 754 2264 760
rect 2283 754 2328 760
rect 1545 748 2328 754
rect 2347 748 2431 806
rect 2432 796 2444 822
rect 2454 850 2500 865
rect 2507 850 2511 865
rect 2532 876 4597 897
rect 2532 870 4462 876
rect 2532 859 2595 870
rect 2599 862 4462 870
rect 2599 859 4226 862
rect 2532 858 4226 859
rect 4236 858 4245 862
rect 2561 850 2595 858
rect 2599 850 4226 858
rect 2454 837 2543 850
rect 2565 846 2597 850
rect 2576 837 2597 846
rect 2454 830 2597 837
rect 2598 830 4226 850
rect 2454 818 2519 830
rect 2525 824 2597 830
rect 2599 824 4226 830
rect 4244 824 4245 858
rect 4266 842 4462 862
rect 4480 873 4597 876
rect 4641 891 4663 905
rect 4679 891 4685 897
rect 4725 894 4763 929
rect 4707 891 4763 894
rect 4641 873 4657 891
rect 4660 873 4663 891
rect 4480 854 4663 873
rect 4675 857 4685 891
rect 4691 873 4763 891
rect 4825 886 5294 939
rect 5313 952 5369 956
rect 5379 952 5381 956
rect 5313 901 5401 952
rect 5455 935 5559 969
rect 5455 919 5513 935
rect 5529 919 5559 935
rect 5595 926 5621 1007
rect 5629 1020 5805 1062
rect 5809 1045 6085 1079
rect 6108 1068 6149 1079
rect 6119 1056 6149 1068
rect 6153 1115 7283 1124
rect 6153 1113 6812 1115
rect 6153 1059 6806 1113
rect 6880 1059 6914 1115
rect 6933 1059 6967 1115
rect 6997 1113 7001 1115
rect 7013 1113 7283 1115
rect 6997 1098 7283 1113
rect 7013 1060 7093 1098
rect 7123 1090 7181 1098
rect 7105 1060 7181 1090
rect 7013 1059 7035 1060
rect 7105 1059 7135 1060
rect 6153 1056 6847 1059
rect 6108 1045 6847 1056
rect 5809 1020 5839 1045
rect 5851 1024 5864 1045
rect 5851 1020 5884 1024
rect 5897 1020 5927 1045
rect 5930 1020 6085 1045
rect 5629 942 5743 1020
rect 5784 1009 5930 1020
rect 5763 963 5930 1009
rect 5933 1011 5973 1020
rect 5933 1008 5952 1011
rect 5763 942 5797 963
rect 5817 959 5830 963
rect 5842 954 5885 963
rect 5905 959 5918 963
rect 5809 942 5912 954
rect 5629 931 5716 942
rect 5790 931 5797 942
rect 5800 931 5912 942
rect 5933 942 5956 1008
rect 5933 935 5952 942
rect 5939 931 5952 935
rect 5964 931 5973 1011
rect 5985 1016 6085 1020
rect 6153 1027 6847 1045
rect 6880 1035 7139 1059
rect 6153 1025 6880 1027
rect 6885 1025 7139 1035
rect 6153 1016 6823 1025
rect 5985 973 6823 1016
rect 6835 973 6857 997
rect 6880 981 6914 1025
rect 6933 981 6967 1025
rect 7079 1022 7139 1025
rect 7075 991 7141 1022
rect 7249 1006 7283 1098
rect 7302 1215 7724 1268
rect 7735 1292 7983 1294
rect 7989 1292 8021 1326
rect 7302 1045 7716 1215
rect 7302 1009 7705 1045
rect 7302 1006 7336 1009
rect 7404 1007 7462 1009
rect 7474 1007 7550 1009
rect 7474 1006 7504 1007
rect 7001 985 7021 991
rect 7079 988 7091 991
rect 7105 988 7141 991
rect 7001 981 7031 985
rect 7079 982 7139 988
rect 6880 973 6967 981
rect 5985 956 6857 973
rect 6900 963 6967 973
rect 6981 963 7031 981
rect 6900 957 7031 963
rect 5985 948 6229 956
rect 6253 948 6317 956
rect 5985 936 6086 948
rect 5985 931 6119 936
rect 5629 930 6119 931
rect 5498 904 5513 919
rect 5313 886 5413 901
rect 4825 876 5288 886
rect 4691 864 4813 873
rect 4691 857 4725 864
rect 4679 854 4685 857
rect 4480 851 4685 854
rect 4266 830 4457 842
rect 4480 836 4681 851
rect 4480 830 4578 836
rect 4266 826 4357 830
rect 4360 826 4578 830
rect 4266 824 4346 826
rect 4360 824 4440 826
rect 4444 824 4578 826
rect 4581 824 4681 836
rect 2525 818 4444 824
rect 2460 816 4444 818
rect 2460 809 2531 816
rect 2460 803 2551 809
rect 2460 796 2553 803
rect 2576 796 2597 816
rect 2599 812 4444 816
rect 2599 796 2606 812
rect 2616 796 4444 812
rect 2466 792 4444 796
rect 2466 790 4440 792
rect 4480 790 4578 824
rect 4641 823 4681 824
rect 4849 850 5288 876
rect 5313 852 5328 886
rect 5342 874 5413 886
rect 5467 874 5501 901
rect 5342 867 5401 874
rect 5629 867 5716 930
rect 5790 926 5797 930
rect 5839 922 5889 930
rect 5828 916 5889 922
rect 5824 892 5890 916
rect 5897 904 5927 930
rect 5939 926 5952 930
rect 5964 926 5973 930
rect 5828 882 5889 892
rect 5828 876 5886 882
rect 5345 862 5513 867
rect 5518 862 5570 867
rect 5646 862 5716 867
rect 5998 863 6032 930
rect 6051 870 6119 930
rect 6153 922 6317 948
rect 6153 917 6295 922
rect 6153 910 6299 917
rect 6161 879 6195 910
rect 6237 886 6241 910
rect 6249 897 6281 901
rect 6201 879 6225 886
rect 6161 870 6225 879
rect 6051 863 6086 870
rect 6193 869 6225 870
rect 6227 879 6243 886
rect 6249 879 6283 897
rect 6227 870 6283 879
rect 6227 869 6259 870
rect 6193 863 6207 869
rect 6237 863 6259 869
rect 6295 863 6363 910
rect 6367 863 6401 956
rect 4849 823 4936 850
rect 4617 820 4681 821
rect 2466 788 4578 790
rect 2466 782 2553 788
rect 2599 787 4578 788
rect 4623 819 4681 820
rect 4735 819 4769 821
rect 4623 798 4693 819
rect 4623 790 4650 798
rect 4651 796 4693 798
rect 4679 790 4693 796
rect 4735 790 4781 819
rect 4623 787 4693 790
rect 4723 787 4781 790
rect 4849 787 4947 823
rect 2466 774 2555 782
rect 2599 780 4947 787
rect 2599 774 4226 780
rect 4294 778 4352 780
rect 4382 778 4428 780
rect 4294 774 4428 778
rect 2466 760 2576 774
rect 2599 764 4428 774
rect 2466 753 2597 760
rect 2466 748 2576 753
rect 2599 748 4390 764
rect 4394 748 4428 764
rect 58 737 1456 748
rect 128 724 1456 737
rect 142 716 1456 724
rect 142 715 714 716
rect 768 715 1456 716
rect 1458 737 4428 748
rect 1458 729 1819 737
rect 1827 736 4428 737
rect 4480 774 4947 780
rect 5004 774 5005 850
rect 5010 848 5176 850
rect 5027 836 5176 848
rect 5027 825 5172 836
rect 5184 825 5187 850
rect 5199 825 5267 850
rect 5027 824 5267 825
rect 5027 798 5056 824
rect 5065 820 5099 824
rect 5031 796 5056 798
rect 5104 805 5144 824
rect 5031 786 5050 796
rect 5104 786 5150 805
rect 5153 796 5172 824
rect 5184 820 5187 824
rect 5218 801 5221 824
rect 5111 782 5150 786
rect 4480 770 5005 774
rect 5016 770 5050 782
rect 5104 774 5150 782
rect 5218 790 5229 801
rect 5241 790 5252 801
rect 5277 797 5288 850
rect 5345 834 5369 862
rect 5351 796 5369 834
rect 5379 796 5397 862
rect 5425 836 5455 862
rect 5518 856 5716 862
rect 5529 844 5716 856
rect 5518 833 5716 844
rect 5646 832 5716 833
rect 5646 802 5699 832
rect 5705 821 5716 832
rect 6003 802 6032 863
rect 5646 797 6032 802
rect 5218 774 5252 790
rect 5682 780 6032 797
rect 6037 858 6295 863
rect 6037 829 6086 858
rect 6119 832 6149 858
rect 6157 840 6259 858
rect 6157 829 6270 840
rect 6352 829 6401 863
rect 6037 774 6085 829
rect 6169 824 6223 829
rect 6237 824 6259 829
rect 6169 823 6259 824
rect 6169 813 6207 823
rect 6237 813 6259 823
rect 6169 796 6195 813
rect 6353 810 6401 829
rect 6420 810 6454 956
rect 6522 933 6857 956
rect 6528 903 6857 933
rect 6613 898 6690 903
rect 6713 898 6857 903
rect 6901 939 6914 957
rect 6931 939 7031 957
rect 7105 972 7139 982
rect 7105 963 7116 972
rect 7124 963 7139 972
rect 6901 920 7047 939
rect 7105 920 7139 963
rect 7158 972 7175 1006
rect 7249 982 7508 1006
rect 7192 972 7249 974
rect 7254 972 7508 982
rect 7158 920 7192 972
rect 7268 938 7283 972
rect 6901 910 7187 920
rect 6613 887 6668 898
rect 6736 887 6823 898
rect 6613 886 6823 887
rect 6837 886 6847 898
rect 6901 891 7192 910
rect 6903 889 6913 891
rect 6933 886 7192 891
rect 7266 886 7283 938
rect 7302 910 7336 972
rect 7448 969 7508 972
rect 7618 989 7705 1009
rect 7735 1026 7769 1292
rect 7849 1284 7895 1292
rect 7849 1258 7883 1284
rect 7931 1266 7983 1292
rect 7795 1232 7883 1258
rect 7937 1232 7983 1266
rect 7987 1232 8021 1292
rect 8023 1281 8121 1619
rect 8409 1604 8480 1619
rect 8409 1487 8479 1604
rect 8591 1536 8649 1542
rect 8591 1502 8603 1536
rect 8591 1496 8649 1502
rect 8222 1481 8280 1487
rect 8222 1447 8234 1481
rect 8222 1441 8280 1447
rect 8392 1413 8479 1487
rect 9895 1419 9930 1453
rect 8166 1397 8224 1411
rect 8166 1377 8190 1397
rect 8278 1377 8312 1411
rect 8178 1343 8324 1377
rect 8392 1360 8490 1413
rect 9896 1400 9930 1419
rect 8178 1319 8192 1343
rect 8023 1232 8138 1281
rect 8234 1247 8296 1281
rect 8262 1241 8296 1247
rect 8392 1241 8831 1360
rect 9211 1307 9246 1325
rect 9175 1292 9246 1307
rect 7791 1198 7983 1232
rect 7837 1190 7897 1198
rect 7837 1175 7894 1190
rect 7953 1175 7983 1198
rect 7835 1171 7883 1175
rect 7895 1174 7921 1175
rect 7835 1162 7861 1171
rect 7895 1162 7903 1174
rect 7953 1171 7971 1175
rect 7785 1143 7803 1147
rect 7835 1144 7907 1162
rect 7859 1143 7907 1144
rect 7773 1026 7823 1143
rect 7859 1128 7919 1143
rect 7877 1078 7919 1128
rect 7927 1094 7941 1128
rect 7904 1063 7919 1078
rect 7873 1026 7907 1060
rect 7987 1026 8021 1230
rect 8040 1109 8138 1232
rect 8218 1179 8252 1207
rect 8392 1179 8406 1241
rect 8206 1145 8352 1179
rect 8218 1109 8252 1145
rect 8051 1044 8138 1109
rect 8250 1075 8308 1081
rect 8250 1046 8262 1075
rect 8409 1056 8831 1241
rect 8842 1237 8877 1271
rect 8250 1044 8284 1046
rect 8051 1041 8284 1044
rect 8051 1035 8308 1041
rect 8051 1026 8282 1035
rect 7735 1007 7759 1026
rect 7773 1008 8021 1026
rect 8068 1008 8282 1026
rect 7773 1007 8282 1008
rect 7735 992 8282 1007
rect 7773 989 7831 992
rect 7861 989 7931 992
rect 7618 974 7931 989
rect 7987 974 8282 992
rect 7444 938 7510 969
rect 7448 935 7460 938
rect 7474 935 7510 938
rect 7448 929 7508 935
rect 7474 919 7508 929
rect 7474 910 7485 919
rect 7493 910 7508 919
rect 7302 904 7362 910
rect 7300 901 7336 904
rect 6522 870 6537 885
rect 6522 857 6580 870
rect 6656 857 6668 886
rect 6520 840 6580 857
rect 6530 820 6580 840
rect 6736 810 6823 886
rect 6979 885 7029 886
rect 6897 873 6913 885
rect 6933 873 6949 885
rect 6897 865 6949 873
rect 6979 865 7037 885
rect 6897 863 6913 865
rect 6933 861 6949 865
rect 6985 863 7037 865
rect 6989 861 7037 863
rect 6169 795 6283 796
rect 6353 790 6364 801
rect 6372 790 6401 810
rect 5104 770 5288 774
rect 5646 772 6085 774
rect 4480 760 5288 770
rect 4480 748 4578 760
rect 4595 753 5288 760
rect 4635 748 4681 753
rect 4735 748 4769 753
rect 4849 748 5288 753
rect 5632 761 6085 772
rect 6147 761 6195 782
rect 6229 761 6305 782
rect 6353 774 6401 790
rect 6406 802 6455 810
rect 6406 790 6502 802
rect 6551 799 6823 810
rect 6406 787 6513 790
rect 6562 788 6823 799
rect 6891 795 6931 802
rect 6997 795 7037 802
rect 6562 787 6722 788
rect 6406 776 6516 787
rect 6551 776 6722 787
rect 6753 782 6823 788
rect 6406 774 6454 776
rect 6353 761 6485 774
rect 6588 766 6722 774
rect 6736 770 6823 782
rect 5632 760 6485 761
rect 6562 760 6722 766
rect 5632 748 6071 760
rect 6147 748 6305 760
rect 6353 748 6485 760
rect 6588 748 6722 760
rect 6753 748 6823 770
rect 6947 757 6981 782
rect 1827 729 4440 736
rect 1458 728 4440 729
rect 1458 715 1948 728
rect 1972 725 4440 728
rect 1961 720 4440 725
rect 1961 715 2162 720
rect 2168 715 4440 720
rect 142 714 4440 715
rect 282 674 300 708
rect 304 702 362 714
rect 392 702 450 714
rect 480 702 538 714
rect 568 702 626 714
rect 656 702 714 714
rect 768 704 1210 714
rect 771 672 1210 704
rect 1222 702 1264 714
rect 1318 702 1368 714
rect 1222 700 1280 702
rect 1310 700 1432 702
rect 1234 696 1244 700
rect 192 656 392 672
rect 762 652 1210 672
rect 771 648 1210 652
rect 1492 648 1526 714
rect 771 631 1228 648
rect 1269 637 1321 648
rect 1357 643 1473 648
rect 1421 637 1473 643
rect 1176 630 1228 631
rect 1280 630 1310 637
rect 1432 630 1462 637
rect 1510 630 1526 648
rect 1545 630 1579 714
rect 1610 630 1613 714
rect 1663 713 1698 714
rect 1705 713 1790 714
rect 1663 708 1790 713
rect 1669 703 1744 708
rect 1669 697 1749 703
rect 1760 697 1790 708
rect 1687 663 1790 697
rect 1861 708 1948 714
rect 1861 698 1895 708
rect 1687 647 1753 663
rect 1760 647 1790 663
rect 1832 682 1854 688
rect 1861 682 1898 698
rect 1832 676 1898 682
rect 1832 672 1854 676
rect 1861 672 1898 676
rect 1914 672 1948 708
rect 2016 691 2017 714
rect 2104 706 2106 714
rect 2104 703 2116 706
rect 2104 691 2121 703
rect 2190 700 2216 714
rect 1832 668 1972 672
rect 1729 630 1744 647
rect 1176 614 1579 630
rect 1082 600 1208 608
rect 1510 600 1579 614
rect 1598 600 1656 630
rect 1686 600 1744 630
rect 1804 604 1826 660
rect 1832 632 1898 668
rect 1861 630 1895 632
rect 1914 630 1948 668
rect 1510 585 1525 600
rect 1545 595 1579 600
rect 1610 595 1613 600
rect 1729 595 1744 600
rect 1861 600 1948 630
rect 1861 595 1895 600
rect 1545 590 1872 595
rect 1880 590 1895 595
rect 1545 589 1895 590
rect 1545 561 1744 589
rect 1749 584 1895 589
rect 1760 572 1895 584
rect 1749 561 1895 572
rect 1914 590 1948 600
rect 58 532 86 536
rect 1914 527 1929 590
rect 1937 589 1948 590
rect 2032 576 2048 678
rect 2060 644 2118 650
rect 2060 610 2076 644
rect 2060 604 2118 610
rect 2230 600 2264 714
rect 2056 594 2122 596
rect 2230 589 2241 600
rect 1961 531 2131 542
rect 2163 531 2215 542
rect 1914 519 1928 527
rect 1972 524 2120 531
rect 2090 519 2120 524
rect 2174 519 2204 531
rect 1914 508 1939 519
rect 2079 508 2131 519
rect 2163 508 2215 519
rect 2249 508 2264 600
rect 2283 696 2324 714
rect 2347 712 2431 714
rect 2466 712 2519 714
rect 2347 701 2381 712
rect 2397 701 2431 712
rect 2432 701 2437 708
rect 2460 701 2465 708
rect 2485 701 2519 712
rect 2599 713 4440 714
rect 4446 713 4478 736
rect 2599 704 4478 713
rect 2599 702 4181 704
rect 4192 702 4478 704
rect 2599 701 4226 702
rect 2347 700 4226 701
rect 2283 652 2317 696
rect 2347 672 2371 700
rect 2385 678 4226 700
rect 4294 692 4352 702
rect 2385 672 3640 678
rect 3644 672 3704 678
rect 2347 667 3694 672
rect 2283 630 2298 652
rect 2313 641 2317 652
rect 2397 650 2443 667
rect 2409 645 2443 650
rect 2502 645 2525 654
rect 2599 652 3694 667
rect 2599 650 3586 652
rect 3592 650 3660 652
rect 2306 630 2317 641
rect 2385 638 2443 645
rect 2473 638 2531 645
rect 2599 644 3660 650
rect 2283 508 2317 630
rect 2599 635 3638 644
rect 2401 576 2412 625
rect 2530 610 2553 626
rect 2425 568 2426 598
rect 2429 591 2487 597
rect 2429 568 2441 591
rect 2425 541 2491 568
rect 2599 544 3586 635
rect 3596 594 3638 635
rect 3646 610 3660 644
rect 3623 579 3638 594
rect 2599 534 3002 544
rect 2426 523 2492 526
rect 72 504 86 508
rect 2283 498 2298 508
rect 282 244 300 480
rect 1964 472 2510 498
rect 2599 489 2606 534
rect 2565 478 2606 489
rect 310 272 328 452
rect 2247 430 2510 472
rect 2576 466 2606 478
rect 2616 504 3002 534
rect 2616 466 2686 504
rect 2798 498 2856 504
rect 2968 498 3002 504
rect 2565 455 2686 466
rect 2308 421 2342 430
rect 2396 421 2430 430
rect 2442 426 2510 430
rect 2616 436 2686 455
rect 2968 455 2982 498
rect 2987 455 3002 498
rect 2968 436 3002 455
rect 2616 426 2705 436
rect 2753 434 2881 436
rect 2442 425 2705 426
rect 2442 419 2694 425
rect 1598 394 1640 418
rect 2652 413 2694 419
rect 2750 416 2884 434
rect 2907 416 3002 436
rect 2652 412 2705 413
rect 2750 412 3002 416
rect 2652 408 3002 412
rect 3021 542 3550 544
rect 3592 542 3626 576
rect 3706 542 3740 678
rect 3021 525 3740 542
rect 3021 424 3055 525
rect 3123 523 3173 525
rect 3211 523 3269 525
rect 3128 501 3158 523
rect 3181 501 3200 523
rect 3216 501 3246 523
rect 3163 498 3200 501
rect 3082 476 3089 480
rect 3163 476 3238 498
rect 2652 402 3004 408
rect 1626 366 1640 390
rect 1802 380 1840 390
rect 288 206 300 244
rect 316 206 328 272
rect 1802 244 1826 380
rect 2784 368 2850 400
rect 2987 374 3004 402
rect 1830 352 1868 362
rect 1830 272 1854 352
rect 3021 349 3038 424
rect 3045 383 3055 424
rect 3070 383 3109 476
rect 3158 461 3251 476
rect 3163 451 3251 461
rect 3163 435 3216 451
rect 3258 417 3263 480
rect 3337 395 3371 525
rect 3337 391 3358 395
rect 3337 383 3371 391
rect 3070 349 3304 383
rect 3358 349 3371 383
rect 3170 292 3204 349
rect 3390 330 3424 525
rect 3454 508 3458 525
rect 3470 508 3740 525
rect 3470 442 3492 508
rect 3498 470 3550 508
rect 3536 432 3594 438
rect 3536 398 3548 432
rect 3573 398 3594 432
rect 3536 392 3594 398
rect 3601 364 3622 466
rect 3706 392 3740 508
rect 3390 301 3504 330
rect 3509 319 3561 330
rect 3520 307 3550 319
rect 3390 296 3457 301
rect 3509 296 3561 307
rect 3725 296 3740 392
rect 3759 672 4226 678
rect 4228 672 4352 692
rect 4382 672 4440 702
rect 3759 630 4181 672
rect 4192 630 4226 672
rect 4294 668 4340 672
rect 4252 642 4340 668
rect 4394 642 4440 672
rect 4444 642 4478 702
rect 4480 735 5288 748
rect 5648 746 6401 748
rect 5730 736 5956 746
rect 6003 736 6401 746
rect 5668 735 6401 736
rect 4480 727 6401 735
rect 4480 715 6071 727
rect 6085 715 6387 727
rect 6406 715 6485 748
rect 4480 714 6485 715
rect 6614 737 7008 748
rect 6614 725 6997 737
rect 6614 723 7008 725
rect 6614 714 7017 723
rect 7105 717 7139 886
rect 4480 691 4578 714
rect 4651 708 4793 714
rect 4679 691 4737 697
rect 4480 642 4595 691
rect 4675 685 4765 691
rect 4675 680 4769 685
rect 4691 672 4753 680
rect 4248 630 4440 642
rect 4444 630 4478 640
rect 4497 630 4595 642
rect 4675 651 4769 672
rect 4849 651 5288 714
rect 5632 702 5703 714
rect 5632 681 5702 702
rect 4675 641 4721 651
rect 3759 608 4595 630
rect 4671 613 4721 641
rect 3759 455 4173 608
rect 3759 419 4162 455
rect 3759 296 3793 419
rect 3905 379 3963 385
rect 3905 345 3917 379
rect 3905 339 3963 345
rect 1808 206 1826 244
rect 1836 206 1854 272
rect 3759 262 3774 296
rect 4092 243 4162 419
rect 4192 436 4226 608
rect 4294 600 4354 608
rect 4382 600 4440 608
rect 4294 585 4351 600
rect 4394 597 4440 600
rect 4410 585 4440 597
rect 4292 581 4340 585
rect 4352 584 4378 585
rect 4292 572 4318 581
rect 4352 572 4360 584
rect 4410 581 4428 585
rect 4242 553 4260 557
rect 4292 554 4364 572
rect 4316 553 4364 554
rect 4230 436 4280 553
rect 4316 538 4376 553
rect 4334 488 4376 538
rect 4384 504 4398 538
rect 4361 473 4376 488
rect 4330 436 4364 470
rect 4444 436 4478 608
rect 4497 519 4595 608
rect 4663 600 4721 613
rect 4751 650 4769 651
rect 4751 613 4801 650
rect 4849 630 4860 641
rect 4866 630 5288 651
rect 4751 600 4809 613
rect 4663 589 4709 600
rect 4794 589 4809 600
rect 4849 600 5288 630
rect 4849 589 4863 600
rect 4663 555 4809 589
rect 4675 519 4709 555
rect 4508 436 4595 519
rect 4707 485 4765 491
rect 4707 451 4719 485
rect 4866 466 5288 600
rect 5299 680 5702 681
rect 5299 647 5334 680
rect 4707 445 4765 451
rect 4192 402 4216 436
rect 4230 402 4478 436
rect 4274 326 4332 332
rect 4274 292 4286 326
rect 4274 286 4332 292
rect 4444 286 4478 402
rect 4525 402 4595 436
rect 4525 366 4578 402
rect 4896 349 4911 466
rect 4930 349 4964 466
rect 5076 432 5134 438
rect 5076 398 5088 432
rect 5076 392 5134 398
rect 4930 315 4945 349
rect 5265 296 5280 466
rect 5299 296 5333 647
rect 5615 630 5626 641
rect 5632 630 5702 680
rect 5399 600 5549 630
rect 5615 600 5702 630
rect 5615 589 5626 600
rect 5445 579 5503 585
rect 5445 545 5457 579
rect 5445 539 5503 545
rect 5445 379 5503 385
rect 5445 345 5457 379
rect 5445 339 5503 345
rect 5299 262 5314 296
rect 5632 243 5702 600
rect 5814 634 5872 640
rect 5814 600 5826 634
rect 5984 630 5995 641
rect 6003 630 6018 714
rect 5984 600 6018 630
rect 5814 594 5872 600
rect 5984 589 5995 600
rect 5814 326 5872 332
rect 5814 292 5826 326
rect 5814 286 5872 292
rect 4092 207 4145 243
rect 5632 207 5685 243
rect 6003 203 6018 600
rect 6037 203 6071 714
rect 6151 680 6185 684
rect 6239 680 6273 684
rect 6139 630 6154 645
rect 6270 630 6285 645
rect 6139 600 6197 630
rect 6227 600 6285 630
rect 6139 585 6154 600
rect 6270 585 6285 600
rect 6353 630 6364 641
rect 6372 630 6387 714
rect 6353 600 6387 630
rect 6353 589 6364 600
rect 6183 273 6241 279
rect 6183 256 6195 273
rect 6372 256 6387 600
rect 6406 674 6441 714
rect 6464 697 6516 708
rect 6537 697 6722 708
rect 6475 685 6505 697
rect 6548 685 6722 697
rect 6464 681 6516 685
rect 6537 681 6722 685
rect 6464 680 6722 681
rect 6464 674 6708 680
rect 6753 674 6823 714
rect 6406 256 6440 674
rect 6508 585 6520 627
rect 6753 621 6810 674
rect 7124 621 7139 717
rect 7158 621 7192 886
rect 7300 870 7366 901
rect 7302 867 7362 870
rect 7474 867 7508 910
rect 7527 919 7544 953
rect 7618 932 7930 974
rect 7618 929 7913 932
rect 7561 919 7618 921
rect 7623 919 7913 929
rect 7527 867 7561 919
rect 7635 912 7913 919
rect 7272 857 7556 867
rect 7272 836 7561 857
rect 7302 833 7561 836
rect 7302 808 7318 832
rect 7348 808 7406 832
rect 7304 704 7362 710
rect 7304 670 7316 704
rect 7304 664 7362 670
rect 7474 664 7508 833
rect 6753 585 6792 621
rect 7158 587 7173 621
rect 7493 568 7508 664
rect 7527 568 7561 833
rect 7635 744 7930 912
rect 7987 876 8021 974
rect 8068 912 8282 974
rect 8439 939 8454 1056
rect 8473 939 8507 1056
rect 8619 1022 8677 1028
rect 8619 988 8631 1022
rect 8619 982 8677 988
rect 8042 906 8282 912
rect 8002 825 8021 876
rect 8038 872 8059 906
rect 8068 903 8282 906
rect 8473 905 8488 939
rect 8808 938 8823 1056
rect 8842 938 8876 1237
rect 8988 1169 9046 1175
rect 8988 1135 9000 1169
rect 8988 1129 9046 1135
rect 8988 969 9046 975
rect 8988 940 9000 969
rect 8988 938 9022 940
rect 8598 935 9022 938
rect 8598 929 9046 935
rect 8598 901 9020 929
rect 8212 883 8246 901
rect 8473 886 9020 901
rect 8042 866 8100 872
rect 8212 847 8282 883
rect 8598 850 9020 886
rect 7998 780 8021 825
rect 8229 813 8300 847
rect 7673 651 7731 657
rect 7673 617 7685 651
rect 7673 611 7731 617
rect 7527 534 7542 568
rect 6722 505 6756 523
rect 7860 515 7930 744
rect 8042 598 8100 604
rect 8042 564 8054 598
rect 8042 558 8100 564
rect 6722 469 6792 505
rect 7860 479 7913 515
rect 8229 472 8299 813
rect 8411 745 8469 751
rect 8411 711 8423 745
rect 8411 705 8469 711
rect 8411 545 8469 551
rect 8411 511 8423 545
rect 8411 505 8469 511
rect 6739 435 6810 469
rect 7090 435 7125 469
rect 7896 462 8299 472
rect 6739 256 6809 435
rect 7091 416 7125 435
rect 6921 367 6979 373
rect 6921 333 6933 367
rect 6921 327 6979 333
rect 6116 203 6809 256
rect 5747 154 6809 203
rect 3573 -120 3586 136
rect 3601 -92 3614 108
rect 6001 101 6809 154
rect 6921 167 6979 173
rect 6921 133 6933 167
rect 6921 127 6979 133
rect 6370 84 6809 101
rect 6370 73 6792 84
rect 7110 73 7125 416
rect 6370 65 6809 73
rect 7091 65 7125 73
rect 6370 48 7125 65
rect 6775 31 7125 48
rect 7144 382 7179 416
rect 7459 382 7494 416
rect 7882 399 7917 417
rect 7144 72 7178 382
rect 7460 363 7494 382
rect 7846 384 7917 399
rect 8229 409 8286 462
rect 8598 409 8668 850
rect 8806 806 9020 850
rect 8780 800 9020 806
rect 8780 766 8792 800
rect 8806 797 9020 800
rect 9175 833 9245 1292
rect 9357 1224 9415 1230
rect 9357 1190 9369 1224
rect 9357 1184 9415 1190
rect 9357 916 9415 922
rect 9357 882 9369 916
rect 9357 876 9415 882
rect 9175 797 9228 833
rect 9175 795 9274 797
rect 9434 796 9465 814
rect 9546 796 9561 1326
rect 9580 796 9614 1380
rect 9726 1351 9784 1357
rect 9726 1317 9738 1351
rect 9726 1311 9784 1317
rect 9726 863 9784 869
rect 9726 834 9738 863
rect 9726 830 9760 834
rect 9722 829 9760 830
rect 9726 823 9784 829
rect 8950 777 8984 795
rect 9175 780 9407 795
rect 9468 780 9499 796
rect 9614 795 9722 796
rect 9175 777 9274 780
rect 9372 777 9407 780
rect 8780 760 8838 766
rect 8950 741 9020 777
rect 9175 762 9407 777
rect 9614 762 9688 795
rect 9175 744 9406 762
rect 8967 707 9038 741
rect 8780 492 8838 498
rect 8780 458 8792 492
rect 8780 452 8838 458
rect 7290 314 7348 320
rect 7290 280 7302 314
rect 7290 274 7348 280
rect 7290 114 7348 120
rect 7290 106 7302 114
rect 7286 80 7352 106
rect 7290 74 7348 80
rect 7144 66 7179 72
rect 7252 66 7386 72
rect 7144 38 7460 66
rect 6775 2 7125 19
rect 6739 -3 7125 2
rect 6739 -15 6810 -3
rect 6406 -68 6441 -34
rect 6037 -121 6072 -87
rect 288 -194 300 -156
rect 282 -430 300 -194
rect 316 -222 328 -156
rect 1808 -220 1826 -156
rect 1836 -220 1854 -156
rect 4128 -157 4163 -140
rect 5668 -157 5703 -140
rect 4092 -174 4163 -157
rect 5632 -174 5703 -157
rect 310 -402 328 -222
rect 3759 -227 3794 -193
rect 2606 -301 2664 -298
rect 1626 -340 1640 -316
rect 1598 -368 1640 -344
rect 2179 -354 2442 -301
rect 2518 -308 2664 -301
rect 2694 -308 2752 -298
rect 3170 -299 3204 -242
rect 3390 -251 3457 -246
rect 3390 -280 3504 -251
rect 3509 -257 3561 -246
rect 3520 -269 3550 -257
rect 3509 -280 3561 -269
rect 2784 -350 2850 -318
rect 2987 -352 3004 -324
rect 2032 -369 2442 -354
rect 2652 -363 2705 -352
rect 2750 -358 3004 -352
rect 2652 -369 2694 -363
rect 2032 -379 2247 -369
rect 2296 -379 2354 -369
rect 2384 -379 2510 -369
rect 2032 -380 2510 -379
rect 2616 -375 2694 -369
rect 2750 -366 3002 -358
rect 2308 -384 2342 -380
rect 2396 -384 2430 -380
rect 2616 -386 2705 -375
rect 2750 -384 2884 -366
rect 2938 -374 3002 -366
rect 2952 -375 2982 -374
rect 2941 -386 2982 -375
rect 2616 -405 2686 -386
rect 2283 -410 2464 -405
rect 2283 -418 2492 -410
rect 2565 -416 2686 -405
rect 2283 -439 2318 -418
rect 2354 -428 2384 -418
rect 2343 -432 2384 -428
rect 2426 -428 2492 -418
rect 2576 -428 2606 -416
rect 2426 -432 2503 -428
rect 2343 -439 2503 -432
rect 2565 -439 2606 -428
rect 1914 -469 1939 -458
rect 2079 -469 2131 -458
rect 2163 -469 2215 -458
rect 1914 -477 1928 -469
rect 2090 -474 2120 -469
rect 1545 -545 1744 -511
rect 1749 -522 1895 -511
rect 1760 -534 1895 -522
rect 1749 -540 1895 -534
rect 1749 -545 1801 -540
rect 1880 -545 1895 -540
rect 1176 -581 1228 -564
rect 1269 -571 1401 -564
rect 1269 -575 1321 -571
rect 1421 -575 1473 -564
rect 771 -596 1228 -581
rect 1280 -587 1310 -575
rect 1432 -587 1462 -575
rect 1269 -596 1321 -587
rect 1421 -593 1473 -587
rect 1357 -596 1473 -593
rect 1510 -596 1526 -564
rect 771 -598 1526 -596
rect 282 -648 300 -624
rect 114 -674 162 -648
rect 192 -674 304 -648
rect 316 -652 350 -640
rect 310 -668 350 -652
rect 316 -674 350 -668
rect 404 -670 438 -640
rect 492 -670 526 -640
rect 534 -648 580 -640
rect 614 -648 668 -640
rect 534 -664 668 -648
rect 692 -664 702 -640
rect 534 -670 702 -664
rect 771 -670 1210 -598
rect 1234 -650 1244 -646
rect 1300 -650 1356 -632
rect 1410 -650 1418 -646
rect 404 -674 714 -670
rect 768 -674 1210 -670
rect 128 -687 1210 -674
rect 58 -708 1210 -687
rect 58 -822 472 -708
rect 492 -724 506 -708
rect 699 -724 714 -709
rect 480 -754 538 -724
rect 568 -738 626 -724
rect 656 -725 714 -724
rect 630 -738 714 -725
rect 562 -754 714 -738
rect 492 -796 506 -754
rect 562 -756 580 -754
rect 620 -756 680 -754
rect 562 -766 626 -756
rect 630 -766 680 -756
rect 562 -772 680 -766
rect 699 -769 714 -754
rect 580 -796 680 -772
rect 492 -820 526 -796
rect 492 -822 506 -820
rect 518 -822 526 -820
rect 580 -806 702 -796
rect 580 -822 626 -806
rect 634 -812 642 -806
rect 662 -820 702 -806
rect 662 -822 680 -820
rect 58 -832 714 -822
rect 754 -832 1210 -708
rect 1222 -709 1264 -650
rect 1300 -662 1418 -650
rect 1300 -666 1444 -662
rect 1318 -700 1444 -666
rect 1222 -719 1268 -709
rect 1318 -716 1368 -700
rect 1376 -706 1380 -700
rect 1222 -830 1274 -719
rect 1290 -747 1302 -743
rect 1284 -748 1302 -747
rect 1322 -747 1366 -716
rect 1404 -734 1408 -700
rect 1378 -747 1390 -743
rect 1280 -759 1310 -748
rect 1322 -759 1362 -747
rect 1284 -818 1362 -759
rect 1284 -830 1324 -818
rect 58 -915 472 -832
rect 23 -1083 27 -915
rect 47 -926 472 -915
rect 56 -938 472 -926
rect 47 -949 472 -938
rect 35 -950 472 -949
rect 492 -834 506 -832
rect 518 -834 532 -832
rect 598 -834 626 -832
rect 662 -834 708 -832
rect 492 -858 532 -834
rect 552 -853 560 -849
rect 580 -853 626 -834
rect 640 -853 648 -849
rect 668 -853 708 -834
rect 492 -950 506 -858
rect 514 -860 532 -858
rect 514 -894 526 -860
rect 540 -893 708 -853
rect 714 -893 1210 -832
rect 1234 -834 1244 -830
rect 1256 -834 1268 -830
rect 514 -922 532 -894
rect 514 -950 526 -922
rect 540 -950 1210 -893
rect 1280 -912 1324 -830
rect 1344 -830 1362 -818
rect 1368 -759 1398 -747
rect 1410 -759 1444 -700
rect 1368 -818 1444 -759
rect 1344 -858 1356 -830
rect 1368 -841 1412 -818
rect 1368 -886 1424 -841
rect 1278 -913 1324 -912
rect 1378 -901 1424 -886
rect 1378 -913 1412 -901
rect 1278 -927 1336 -913
rect 1366 -927 1424 -913
rect 1336 -928 1352 -927
rect 35 -990 718 -950
rect 720 -976 742 -950
rect 754 -963 1210 -950
rect 1334 -963 1368 -942
rect 1492 -944 1526 -598
rect 1545 -687 1579 -545
rect 1610 -687 1613 -545
rect 1669 -592 1698 -579
rect 1737 -582 1744 -566
rect 1650 -597 1698 -592
rect 1729 -597 1744 -582
rect 1760 -592 1790 -555
rect 1804 -592 1826 -554
rect 1650 -610 1744 -597
rect 1749 -610 1826 -592
rect 1669 -613 1744 -610
rect 1760 -613 1790 -610
rect 1687 -620 1790 -613
rect 1832 -620 1854 -582
rect 1650 -638 1854 -620
rect 1861 -598 1895 -545
rect 1914 -540 1929 -477
rect 1972 -481 2120 -474
rect 2174 -481 2204 -469
rect 1961 -492 2131 -481
rect 2163 -492 2215 -481
rect 2014 -504 2120 -502
rect 1914 -582 1948 -540
rect 1861 -632 1898 -598
rect 1914 -618 1932 -582
rect 1937 -618 1948 -607
rect 1687 -647 1790 -638
rect 1625 -668 1644 -656
rect 1687 -663 1744 -647
rect 1760 -663 1790 -647
rect 1621 -687 1644 -668
rect 1698 -678 1744 -663
rect 1698 -687 1735 -678
rect 1861 -687 1895 -632
rect 1914 -674 1948 -618
rect 2032 -628 2048 -526
rect 2060 -560 2118 -554
rect 2249 -560 2264 -458
rect 2060 -594 2076 -560
rect 2060 -600 2118 -594
rect 2116 -641 2150 -636
rect 2016 -670 2017 -641
rect 2104 -650 2162 -641
rect 2248 -650 2264 -560
rect 2028 -670 2062 -653
rect 2104 -656 2150 -650
rect 2104 -670 2106 -656
rect 2116 -670 2150 -656
rect 2190 -670 2216 -650
rect 2230 -670 2264 -650
rect 2283 -560 2317 -439
rect 2383 -462 2492 -449
rect 2383 -491 2384 -462
rect 2426 -476 2492 -462
rect 2599 -484 2606 -439
rect 2616 -454 2686 -416
rect 2794 -448 2832 -442
rect 2968 -448 2982 -386
rect 2987 -448 3002 -374
rect 2794 -454 2856 -448
rect 2968 -454 3002 -448
rect 2616 -484 3002 -454
rect 2283 -563 2298 -560
rect 2283 -646 2317 -563
rect 2401 -575 2412 -526
rect 2425 -548 2426 -491
rect 2599 -494 3002 -484
rect 3021 -374 3038 -299
rect 3070 -333 3304 -299
rect 3358 -308 3371 -299
rect 3390 -308 3424 -280
rect 3358 -329 3424 -308
rect 3358 -333 3371 -329
rect 3390 -330 3424 -329
rect 3045 -374 3055 -333
rect 3021 -475 3055 -374
rect 3070 -419 3109 -333
rect 3337 -341 3371 -333
rect 3378 -341 3424 -330
rect 3337 -345 3358 -341
rect 3145 -376 3170 -367
rect 3141 -380 3204 -376
rect 3213 -380 3251 -363
rect 3141 -414 3251 -380
rect 3158 -419 3251 -414
rect 3258 -419 3263 -367
rect 3070 -426 3128 -419
rect 3158 -426 3304 -419
rect 3337 -426 3371 -345
rect 3082 -430 3089 -426
rect 3163 -435 3216 -426
rect 3224 -435 3229 -426
rect 3258 -430 3263 -426
rect 3163 -451 3200 -435
rect 3181 -473 3200 -451
rect 3216 -473 3246 -451
rect 3123 -475 3173 -473
rect 3211 -475 3261 -473
rect 3356 -475 3371 -426
rect 3390 -475 3424 -341
rect 3536 -348 3594 -342
rect 3536 -382 3548 -348
rect 3573 -382 3594 -348
rect 3536 -388 3594 -382
rect 3470 -458 3492 -392
rect 3601 -416 3622 -314
rect 3725 -342 3740 -246
rect 3498 -458 3550 -420
rect 3592 -458 3626 -424
rect 3706 -458 3740 -342
rect 3454 -475 3458 -458
rect 3470 -475 3740 -458
rect 3021 -492 3740 -475
rect 3021 -494 3550 -492
rect 2429 -507 2487 -501
rect 2429 -541 2441 -507
rect 2599 -518 3586 -494
rect 2599 -522 3608 -518
rect 2429 -547 2487 -541
rect 2599 -544 3620 -522
rect 3623 -544 3638 -529
rect 2599 -554 3638 -544
rect 2599 -560 3646 -554
rect 2530 -576 2553 -560
rect 2485 -588 2519 -583
rect 2385 -593 2443 -588
rect 2409 -600 2443 -593
rect 2397 -617 2443 -600
rect 2485 -604 2525 -588
rect 2599 -600 3638 -560
rect 3646 -588 3660 -560
rect 2485 -617 2519 -604
rect 2599 -617 3586 -600
rect 3592 -604 3640 -600
rect 3596 -610 3640 -604
rect 2347 -622 3586 -617
rect 2283 -670 2324 -646
rect 2347 -650 2371 -622
rect 2385 -628 3586 -622
rect 3614 -628 3640 -610
rect 3706 -628 3740 -492
rect 3759 -369 3793 -227
rect 3905 -295 3963 -289
rect 3905 -329 3917 -295
rect 3905 -335 3963 -329
rect 4092 -369 4162 -174
rect 5299 -227 5334 -193
rect 4274 -242 4332 -236
rect 4274 -276 4286 -242
rect 4274 -282 4332 -276
rect 4330 -352 4364 -318
rect 4444 -352 4478 -236
rect 4930 -280 4965 -246
rect 4561 -316 4596 -299
rect 3759 -405 4162 -369
rect 4192 -386 4227 -352
rect 4230 -386 4478 -352
rect 4525 -333 4596 -316
rect 4525 -386 4595 -333
rect 3759 -575 4173 -405
rect 3759 -628 4181 -575
rect 2385 -650 4181 -628
rect 2347 -651 4181 -650
rect 2347 -662 2381 -651
rect 2397 -662 2431 -651
rect 1914 -687 1960 -674
rect 1978 -678 2013 -670
rect 2016 -678 2162 -670
rect 1978 -687 2162 -678
rect 1545 -704 2162 -687
rect 2190 -704 2328 -670
rect 1545 -944 2012 -704
rect 2014 -809 2062 -704
rect 2104 -738 2106 -704
rect 2190 -725 2216 -704
rect 2190 -738 2217 -725
rect 2102 -772 2116 -738
rect 2147 -756 2162 -741
rect 2104 -806 2106 -772
rect 2120 -806 2162 -756
rect 2168 -772 2182 -766
rect 2164 -806 2186 -772
rect 2190 -799 2220 -738
rect 2230 -799 2264 -704
rect 2014 -821 2048 -809
rect 2104 -821 2162 -806
rect 2014 -858 2060 -821
rect 2116 -825 2164 -821
rect 2138 -834 2164 -825
rect 2190 -830 2278 -799
rect 2202 -834 2264 -830
rect 2092 -853 2164 -834
rect 2180 -853 2214 -849
rect 2014 -862 2048 -858
rect 2080 -862 2140 -853
rect 2174 -858 2226 -853
rect 2060 -868 2140 -862
rect 2180 -868 2226 -858
rect 2056 -902 2140 -868
rect 2056 -908 2122 -902
rect 2056 -918 2076 -908
rect 2080 -918 2122 -908
rect 2080 -922 2106 -918
rect 2032 -928 2106 -922
rect 2196 -928 2226 -868
rect 2032 -936 2138 -928
rect 1492 -958 2012 -944
rect 1492 -963 1526 -958
rect 1545 -961 2012 -958
rect 754 -976 1536 -963
rect 1573 -970 2012 -961
rect 2080 -958 2138 -936
rect 2168 -958 2226 -928
rect 2080 -970 2095 -958
rect 2180 -970 2226 -958
rect 2230 -970 2264 -834
rect 2283 -917 2328 -704
rect 2347 -756 2431 -662
rect 2347 -781 2412 -756
rect 2432 -768 2437 -651
rect 2455 -662 2473 -651
rect 2485 -662 2519 -651
rect 2599 -654 4181 -651
rect 4192 -652 4226 -386
rect 4230 -503 4280 -386
rect 4316 -454 4330 -420
rect 4361 -438 4376 -423
rect 4334 -488 4376 -438
rect 4384 -488 4398 -454
rect 4319 -503 4376 -488
rect 4242 -507 4260 -503
rect 4330 -507 4378 -503
rect 4352 -516 4378 -507
rect 4306 -524 4378 -516
rect 4286 -535 4378 -524
rect 4410 -535 4428 -531
rect 4286 -550 4354 -535
rect 4294 -558 4354 -550
rect 4410 -558 4440 -535
rect 4259 -569 4440 -558
rect 4270 -581 4440 -569
rect 4259 -592 4440 -581
rect 4444 -590 4478 -386
rect 4508 -469 4595 -386
rect 4707 -401 4765 -395
rect 4707 -435 4719 -401
rect 4896 -416 4911 -299
rect 4930 -416 4964 -280
rect 5076 -348 5134 -342
rect 5076 -382 5088 -348
rect 5076 -388 5134 -382
rect 5144 -416 5169 -392
rect 5265 -416 5280 -246
rect 4707 -441 4765 -435
rect 4497 -592 4595 -469
rect 4675 -505 4709 -469
rect 4663 -539 4809 -505
rect 4675 -567 4709 -539
rect 4849 -563 4863 -539
rect 4294 -615 4340 -592
rect 4306 -644 4340 -615
rect 4394 -626 4440 -592
rect 4306 -652 4352 -644
rect 4388 -652 4440 -626
rect 4444 -652 4478 -592
rect 4192 -654 4440 -652
rect 2460 -768 2465 -662
rect 2466 -688 2519 -662
rect 2466 -738 2531 -688
rect 2539 -738 2553 -719
rect 2466 -753 2553 -738
rect 2466 -759 2551 -753
rect 2466 -766 2531 -759
rect 2576 -766 2597 -661
rect 2466 -768 2597 -766
rect 2347 -818 2418 -781
rect 2454 -800 2512 -768
rect 2525 -769 2597 -768
rect 2599 -686 4440 -654
rect 4446 -686 4478 -652
rect 4480 -641 4595 -592
rect 4866 -601 5288 -416
rect 4691 -635 4753 -601
rect 4691 -641 4725 -635
rect 2599 -740 4226 -686
rect 4306 -694 4428 -686
rect 4306 -710 4352 -694
rect 4360 -700 4368 -694
rect 4324 -740 4352 -710
rect 4388 -728 4428 -694
rect 4366 -740 4374 -737
rect 4394 -740 4428 -728
rect 2525 -787 2579 -769
rect 2576 -796 2579 -787
rect 2599 -774 4440 -740
rect 4446 -774 4478 -740
rect 2565 -800 2583 -796
rect 2454 -801 2511 -800
rect 2429 -815 2446 -809
rect 2450 -812 2511 -801
rect 2561 -810 2595 -800
rect 2454 -815 2511 -812
rect 2347 -917 2381 -818
rect 2391 -830 2418 -818
rect 2425 -818 2511 -815
rect 2534 -812 2595 -810
rect 2391 -834 2412 -830
rect 2425 -849 2509 -818
rect 2534 -844 2549 -812
rect 2561 -815 2595 -812
rect 2565 -828 2595 -815
rect 2429 -855 2495 -849
rect 2449 -860 2495 -855
rect 2401 -865 2495 -860
rect 2401 -880 2464 -865
rect 2401 -883 2455 -880
rect 2552 -883 2595 -828
rect 2549 -917 2595 -883
rect 2599 -917 4226 -774
rect 4266 -808 4346 -774
rect 4252 -842 4354 -808
rect 2283 -922 2595 -917
rect 2598 -922 4226 -917
rect 4266 -876 4354 -842
rect 4266 -883 4346 -876
rect 4266 -885 4324 -883
rect 4332 -885 4346 -883
rect 4266 -895 4346 -885
rect 4360 -883 4440 -774
rect 4360 -895 4400 -883
rect 4410 -895 4440 -883
rect 4266 -899 4340 -895
rect 4354 -899 4428 -895
rect 4266 -908 4324 -899
rect 4354 -908 4412 -899
rect 4266 -919 4412 -908
rect 2283 -951 4226 -922
rect 4242 -921 4412 -919
rect 4242 -923 4276 -921
rect 4278 -923 4312 -921
rect 1573 -976 2226 -970
rect 2249 -976 2264 -970
rect 2294 -976 2328 -951
rect 2347 -976 2381 -951
rect 2461 -968 2495 -951
rect 2549 -968 2583 -951
rect 2616 -976 4226 -951
rect 732 -985 762 -976
rect 771 -982 4226 -976
rect 4230 -925 4312 -923
rect 4316 -923 4364 -921
rect 4366 -923 4400 -921
rect 4316 -925 4400 -923
rect 4230 -949 4282 -925
rect 4316 -936 4376 -925
rect 4444 -933 4478 -774
rect 4316 -942 4396 -936
rect 4230 -950 4280 -949
rect 4230 -959 4276 -950
rect 4324 -952 4400 -942
rect 771 -985 4198 -982
rect 4230 -984 4271 -959
rect 4272 -984 4276 -959
rect 4318 -959 4400 -952
rect 35 -1002 714 -990
rect 35 -1010 708 -1002
rect 725 -1008 4198 -985
rect 725 -1010 4181 -1008
rect 35 -1028 472 -1010
rect 540 -1022 656 -1010
rect 671 -1022 686 -1010
rect 35 -1052 534 -1028
rect 540 -1033 686 -1022
rect 708 -1022 1536 -1010
rect 1573 -1011 2226 -1010
rect 1568 -1022 2226 -1011
rect 2227 -1022 2238 -1011
rect 708 -1031 2238 -1022
rect 548 -1052 598 -1033
rect 708 -1052 2012 -1031
rect 2080 -1033 2138 -1031
rect 2168 -1033 2238 -1031
rect 2092 -1037 2126 -1033
rect 2180 -1037 2238 -1033
rect 23 -1094 34 -1083
rect 35 -1094 472 -1052
rect 534 -1071 614 -1052
rect 550 -1072 598 -1071
rect 558 -1086 584 -1072
rect 600 -1080 614 -1071
rect 596 -1084 622 -1080
rect 596 -1088 630 -1084
rect 16 -1114 472 -1094
rect 580 -1114 646 -1088
rect 708 -1111 1553 -1052
rect 1573 -1058 2012 -1052
rect 2204 -1052 2238 -1037
rect 2204 -1058 2215 -1052
rect 1573 -1063 2215 -1058
rect 2227 -1058 2238 -1052
rect 2283 -1022 2328 -1010
rect 2347 -1022 2577 -1010
rect 2616 -1022 4181 -1010
rect 2283 -1039 4181 -1022
rect 2227 -1063 2264 -1058
rect 1573 -1083 2208 -1063
rect 1573 -1092 2215 -1083
rect 1573 -1111 2012 -1092
rect 2120 -1094 2138 -1092
rect 0 -1182 472 -1114
rect 626 -1122 662 -1114
rect 610 -1129 676 -1122
rect 594 -1133 676 -1129
rect 494 -1139 552 -1133
rect 494 -1182 495 -1139
rect 538 -1145 552 -1142
rect 506 -1148 552 -1145
rect 500 -1150 552 -1148
rect 582 -1148 676 -1133
rect 582 -1150 662 -1148
rect 674 -1150 676 -1148
rect 708 -1124 2012 -1111
rect 708 -1150 1554 -1124
rect 1573 -1150 2012 -1124
rect 2030 -1102 2096 -1099
rect 2120 -1102 2130 -1094
rect 2030 -1112 2164 -1102
rect 2170 -1112 2186 -1092
rect 2030 -1114 2186 -1112
rect 2204 -1093 2220 -1092
rect 2204 -1094 2238 -1093
rect 2249 -1094 2264 -1063
rect 2030 -1124 2164 -1114
rect 2030 -1126 2096 -1124
rect 2120 -1126 2164 -1124
rect 2030 -1130 2164 -1126
rect 2204 -1122 2264 -1094
rect 2283 -1122 2328 -1039
rect 2347 -1122 2381 -1039
rect 2505 -1048 2539 -1039
rect 2383 -1052 2533 -1049
rect 2489 -1077 2555 -1052
rect 2599 -1079 4181 -1039
rect 4203 -1044 4226 -984
rect 4230 -985 4280 -984
rect 4306 -985 4310 -968
rect 4318 -974 4376 -959
rect 4384 -974 4398 -959
rect 4318 -976 4398 -974
rect 4318 -985 4390 -976
rect 4446 -985 4478 -933
rect 4480 -979 4578 -641
rect 4581 -679 4595 -641
rect 4623 -691 4681 -669
rect 4623 -703 4649 -691
rect 4735 -703 4769 -669
rect 4635 -737 4781 -703
rect 4849 -720 5288 -601
rect 5299 -597 5333 -227
rect 5445 -295 5503 -289
rect 5445 -329 5457 -295
rect 5445 -335 5503 -329
rect 5445 -495 5503 -489
rect 5445 -529 5457 -495
rect 5445 -535 5503 -529
rect 5299 -631 5334 -597
rect 5632 -631 5702 -174
rect 5814 -242 5872 -236
rect 5814 -276 5826 -242
rect 5814 -282 5872 -276
rect 5814 -550 5872 -544
rect 5814 -584 5826 -550
rect 5814 -590 5872 -584
rect 5632 -667 5685 -631
rect 6003 -686 6018 -140
rect 6037 -686 6071 -121
rect 6183 -189 6241 -183
rect 6183 -223 6195 -189
rect 6183 -229 6241 -223
rect 6183 -677 6241 -671
rect 6037 -707 6052 -686
rect 4849 -773 4947 -720
rect 4679 -807 4737 -801
rect 4679 -841 4691 -807
rect 4679 -847 4737 -841
rect 4849 -847 4936 -773
rect 5141 -815 5144 -720
rect 5169 -820 5172 -720
rect 5632 -722 6057 -707
rect 6183 -711 6195 -677
rect 6183 -717 6241 -711
rect 6372 -794 6387 -87
rect 6406 -726 6440 -68
rect 6552 -136 6610 -130
rect 6552 -170 6564 -136
rect 6552 -176 6610 -170
rect 6739 -385 6809 -15
rect 6921 -83 6979 -77
rect 6921 -117 6933 -83
rect 6921 -123 6979 -117
rect 6921 -283 6979 -277
rect 6921 -317 6933 -283
rect 6921 -323 6979 -317
rect 6739 -419 6810 -385
rect 7110 -400 7125 -3
rect 7144 12 7178 38
rect 7144 4 7460 12
rect 7144 -22 7179 4
rect 7252 -22 7386 4
rect 7144 -332 7178 -22
rect 7290 -30 7348 -24
rect 7286 -56 7352 -30
rect 7290 -64 7302 -56
rect 7290 -70 7348 -64
rect 7290 -230 7348 -224
rect 7290 -264 7302 -230
rect 7290 -270 7348 -264
rect 7144 -366 7179 -332
rect 7479 -347 7494 363
rect 7513 329 7548 363
rect 7513 125 7547 329
rect 7846 267 7916 384
rect 8229 373 8268 409
rect 8598 373 8651 409
rect 8967 391 9037 707
rect 9149 639 9207 645
rect 9149 605 9161 639
rect 9149 599 9207 605
rect 9149 439 9207 445
rect 9336 444 9406 744
rect 9614 734 9688 761
rect 9580 728 9602 732
rect 9614 728 9756 734
rect 9580 727 9614 728
rect 9676 727 9756 728
rect 9915 727 9930 1400
rect 9949 1366 9984 1400
rect 9949 727 9983 1366
rect 10095 1298 10153 1304
rect 10095 1264 10107 1298
rect 10095 1258 10153 1264
rect 10265 1095 10299 1113
rect 10265 1059 10335 1095
rect 10282 1025 10353 1059
rect 10633 1025 10668 1059
rect 10095 810 10153 816
rect 10095 776 10107 810
rect 10095 770 10153 776
rect 9518 694 9576 700
rect 9518 660 9530 694
rect 9564 693 9580 694
rect 9949 693 9964 727
rect 9518 654 9576 660
rect 9913 638 10012 691
rect 10282 674 10352 1025
rect 10634 1006 10668 1025
rect 10464 957 10522 963
rect 10464 923 10476 957
rect 10464 917 10522 923
rect 10464 757 10522 763
rect 10464 723 10476 757
rect 10464 717 10522 723
rect 10282 638 10335 674
rect 10653 621 10668 1006
rect 10687 972 10722 1006
rect 11002 972 11018 1006
rect 10687 621 10721 972
rect 11003 953 11018 972
rect 10833 904 10891 910
rect 10833 870 10845 904
rect 10833 864 10891 870
rect 10833 704 10891 710
rect 10833 670 10845 704
rect 10833 664 10891 670
rect 10687 587 10702 621
rect 11389 479 11442 989
rect 9149 405 9161 439
rect 9149 399 9207 405
rect 8950 390 9037 391
rect 9319 390 9406 444
rect 9474 433 9514 444
rect 9580 433 9620 444
rect 11758 426 11811 883
rect 9496 390 9598 420
rect 8935 366 9037 390
rect 8634 356 9037 366
rect 9322 356 9407 390
rect 9492 356 9602 390
rect 12127 373 12180 883
rect 8028 316 8086 322
rect 8028 282 8040 316
rect 8198 293 8232 322
rect 8620 293 8655 311
rect 8028 276 8086 282
rect 7659 261 7717 267
rect 7659 227 7671 261
rect 7659 221 7717 227
rect 7829 178 7916 267
rect 8198 257 8268 293
rect 7996 178 8030 212
rect 8084 178 8118 212
rect 8198 197 8286 257
rect 8347 197 8505 257
rect 8584 250 8655 293
rect 8716 250 8874 312
rect 8953 303 9024 356
rect 9085 303 9257 337
rect 9322 303 9406 356
rect 9518 352 9530 356
rect 9518 346 9576 352
rect 9514 336 9580 346
rect 7627 125 7661 159
rect 7715 125 7749 159
rect 7829 144 7917 178
rect 7978 144 8130 178
rect 8136 144 8152 178
rect 7513 91 7548 125
rect 7615 99 7761 125
rect 7767 111 7783 125
rect 7624 95 7752 99
rect 7621 91 7755 95
rect 7513 -41 7547 91
rect 7655 27 7721 61
rect 7655 -11 7721 23
rect 7829 0 7916 144
rect 8002 92 8030 114
rect 8074 92 8121 123
rect 8002 85 8042 92
rect 8072 85 8121 92
rect 8002 67 8121 85
rect 8009 55 8121 67
rect 7992 42 8122 55
rect 8024 36 8090 42
rect 8024 26 8042 36
rect 8072 26 8090 36
rect 8028 8 8086 14
rect 7513 -75 7548 -41
rect 7621 -45 7755 -41
rect 7662 -49 7714 -45
rect 7615 -75 7761 -49
rect 7513 -279 7547 -75
rect 7846 -94 7916 0
rect 7992 -5 8122 8
rect 8009 -17 8121 -5
rect 8002 -26 8121 -17
rect 8002 -42 8042 -26
rect 8072 -42 8112 -26
rect 8002 -64 8030 -42
rect 8084 -64 8112 -42
rect 7846 -128 7917 -94
rect 7984 -128 8130 -94
rect 7659 -177 7717 -171
rect 7659 -211 7671 -177
rect 7659 -217 7717 -211
rect 7513 -313 7548 -279
rect 7846 -313 7916 -128
rect 7996 -189 8030 -128
rect 8084 -189 8118 -128
rect 8198 -147 8285 197
rect 8584 161 8654 250
rect 8953 216 9023 303
rect 9322 260 9393 303
rect 9504 288 9562 294
rect 9504 284 9516 288
rect 9489 273 9577 284
rect 9500 261 9566 273
rect 9406 260 9660 261
rect 9674 260 9708 294
rect 9322 250 9708 260
rect 9322 241 9392 250
rect 9504 248 9562 250
rect 8778 167 8812 210
rect 8409 129 8443 155
rect 8361 89 8491 129
rect 8361 83 8411 89
rect 8365 79 8411 83
rect 8441 83 8491 89
rect 8441 79 8487 83
rect 8365 61 8405 79
rect 8447 61 8487 79
rect 8365 0 8399 61
rect 8453 0 8487 61
rect 8371 -11 8481 -7
rect 8365 -33 8487 -11
rect 8361 -39 8411 -33
rect 8441 -39 8491 -33
rect 8361 -79 8491 -39
rect 8409 -105 8443 -79
rect 8567 -111 8654 161
rect 8762 148 8828 167
rect 8936 151 9023 216
rect 9135 235 9193 241
rect 9135 201 9147 235
rect 9305 206 9392 241
rect 9135 195 9193 201
rect 9305 172 9393 206
rect 9460 172 9606 206
rect 9103 151 9137 167
rect 9191 151 9225 167
rect 8766 142 8824 148
rect 8734 129 8768 133
rect 8822 129 8856 133
rect 8734 117 8780 129
rect 8810 117 8856 129
rect 8734 114 8774 117
rect 8816 114 8856 117
rect 8734 -51 8768 114
rect 8822 -51 8856 114
rect 8734 -67 8856 -51
rect 8936 117 9024 151
rect 9091 117 9237 151
rect 8936 -67 9023 117
rect 9103 87 9137 117
rect 9191 87 9225 117
rect 9103 73 9225 87
rect 9103 69 9137 73
rect 9191 69 9225 73
rect 9135 49 9193 55
rect 9131 35 9197 49
rect 9147 15 9181 35
rect 9131 1 9197 15
rect 9135 -5 9193 1
rect 9103 -23 9137 -19
rect 9191 -23 9225 -19
rect 9103 -30 9149 -23
rect 9179 -30 9225 -23
rect 9103 -33 9143 -30
rect 9185 -33 9225 -30
rect 9103 -67 9137 -33
rect 9191 -67 9225 -33
rect 8731 -79 8859 -67
rect 8734 -83 8768 -79
rect 8822 -83 8856 -79
rect 8766 -98 8824 -92
rect 8198 -207 8286 -147
rect 8347 -207 8505 -147
rect 8584 -200 8654 -111
rect 8762 -117 8828 -98
rect 8936 -101 9024 -67
rect 9091 -101 9237 -67
rect 9243 -101 9259 -67
rect 8778 -160 8812 -117
rect 8936 -166 9023 -101
rect 9305 -122 9392 172
rect 9478 120 9506 142
rect 9550 120 9597 151
rect 9478 104 9518 120
rect 9548 104 9597 120
rect 9478 77 9597 104
rect 9460 27 9606 77
rect 9466 -1 9512 23
rect 9550 -1 9600 23
rect 9478 -4 9506 -1
rect 9550 -4 9597 -1
rect 9478 -20 9518 -4
rect 9548 -20 9597 -4
rect 9478 -54 9597 -20
rect 9478 -70 9518 -54
rect 9548 -70 9588 -54
rect 9478 -88 9506 -70
rect 9472 -122 9506 -88
rect 9560 -88 9588 -70
rect 9560 -122 9594 -88
rect 8584 -207 8655 -200
rect 8028 -232 8086 -226
rect 8028 -266 8040 -232
rect 8198 -243 8268 -207
rect 8584 -243 8637 -207
rect 8028 -272 8086 -266
rect 8198 -272 8232 -243
rect 8716 -262 8874 -200
rect 8953 -253 9023 -166
rect 9135 -151 9193 -145
rect 9135 -185 9147 -151
rect 9305 -156 9393 -122
rect 9460 -156 9606 -122
rect 9612 -145 9628 -122
rect 9135 -191 9193 -185
rect 9305 -191 9392 -156
rect 8953 -262 9024 -253
rect 8953 -298 9006 -262
rect 9322 -287 9392 -191
rect 9504 -204 9562 -198
rect 9504 -238 9516 -204
rect 9504 -244 9562 -238
rect 9674 -244 9708 250
rect 7846 -349 7899 -313
rect 9322 -323 9375 -287
rect 6739 -455 6792 -419
rect 6552 -624 6610 -618
rect 6552 -658 6564 -624
rect 6589 -658 6610 -624
rect 6552 -664 6610 -658
rect 6617 -692 6638 -626
rect 6406 -760 6441 -726
rect 6603 -796 6792 -739
rect 6001 -813 6057 -796
rect 4866 -943 4936 -847
rect 6001 -849 6423 -813
rect 5048 -862 5106 -856
rect 5048 -896 5060 -862
rect 5048 -902 5106 -896
rect 4866 -945 4919 -943
rect 4866 -963 4936 -945
rect 5048 -963 5083 -945
rect 4866 -964 5083 -963
rect 5122 -964 5302 -944
rect 4866 -978 5302 -964
rect 5363 -978 5398 -944
rect 4480 -982 4542 -979
rect 4480 -985 4532 -982
rect 2409 -1107 2475 -1095
rect 2599 -1096 4223 -1079
rect 4230 -1096 4578 -985
rect 4866 -998 5156 -978
rect 5364 -997 5398 -978
rect 4679 -1020 4694 -999
rect 4866 -1002 5082 -998
rect 4713 -1020 5082 -1002
rect 4623 -1021 5082 -1020
rect 4605 -1055 5082 -1021
rect 5383 -1040 5398 -997
rect 4606 -1056 5082 -1055
rect 2599 -1104 4578 -1096
rect 2409 -1112 2441 -1107
rect 2599 -1111 4181 -1104
rect 2409 -1122 2475 -1112
rect 2599 -1122 4191 -1111
rect 2030 -1133 2140 -1130
rect 2038 -1150 2140 -1133
rect 2204 -1150 4191 -1122
rect 4237 -1114 4578 -1104
rect 4623 -1114 5082 -1056
rect 4237 -1150 5082 -1114
rect 5162 -1150 5196 -1116
rect 5250 -1150 5284 -1116
rect 5364 -1150 5398 -1040
rect 5417 -1031 5452 -997
rect 5417 -1150 5451 -1031
rect 7208 -1063 7243 -1029
rect 5563 -1099 5621 -1093
rect 5563 -1112 5575 -1099
rect 5563 -1114 5609 -1112
rect 5563 -1116 5621 -1114
rect 5559 -1133 5625 -1116
rect 5733 -1122 5767 -1093
rect 6119 -1122 6330 -1067
rect 7209 -1082 7243 -1063
rect 5563 -1139 5621 -1133
rect 5535 -1150 5649 -1142
rect 5733 -1150 6076 -1122
rect 500 -1182 6076 -1150
rect 0 -1193 491 -1182
rect 494 -1184 6076 -1182
rect 0 -1196 480 -1193
rect 494 -1196 692 -1184
rect 0 -1197 481 -1196
rect 0 -1224 426 -1197
rect 438 -1198 481 -1197
rect 491 -1198 692 -1196
rect 708 -1190 4191 -1184
rect 708 -1196 4162 -1190
rect 708 -1197 3012 -1196
rect 708 -1198 1885 -1197
rect 438 -1202 1885 -1198
rect 1888 -1202 1948 -1197
rect 438 -1216 1948 -1202
rect 1978 -1216 3012 -1197
rect 463 -1224 481 -1216
rect 0 -1238 481 -1224
rect 491 -1224 552 -1216
rect 491 -1238 588 -1224
rect 0 -1248 426 -1238
rect 492 -1246 552 -1238
rect 594 -1246 640 -1216
rect 708 -1224 1948 -1216
rect 689 -1238 1948 -1224
rect 655 -1246 662 -1238
rect 492 -1248 580 -1246
rect 594 -1248 668 -1246
rect 0 -1250 438 -1248
rect 492 -1250 702 -1248
rect 0 -1252 426 -1250
rect 492 -1252 580 -1250
rect 0 -1266 444 -1252
rect 486 -1264 588 -1252
rect 594 -1264 668 -1250
rect 486 -1266 668 -1264
rect 0 -1287 426 -1266
rect 492 -1270 668 -1266
rect 674 -1252 702 -1250
rect 708 -1252 1948 -1238
rect 674 -1266 1948 -1252
rect 674 -1270 702 -1266
rect 708 -1270 1948 -1266
rect 438 -1287 1948 -1270
rect 0 -1304 1948 -1287
rect 0 -1376 472 -1304
rect 492 -1326 526 -1304
rect 533 -1313 546 -1304
rect 561 -1313 634 -1304
rect 533 -1317 540 -1313
rect 561 -1317 628 -1313
rect 561 -1326 614 -1317
rect 649 -1325 702 -1304
rect 0 -1408 485 -1376
rect 492 -1408 532 -1326
rect 561 -1341 618 -1326
rect 534 -1354 538 -1344
rect 534 -1360 560 -1354
rect 567 -1356 618 -1341
rect 567 -1360 626 -1356
rect 534 -1366 626 -1360
rect 630 -1366 702 -1325
rect 534 -1394 702 -1366
rect 534 -1400 560 -1394
rect 567 -1399 702 -1394
rect 708 -1326 1948 -1304
rect 1990 -1230 2036 -1216
rect 2042 -1230 2124 -1216
rect 1990 -1237 2124 -1230
rect 2130 -1237 3012 -1216
rect 1990 -1238 3012 -1237
rect 1990 -1241 2150 -1238
rect 1990 -1248 2156 -1241
rect 2159 -1248 2162 -1241
rect 1990 -1264 2177 -1248
rect 1990 -1289 2002 -1264
rect 1990 -1298 2005 -1289
rect 2010 -1298 2177 -1264
rect 1990 -1300 2062 -1298
rect 2090 -1300 2177 -1298
rect 1990 -1304 2072 -1300
rect 708 -1330 1953 -1326
rect 1990 -1330 2068 -1304
rect 2084 -1316 2177 -1300
rect 2084 -1330 2162 -1316
rect 708 -1399 1959 -1330
rect 1982 -1345 1987 -1341
rect 1976 -1346 1987 -1345
rect 2002 -1345 2068 -1330
rect 2070 -1332 2162 -1330
rect 2002 -1346 2062 -1345
rect 2070 -1346 2150 -1332
rect 1971 -1357 1995 -1346
rect 2002 -1348 2150 -1346
rect 2007 -1357 2104 -1348
rect 534 -1408 538 -1400
rect 567 -1406 1959 -1399
rect 0 -1432 540 -1408
rect 567 -1412 642 -1406
rect 567 -1418 628 -1412
rect 649 -1418 1959 -1406
rect 0 -1457 476 -1432
rect 0 -1462 472 -1457
rect 480 -1462 530 -1432
rect 552 -1448 628 -1418
rect 640 -1432 1959 -1418
rect 640 -1436 702 -1432
rect 640 -1448 701 -1436
rect 552 -1449 567 -1448
rect 552 -1453 560 -1449
rect 568 -1453 581 -1448
rect 586 -1452 614 -1448
rect 598 -1453 614 -1452
rect 640 -1449 655 -1448
rect 640 -1453 648 -1449
rect 674 -1452 689 -1448
rect 540 -1458 583 -1453
rect 540 -1460 567 -1458
rect 533 -1462 567 -1460
rect 568 -1462 583 -1458
rect 606 -1462 614 -1453
rect 628 -1462 671 -1453
rect 683 -1462 686 -1453
rect 708 -1462 1959 -1432
rect 0 -1470 1959 -1462
rect 0 -1486 472 -1470
rect 480 -1473 530 -1470
rect 533 -1473 1959 -1470
rect 488 -1486 506 -1473
rect 533 -1476 1219 -1473
rect 540 -1486 1219 -1476
rect 0 -1496 686 -1486
rect 706 -1496 1219 -1486
rect 0 -1540 472 -1496
rect 552 -1540 586 -1496
rect 593 -1540 598 -1496
rect 628 -1508 656 -1496
rect 671 -1508 686 -1496
rect 628 -1538 686 -1508
rect 640 -1540 686 -1538
rect 725 -1540 1219 -1496
rect 0 -1553 1219 -1540
rect 1239 -1553 1244 -1473
rect 1250 -1481 1356 -1473
rect 1421 -1481 1424 -1473
rect 1250 -1500 1424 -1481
rect 1250 -1516 1336 -1500
rect 1250 -1538 1279 -1516
rect 1284 -1527 1336 -1516
rect 1342 -1527 1424 -1500
rect 1446 -1475 1959 -1473
rect 1976 -1360 2062 -1357
rect 2070 -1360 2104 -1357
rect 2116 -1360 2150 -1348
rect 1976 -1406 2150 -1360
rect 2159 -1406 2162 -1332
rect 1976 -1421 2162 -1406
rect 2184 -1350 3012 -1238
rect 3021 -1264 3055 -1196
rect 3057 -1211 3091 -1196
rect 3119 -1207 3145 -1196
rect 3119 -1210 3169 -1207
rect 3223 -1210 3257 -1196
rect 3119 -1211 3181 -1210
rect 3211 -1211 3269 -1210
rect 3328 -1211 4162 -1196
rect 3057 -1227 4162 -1211
rect 4237 -1202 5414 -1184
rect 5417 -1202 5451 -1184
rect 5493 -1196 5665 -1184
rect 3057 -1245 4169 -1227
rect 3123 -1253 3181 -1245
rect 3211 -1253 3269 -1245
rect 3328 -1252 4169 -1245
rect 3135 -1257 3169 -1253
rect 3223 -1257 3257 -1253
rect 3328 -1263 4183 -1252
rect 3328 -1264 4172 -1263
rect 3021 -1268 4172 -1264
rect 4184 -1268 4191 -1238
rect 4237 -1252 5451 -1202
rect 5531 -1222 5565 -1196
rect 5619 -1217 5653 -1196
rect 5589 -1222 5653 -1217
rect 5713 -1212 5719 -1196
rect 5733 -1212 6076 -1184
rect 5589 -1230 5636 -1222
rect 4224 -1268 5451 -1252
rect 5521 -1264 5531 -1230
rect 5571 -1238 5639 -1230
rect 5539 -1258 5577 -1248
rect 5589 -1258 5639 -1238
rect 3021 -1279 5451 -1268
rect 3021 -1326 3036 -1279
rect 3101 -1291 3291 -1279
rect 3328 -1286 5451 -1279
rect 3152 -1298 3240 -1291
rect 3328 -1301 4163 -1286
rect 3021 -1331 3055 -1326
rect 3163 -1341 3229 -1308
rect 3328 -1326 4145 -1301
rect 4150 -1313 4163 -1301
rect 4150 -1317 4157 -1313
rect 1976 -1425 2138 -1421
rect 1976 -1468 2116 -1425
rect 2184 -1447 3029 -1350
rect 3328 -1357 4147 -1326
rect 4178 -1339 4195 -1286
rect 4178 -1341 4191 -1339
rect 4184 -1351 4191 -1341
rect 3153 -1366 3187 -1359
rect 3043 -1427 3297 -1393
rect 3328 -1407 3955 -1357
rect 4045 -1360 4049 -1357
rect 3971 -1392 3981 -1376
rect 3966 -1407 3981 -1392
rect 4062 -1387 4083 -1357
rect 4084 -1387 4147 -1357
rect 4203 -1387 4230 -1286
rect 4237 -1387 5451 -1286
rect 5539 -1266 5639 -1258
rect 5650 -1266 5665 -1251
rect 5519 -1298 5534 -1289
rect 5539 -1298 5665 -1266
rect 5519 -1302 5577 -1298
rect 5619 -1300 5665 -1298
rect 5585 -1302 5601 -1300
rect 5519 -1304 5601 -1302
rect 5477 -1330 5482 -1326
rect 5519 -1330 5577 -1304
rect 5477 -1342 5488 -1330
rect 4062 -1394 5451 -1387
rect 3328 -1410 3981 -1407
rect 3109 -1438 3143 -1434
rect 3197 -1438 3231 -1434
rect 1976 -1475 2047 -1468
rect 1446 -1498 2047 -1475
rect 1446 -1509 2016 -1498
rect 2022 -1509 2047 -1498
rect 2056 -1502 2138 -1468
rect 2058 -1509 2116 -1502
rect 1446 -1510 2158 -1509
rect 1290 -1531 1307 -1527
rect 1252 -1553 1279 -1538
rect 1336 -1550 1366 -1527
rect 1373 -1528 1408 -1527
rect 1373 -1550 1439 -1528
rect 1336 -1553 1439 -1550
rect 1446 -1543 1909 -1510
rect 1948 -1516 1953 -1510
rect 1965 -1516 2158 -1510
rect 2184 -1516 2218 -1447
rect 2221 -1516 3029 -1447
rect 3097 -1452 3155 -1438
rect 3185 -1452 3243 -1438
rect 3109 -1461 3143 -1452
rect 3197 -1461 3231 -1452
rect 1948 -1525 2787 -1516
rect 1948 -1536 2010 -1525
rect 2022 -1532 2070 -1525
rect 2017 -1536 2070 -1532
rect 2076 -1536 2787 -1525
rect 1948 -1543 2787 -1536
rect 1446 -1553 1902 -1543
rect 0 -1574 1902 -1553
rect 0 -1576 472 -1574
rect 552 -1576 586 -1574
rect 593 -1576 598 -1574
rect 640 -1576 674 -1574
rect 681 -1576 1902 -1574
rect 0 -1587 1902 -1576
rect 1914 -1553 1953 -1543
rect 1914 -1570 1948 -1553
rect 1968 -1556 2094 -1543
rect 1992 -1570 2094 -1556
rect 2117 -1570 2118 -1543
rect 2184 -1570 2218 -1543
rect 2221 -1547 2787 -1543
rect 2221 -1553 2830 -1547
rect 2221 -1570 2787 -1553
rect 1914 -1577 2787 -1570
rect 1914 -1581 2168 -1577
rect 1914 -1582 1956 -1581
rect 1965 -1582 1995 -1581
rect 1914 -1587 1995 -1582
rect 2010 -1587 2168 -1581
rect 0 -1604 2168 -1587
rect 2184 -1604 2218 -1577
rect 2221 -1587 2787 -1577
rect 2221 -1604 2547 -1587
rect 0 -1610 2147 -1604
rect 0 -1666 472 -1610
rect 496 -1618 617 -1610
rect 540 -1633 617 -1618
rect 660 -1629 686 -1610
rect 628 -1633 686 -1629
rect 694 -1612 2158 -1610
rect 2184 -1612 2547 -1604
rect 694 -1620 1936 -1612
rect 1999 -1620 2158 -1612
rect 694 -1621 2158 -1620
rect 694 -1623 1908 -1621
rect 2117 -1622 2118 -1621
rect 694 -1633 1885 -1623
rect 552 -1636 586 -1633
rect 524 -1637 586 -1636
rect 524 -1642 567 -1637
rect 520 -1654 586 -1642
rect 518 -1661 586 -1654
rect 35 -1696 43 -1666
rect 14 -1704 43 -1696
rect 69 -1704 103 -1666
rect 123 -1679 137 -1675
rect 211 -1679 245 -1675
rect 111 -1694 139 -1679
rect 199 -1690 257 -1679
rect 111 -1704 137 -1694
rect 199 -1704 245 -1690
rect 342 -1693 472 -1666
rect 520 -1662 586 -1661
rect 593 -1662 628 -1633
rect 660 -1637 674 -1633
rect 694 -1636 708 -1633
rect 711 -1636 1885 -1633
rect 520 -1664 628 -1662
rect 694 -1654 1885 -1636
rect 694 -1655 842 -1654
rect 890 -1655 1885 -1654
rect 520 -1671 586 -1664
rect 520 -1692 538 -1674
rect 546 -1676 586 -1671
rect 601 -1674 612 -1664
rect 568 -1680 580 -1676
rect 568 -1685 620 -1680
rect 568 -1692 646 -1685
rect 325 -1704 472 -1693
rect -14 -1751 472 -1704
rect 488 -1716 538 -1696
rect 580 -1714 646 -1692
rect 580 -1716 648 -1714
rect 491 -1723 538 -1716
rect 585 -1719 648 -1716
rect 580 -1723 648 -1719
rect 480 -1728 648 -1723
rect 480 -1732 670 -1728
rect 677 -1730 688 -1674
rect 694 -1704 824 -1655
rect 973 -1704 997 -1655
rect 999 -1657 1885 -1655
rect 1895 -1657 1908 -1623
rect 2218 -1626 2547 -1612
rect 2221 -1631 2547 -1626
rect 2184 -1642 2195 -1631
rect 2213 -1632 2547 -1631
rect 2213 -1642 2224 -1632
rect 999 -1674 1908 -1657
rect 2117 -1674 2124 -1642
rect 2184 -1674 2224 -1642
rect 2322 -1657 2547 -1632
rect 2590 -1632 2787 -1587
rect 2590 -1639 2801 -1632
rect 2959 -1639 3029 -1516
rect 3328 -1463 3407 -1410
rect 3516 -1423 3981 -1410
rect 3516 -1457 4003 -1423
rect 4049 -1447 5451 -1394
rect 5473 -1447 5488 -1342
rect 5511 -1345 5516 -1341
rect 5505 -1346 5516 -1345
rect 5531 -1345 5577 -1330
rect 5613 -1313 5665 -1300
rect 5672 -1313 5688 -1282
rect 5613 -1316 5688 -1313
rect 5613 -1332 5665 -1316
rect 5599 -1345 5604 -1341
rect 5500 -1357 5524 -1346
rect 5531 -1348 5576 -1345
rect 5593 -1346 5604 -1345
rect 5588 -1347 5607 -1346
rect 5619 -1347 5665 -1332
rect 5713 -1347 6076 -1212
rect 5536 -1357 5576 -1348
rect 3516 -1462 3981 -1457
rect 4049 -1462 5488 -1447
rect 3141 -1566 3199 -1560
rect 3328 -1565 3398 -1463
rect 3516 -1473 5488 -1462
rect 3516 -1479 4857 -1473
rect 3566 -1502 3611 -1479
rect 3665 -1502 3787 -1479
rect 3841 -1502 3881 -1479
rect 3921 -1491 4857 -1479
rect 3921 -1496 3981 -1491
rect 4017 -1493 4857 -1491
rect 4860 -1493 4867 -1473
rect 4975 -1474 5488 -1473
rect 5505 -1360 5576 -1357
rect 5578 -1360 6076 -1347
rect 5505 -1391 5570 -1360
rect 5577 -1370 5645 -1360
rect 5646 -1364 6076 -1360
rect 6119 -1137 6190 -1122
rect 7039 -1131 7097 -1125
rect 6119 -1364 6189 -1137
rect 7039 -1165 7051 -1131
rect 7039 -1171 7097 -1165
rect 6301 -1205 6359 -1199
rect 6301 -1239 6313 -1205
rect 6471 -1228 6505 -1210
rect 6893 -1228 6927 -1210
rect 6301 -1245 6359 -1239
rect 6471 -1264 6541 -1228
rect 5646 -1370 6189 -1364
rect 5577 -1373 6189 -1370
rect 5576 -1381 6189 -1373
rect 5576 -1391 5645 -1381
rect 5505 -1409 5645 -1391
rect 5713 -1400 6189 -1381
rect 6488 -1298 6559 -1264
rect 5505 -1457 5646 -1409
rect 5713 -1434 6201 -1400
rect 6257 -1434 6297 -1400
rect 5713 -1449 6189 -1434
rect 5505 -1474 5576 -1457
rect 4975 -1493 5576 -1474
rect 4017 -1496 5576 -1493
rect 3566 -1514 3600 -1502
rect 3680 -1514 3714 -1502
rect 3534 -1529 3600 -1514
rect 3608 -1529 3612 -1514
rect 3534 -1561 3612 -1529
rect 3141 -1588 3153 -1566
rect 3141 -1606 3199 -1588
rect 3113 -1634 3227 -1616
rect 3311 -1619 3398 -1565
rect 3466 -1572 3506 -1565
rect 3554 -1585 3615 -1561
rect 3554 -1596 3635 -1585
rect 3554 -1610 3604 -1596
rect 3510 -1619 3568 -1613
rect 2590 -1649 3029 -1639
rect 2590 -1657 2801 -1649
rect 2513 -1666 2547 -1657
rect 2576 -1666 2801 -1657
rect 999 -1685 1936 -1674
rect 2005 -1684 2093 -1674
rect 1967 -1685 2093 -1684
rect 2106 -1676 2224 -1674
rect 2106 -1685 2147 -1676
rect 2213 -1683 2224 -1676
rect 999 -1686 1925 -1685
rect 1967 -1686 2082 -1685
rect 2117 -1686 2147 -1685
rect 2190 -1686 2224 -1683
rect 999 -1691 2224 -1686
rect 999 -1704 1539 -1691
rect 694 -1712 1539 -1704
rect 1585 -1712 1589 -1691
rect 477 -1740 538 -1732
rect 568 -1740 670 -1732
rect 694 -1740 1607 -1712
rect 1619 -1717 1653 -1706
rect 1665 -1717 1695 -1691
rect 1715 -1706 1737 -1691
rect 1707 -1717 1741 -1706
rect 1821 -1712 1855 -1691
rect 1868 -1708 2224 -1691
rect 1753 -1717 1855 -1712
rect 1613 -1718 1665 -1717
rect 1616 -1729 1665 -1718
rect 1619 -1732 1665 -1729
rect 1700 -1732 1855 -1717
rect 1619 -1740 1661 -1732
rect 1707 -1740 1749 -1732
rect 1753 -1740 1855 -1732
rect 1874 -1740 1908 -1708
rect 1967 -1723 2082 -1708
rect 1967 -1734 2033 -1723
rect 2117 -1739 2124 -1708
rect 2190 -1712 2224 -1708
rect 2576 -1712 2787 -1666
rect 2959 -1702 3016 -1649
rect 3314 -1653 3399 -1619
rect 3495 -1630 3669 -1619
rect 3506 -1642 3572 -1630
rect 3623 -1642 3653 -1630
rect 3699 -1638 3714 -1514
rect 3495 -1653 3583 -1642
rect 3612 -1653 3664 -1642
rect 3314 -1702 3398 -1653
rect 3510 -1659 3568 -1653
rect 3506 -1669 3572 -1663
rect 3685 -1666 3714 -1638
rect 3733 -1514 3767 -1502
rect 3685 -1672 3719 -1666
rect 3733 -1672 3748 -1514
rect 3765 -1635 3767 -1533
rect 3835 -1536 3844 -1514
rect 3847 -1520 3881 -1502
rect 4049 -1508 5576 -1496
rect 4049 -1509 5451 -1508
rect 5477 -1509 5576 -1508
rect 5578 -1509 5646 -1457
rect 5720 -1499 6189 -1449
rect 6263 -1466 6297 -1434
rect 6275 -1496 6297 -1475
rect 4049 -1510 5687 -1509
rect 3847 -1536 3894 -1520
rect 3799 -1601 3801 -1567
rect 3835 -1601 3894 -1536
rect 4049 -1538 5436 -1510
rect 5477 -1520 5687 -1510
rect 5477 -1532 5676 -1520
rect 5738 -1530 6189 -1499
rect 5680 -1532 6189 -1530
rect 4049 -1543 5432 -1538
rect 5477 -1542 6189 -1532
rect 3778 -1644 3801 -1615
rect 3806 -1616 3829 -1615
rect 3787 -1666 3801 -1644
rect 3815 -1666 3829 -1616
rect 3835 -1617 3865 -1601
rect 3923 -1610 3941 -1567
rect 4049 -1576 5431 -1543
rect 5477 -1553 5482 -1542
rect 5483 -1543 6189 -1542
rect 5521 -1570 5566 -1543
rect 5521 -1572 5535 -1570
rect 3835 -1618 3850 -1617
rect 3923 -1618 3956 -1610
rect 3835 -1625 3875 -1618
rect 3923 -1625 3981 -1618
rect 4049 -1626 5417 -1576
rect 5420 -1582 5431 -1576
rect 4049 -1629 5414 -1626
rect 5424 -1629 5431 -1582
rect 5525 -1606 5535 -1572
rect 5539 -1572 5566 -1570
rect 5578 -1572 5623 -1543
rect 5539 -1577 5623 -1572
rect 5539 -1606 5566 -1577
rect 5525 -1612 5566 -1606
rect 5578 -1606 5623 -1577
rect 4049 -1634 5479 -1629
rect 3685 -1688 3748 -1672
rect 3767 -1672 3867 -1666
rect 3879 -1672 3937 -1666
rect 3767 -1683 3952 -1672
rect 3767 -1688 3867 -1683
rect 3685 -1692 3867 -1688
rect 2034 -1740 2064 -1739
rect 2190 -1740 2533 -1712
rect 477 -1751 2533 -1740
rect -14 -1774 2533 -1751
rect -14 -1782 538 -1774
rect 569 -1782 635 -1774
rect 694 -1780 1871 -1774
rect 1874 -1780 1925 -1774
rect 1950 -1775 2147 -1774
rect 1950 -1780 2158 -1775
rect 694 -1782 2158 -1780
rect -14 -1784 2158 -1782
rect -14 -1786 2170 -1784
rect -14 -1816 1917 -1786
rect -14 -1819 538 -1816
rect -14 -1908 412 -1819
rect 424 -1908 446 -1819
rect 449 -1828 467 -1819
rect 449 -1856 464 -1828
rect 454 -1897 464 -1856
rect 458 -1908 464 -1897
rect 470 -1882 538 -1819
rect 580 -1817 614 -1816
rect 580 -1828 626 -1817
rect 546 -1857 561 -1828
rect 574 -1857 626 -1828
rect 546 -1858 626 -1857
rect 641 -1858 648 -1828
rect 694 -1852 1917 -1816
rect 1937 -1792 1942 -1786
rect 1954 -1792 1971 -1786
rect 1937 -1812 1971 -1792
rect 553 -1859 620 -1858
rect 542 -1870 620 -1859
rect 553 -1875 620 -1870
rect 635 -1864 648 -1858
rect 660 -1858 675 -1854
rect 694 -1858 1925 -1852
rect 660 -1864 687 -1858
rect 635 -1875 687 -1864
rect 553 -1882 687 -1875
rect 470 -1908 687 -1882
rect -14 -1909 687 -1908
rect -14 -2014 412 -1909
rect 424 -1913 446 -1909
rect 515 -1916 516 -1909
rect 527 -1916 687 -1909
rect 502 -1950 687 -1916
rect 515 -1964 687 -1950
rect 515 -1976 675 -1964
rect 520 -1984 604 -1976
rect 439 -2010 444 -1997
rect 520 -2000 599 -1984
rect 541 -2004 556 -2000
rect 463 -2010 481 -2004
rect 491 -2010 556 -2004
rect 573 -2010 599 -2000
rect 615 -2004 621 -1976
rect 660 -2010 675 -1976
rect 677 -2010 687 -1964
rect -14 -2018 428 -2014
rect 481 -2018 599 -2010
rect -14 -2047 444 -2018
rect 481 -2040 509 -2018
rect 541 -2038 599 -2018
rect 629 -2038 687 -2010
rect 694 -1866 1908 -1858
rect 1909 -1866 1925 -1858
rect 1937 -1866 1942 -1812
rect 1950 -1828 1971 -1812
rect 1976 -1820 1983 -1786
rect 1988 -1812 2022 -1786
rect 2076 -1807 2110 -1786
rect 2046 -1812 2110 -1807
rect 1988 -1820 2009 -1812
rect 2046 -1820 2093 -1812
rect 1976 -1828 2009 -1820
rect 2028 -1828 2096 -1820
rect 1950 -1838 2009 -1828
rect 2046 -1830 2096 -1828
rect 2117 -1824 2170 -1786
rect 2117 -1828 2173 -1824
rect 2117 -1830 2170 -1828
rect 2190 -1830 2533 -1774
rect 1950 -1848 2034 -1838
rect 2046 -1848 2533 -1830
rect 1950 -1856 2533 -1848
rect 1950 -1858 1971 -1856
rect 1954 -1866 1971 -1858
rect 1976 -1866 1983 -1856
rect 694 -1870 1983 -1866
rect 694 -2010 1908 -1870
rect 1909 -1894 1925 -1870
rect 1937 -1874 1942 -1870
rect 1954 -1874 1971 -1870
rect 1988 -1879 2533 -1856
rect 1976 -1888 2533 -1879
rect 1954 -1894 1971 -1890
rect 1951 -1896 1971 -1894
rect 1934 -1932 1939 -1916
rect 1930 -2010 1939 -1932
rect 1954 -1931 1971 -1896
rect 1976 -1892 2034 -1888
rect 2037 -1892 2058 -1890
rect 1976 -1894 2058 -1892
rect 1976 -1920 2034 -1894
rect 2059 -1906 2533 -1888
rect 2059 -1920 2145 -1906
rect 1954 -1935 1973 -1931
rect 1982 -1935 2034 -1920
rect 2056 -1922 2145 -1920
rect 2056 -1930 2139 -1922
rect 2056 -1935 2122 -1930
rect 1968 -1936 1973 -1935
rect 1957 -1947 1981 -1936
rect 1988 -1938 2033 -1935
rect 2050 -1936 2122 -1935
rect 1993 -1947 2033 -1938
rect 2045 -1941 2122 -1936
rect 2153 -1941 2533 -1906
rect 2045 -1942 2533 -1941
rect 2045 -1947 2064 -1942
rect 2088 -1947 2122 -1942
rect 1968 -1950 2033 -1947
rect 2050 -1950 2122 -1947
rect 2159 -1950 2533 -1942
rect 1968 -1981 2027 -1950
rect 2034 -1963 2039 -1950
rect 2044 -1963 2102 -1950
rect 2033 -1976 2102 -1963
rect 2125 -1970 2159 -1950
rect 2033 -1981 2159 -1976
rect 1968 -1984 2159 -1981
rect 1968 -1991 2039 -1984
rect 2044 -1991 2102 -1984
rect 1968 -2004 2102 -1991
rect -14 -2052 412 -2047
rect 463 -2052 481 -2040
rect -14 -2069 481 -2052
rect 37 -2085 344 -2069
rect 356 -2085 481 -2069
rect 37 -2086 481 -2085
rect 463 -2092 481 -2086
rect 491 -2092 509 -2040
rect 553 -2042 587 -2038
rect 629 -2052 679 -2038
rect 694 -2040 1951 -2010
rect 1968 -2012 2159 -2004
rect 1968 -2026 2102 -2012
rect 2170 -2026 2533 -1950
rect 1968 -2031 2103 -2026
rect 694 -2052 1939 -2040
rect 1968 -2047 2039 -2031
rect 2044 -2047 2103 -2031
rect 1968 -2052 2027 -2047
rect 2056 -2052 2103 -2047
rect 2133 -2052 2533 -2026
rect 519 -2063 2533 -2052
rect 519 -2071 1355 -2063
rect 1398 -2071 2533 -2063
rect 519 -2076 2533 -2071
rect 535 -2086 2533 -2076
rect 711 -2122 1150 -2086
rect 477 -2158 1150 -2122
rect 1236 -2121 1271 -2086
rect 1274 -2090 1297 -2086
rect 1317 -2102 1324 -2086
rect 1393 -2088 1922 -2086
rect 1930 -2088 2027 -2086
rect 1393 -2092 1908 -2088
rect 1432 -2099 1908 -2092
rect 1934 -2099 2002 -2088
rect 2022 -2092 2027 -2088
rect 2056 -2092 2102 -2086
rect 2022 -2099 2033 -2092
rect 2050 -2099 2102 -2092
rect 1432 -2100 2170 -2099
rect 1359 -2106 1366 -2102
rect 1393 -2118 1425 -2102
rect 1359 -2120 1425 -2118
rect 1236 -2128 1259 -2121
rect 1375 -2124 1425 -2120
rect 1359 -2152 1425 -2124
rect 1432 -2128 1893 -2100
rect 1934 -2115 2170 -2100
rect 1934 -2120 1981 -2115
rect 1432 -2133 1889 -2128
rect 1432 -2158 1888 -2133
rect 1934 -2143 1939 -2120
rect 1951 -2122 1981 -2120
rect 2014 -2120 2056 -2115
rect 2090 -2120 2170 -2115
rect 2014 -2122 2044 -2120
rect 2103 -2122 2133 -2120
rect 1940 -2124 1992 -2122
rect 2003 -2124 2055 -2122
rect 1940 -2128 2084 -2124
rect 2092 -2128 2144 -2122
rect 1940 -2133 2144 -2128
rect 2204 -2133 2533 -2086
rect 1954 -2146 1981 -2133
rect 2014 -2146 2023 -2133
rect 477 -2175 1271 -2158
rect 1276 -2169 1888 -2158
rect 235 -2234 258 -2205
rect 263 -2206 286 -2205
rect 244 -2278 258 -2234
rect 240 -2282 258 -2278
rect 272 -2306 286 -2206
rect 477 -2244 721 -2175
rect 1082 -2226 1083 -2175
rect 1116 -2192 1271 -2175
rect 1287 -2181 1317 -2169
rect 1325 -2181 1888 -2169
rect 1276 -2186 1888 -2181
rect 1276 -2192 1328 -2186
rect 1449 -2245 1888 -2186
rect 1996 -2162 2023 -2146
rect 1996 -2167 2062 -2162
rect 1996 -2202 2023 -2167
rect 2103 -2212 2104 -2133
rect 1449 -2281 1871 -2245
rect 1881 -2264 1888 -2245
rect 2170 -2232 2181 -2221
rect 2193 -2232 2204 -2221
rect 2207 -2222 2533 -2133
rect 2576 -1727 2647 -1712
rect 2576 -2186 2646 -1727
rect 2959 -1738 2998 -1702
rect 3314 -1738 3381 -1702
rect 3685 -1712 3748 -1692
rect 3543 -1715 3645 -1712
rect 3666 -1715 3748 -1712
rect 3496 -1721 3645 -1715
rect 3481 -1732 3611 -1721
rect 3612 -1732 3664 -1721
rect 3492 -1734 3611 -1732
rect 3618 -1734 3653 -1732
rect 3685 -1734 3748 -1715
rect 3767 -1695 3867 -1692
rect 3875 -1695 3941 -1683
rect 3767 -1706 3952 -1695
rect 3767 -1716 3867 -1706
rect 3879 -1712 3937 -1706
rect 3752 -1720 3867 -1716
rect 3767 -1734 3867 -1720
rect 3875 -1722 3911 -1716
rect 3492 -1740 3787 -1734
rect 3492 -1744 3767 -1740
rect 3481 -1748 3767 -1744
rect 3398 -1755 3767 -1748
rect 3799 -1751 3867 -1734
rect 3953 -1740 3965 -1638
rect 4049 -1654 5414 -1634
rect 4009 -1706 4046 -1705
rect 4035 -1716 4046 -1706
rect 4049 -1712 4136 -1654
rect 4204 -1672 4236 -1654
rect 4204 -1675 4250 -1672
rect 4204 -1687 4251 -1675
rect 4206 -1709 4236 -1687
rect 4262 -1709 4278 -1687
rect 4064 -1716 4136 -1712
rect 4035 -1746 4136 -1716
rect 4035 -1751 4046 -1746
rect 4064 -1751 4136 -1746
rect 3496 -1761 3554 -1755
rect 3565 -1780 3594 -1755
rect 3665 -1774 3767 -1755
rect 3785 -1768 3867 -1751
rect 3911 -1768 4136 -1751
rect 4148 -1765 4170 -1732
rect 3785 -1774 4136 -1768
rect 2758 -1795 2816 -1789
rect 2758 -1829 2770 -1795
rect 2928 -1818 2962 -1800
rect 3350 -1818 3384 -1800
rect 2758 -1835 2816 -1829
rect 2928 -1854 2998 -1818
rect 2945 -1888 3016 -1854
rect 2758 -2103 2816 -2097
rect 2758 -2137 2770 -2103
rect 2758 -2143 2816 -2137
rect 2576 -2222 2629 -2186
rect 2170 -2264 2204 -2232
rect 1881 -2275 1922 -2264
rect 2092 -2266 2204 -2264
rect 1881 -2287 1911 -2275
rect 1870 -2288 1911 -2287
rect 1953 -2287 2019 -2274
rect 2092 -2275 2133 -2266
rect 2103 -2287 2133 -2275
rect 2193 -2277 2204 -2266
rect 2576 -2256 2787 -2222
rect 2945 -2239 3015 -1888
rect 3127 -1956 3185 -1950
rect 3127 -1990 3139 -1956
rect 3127 -1996 3185 -1990
rect 3127 -2156 3185 -2150
rect 3127 -2190 3139 -2156
rect 3127 -2196 3185 -2190
rect 2576 -2275 2753 -2256
rect 2945 -2275 2998 -2239
rect 1953 -2288 2030 -2287
rect 1870 -2298 2030 -2288
rect 2092 -2298 2144 -2287
rect 3314 -2292 3384 -1818
rect 3565 -1902 3620 -1780
rect 3665 -1808 4136 -1774
rect 4244 -1775 4278 -1709
rect 3665 -1902 3753 -1808
rect 3767 -1819 4123 -1808
rect 3767 -1824 3911 -1819
rect 3767 -1855 3909 -1824
rect 3947 -1831 3951 -1819
rect 3953 -1833 3987 -1819
rect 3999 -1832 4123 -1819
rect 4230 -1827 4356 -1824
rect 4418 -1827 4452 -1654
rect 4471 -1827 4486 -1654
rect 4195 -1832 4298 -1827
rect 3921 -1855 3933 -1851
rect 3953 -1855 3989 -1833
rect 3565 -1913 3598 -1902
rect 3666 -1913 3700 -1902
rect 3719 -1913 3753 -1902
rect 3799 -1897 3989 -1855
rect 3999 -1846 4298 -1832
rect 4299 -1838 4351 -1827
rect 4387 -1830 4486 -1827
rect 4502 -1830 4505 -1654
rect 4528 -1657 5414 -1654
rect 5424 -1657 5431 -1634
rect 4528 -1672 5457 -1657
rect 4528 -1674 5454 -1672
rect 5525 -1674 5559 -1612
rect 5578 -1674 5612 -1606
rect 5680 -1627 5691 -1543
rect 5680 -1642 5695 -1627
rect 5713 -1642 5747 -1543
rect 5750 -1615 6189 -1543
rect 6263 -1497 6297 -1496
rect 6263 -1507 6321 -1497
rect 6263 -1513 6359 -1507
rect 6263 -1547 6321 -1513
rect 6263 -1553 6359 -1547
rect 6263 -1563 6321 -1553
rect 6263 -1615 6297 -1563
rect 5750 -1632 6195 -1615
rect 5780 -1642 5826 -1632
rect 5680 -1674 5747 -1642
rect 4528 -1691 5457 -1674
rect 4528 -1706 5226 -1691
rect 4528 -1728 5034 -1706
rect 5056 -1718 5082 -1706
rect 5084 -1718 5110 -1706
rect 5076 -1728 5088 -1726
rect 4528 -1758 5088 -1728
rect 4528 -1778 5034 -1758
rect 4544 -1792 4874 -1778
rect 4544 -1796 4924 -1792
rect 4942 -1793 4997 -1785
rect 5000 -1786 5024 -1778
rect 4668 -1816 4924 -1796
rect 4958 -1816 4994 -1797
rect 5000 -1815 5028 -1786
rect 5036 -1793 5088 -1758
rect 5122 -1780 5148 -1776
rect 5102 -1793 5148 -1780
rect 4668 -1818 4675 -1816
rect 4787 -1820 4821 -1816
rect 4840 -1820 4874 -1816
rect 4387 -1838 4428 -1830
rect 4310 -1846 4340 -1838
rect 4398 -1846 4428 -1838
rect 4437 -1842 4505 -1830
rect 4471 -1846 4505 -1842
rect 4696 -1844 4896 -1820
rect 5008 -1821 5028 -1815
rect 4986 -1831 4994 -1825
rect 5056 -1826 5086 -1793
rect 5108 -1821 5110 -1793
rect 4998 -1831 5086 -1826
rect 4696 -1846 4703 -1844
rect 3999 -1861 4452 -1846
rect 3999 -1897 4105 -1861
rect 4144 -1895 4178 -1882
rect 3799 -1908 3967 -1897
rect 3999 -1898 4069 -1897
rect 3999 -1908 4103 -1898
rect 3799 -1909 4103 -1908
rect 3799 -1913 3867 -1909
rect 3565 -1914 3867 -1913
rect 3501 -2120 3504 -1976
rect 3540 -1982 3559 -1930
rect 3583 -1982 3598 -1967
rect 3529 -2092 3532 -2004
rect 3540 -2012 3598 -1982
rect 3583 -2014 3598 -2012
rect 3552 -2026 3598 -2014
rect 3666 -2026 3700 -1914
rect 3719 -1982 3753 -1914
rect 3719 -2012 3741 -1982
rect 3799 -2004 3801 -1914
rect 3827 -2004 3829 -1914
rect 3887 -2004 3899 -1909
rect 3911 -1935 3941 -1909
rect 3915 -1947 3933 -1935
rect 3915 -2004 3927 -1947
rect 4044 -1964 4103 -1909
rect 4044 -1975 4069 -1964
rect 4105 -1975 4173 -1897
rect 4352 -1924 4386 -1861
rect 4471 -1914 4486 -1846
rect 4502 -1880 4505 -1846
rect 4558 -1880 4748 -1864
rect 4502 -1891 4543 -1880
rect 4558 -1886 4626 -1880
rect 4627 -1886 4714 -1880
rect 4725 -1886 4748 -1880
rect 4502 -1903 4532 -1891
rect 4558 -1898 4748 -1886
rect 4491 -1914 4543 -1903
rect 4567 -1914 4748 -1898
rect 4806 -1914 4821 -1844
rect 4840 -1848 4896 -1844
rect 4906 -1848 4908 -1844
rect 4840 -1899 4928 -1848
rect 4982 -1865 5086 -1831
rect 4982 -1881 5040 -1865
rect 5056 -1881 5086 -1865
rect 5122 -1874 5148 -1793
rect 5156 -1780 5226 -1706
rect 5233 -1712 5243 -1691
rect 5233 -1726 5311 -1712
rect 5233 -1773 5332 -1726
rect 5237 -1780 5332 -1773
rect 5336 -1780 5366 -1691
rect 5378 -1780 5391 -1691
rect 5397 -1698 5457 -1691
rect 5493 -1676 5747 -1674
rect 5768 -1676 5826 -1642
rect 5493 -1697 5676 -1676
rect 5680 -1697 5747 -1676
rect 5493 -1698 5747 -1697
rect 5397 -1708 5747 -1698
rect 5780 -1691 5826 -1676
rect 5780 -1703 5814 -1691
rect 5424 -1712 5457 -1708
rect 5525 -1712 5612 -1708
rect 5424 -1743 5612 -1712
rect 5424 -1780 5454 -1743
rect 5457 -1780 5612 -1743
rect 5156 -1858 5270 -1780
rect 5311 -1791 5457 -1780
rect 5290 -1837 5457 -1791
rect 5460 -1792 5479 -1780
rect 5290 -1858 5324 -1837
rect 5344 -1841 5357 -1837
rect 5369 -1846 5412 -1837
rect 5432 -1841 5445 -1837
rect 5336 -1858 5439 -1846
rect 5156 -1869 5243 -1858
rect 5317 -1869 5324 -1858
rect 5327 -1869 5439 -1858
rect 5460 -1858 5483 -1792
rect 5460 -1865 5479 -1858
rect 5466 -1869 5479 -1865
rect 5491 -1869 5500 -1780
rect 5512 -1784 5612 -1780
rect 5680 -1784 5691 -1708
rect 5780 -1718 5826 -1703
rect 5512 -1798 5691 -1784
rect 5512 -1830 5730 -1798
rect 5734 -1830 5738 -1718
rect 5768 -1750 5826 -1718
rect 5780 -1765 5826 -1750
rect 5780 -1830 5814 -1765
rect 5823 -1810 5826 -1765
rect 5894 -1776 5928 -1632
rect 5947 -1750 5962 -1632
rect 6155 -1649 6195 -1632
rect 6251 -1649 6409 -1615
rect 6488 -1649 6558 -1298
rect 6670 -1366 6728 -1360
rect 6670 -1400 6682 -1366
rect 6670 -1406 6728 -1400
rect 6670 -1566 6728 -1560
rect 6670 -1600 6682 -1566
rect 6670 -1606 6728 -1600
rect 6263 -1705 6297 -1649
rect 6488 -1685 6541 -1649
rect 6524 -1702 6720 -1687
rect 6857 -1702 6927 -1228
rect 7039 -1619 7097 -1613
rect 7039 -1653 7051 -1619
rect 7039 -1659 7097 -1653
rect 6263 -1741 6333 -1705
rect 6857 -1738 6910 -1702
rect 5512 -1852 5756 -1830
rect 5780 -1852 5844 -1830
rect 5870 -1844 5873 -1810
rect 5894 -1844 5938 -1776
rect 5512 -1864 5613 -1852
rect 5512 -1869 5646 -1864
rect 5156 -1870 5646 -1869
rect 5025 -1896 5040 -1881
rect 4840 -1914 4940 -1899
rect 4840 -1948 4855 -1914
rect 4869 -1926 4940 -1914
rect 4994 -1926 5028 -1899
rect 4869 -1933 4928 -1926
rect 5156 -1933 5243 -1870
rect 5317 -1874 5324 -1870
rect 5366 -1878 5416 -1870
rect 5355 -1884 5416 -1878
rect 5351 -1908 5417 -1884
rect 5424 -1896 5454 -1870
rect 5466 -1874 5479 -1870
rect 5491 -1874 5500 -1870
rect 5525 -1883 5534 -1870
rect 5544 -1883 5559 -1870
rect 5355 -1918 5416 -1908
rect 5355 -1924 5413 -1918
rect 4872 -1938 5040 -1933
rect 5045 -1938 5097 -1933
rect 5173 -1938 5243 -1933
rect 5525 -1937 5559 -1883
rect 5578 -1930 5646 -1870
rect 5680 -1878 5844 -1852
rect 5680 -1883 5822 -1878
rect 5680 -1890 5826 -1883
rect 5688 -1921 5722 -1890
rect 5764 -1914 5768 -1890
rect 5776 -1903 5808 -1899
rect 5728 -1921 5752 -1914
rect 5688 -1930 5752 -1921
rect 5578 -1937 5613 -1930
rect 5720 -1931 5752 -1930
rect 5754 -1921 5770 -1914
rect 5776 -1921 5810 -1903
rect 5754 -1930 5810 -1921
rect 5754 -1931 5786 -1930
rect 5720 -1937 5734 -1931
rect 5764 -1937 5786 -1931
rect 5822 -1937 5890 -1890
rect 5894 -1937 5928 -1844
rect 4872 -1966 4896 -1938
rect 4044 -1976 4173 -1975
rect 4035 -2004 4046 -1999
rect 3992 -2010 4010 -2004
rect 4020 -2010 4046 -2004
rect 4052 -2010 4105 -1977
rect 4144 -1980 4178 -1979
rect 4878 -2004 4896 -1966
rect 4906 -2004 4924 -1938
rect 4952 -1964 4982 -1938
rect 5045 -1944 5243 -1938
rect 5056 -1956 5243 -1944
rect 5045 -1967 5243 -1956
rect 5173 -1968 5243 -1967
rect 5173 -1998 5226 -1968
rect 5232 -1979 5243 -1968
rect 5530 -1998 5559 -1937
rect 5173 -2003 5559 -1998
rect 3719 -2026 3753 -2012
rect 4035 -2013 4105 -2010
rect 3552 -2027 3821 -2026
rect 3552 -2052 3586 -2027
rect 3598 -2052 3821 -2027
rect 3833 -2052 3867 -2018
rect 3921 -2052 3955 -2018
rect 3967 -2052 4019 -2026
rect 4035 -2040 4438 -2013
rect 5209 -2020 5559 -2003
rect 5564 -1942 5822 -1937
rect 5564 -1971 5613 -1942
rect 5646 -1968 5676 -1942
rect 5684 -1960 5786 -1942
rect 5684 -1971 5797 -1960
rect 5879 -1971 5928 -1937
rect 5564 -2026 5612 -1971
rect 5696 -1976 5750 -1971
rect 5764 -1976 5786 -1971
rect 5696 -1977 5786 -1976
rect 5696 -1987 5734 -1977
rect 5764 -1987 5786 -1977
rect 5696 -2004 5722 -1987
rect 5880 -1990 5928 -1971
rect 5947 -1990 5981 -1750
rect 6263 -1775 6351 -1741
rect 6631 -1775 6666 -1741
rect 6893 -1755 7089 -1740
rect 7228 -1755 7243 -1082
rect 7262 -1116 7297 -1082
rect 7262 -1755 7296 -1116
rect 7408 -1184 7466 -1178
rect 7408 -1218 7420 -1184
rect 7408 -1224 7466 -1218
rect 7578 -1387 7612 -1369
rect 9422 -1381 9457 -1347
rect 7578 -1423 7648 -1387
rect 9423 -1400 9457 -1381
rect 7595 -1457 7666 -1423
rect 7946 -1457 7981 -1423
rect 7408 -1672 7466 -1666
rect 7408 -1706 7420 -1672
rect 7408 -1712 7466 -1706
rect 6049 -1930 6064 -1915
rect 6074 -1930 6089 -1928
rect 6049 -1943 6089 -1930
rect 6155 -1943 6195 -1936
rect 6047 -1960 6074 -1943
rect 6107 -1960 6116 -1943
rect 6093 -1990 6151 -1984
rect 5696 -2005 5810 -2004
rect 5880 -2010 5891 -1999
rect 5899 -2010 5928 -1990
rect 5173 -2028 5612 -2026
rect 3552 -2085 3624 -2052
rect 3632 -2085 3753 -2052
rect 3799 -2085 3967 -2052
rect 3969 -2085 3989 -2052
rect 3992 -2085 4019 -2052
rect 3552 -2086 4019 -2085
rect 4020 -2047 4404 -2040
rect 4020 -2052 4122 -2047
rect 4427 -2051 4438 -2040
rect 5159 -2039 5612 -2028
rect 5674 -2039 5722 -2018
rect 5756 -2039 5832 -2018
rect 5880 -2026 5928 -2010
rect 5933 -1998 5982 -1990
rect 5933 -2010 6029 -1998
rect 6078 -2001 6166 -1990
rect 5933 -2013 6040 -2010
rect 5933 -2024 6043 -2013
rect 5933 -2026 5981 -2024
rect 5880 -2039 6012 -2026
rect 5159 -2040 6012 -2039
rect 5159 -2052 5598 -2040
rect 5674 -2052 5832 -2040
rect 5880 -2052 6012 -2040
rect 6065 -2052 6074 -2004
rect 6089 -2013 6155 -2001
rect 6078 -2024 6166 -2013
rect 6093 -2030 6151 -2024
rect 6263 -2030 6350 -1775
rect 6632 -1794 6666 -1775
rect 6857 -1791 7071 -1758
rect 7262 -1789 7277 -1755
rect 7595 -1756 7665 -1457
rect 7947 -1476 7981 -1457
rect 7777 -1525 7835 -1519
rect 7777 -1559 7789 -1525
rect 7777 -1565 7835 -1559
rect 7777 -1725 7835 -1719
rect 7777 -1754 7789 -1725
rect 7777 -1756 7811 -1754
rect 7595 -1759 7811 -1756
rect 7595 -1765 7835 -1759
rect 7485 -1792 7516 -1774
rect 6462 -1843 6520 -1837
rect 6462 -1877 6474 -1843
rect 6462 -1883 6520 -1877
rect 6089 -2040 6155 -2034
rect 4020 -2064 4105 -2052
rect 4122 -2064 4404 -2052
rect 5175 -2054 5928 -2052
rect 5257 -2064 5483 -2054
rect 5530 -2064 5928 -2054
rect 4020 -2073 5928 -2064
rect 4020 -2085 5598 -2073
rect 5612 -2085 5914 -2073
rect 5933 -2085 6012 -2052
rect 4020 -2086 6012 -2085
rect 3552 -2124 3586 -2086
rect 3496 -2209 3554 -2203
rect 3496 -2243 3508 -2209
rect 3541 -2243 3554 -2209
rect 3496 -2249 3554 -2243
rect 3569 -2277 3582 -2226
rect 2180 -2298 2204 -2297
rect 240 -2310 286 -2306
rect 1818 -2334 2037 -2302
rect 3314 -2328 3367 -2292
rect 3685 -2345 3700 -2086
rect 3719 -2345 3753 -2086
rect 3992 -2092 4010 -2086
rect 4020 -2092 4122 -2086
rect 4206 -2092 4320 -2086
rect 4038 -2120 4122 -2092
rect 4234 -2115 4292 -2109
rect 4230 -2120 4296 -2115
rect 3865 -2262 3923 -2256
rect 3865 -2296 3877 -2262
rect 3865 -2302 3923 -2296
rect 3719 -2379 3734 -2345
rect 0 -2400 28 -2388
rect 1125 -2406 1167 -2382
rect 4052 -2398 4122 -2120
rect 4234 -2124 4280 -2120
rect 4234 -2149 4246 -2124
rect 4234 -2155 4292 -2149
rect 4234 -2315 4292 -2309
rect 4234 -2349 4246 -2315
rect 4234 -2355 4292 -2349
rect 26 -2428 28 -2416
rect 447 -2476 456 -2422
rect 1153 -2434 1167 -2410
rect 1329 -2420 1367 -2410
rect 501 -2499 510 -2476
rect 1329 -2556 1353 -2420
rect 4052 -2434 4105 -2398
rect 1357 -2448 1395 -2438
rect 1357 -2528 1381 -2448
rect 4423 -2451 4438 -2086
rect 4457 -2100 4492 -2086
rect 4553 -2100 4711 -2086
rect 4772 -2100 4807 -2086
rect 4457 -2451 4491 -2100
rect 4773 -2119 4807 -2100
rect 5159 -2098 5230 -2086
rect 5159 -2119 5229 -2098
rect 4603 -2168 4661 -2162
rect 4603 -2202 4615 -2168
rect 4603 -2208 4661 -2202
rect 4603 -2368 4661 -2362
rect 4603 -2402 4615 -2368
rect 4603 -2408 4661 -2402
rect 4457 -2485 4472 -2451
rect 4792 -2504 4807 -2119
rect 4826 -2120 5229 -2119
rect 4826 -2153 4861 -2120
rect 4826 -2504 4860 -2153
rect 4972 -2221 5030 -2215
rect 4972 -2255 4984 -2221
rect 4972 -2261 5030 -2255
rect 4972 -2421 5030 -2415
rect 4972 -2455 4984 -2421
rect 4972 -2461 5030 -2455
rect 1335 -2594 1353 -2556
rect 1363 -2594 1381 -2528
rect 4826 -2538 4841 -2504
rect 5159 -2557 5229 -2120
rect 5341 -2166 5399 -2160
rect 5341 -2200 5353 -2166
rect 5341 -2206 5399 -2200
rect 5341 -2474 5399 -2468
rect 5341 -2508 5353 -2474
rect 5341 -2514 5399 -2508
rect 5159 -2593 5212 -2557
rect 449 -2600 467 -2594
rect 477 -2600 495 -2594
rect 5530 -2610 5545 -2086
rect 5564 -2610 5598 -2086
rect 5678 -2120 5712 -2116
rect 5766 -2120 5800 -2116
rect 5710 -2527 5768 -2521
rect 5710 -2561 5722 -2527
rect 5710 -2567 5768 -2561
rect 449 -2682 467 -2630
rect 477 -2682 495 -2630
rect 5564 -2644 5579 -2610
rect 5899 -2663 5914 -2086
rect 5933 -2126 5968 -2086
rect 6051 -2092 6074 -2058
rect 6079 -2092 6137 -2086
rect 6064 -2103 6152 -2092
rect 6075 -2115 6141 -2103
rect 6064 -2119 6152 -2115
rect 5981 -2126 6235 -2119
rect 6280 -2126 6350 -2030
rect 6462 -2043 6520 -2037
rect 6462 -2077 6474 -2043
rect 6462 -2083 6520 -2077
rect 5933 -2663 5967 -2126
rect 6079 -2132 6137 -2126
rect 6280 -2179 6337 -2126
rect 6651 -2179 6666 -1794
rect 6685 -1828 6720 -1794
rect 7000 -1828 7035 -1794
rect 7262 -1808 7458 -1793
rect 7519 -1808 7550 -1792
rect 7423 -1811 7458 -1808
rect 6685 -2179 6719 -1828
rect 7001 -1847 7035 -1828
rect 7226 -1826 7458 -1811
rect 7226 -1844 7457 -1826
rect 6831 -1896 6889 -1890
rect 6831 -1930 6843 -1896
rect 6831 -1936 6889 -1930
rect 6831 -2096 6889 -2090
rect 6831 -2130 6843 -2096
rect 6831 -2136 6889 -2130
rect 6280 -2215 6319 -2179
rect 6685 -2213 6700 -2179
rect 7020 -2232 7035 -1847
rect 7054 -1881 7089 -1847
rect 7054 -2232 7088 -1881
rect 7200 -1949 7258 -1943
rect 7200 -1983 7212 -1949
rect 7200 -1989 7258 -1983
rect 7200 -2149 7258 -2143
rect 7200 -2183 7212 -2149
rect 7200 -2189 7258 -2183
rect 7054 -2266 7069 -2232
rect 6249 -2295 6283 -2277
rect 7387 -2285 7457 -1844
rect 7595 -1888 7809 -1765
rect 7966 -1861 7981 -1476
rect 8000 -1510 8035 -1476
rect 8315 -1510 8350 -1476
rect 8738 -1493 8773 -1475
rect 8000 -1861 8034 -1510
rect 8316 -1529 8350 -1510
rect 8702 -1508 8773 -1493
rect 8146 -1578 8204 -1572
rect 8146 -1612 8158 -1578
rect 8146 -1618 8204 -1612
rect 8146 -1778 8204 -1772
rect 8146 -1812 8158 -1778
rect 8146 -1818 8204 -1812
rect 7569 -1894 7809 -1888
rect 7569 -1928 7581 -1894
rect 7595 -1897 7809 -1894
rect 8000 -1895 8015 -1861
rect 8335 -1862 8350 -1529
rect 8369 -1563 8404 -1529
rect 8369 -1862 8403 -1563
rect 8515 -1631 8573 -1625
rect 8515 -1665 8527 -1631
rect 8515 -1671 8573 -1665
rect 8515 -1831 8573 -1825
rect 8515 -1860 8527 -1831
rect 8515 -1862 8549 -1860
rect 8125 -1865 8549 -1862
rect 8125 -1871 8573 -1865
rect 8125 -1899 8547 -1871
rect 7739 -1917 7773 -1899
rect 8000 -1914 8547 -1899
rect 7569 -1934 7627 -1928
rect 7739 -1953 7809 -1917
rect 8125 -1950 8547 -1914
rect 7756 -1987 7827 -1953
rect 7569 -2202 7627 -2196
rect 7569 -2236 7581 -2202
rect 7569 -2242 7627 -2236
rect 6249 -2331 6319 -2295
rect 7387 -2321 7440 -2285
rect 7756 -2328 7826 -1987
rect 7938 -2055 7996 -2049
rect 7938 -2089 7950 -2055
rect 7938 -2095 7996 -2089
rect 7938 -2255 7996 -2249
rect 7938 -2289 7950 -2255
rect 7938 -2295 7996 -2289
rect 6266 -2365 6337 -2331
rect 6617 -2365 6652 -2331
rect 7423 -2338 7826 -2328
rect 6079 -2580 6137 -2574
rect 6079 -2614 6091 -2580
rect 6079 -2620 6137 -2614
rect 5933 -2697 5948 -2663
rect 6266 -2716 6336 -2365
rect 6618 -2384 6652 -2365
rect 6448 -2433 6506 -2427
rect 6448 -2467 6460 -2433
rect 6448 -2473 6506 -2467
rect 6448 -2633 6506 -2627
rect 6448 -2667 6460 -2633
rect 6448 -2673 6506 -2667
rect 6266 -2752 6319 -2716
rect 6637 -2769 6652 -2384
rect 6671 -2418 6706 -2384
rect 6986 -2418 7021 -2384
rect 7409 -2401 7444 -2383
rect 6671 -2769 6705 -2418
rect 6987 -2437 7021 -2418
rect 7373 -2416 7444 -2401
rect 7756 -2391 7813 -2338
rect 8125 -2391 8195 -1950
rect 8333 -1994 8547 -1950
rect 8307 -2000 8547 -1994
rect 8307 -2034 8319 -2000
rect 8333 -2003 8547 -2000
rect 8702 -1967 8772 -1508
rect 8884 -1576 8942 -1570
rect 8884 -1610 8896 -1576
rect 8884 -1616 8942 -1610
rect 8884 -1884 8942 -1878
rect 8884 -1918 8896 -1884
rect 8884 -1924 8942 -1918
rect 8702 -2003 8755 -1967
rect 8702 -2005 8801 -2003
rect 8961 -2004 8992 -1986
rect 9073 -2004 9088 -1474
rect 9107 -2004 9141 -1420
rect 9253 -1449 9311 -1443
rect 9253 -1483 9265 -1449
rect 9253 -1489 9311 -1483
rect 9253 -1937 9311 -1931
rect 9253 -1966 9265 -1937
rect 9253 -1970 9287 -1966
rect 9249 -1971 9287 -1970
rect 9253 -1977 9311 -1971
rect 8477 -2023 8511 -2005
rect 8702 -2020 8934 -2005
rect 8995 -2020 9026 -2004
rect 9141 -2005 9249 -2004
rect 8702 -2023 8801 -2020
rect 8899 -2023 8934 -2020
rect 8307 -2040 8365 -2034
rect 8477 -2059 8547 -2023
rect 8702 -2038 8934 -2023
rect 9141 -2038 9215 -2005
rect 8702 -2056 8933 -2038
rect 8494 -2093 8565 -2059
rect 8307 -2308 8365 -2302
rect 8307 -2342 8319 -2308
rect 8307 -2348 8365 -2342
rect 6817 -2486 6875 -2480
rect 6817 -2520 6829 -2486
rect 6817 -2526 6875 -2520
rect 6817 -2686 6875 -2680
rect 6817 -2720 6829 -2686
rect 6817 -2726 6875 -2720
rect 0 -2800 40 -2788
rect 6671 -2803 6686 -2769
rect 26 -2828 40 -2816
rect 7006 -2822 7021 -2437
rect 7040 -2471 7075 -2437
rect 7040 -2822 7074 -2471
rect 7186 -2539 7244 -2533
rect 7186 -2573 7198 -2539
rect 7186 -2579 7244 -2573
rect 7186 -2739 7244 -2733
rect 7186 -2773 7198 -2739
rect 7186 -2779 7244 -2773
rect 7040 -2856 7055 -2822
rect 7373 -2875 7443 -2416
rect 7756 -2427 7795 -2391
rect 8125 -2427 8178 -2391
rect 8494 -2434 8564 -2093
rect 8676 -2161 8734 -2155
rect 8676 -2195 8688 -2161
rect 8676 -2201 8734 -2195
rect 8676 -2361 8734 -2355
rect 8676 -2395 8688 -2361
rect 8676 -2401 8734 -2395
rect 8161 -2444 8564 -2434
rect 7555 -2484 7613 -2478
rect 7555 -2518 7567 -2484
rect 7725 -2507 7759 -2489
rect 8147 -2507 8182 -2489
rect 7555 -2524 7613 -2518
rect 7725 -2543 7795 -2507
rect 8111 -2522 8182 -2507
rect 8494 -2497 8551 -2444
rect 8863 -2497 8933 -2056
rect 9141 -2066 9215 -2039
rect 9107 -2072 9129 -2068
rect 9141 -2072 9283 -2066
rect 9107 -2073 9141 -2072
rect 9203 -2073 9283 -2072
rect 9442 -2073 9457 -1400
rect 9476 -1434 9511 -1400
rect 9476 -2073 9510 -1434
rect 9622 -1502 9680 -1496
rect 9622 -1536 9634 -1502
rect 9622 -1542 9680 -1536
rect 9792 -1705 9826 -1687
rect 9792 -1741 9862 -1705
rect 9809 -1775 9880 -1741
rect 10160 -1775 10195 -1741
rect 9622 -1990 9680 -1984
rect 9622 -2024 9634 -1990
rect 9622 -2030 9680 -2024
rect 9045 -2106 9103 -2100
rect 9045 -2140 9057 -2106
rect 9091 -2107 9107 -2106
rect 9476 -2107 9491 -2073
rect 9045 -2146 9103 -2140
rect 9440 -2162 9539 -2109
rect 9809 -2126 9879 -1775
rect 10161 -1794 10195 -1775
rect 9991 -1843 10049 -1837
rect 9991 -1877 10003 -1843
rect 9991 -1883 10049 -1877
rect 9991 -2043 10049 -2037
rect 9991 -2077 10003 -2043
rect 9991 -2083 10049 -2077
rect 9809 -2162 9862 -2126
rect 10180 -2179 10195 -1794
rect 10214 -1828 10249 -1794
rect 10529 -1828 10564 -1794
rect 10952 -1811 10987 -1793
rect 10214 -2179 10248 -1828
rect 10530 -1847 10564 -1828
rect 10916 -1826 10987 -1811
rect 10360 -1896 10418 -1890
rect 10360 -1930 10372 -1896
rect 10360 -1936 10418 -1930
rect 10360 -2096 10418 -2090
rect 10360 -2130 10372 -2096
rect 10360 -2136 10418 -2130
rect 10214 -2213 10229 -2179
rect 10549 -2232 10564 -1847
rect 10583 -1881 10618 -1847
rect 10583 -2232 10617 -1881
rect 10729 -1949 10787 -1943
rect 10729 -1983 10741 -1949
rect 10729 -1989 10787 -1983
rect 10729 -2149 10787 -2143
rect 10729 -2183 10741 -2149
rect 10729 -2189 10787 -2183
rect 10583 -2266 10598 -2232
rect 10916 -2285 10986 -1826
rect 10916 -2321 10969 -2285
rect 11285 -2374 11338 -1917
rect 9045 -2414 9103 -2408
rect 9045 -2448 9057 -2414
rect 11654 -2427 11707 -1917
rect 9045 -2454 9103 -2448
rect 12023 -2480 12076 -2023
rect 7742 -2577 7813 -2543
rect 7555 -2792 7613 -2786
rect 7555 -2826 7567 -2792
rect 7555 -2832 7613 -2826
rect 7373 -2911 7426 -2875
rect 7742 -2928 7812 -2577
rect 7924 -2645 7982 -2639
rect 7924 -2679 7936 -2645
rect 7924 -2685 7982 -2679
rect 7924 -2845 7982 -2839
rect 7924 -2879 7936 -2845
rect 7924 -2885 7982 -2879
rect 7742 -2964 7795 -2928
rect 8111 -2981 8181 -2522
rect 8494 -2533 8533 -2497
rect 8863 -2533 8916 -2497
rect 8899 -2550 9249 -2540
rect 8293 -2590 8351 -2584
rect 8293 -2624 8305 -2590
rect 8463 -2613 8497 -2595
rect 8885 -2613 8920 -2595
rect 8293 -2630 8351 -2624
rect 8463 -2649 8533 -2613
rect 8849 -2628 8920 -2613
rect 8480 -2683 8551 -2649
rect 8293 -2898 8351 -2892
rect 8293 -2932 8305 -2898
rect 8293 -2938 8351 -2932
rect 200 -3016 226 -2998
rect 1153 -3010 1353 -2992
rect 8111 -3017 8164 -2981
rect 200 -3044 240 -3026
rect 1167 -3038 1367 -3020
rect 8480 -3034 8550 -2683
rect 8662 -2751 8720 -2745
rect 8662 -2785 8674 -2751
rect 8662 -2791 8720 -2785
rect 8662 -2951 8720 -2945
rect 8662 -2985 8674 -2951
rect 8662 -2991 8720 -2985
rect 8480 -3070 8533 -3034
rect 8849 -3087 8919 -2628
rect 9031 -2696 9089 -2690
rect 9031 -2730 9043 -2696
rect 9031 -2736 9089 -2730
rect 9031 -3004 9089 -2998
rect 9031 -3038 9043 -3004
rect 9031 -3044 9089 -3038
rect 8849 -3123 8902 -3087
rect 0 -3200 40 -3188
rect 26 -3228 40 -3216
rect 26 -3416 226 -3398
rect 1153 -3410 1353 -3392
rect 40 -3444 240 -3426
rect 1167 -3438 1367 -3420
rect 26 -3816 226 -3798
rect 1153 -3810 1353 -3792
rect 40 -3844 240 -3826
rect 1167 -3838 1367 -3820
rect 1153 -4210 1353 -4192
rect 1167 -4238 1367 -4220
<< nwell >>
rect 56 972 3586 1174
rect 3506 544 3586 972
rect 3508 -922 3586 -494
rect 56 -1196 3586 -922
<< poly >>
rect -158 40 -128 1174
rect -86 148 -56 1174
rect 3024 1144 3560 1174
rect 3492 760 3550 788
rect 3426 734 3550 760
rect -86 132 16 148
rect -86 98 -34 132
rect 0 112 16 132
rect 0 98 76 112
rect -86 82 76 98
rect -158 10 70 40
rect -158 -1196 -128 10
rect -86 -48 82 -32
rect -86 -82 -34 -48
rect 0 -62 82 -48
rect 0 -82 16 -62
rect -86 -98 16 -82
rect -86 -1196 -56 -98
rect 3520 -540 3550 734
rect 3520 -556 3586 -540
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 3520 -606 3586 -590
rect 3490 -736 3560 -702
rect 3426 -756 3560 -736
rect 3422 -842 3488 -826
rect 3422 -876 3438 -842
rect 3472 -876 3488 -842
rect 3422 -892 3488 -876
rect 3422 -896 3452 -892
rect 3024 -926 3452 -896
rect 3530 -1196 3560 -756
<< polycont >>
rect -34 98 0 132
rect -34 -82 0 -48
rect 3536 -590 3570 -556
rect 3438 -876 3472 -842
<< locali >>
rect -50 98 -34 132
rect 0 98 16 132
rect -50 -82 -34 -48
rect 0 -82 16 -48
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 3422 -876 3438 -842
rect 3472 -876 3488 -842
<< viali >>
rect -34 98 0 132
rect -34 -82 0 -48
rect 3536 -590 3570 -556
rect 3438 -876 3472 -842
<< metal1 >>
rect 56 972 3586 1174
rect 58 200 3586 206
rect 0 148 3586 200
rect -50 132 3586 148
rect -50 98 -34 132
rect 0 98 3586 132
rect -50 82 3586 98
rect -34 0 3586 82
rect -34 -32 0 0
rect -50 -48 16 -32
rect -50 -82 -34 -48
rect 0 -82 16 -48
rect -50 -98 16 -82
rect 58 -156 3586 0
rect 0 -400 200 -200
rect 3520 -556 3586 -540
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 0 -800 200 -600
rect 3520 -606 3586 -590
rect 3520 -826 3554 -606
rect 3422 -842 3554 -826
rect 3422 -876 3438 -842
rect 3472 -860 3554 -842
rect 3472 -876 3488 -860
rect 3422 -892 3488 -876
rect 56 -1000 3586 -922
rect 0 -1196 3586 -1000
rect 0 -1200 200 -1196
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
<< metal2 >>
rect 2946 364 2998 416
rect 2946 -366 2998 -314
use c1b  c1b_1
timestamp 1624053917
transform 1 0 58 0 -1 -68
box -85 -5128 9686 1784
use c1b  c1b_0
timestamp 1624053917
transform 1 0 58 0 1 118
box -85 -5128 9686 1784
use c1b  x1
timestamp 1624053917
transform 1 0 72 0 1 708
box -85 -5128 9686 1784
use c1b  x2
timestamp 1624053917
transform 1 0 3601 0 1 708
box -85 -5128 9686 1784
<< labels >>
rlabel metal2 2946 364 2998 416 1 b0
rlabel metal2 2946 -366 2998 -314 1 b1
rlabel poly -150 1154 -134 1170 1 clr
rlabel poly -78 1154 -62 1170 1 clk
rlabel metal1 3476 0 3506 58 1 vss
rlabel metal1 924 -996 966 -968 1 vdd
rlabel metal1 3466 992 3496 1050 1 vdd
rlabel poly -78 -54 -62 -38 1 clk
rlabel poly 3540 1152 3552 1168 1 ce
rlabel poly 3538 -916 3554 -874 1 out
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 ce
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 clr
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 b0
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 b1
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 out
port 8 nsew
<< end >>
