magic
tech sky130A
magscale 1 2
timestamp 1616102052
<< nwell >>
rect 428 1004 1392 1008
rect 122 736 1756 1004
rect 120 516 1756 736
rect 120 114 1758 516
rect 120 110 1756 114
<< pwell >>
rect 120 -442 1750 -22
rect 120 -902 1744 -442
<< psubdiff >>
rect 268 -782 292 -602
rect 1632 -782 1656 -602
<< nsubdiff >>
rect 580 958 1320 960
rect 568 928 1328 958
rect 568 832 610 928
rect 1288 832 1328 928
rect 568 792 1328 832
<< psubdiffcont >>
rect 292 -782 1632 -602
<< nsubdiffcont >>
rect 610 832 1288 928
<< poly >>
rect 362 718 392 748
rect 1382 718 1468 730
rect 360 712 1468 718
rect 360 678 1412 712
rect 1446 678 1468 712
rect 360 668 1468 678
rect 362 436 392 668
rect 1382 654 1468 668
rect 636 588 1328 626
rect 638 426 668 588
rect 1290 402 1328 588
rect 266 -68 296 226
rect 362 -70 392 224
rect 638 92 668 228
rect 438 58 668 92
rect 438 24 462 58
rect 496 54 668 58
rect 496 24 514 54
rect 438 8 514 24
rect 458 -78 488 8
rect 734 -24 764 224
rect 916 -24 950 -20
rect 554 -62 952 -24
rect 554 -76 584 -62
rect 266 -444 296 -282
rect 916 -334 950 -62
rect 1294 -80 1324 170
rect 1626 66 1656 166
rect 1478 32 1656 66
rect 1276 -260 1342 -202
rect 1478 -334 1516 32
rect 1626 -82 1656 32
rect 916 -366 1516 -334
rect 1782 -444 1848 -426
rect 266 -452 1848 -444
rect 266 -492 1792 -452
rect 1838 -492 1848 -452
rect 266 -494 1848 -492
rect 1782 -510 1848 -494
<< polycont >>
rect 1412 678 1446 712
rect 462 24 496 58
rect 1792 -492 1838 -452
<< locali >>
rect 1388 716 1464 724
rect 1388 672 1400 716
rect 1450 672 1464 716
rect 1388 662 1464 672
rect 438 62 514 70
rect 438 18 450 62
rect 500 18 514 62
rect 438 8 514 18
rect 1782 -444 1848 -426
rect 1782 -496 1792 -444
rect 1840 -496 1848 -444
rect 1782 -510 1848 -496
rect 276 -782 292 -602
rect 1632 -782 1648 -602
<< viali >>
rect 154 928 1714 970
rect 154 854 610 928
rect 568 832 610 854
rect 610 832 1288 928
rect 1288 854 1714 928
rect 1288 832 1328 854
rect 568 792 1328 832
rect 1400 712 1450 716
rect 1400 678 1412 712
rect 1412 678 1446 712
rect 1446 678 1450 712
rect 1400 672 1450 678
rect 924 108 972 164
rect 92 10 154 72
rect 450 58 500 62
rect 450 24 462 58
rect 462 24 496 58
rect 496 24 500 58
rect 450 18 500 24
rect 1792 -452 1840 -444
rect 1792 -492 1838 -452
rect 1838 -492 1840 -452
rect 1792 -496 1840 -492
rect 292 -782 1632 -602
rect 1774 -754 1828 -688
<< metal1 >>
rect 122 970 1754 1008
rect 122 854 154 970
rect 1714 854 1754 970
rect 122 792 568 854
rect 1328 814 1754 854
rect 1328 792 1340 814
rect 122 786 1340 792
rect 122 784 672 786
rect 314 780 672 784
rect 314 486 348 780
rect 314 388 346 486
rect 502 444 720 486
rect 216 176 250 254
rect 408 176 442 254
rect 500 176 544 444
rect 680 374 720 444
rect 1120 360 1154 786
rect 1382 716 1468 730
rect 1382 672 1400 716
rect 1450 672 1468 716
rect 1382 654 1468 672
rect 1504 658 1538 814
rect 1278 398 1340 452
rect 584 176 624 276
rect 1120 272 1282 360
rect 776 176 816 272
rect 216 116 544 176
rect 216 114 250 116
rect 408 114 442 116
rect 500 112 544 116
rect 582 164 978 176
rect 582 108 924 164
rect 972 108 978 164
rect 582 102 978 108
rect 80 72 166 78
rect 80 10 92 72
rect 154 64 166 72
rect 438 64 514 70
rect 154 62 514 64
rect 154 24 450 62
rect 154 10 166 24
rect 80 4 166 10
rect 438 18 450 24
rect 500 18 514 62
rect 438 8 514 18
rect 916 -28 978 102
rect 400 -58 978 -28
rect 1342 70 1376 242
rect 1406 70 1446 654
rect 1504 510 1540 658
rect 1506 354 1540 510
rect 1608 398 1674 452
rect 1506 278 1610 354
rect 1506 276 1540 278
rect 1342 10 1446 70
rect 1666 56 1706 240
rect 402 -102 446 -58
rect 218 -438 248 -154
rect 602 -416 632 -152
rect 1164 -172 1272 -114
rect 1342 -166 1376 10
rect 1666 4 1846 56
rect 216 -458 248 -438
rect 216 -584 246 -458
rect 596 -584 634 -416
rect 1166 -436 1200 -172
rect 1544 -184 1612 -116
rect 1276 -264 1342 -206
rect 1162 -584 1200 -436
rect 1544 -454 1578 -184
rect 1666 -196 1706 4
rect 1608 -228 1674 -226
rect 1608 -280 1730 -228
rect 1542 -584 1580 -454
rect 216 -602 1670 -584
rect 216 -782 292 -602
rect 1632 -782 1670 -602
rect 1700 -688 1730 -280
rect 1792 -426 1842 4
rect 1782 -444 1848 -426
rect 1782 -496 1792 -444
rect 1840 -496 1848 -444
rect 1782 -510 1848 -496
rect 1768 -688 1834 -676
rect 1700 -754 1774 -688
rect 1828 -754 1834 -688
rect 1768 -766 1834 -754
rect 216 -798 1670 -782
rect 218 -810 1670 -798
rect 1542 -820 1580 -810
use sky130_fd_pr__pfet_01v8_5YQHKB  sky130_fd_pr__pfet_01v8_5YQHKB_0
timestamp 1615740176
transform 1 0 267 0 1 136
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_A66TXA  sky130_fd_pr__pfet_01v8_A66TXA_1
timestamp 1615743317
transform 1 0 1641 0 1 304
box -109 -188 109 154
use sky130_fd_pr__nfet_01v8_J6Z6BK  sky130_fd_pr__nfet_01v8_J6Z6BK_1
timestamp 1615743317
transform 1 0 1641 0 1 -182
box -73 -102 73 102
use sky130_fd_pr__nfet_01v8_J6Z6BK  sky130_fd_pr__nfet_01v8_J6Z6BK_0
timestamp 1615743317
transform 1 0 1309 0 1 -164
box -73 -102 73 102
use sky130_fd_pr__pfet_01v8_A66TXA  sky130_fd_pr__pfet_01v8_A66TXA_0
timestamp 1615743317
transform 1 0 1309 0 1 306
box -109 -188 109 154
use sky130_fd_pr__pfet_01v8_5A4GFE  sky130_fd_pr__pfet_01v8_5A4GFE_0
timestamp 1615743317
transform 1 0 329 0 1 326
box -253 -210 251 192
use sky130_fd_pr__pfet_01v8_5A4GFE  sky130_fd_pr__pfet_01v8_5A4GFE_1
timestamp 1615743317
transform 1 0 701 0 1 324
box -253 -210 251 192
use sky130_fd_pr__nfet_01v8_66KVP3  sky130_fd_pr__nfet_01v8_66KVP3_0
timestamp 1615743317
transform 1 0 425 0 1 -180
box -221 -116 221 118
<< labels >>
rlabel viali 924 108 972 164 1 Z
rlabel nwell 590 814 1298 930 1 vdd
rlabel viali 92 10 154 72 1 A
rlabel pwell 312 -730 1524 -622 1 vss
rlabel viali 1774 -754 1828 -688 1 vin
<< end >>
