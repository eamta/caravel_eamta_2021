magic
tech sky130A
magscale 1 2
timestamp 1615949206
<< metal1 >>
rect 2022 2721 2328 2732
rect 2022 2618 2043 2721
rect 2163 2618 2192 2721
rect 2312 2618 2328 2721
rect 2022 2488 2328 2618
rect 1812 2442 2538 2488
rect 1756 645 1804 2410
rect 1953 870 2000 2442
rect 2152 645 2200 2410
rect 2350 870 2397 2442
rect 2548 645 2596 2410
<< via1 >>
rect 2043 2618 2163 2721
rect 2192 2618 2312 2721
<< metal2 >>
rect 2043 2721 2163 2731
rect 2043 2608 2163 2618
rect 2192 2721 2312 2731
rect 2192 2608 2312 2618
use sky130_fd_pr__nfet_01v8_MXMZMC  sky130_fd_pr__nfet_01v8_MXMZMC_0
timestamp 1615949206
transform 1 0 2175 0 1 1671
box -563 -949 563 949
<< end >>
