magic
tech sky130A
magscale 1 2
timestamp 1615997521
<< nwell >>
rect -3517 -884 3517 884
<< pmoslvt >>
rect -3321 -664 -3111 736
rect -3053 -664 -2843 736
rect -2785 -664 -2575 736
rect -2517 -664 -2307 736
rect -2249 -664 -2039 736
rect -1981 -664 -1771 736
rect -1713 -664 -1503 736
rect -1445 -664 -1235 736
rect -1177 -664 -967 736
rect -909 -664 -699 736
rect -641 -664 -431 736
rect -373 -664 -163 736
rect -105 -664 105 736
rect 163 -664 373 736
rect 431 -664 641 736
rect 699 -664 909 736
rect 967 -664 1177 736
rect 1235 -664 1445 736
rect 1503 -664 1713 736
rect 1771 -664 1981 736
rect 2039 -664 2249 736
rect 2307 -664 2517 736
rect 2575 -664 2785 736
rect 2843 -664 3053 736
rect 3111 -664 3321 736
<< pdiff >>
rect -3379 724 -3321 736
rect -3379 -652 -3367 724
rect -3333 -652 -3321 724
rect -3379 -664 -3321 -652
rect -3111 724 -3053 736
rect -3111 -652 -3099 724
rect -3065 -652 -3053 724
rect -3111 -664 -3053 -652
rect -2843 724 -2785 736
rect -2843 -652 -2831 724
rect -2797 -652 -2785 724
rect -2843 -664 -2785 -652
rect -2575 724 -2517 736
rect -2575 -652 -2563 724
rect -2529 -652 -2517 724
rect -2575 -664 -2517 -652
rect -2307 724 -2249 736
rect -2307 -652 -2295 724
rect -2261 -652 -2249 724
rect -2307 -664 -2249 -652
rect -2039 724 -1981 736
rect -2039 -652 -2027 724
rect -1993 -652 -1981 724
rect -2039 -664 -1981 -652
rect -1771 724 -1713 736
rect -1771 -652 -1759 724
rect -1725 -652 -1713 724
rect -1771 -664 -1713 -652
rect -1503 724 -1445 736
rect -1503 -652 -1491 724
rect -1457 -652 -1445 724
rect -1503 -664 -1445 -652
rect -1235 724 -1177 736
rect -1235 -652 -1223 724
rect -1189 -652 -1177 724
rect -1235 -664 -1177 -652
rect -967 724 -909 736
rect -967 -652 -955 724
rect -921 -652 -909 724
rect -967 -664 -909 -652
rect -699 724 -641 736
rect -699 -652 -687 724
rect -653 -652 -641 724
rect -699 -664 -641 -652
rect -431 724 -373 736
rect -431 -652 -419 724
rect -385 -652 -373 724
rect -431 -664 -373 -652
rect -163 724 -105 736
rect -163 -652 -151 724
rect -117 -652 -105 724
rect -163 -664 -105 -652
rect 105 724 163 736
rect 105 -652 117 724
rect 151 -652 163 724
rect 105 -664 163 -652
rect 373 724 431 736
rect 373 -652 385 724
rect 419 -652 431 724
rect 373 -664 431 -652
rect 641 724 699 736
rect 641 -652 653 724
rect 687 -652 699 724
rect 641 -664 699 -652
rect 909 724 967 736
rect 909 -652 921 724
rect 955 -652 967 724
rect 909 -664 967 -652
rect 1177 724 1235 736
rect 1177 -652 1189 724
rect 1223 -652 1235 724
rect 1177 -664 1235 -652
rect 1445 724 1503 736
rect 1445 -652 1457 724
rect 1491 -652 1503 724
rect 1445 -664 1503 -652
rect 1713 724 1771 736
rect 1713 -652 1725 724
rect 1759 -652 1771 724
rect 1713 -664 1771 -652
rect 1981 724 2039 736
rect 1981 -652 1993 724
rect 2027 -652 2039 724
rect 1981 -664 2039 -652
rect 2249 724 2307 736
rect 2249 -652 2261 724
rect 2295 -652 2307 724
rect 2249 -664 2307 -652
rect 2517 724 2575 736
rect 2517 -652 2529 724
rect 2563 -652 2575 724
rect 2517 -664 2575 -652
rect 2785 724 2843 736
rect 2785 -652 2797 724
rect 2831 -652 2843 724
rect 2785 -664 2843 -652
rect 3053 724 3111 736
rect 3053 -652 3065 724
rect 3099 -652 3111 724
rect 3053 -664 3111 -652
rect 3321 724 3379 736
rect 3321 -652 3333 724
rect 3367 -652 3379 724
rect 3321 -664 3379 -652
<< pdiffc >>
rect -3367 -652 -3333 724
rect -3099 -652 -3065 724
rect -2831 -652 -2797 724
rect -2563 -652 -2529 724
rect -2295 -652 -2261 724
rect -2027 -652 -1993 724
rect -1759 -652 -1725 724
rect -1491 -652 -1457 724
rect -1223 -652 -1189 724
rect -955 -652 -921 724
rect -687 -652 -653 724
rect -419 -652 -385 724
rect -151 -652 -117 724
rect 117 -652 151 724
rect 385 -652 419 724
rect 653 -652 687 724
rect 921 -652 955 724
rect 1189 -652 1223 724
rect 1457 -652 1491 724
rect 1725 -652 1759 724
rect 1993 -652 2027 724
rect 2261 -652 2295 724
rect 2529 -652 2563 724
rect 2797 -652 2831 724
rect 3065 -652 3099 724
rect 3333 -652 3367 724
<< nsubdiff >>
rect -3481 814 -3385 848
rect 3385 814 3481 848
rect -3481 751 -3447 814
rect 3447 751 3481 814
rect -3481 -814 -3447 -751
rect 3447 -814 3481 -751
rect -3481 -848 -3385 -814
rect 3385 -848 3481 -814
<< nsubdiffcont >>
rect -3385 814 3385 848
rect -3481 -751 -3447 751
rect 3447 -751 3481 751
rect -3385 -848 3385 -814
<< poly >>
rect -3321 736 -3111 762
rect -3053 736 -2843 762
rect -2785 736 -2575 762
rect -2517 736 -2307 762
rect -2249 736 -2039 762
rect -1981 736 -1771 762
rect -1713 736 -1503 762
rect -1445 736 -1235 762
rect -1177 736 -967 762
rect -909 736 -699 762
rect -641 736 -431 762
rect -373 736 -163 762
rect -105 736 105 762
rect 163 736 373 762
rect 431 736 641 762
rect 699 736 909 762
rect 967 736 1177 762
rect 1235 736 1445 762
rect 1503 736 1713 762
rect 1771 736 1981 762
rect 2039 736 2249 762
rect 2307 736 2517 762
rect 2575 736 2785 762
rect 2843 736 3053 762
rect 3111 736 3321 762
rect -3321 -711 -3111 -664
rect -3321 -745 -3305 -711
rect -3127 -745 -3111 -711
rect -3321 -761 -3111 -745
rect -3053 -711 -2843 -664
rect -3053 -745 -3037 -711
rect -2859 -745 -2843 -711
rect -3053 -761 -2843 -745
rect -2785 -711 -2575 -664
rect -2785 -745 -2769 -711
rect -2591 -745 -2575 -711
rect -2785 -761 -2575 -745
rect -2517 -711 -2307 -664
rect -2517 -745 -2501 -711
rect -2323 -745 -2307 -711
rect -2517 -761 -2307 -745
rect -2249 -711 -2039 -664
rect -2249 -745 -2233 -711
rect -2055 -745 -2039 -711
rect -2249 -761 -2039 -745
rect -1981 -711 -1771 -664
rect -1981 -745 -1965 -711
rect -1787 -745 -1771 -711
rect -1981 -761 -1771 -745
rect -1713 -711 -1503 -664
rect -1713 -745 -1697 -711
rect -1519 -745 -1503 -711
rect -1713 -761 -1503 -745
rect -1445 -711 -1235 -664
rect -1445 -745 -1429 -711
rect -1251 -745 -1235 -711
rect -1445 -761 -1235 -745
rect -1177 -711 -967 -664
rect -1177 -745 -1161 -711
rect -983 -745 -967 -711
rect -1177 -761 -967 -745
rect -909 -711 -699 -664
rect -909 -745 -893 -711
rect -715 -745 -699 -711
rect -909 -761 -699 -745
rect -641 -711 -431 -664
rect -641 -745 -625 -711
rect -447 -745 -431 -711
rect -641 -761 -431 -745
rect -373 -711 -163 -664
rect -373 -745 -357 -711
rect -179 -745 -163 -711
rect -373 -761 -163 -745
rect -105 -711 105 -664
rect -105 -745 -89 -711
rect 89 -745 105 -711
rect -105 -761 105 -745
rect 163 -711 373 -664
rect 163 -745 179 -711
rect 357 -745 373 -711
rect 163 -761 373 -745
rect 431 -711 641 -664
rect 431 -745 447 -711
rect 625 -745 641 -711
rect 431 -761 641 -745
rect 699 -711 909 -664
rect 699 -745 715 -711
rect 893 -745 909 -711
rect 699 -761 909 -745
rect 967 -711 1177 -664
rect 967 -745 983 -711
rect 1161 -745 1177 -711
rect 967 -761 1177 -745
rect 1235 -711 1445 -664
rect 1235 -745 1251 -711
rect 1429 -745 1445 -711
rect 1235 -761 1445 -745
rect 1503 -711 1713 -664
rect 1503 -745 1519 -711
rect 1697 -745 1713 -711
rect 1503 -761 1713 -745
rect 1771 -711 1981 -664
rect 1771 -745 1787 -711
rect 1965 -745 1981 -711
rect 1771 -761 1981 -745
rect 2039 -711 2249 -664
rect 2039 -745 2055 -711
rect 2233 -745 2249 -711
rect 2039 -761 2249 -745
rect 2307 -711 2517 -664
rect 2307 -745 2323 -711
rect 2501 -745 2517 -711
rect 2307 -761 2517 -745
rect 2575 -711 2785 -664
rect 2575 -745 2591 -711
rect 2769 -745 2785 -711
rect 2575 -761 2785 -745
rect 2843 -711 3053 -664
rect 2843 -745 2859 -711
rect 3037 -745 3053 -711
rect 2843 -761 3053 -745
rect 3111 -711 3321 -664
rect 3111 -745 3127 -711
rect 3305 -745 3321 -711
rect 3111 -761 3321 -745
<< polycont >>
rect -3305 -745 -3127 -711
rect -3037 -745 -2859 -711
rect -2769 -745 -2591 -711
rect -2501 -745 -2323 -711
rect -2233 -745 -2055 -711
rect -1965 -745 -1787 -711
rect -1697 -745 -1519 -711
rect -1429 -745 -1251 -711
rect -1161 -745 -983 -711
rect -893 -745 -715 -711
rect -625 -745 -447 -711
rect -357 -745 -179 -711
rect -89 -745 89 -711
rect 179 -745 357 -711
rect 447 -745 625 -711
rect 715 -745 893 -711
rect 983 -745 1161 -711
rect 1251 -745 1429 -711
rect 1519 -745 1697 -711
rect 1787 -745 1965 -711
rect 2055 -745 2233 -711
rect 2323 -745 2501 -711
rect 2591 -745 2769 -711
rect 2859 -745 3037 -711
rect 3127 -745 3305 -711
<< locali >>
rect -3481 814 -3385 848
rect 3385 814 3481 848
rect -3481 751 -3447 814
rect 3447 751 3481 814
rect -3367 724 -3333 740
rect -3367 -668 -3333 -652
rect -3099 724 -3065 740
rect -3099 -668 -3065 -652
rect -2831 724 -2797 740
rect -2831 -668 -2797 -652
rect -2563 724 -2529 740
rect -2563 -668 -2529 -652
rect -2295 724 -2261 740
rect -2295 -668 -2261 -652
rect -2027 724 -1993 740
rect -2027 -668 -1993 -652
rect -1759 724 -1725 740
rect -1759 -668 -1725 -652
rect -1491 724 -1457 740
rect -1491 -668 -1457 -652
rect -1223 724 -1189 740
rect -1223 -668 -1189 -652
rect -955 724 -921 740
rect -955 -668 -921 -652
rect -687 724 -653 740
rect -687 -668 -653 -652
rect -419 724 -385 740
rect -419 -668 -385 -652
rect -151 724 -117 740
rect -151 -668 -117 -652
rect 117 724 151 740
rect 117 -668 151 -652
rect 385 724 419 740
rect 385 -668 419 -652
rect 653 724 687 740
rect 653 -668 687 -652
rect 921 724 955 740
rect 921 -668 955 -652
rect 1189 724 1223 740
rect 1189 -668 1223 -652
rect 1457 724 1491 740
rect 1457 -668 1491 -652
rect 1725 724 1759 740
rect 1725 -668 1759 -652
rect 1993 724 2027 740
rect 1993 -668 2027 -652
rect 2261 724 2295 740
rect 2261 -668 2295 -652
rect 2529 724 2563 740
rect 2529 -668 2563 -652
rect 2797 724 2831 740
rect 2797 -668 2831 -652
rect 3065 724 3099 740
rect 3065 -668 3099 -652
rect 3333 724 3367 740
rect 3333 -668 3367 -652
rect -3321 -745 -3305 -711
rect -3127 -745 -3111 -711
rect -3053 -745 -3037 -711
rect -2859 -745 -2843 -711
rect -2785 -745 -2769 -711
rect -2591 -745 -2575 -711
rect -2517 -745 -2501 -711
rect -2323 -745 -2307 -711
rect -2249 -745 -2233 -711
rect -2055 -745 -2039 -711
rect -1981 -745 -1965 -711
rect -1787 -745 -1771 -711
rect -1713 -745 -1697 -711
rect -1519 -745 -1503 -711
rect -1445 -745 -1429 -711
rect -1251 -745 -1235 -711
rect -1177 -745 -1161 -711
rect -983 -745 -967 -711
rect -909 -745 -893 -711
rect -715 -745 -699 -711
rect -641 -745 -625 -711
rect -447 -745 -431 -711
rect -373 -745 -357 -711
rect -179 -745 -163 -711
rect -105 -745 -89 -711
rect 89 -745 105 -711
rect 163 -745 179 -711
rect 357 -745 373 -711
rect 431 -745 447 -711
rect 625 -745 641 -711
rect 699 -745 715 -711
rect 893 -745 909 -711
rect 967 -745 983 -711
rect 1161 -745 1177 -711
rect 1235 -745 1251 -711
rect 1429 -745 1445 -711
rect 1503 -745 1519 -711
rect 1697 -745 1713 -711
rect 1771 -745 1787 -711
rect 1965 -745 1981 -711
rect 2039 -745 2055 -711
rect 2233 -745 2249 -711
rect 2307 -745 2323 -711
rect 2501 -745 2517 -711
rect 2575 -745 2591 -711
rect 2769 -745 2785 -711
rect 2843 -745 2859 -711
rect 3037 -745 3053 -711
rect 3111 -745 3127 -711
rect 3305 -745 3321 -711
rect -3481 -814 -3447 -751
rect 3447 -814 3481 -751
rect -3481 -848 -3385 -814
rect 3385 -848 3481 -814
<< viali >>
rect -3367 -652 -3333 724
rect -3099 -652 -3065 724
rect -2831 -652 -2797 724
rect -2563 -652 -2529 724
rect -2295 -652 -2261 724
rect -2027 -652 -1993 724
rect -1759 -652 -1725 724
rect -1491 -652 -1457 724
rect -1223 -652 -1189 724
rect -955 -652 -921 724
rect -687 -652 -653 724
rect -419 -652 -385 724
rect -151 -652 -117 724
rect 117 -652 151 724
rect 385 -652 419 724
rect 653 -652 687 724
rect 921 -652 955 724
rect 1189 -652 1223 724
rect 1457 -652 1491 724
rect 1725 -652 1759 724
rect 1993 -652 2027 724
rect 2261 -652 2295 724
rect 2529 -652 2563 724
rect 2797 -652 2831 724
rect 3065 -652 3099 724
rect 3333 -652 3367 724
rect -3305 -745 -3127 -711
rect -3037 -745 -2859 -711
rect -2769 -745 -2591 -711
rect -2501 -745 -2323 -711
rect -2233 -745 -2055 -711
rect -1965 -745 -1787 -711
rect -1697 -745 -1519 -711
rect -1429 -745 -1251 -711
rect -1161 -745 -983 -711
rect -893 -745 -715 -711
rect -625 -745 -447 -711
rect -357 -745 -179 -711
rect -89 -745 89 -711
rect 179 -745 357 -711
rect 447 -745 625 -711
rect 715 -745 893 -711
rect 983 -745 1161 -711
rect 1251 -745 1429 -711
rect 1519 -745 1697 -711
rect 1787 -745 1965 -711
rect 2055 -745 2233 -711
rect 2323 -745 2501 -711
rect 2591 -745 2769 -711
rect 2859 -745 3037 -711
rect 3127 -745 3305 -711
<< metal1 >>
rect -3373 724 -3327 736
rect -3373 -652 -3367 724
rect -3333 -652 -3327 724
rect -3373 -664 -3327 -652
rect -3105 724 -3059 736
rect -3105 -652 -3099 724
rect -3065 -652 -3059 724
rect -3105 -664 -3059 -652
rect -2837 724 -2791 736
rect -2837 -652 -2831 724
rect -2797 -652 -2791 724
rect -2837 -664 -2791 -652
rect -2569 724 -2523 736
rect -2569 -652 -2563 724
rect -2529 -652 -2523 724
rect -2569 -664 -2523 -652
rect -2301 724 -2255 736
rect -2301 -652 -2295 724
rect -2261 -652 -2255 724
rect -2301 -664 -2255 -652
rect -2033 724 -1987 736
rect -2033 -652 -2027 724
rect -1993 -652 -1987 724
rect -2033 -664 -1987 -652
rect -1765 724 -1719 736
rect -1765 -652 -1759 724
rect -1725 -652 -1719 724
rect -1765 -664 -1719 -652
rect -1497 724 -1451 736
rect -1497 -652 -1491 724
rect -1457 -652 -1451 724
rect -1497 -664 -1451 -652
rect -1229 724 -1183 736
rect -1229 -652 -1223 724
rect -1189 -652 -1183 724
rect -1229 -664 -1183 -652
rect -961 724 -915 736
rect -961 -652 -955 724
rect -921 -652 -915 724
rect -961 -664 -915 -652
rect -693 724 -647 736
rect -693 -652 -687 724
rect -653 -652 -647 724
rect -693 -664 -647 -652
rect -425 724 -379 736
rect -425 -652 -419 724
rect -385 -652 -379 724
rect -425 -664 -379 -652
rect -157 724 -111 736
rect -157 -652 -151 724
rect -117 -652 -111 724
rect -157 -664 -111 -652
rect 111 724 157 736
rect 111 -652 117 724
rect 151 -652 157 724
rect 111 -664 157 -652
rect 379 724 425 736
rect 379 -652 385 724
rect 419 -652 425 724
rect 379 -664 425 -652
rect 647 724 693 736
rect 647 -652 653 724
rect 687 -652 693 724
rect 647 -664 693 -652
rect 915 724 961 736
rect 915 -652 921 724
rect 955 -652 961 724
rect 915 -664 961 -652
rect 1183 724 1229 736
rect 1183 -652 1189 724
rect 1223 -652 1229 724
rect 1183 -664 1229 -652
rect 1451 724 1497 736
rect 1451 -652 1457 724
rect 1491 -652 1497 724
rect 1451 -664 1497 -652
rect 1719 724 1765 736
rect 1719 -652 1725 724
rect 1759 -652 1765 724
rect 1719 -664 1765 -652
rect 1987 724 2033 736
rect 1987 -652 1993 724
rect 2027 -652 2033 724
rect 1987 -664 2033 -652
rect 2255 724 2301 736
rect 2255 -652 2261 724
rect 2295 -652 2301 724
rect 2255 -664 2301 -652
rect 2523 724 2569 736
rect 2523 -652 2529 724
rect 2563 -652 2569 724
rect 2523 -664 2569 -652
rect 2791 724 2837 736
rect 2791 -652 2797 724
rect 2831 -652 2837 724
rect 2791 -664 2837 -652
rect 3059 724 3105 736
rect 3059 -652 3065 724
rect 3099 -652 3105 724
rect 3059 -664 3105 -652
rect 3327 724 3373 736
rect 3327 -652 3333 724
rect 3367 -652 3373 724
rect 3327 -664 3373 -652
rect -3317 -711 -3115 -705
rect -3317 -745 -3305 -711
rect -3127 -745 -3115 -711
rect -3317 -751 -3115 -745
rect -3049 -711 -2847 -705
rect -3049 -745 -3037 -711
rect -2859 -745 -2847 -711
rect -3049 -751 -2847 -745
rect -2781 -711 -2579 -705
rect -2781 -745 -2769 -711
rect -2591 -745 -2579 -711
rect -2781 -751 -2579 -745
rect -2513 -711 -2311 -705
rect -2513 -745 -2501 -711
rect -2323 -745 -2311 -711
rect -2513 -751 -2311 -745
rect -2245 -711 -2043 -705
rect -2245 -745 -2233 -711
rect -2055 -745 -2043 -711
rect -2245 -751 -2043 -745
rect -1977 -711 -1775 -705
rect -1977 -745 -1965 -711
rect -1787 -745 -1775 -711
rect -1977 -751 -1775 -745
rect -1709 -711 -1507 -705
rect -1709 -745 -1697 -711
rect -1519 -745 -1507 -711
rect -1709 -751 -1507 -745
rect -1441 -711 -1239 -705
rect -1441 -745 -1429 -711
rect -1251 -745 -1239 -711
rect -1441 -751 -1239 -745
rect -1173 -711 -971 -705
rect -1173 -745 -1161 -711
rect -983 -745 -971 -711
rect -1173 -751 -971 -745
rect -905 -711 -703 -705
rect -905 -745 -893 -711
rect -715 -745 -703 -711
rect -905 -751 -703 -745
rect -637 -711 -435 -705
rect -637 -745 -625 -711
rect -447 -745 -435 -711
rect -637 -751 -435 -745
rect -369 -711 -167 -705
rect -369 -745 -357 -711
rect -179 -745 -167 -711
rect -369 -751 -167 -745
rect -101 -711 101 -705
rect -101 -745 -89 -711
rect 89 -745 101 -711
rect -101 -751 101 -745
rect 167 -711 369 -705
rect 167 -745 179 -711
rect 357 -745 369 -711
rect 167 -751 369 -745
rect 435 -711 637 -705
rect 435 -745 447 -711
rect 625 -745 637 -711
rect 435 -751 637 -745
rect 703 -711 905 -705
rect 703 -745 715 -711
rect 893 -745 905 -711
rect 703 -751 905 -745
rect 971 -711 1173 -705
rect 971 -745 983 -711
rect 1161 -745 1173 -711
rect 971 -751 1173 -745
rect 1239 -711 1441 -705
rect 1239 -745 1251 -711
rect 1429 -745 1441 -711
rect 1239 -751 1441 -745
rect 1507 -711 1709 -705
rect 1507 -745 1519 -711
rect 1697 -745 1709 -711
rect 1507 -751 1709 -745
rect 1775 -711 1977 -705
rect 1775 -745 1787 -711
rect 1965 -745 1977 -711
rect 1775 -751 1977 -745
rect 2043 -711 2245 -705
rect 2043 -745 2055 -711
rect 2233 -745 2245 -711
rect 2043 -751 2245 -745
rect 2311 -711 2513 -705
rect 2311 -745 2323 -711
rect 2501 -745 2513 -711
rect 2311 -751 2513 -745
rect 2579 -711 2781 -705
rect 2579 -745 2591 -711
rect 2769 -745 2781 -711
rect 2579 -751 2781 -745
rect 2847 -711 3049 -705
rect 2847 -745 2859 -711
rect 3037 -745 3049 -711
rect 2847 -751 3049 -745
rect 3115 -711 3317 -705
rect 3115 -745 3127 -711
rect 3305 -745 3317 -711
rect 3115 -751 3317 -745
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -3464 -831 3464 831
string parameters w 7 l 1.05 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
