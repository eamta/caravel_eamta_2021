magic
tech sky130A
magscale 1 2
timestamp 1622937437
<< error_p >>
rect -845 1947 -787 1953
rect -653 1947 -595 1953
rect -461 1947 -403 1953
rect -269 1947 -211 1953
rect -77 1947 -19 1953
rect 115 1947 173 1953
rect 307 1947 365 1953
rect 499 1947 557 1953
rect 691 1947 749 1953
rect 883 1947 941 1953
rect -845 1913 -833 1947
rect -653 1913 -641 1947
rect -461 1913 -449 1947
rect -269 1913 -257 1947
rect -77 1913 -65 1947
rect 115 1913 127 1947
rect 307 1913 319 1947
rect 499 1913 511 1947
rect 691 1913 703 1947
rect 883 1913 895 1947
rect -845 1907 -787 1913
rect -653 1907 -595 1913
rect -461 1907 -403 1913
rect -269 1907 -211 1913
rect -77 1907 -19 1913
rect 115 1907 173 1913
rect 307 1907 365 1913
rect 499 1907 557 1913
rect 691 1907 749 1913
rect 883 1907 941 1913
rect -941 -1913 -883 -1907
rect -749 -1913 -691 -1907
rect -557 -1913 -499 -1907
rect -365 -1913 -307 -1907
rect -173 -1913 -115 -1907
rect 19 -1913 77 -1907
rect 211 -1913 269 -1907
rect 403 -1913 461 -1907
rect 595 -1913 653 -1907
rect 787 -1913 845 -1907
rect -941 -1947 -929 -1913
rect -749 -1947 -737 -1913
rect -557 -1947 -545 -1913
rect -365 -1947 -353 -1913
rect -173 -1947 -161 -1913
rect 19 -1947 31 -1913
rect 211 -1947 223 -1913
rect 403 -1947 415 -1913
rect 595 -1947 607 -1913
rect 787 -1947 799 -1913
rect -941 -1953 -883 -1947
rect -749 -1953 -691 -1947
rect -557 -1953 -499 -1947
rect -365 -1953 -307 -1947
rect -173 -1953 -115 -1947
rect 19 -1953 77 -1947
rect 211 -1953 269 -1947
rect 403 -1953 461 -1947
rect 595 -1953 653 -1947
rect 787 -1953 845 -1947
<< pwell >>
rect -1127 -2085 1127 2085
<< nmos >>
rect -927 -1875 -897 1875
rect -831 -1875 -801 1875
rect -735 -1875 -705 1875
rect -639 -1875 -609 1875
rect -543 -1875 -513 1875
rect -447 -1875 -417 1875
rect -351 -1875 -321 1875
rect -255 -1875 -225 1875
rect -159 -1875 -129 1875
rect -63 -1875 -33 1875
rect 33 -1875 63 1875
rect 129 -1875 159 1875
rect 225 -1875 255 1875
rect 321 -1875 351 1875
rect 417 -1875 447 1875
rect 513 -1875 543 1875
rect 609 -1875 639 1875
rect 705 -1875 735 1875
rect 801 -1875 831 1875
rect 897 -1875 927 1875
<< ndiff >>
rect -989 1863 -927 1875
rect -989 -1863 -977 1863
rect -943 -1863 -927 1863
rect -989 -1875 -927 -1863
rect -897 1863 -831 1875
rect -897 -1863 -881 1863
rect -847 -1863 -831 1863
rect -897 -1875 -831 -1863
rect -801 1863 -735 1875
rect -801 -1863 -785 1863
rect -751 -1863 -735 1863
rect -801 -1875 -735 -1863
rect -705 1863 -639 1875
rect -705 -1863 -689 1863
rect -655 -1863 -639 1863
rect -705 -1875 -639 -1863
rect -609 1863 -543 1875
rect -609 -1863 -593 1863
rect -559 -1863 -543 1863
rect -609 -1875 -543 -1863
rect -513 1863 -447 1875
rect -513 -1863 -497 1863
rect -463 -1863 -447 1863
rect -513 -1875 -447 -1863
rect -417 1863 -351 1875
rect -417 -1863 -401 1863
rect -367 -1863 -351 1863
rect -417 -1875 -351 -1863
rect -321 1863 -255 1875
rect -321 -1863 -305 1863
rect -271 -1863 -255 1863
rect -321 -1875 -255 -1863
rect -225 1863 -159 1875
rect -225 -1863 -209 1863
rect -175 -1863 -159 1863
rect -225 -1875 -159 -1863
rect -129 1863 -63 1875
rect -129 -1863 -113 1863
rect -79 -1863 -63 1863
rect -129 -1875 -63 -1863
rect -33 1863 33 1875
rect -33 -1863 -17 1863
rect 17 -1863 33 1863
rect -33 -1875 33 -1863
rect 63 1863 129 1875
rect 63 -1863 79 1863
rect 113 -1863 129 1863
rect 63 -1875 129 -1863
rect 159 1863 225 1875
rect 159 -1863 175 1863
rect 209 -1863 225 1863
rect 159 -1875 225 -1863
rect 255 1863 321 1875
rect 255 -1863 271 1863
rect 305 -1863 321 1863
rect 255 -1875 321 -1863
rect 351 1863 417 1875
rect 351 -1863 367 1863
rect 401 -1863 417 1863
rect 351 -1875 417 -1863
rect 447 1863 513 1875
rect 447 -1863 463 1863
rect 497 -1863 513 1863
rect 447 -1875 513 -1863
rect 543 1863 609 1875
rect 543 -1863 559 1863
rect 593 -1863 609 1863
rect 543 -1875 609 -1863
rect 639 1863 705 1875
rect 639 -1863 655 1863
rect 689 -1863 705 1863
rect 639 -1875 705 -1863
rect 735 1863 801 1875
rect 735 -1863 751 1863
rect 785 -1863 801 1863
rect 735 -1875 801 -1863
rect 831 1863 897 1875
rect 831 -1863 847 1863
rect 881 -1863 897 1863
rect 831 -1875 897 -1863
rect 927 1863 989 1875
rect 927 -1863 943 1863
rect 977 -1863 989 1863
rect 927 -1875 989 -1863
<< ndiffc >>
rect -977 -1863 -943 1863
rect -881 -1863 -847 1863
rect -785 -1863 -751 1863
rect -689 -1863 -655 1863
rect -593 -1863 -559 1863
rect -497 -1863 -463 1863
rect -401 -1863 -367 1863
rect -305 -1863 -271 1863
rect -209 -1863 -175 1863
rect -113 -1863 -79 1863
rect -17 -1863 17 1863
rect 79 -1863 113 1863
rect 175 -1863 209 1863
rect 271 -1863 305 1863
rect 367 -1863 401 1863
rect 463 -1863 497 1863
rect 559 -1863 593 1863
rect 655 -1863 689 1863
rect 751 -1863 785 1863
rect 847 -1863 881 1863
rect 943 -1863 977 1863
<< psubdiff >>
rect -1091 2015 -995 2049
rect 995 2015 1091 2049
rect -1091 1953 -1057 2015
rect 1057 1953 1091 2015
rect -1091 -2015 -1057 -1953
rect 1057 -2015 1091 -1953
rect -1091 -2049 -995 -2015
rect 995 -2049 1091 -2015
<< psubdiffcont >>
rect -995 2015 995 2049
rect -1091 -1953 -1057 1953
rect 1057 -1953 1091 1953
rect -995 -2049 995 -2015
<< poly >>
rect -849 1947 -783 1963
rect -849 1913 -833 1947
rect -799 1913 -783 1947
rect -927 1875 -897 1901
rect -849 1897 -783 1913
rect -657 1947 -591 1963
rect -657 1913 -641 1947
rect -607 1913 -591 1947
rect -831 1875 -801 1897
rect -735 1875 -705 1901
rect -657 1897 -591 1913
rect -465 1947 -399 1963
rect -465 1913 -449 1947
rect -415 1913 -399 1947
rect -639 1875 -609 1897
rect -543 1875 -513 1901
rect -465 1897 -399 1913
rect -273 1947 -207 1963
rect -273 1913 -257 1947
rect -223 1913 -207 1947
rect -447 1875 -417 1897
rect -351 1875 -321 1901
rect -273 1897 -207 1913
rect -81 1947 -15 1963
rect -81 1913 -65 1947
rect -31 1913 -15 1947
rect -255 1875 -225 1897
rect -159 1875 -129 1901
rect -81 1897 -15 1913
rect 111 1947 177 1963
rect 111 1913 127 1947
rect 161 1913 177 1947
rect -63 1875 -33 1897
rect 33 1875 63 1901
rect 111 1897 177 1913
rect 303 1947 369 1963
rect 303 1913 319 1947
rect 353 1913 369 1947
rect 129 1875 159 1897
rect 225 1875 255 1901
rect 303 1897 369 1913
rect 495 1947 561 1963
rect 495 1913 511 1947
rect 545 1913 561 1947
rect 321 1875 351 1897
rect 417 1875 447 1901
rect 495 1897 561 1913
rect 687 1947 753 1963
rect 687 1913 703 1947
rect 737 1913 753 1947
rect 513 1875 543 1897
rect 609 1875 639 1901
rect 687 1897 753 1913
rect 879 1947 945 1963
rect 879 1913 895 1947
rect 929 1913 945 1947
rect 705 1875 735 1897
rect 801 1875 831 1901
rect 879 1897 945 1913
rect 897 1875 927 1897
rect -927 -1897 -897 -1875
rect -945 -1913 -879 -1897
rect -831 -1901 -801 -1875
rect -735 -1897 -705 -1875
rect -945 -1947 -929 -1913
rect -895 -1947 -879 -1913
rect -945 -1963 -879 -1947
rect -753 -1913 -687 -1897
rect -639 -1901 -609 -1875
rect -543 -1897 -513 -1875
rect -753 -1947 -737 -1913
rect -703 -1947 -687 -1913
rect -753 -1963 -687 -1947
rect -561 -1913 -495 -1897
rect -447 -1901 -417 -1875
rect -351 -1897 -321 -1875
rect -561 -1947 -545 -1913
rect -511 -1947 -495 -1913
rect -561 -1963 -495 -1947
rect -369 -1913 -303 -1897
rect -255 -1901 -225 -1875
rect -159 -1897 -129 -1875
rect -369 -1947 -353 -1913
rect -319 -1947 -303 -1913
rect -369 -1963 -303 -1947
rect -177 -1913 -111 -1897
rect -63 -1901 -33 -1875
rect 33 -1897 63 -1875
rect -177 -1947 -161 -1913
rect -127 -1947 -111 -1913
rect -177 -1963 -111 -1947
rect 15 -1913 81 -1897
rect 129 -1901 159 -1875
rect 225 -1897 255 -1875
rect 15 -1947 31 -1913
rect 65 -1947 81 -1913
rect 15 -1963 81 -1947
rect 207 -1913 273 -1897
rect 321 -1901 351 -1875
rect 417 -1897 447 -1875
rect 207 -1947 223 -1913
rect 257 -1947 273 -1913
rect 207 -1963 273 -1947
rect 399 -1913 465 -1897
rect 513 -1901 543 -1875
rect 609 -1897 639 -1875
rect 399 -1947 415 -1913
rect 449 -1947 465 -1913
rect 399 -1963 465 -1947
rect 591 -1913 657 -1897
rect 705 -1901 735 -1875
rect 801 -1897 831 -1875
rect 591 -1947 607 -1913
rect 641 -1947 657 -1913
rect 591 -1963 657 -1947
rect 783 -1913 849 -1897
rect 897 -1901 927 -1875
rect 783 -1947 799 -1913
rect 833 -1947 849 -1913
rect 783 -1963 849 -1947
<< polycont >>
rect -833 1913 -799 1947
rect -641 1913 -607 1947
rect -449 1913 -415 1947
rect -257 1913 -223 1947
rect -65 1913 -31 1947
rect 127 1913 161 1947
rect 319 1913 353 1947
rect 511 1913 545 1947
rect 703 1913 737 1947
rect 895 1913 929 1947
rect -929 -1947 -895 -1913
rect -737 -1947 -703 -1913
rect -545 -1947 -511 -1913
rect -353 -1947 -319 -1913
rect -161 -1947 -127 -1913
rect 31 -1947 65 -1913
rect 223 -1947 257 -1913
rect 415 -1947 449 -1913
rect 607 -1947 641 -1913
rect 799 -1947 833 -1913
<< locali >>
rect -1091 2015 -995 2049
rect 995 2015 1091 2049
rect -1091 1953 -1057 2015
rect 1057 1953 1091 2015
rect -849 1913 -833 1947
rect -799 1913 -783 1947
rect -657 1913 -641 1947
rect -607 1913 -591 1947
rect -465 1913 -449 1947
rect -415 1913 -399 1947
rect -273 1913 -257 1947
rect -223 1913 -207 1947
rect -81 1913 -65 1947
rect -31 1913 -15 1947
rect 111 1913 127 1947
rect 161 1913 177 1947
rect 303 1913 319 1947
rect 353 1913 369 1947
rect 495 1913 511 1947
rect 545 1913 561 1947
rect 687 1913 703 1947
rect 737 1913 753 1947
rect 879 1913 895 1947
rect 929 1913 945 1947
rect -977 1863 -943 1879
rect -977 -1879 -943 -1863
rect -881 1863 -847 1879
rect -881 -1879 -847 -1863
rect -785 1863 -751 1879
rect -785 -1879 -751 -1863
rect -689 1863 -655 1879
rect -689 -1879 -655 -1863
rect -593 1863 -559 1879
rect -593 -1879 -559 -1863
rect -497 1863 -463 1879
rect -497 -1879 -463 -1863
rect -401 1863 -367 1879
rect -401 -1879 -367 -1863
rect -305 1863 -271 1879
rect -305 -1879 -271 -1863
rect -209 1863 -175 1879
rect -209 -1879 -175 -1863
rect -113 1863 -79 1879
rect -113 -1879 -79 -1863
rect -17 1863 17 1879
rect -17 -1879 17 -1863
rect 79 1863 113 1879
rect 79 -1879 113 -1863
rect 175 1863 209 1879
rect 175 -1879 209 -1863
rect 271 1863 305 1879
rect 271 -1879 305 -1863
rect 367 1863 401 1879
rect 367 -1879 401 -1863
rect 463 1863 497 1879
rect 463 -1879 497 -1863
rect 559 1863 593 1879
rect 559 -1879 593 -1863
rect 655 1863 689 1879
rect 655 -1879 689 -1863
rect 751 1863 785 1879
rect 751 -1879 785 -1863
rect 847 1863 881 1879
rect 847 -1879 881 -1863
rect 943 1863 977 1879
rect 943 -1879 977 -1863
rect -945 -1947 -929 -1913
rect -895 -1947 -879 -1913
rect -753 -1947 -737 -1913
rect -703 -1947 -687 -1913
rect -561 -1947 -545 -1913
rect -511 -1947 -495 -1913
rect -369 -1947 -353 -1913
rect -319 -1947 -303 -1913
rect -177 -1947 -161 -1913
rect -127 -1947 -111 -1913
rect 15 -1947 31 -1913
rect 65 -1947 81 -1913
rect 207 -1947 223 -1913
rect 257 -1947 273 -1913
rect 399 -1947 415 -1913
rect 449 -1947 465 -1913
rect 591 -1947 607 -1913
rect 641 -1947 657 -1913
rect 783 -1947 799 -1913
rect 833 -1947 849 -1913
rect -1091 -2015 -1057 -1953
rect 1057 -2015 1091 -1953
rect -1091 -2049 -995 -2015
rect 995 -2049 1091 -2015
<< viali >>
rect -833 1913 -799 1947
rect -641 1913 -607 1947
rect -449 1913 -415 1947
rect -257 1913 -223 1947
rect -65 1913 -31 1947
rect 127 1913 161 1947
rect 319 1913 353 1947
rect 511 1913 545 1947
rect 703 1913 737 1947
rect 895 1913 929 1947
rect -977 -1863 -943 1863
rect -881 -1863 -847 1863
rect -785 -1863 -751 1863
rect -689 -1863 -655 1863
rect -593 -1863 -559 1863
rect -497 -1863 -463 1863
rect -401 -1863 -367 1863
rect -305 -1863 -271 1863
rect -209 -1863 -175 1863
rect -113 -1863 -79 1863
rect -17 -1863 17 1863
rect 79 -1863 113 1863
rect 175 -1863 209 1863
rect 271 -1863 305 1863
rect 367 -1863 401 1863
rect 463 -1863 497 1863
rect 559 -1863 593 1863
rect 655 -1863 689 1863
rect 751 -1863 785 1863
rect 847 -1863 881 1863
rect 943 -1863 977 1863
rect -929 -1947 -895 -1913
rect -737 -1947 -703 -1913
rect -545 -1947 -511 -1913
rect -353 -1947 -319 -1913
rect -161 -1947 -127 -1913
rect 31 -1947 65 -1913
rect 223 -1947 257 -1913
rect 415 -1947 449 -1913
rect 607 -1947 641 -1913
rect 799 -1947 833 -1913
<< metal1 >>
rect -845 1947 -787 1953
rect -845 1913 -833 1947
rect -799 1913 -787 1947
rect -845 1907 -787 1913
rect -653 1947 -595 1953
rect -653 1913 -641 1947
rect -607 1913 -595 1947
rect -653 1907 -595 1913
rect -461 1947 -403 1953
rect -461 1913 -449 1947
rect -415 1913 -403 1947
rect -461 1907 -403 1913
rect -269 1947 -211 1953
rect -269 1913 -257 1947
rect -223 1913 -211 1947
rect -269 1907 -211 1913
rect -77 1947 -19 1953
rect -77 1913 -65 1947
rect -31 1913 -19 1947
rect -77 1907 -19 1913
rect 115 1947 173 1953
rect 115 1913 127 1947
rect 161 1913 173 1947
rect 115 1907 173 1913
rect 307 1947 365 1953
rect 307 1913 319 1947
rect 353 1913 365 1947
rect 307 1907 365 1913
rect 499 1947 557 1953
rect 499 1913 511 1947
rect 545 1913 557 1947
rect 499 1907 557 1913
rect 691 1947 749 1953
rect 691 1913 703 1947
rect 737 1913 749 1947
rect 691 1907 749 1913
rect 883 1947 941 1953
rect 883 1913 895 1947
rect 929 1913 941 1947
rect 883 1907 941 1913
rect -983 1863 -937 1875
rect -983 -1863 -977 1863
rect -943 -1863 -937 1863
rect -983 -1875 -937 -1863
rect -887 1863 -841 1875
rect -887 -1863 -881 1863
rect -847 -1863 -841 1863
rect -887 -1875 -841 -1863
rect -791 1863 -745 1875
rect -791 -1863 -785 1863
rect -751 -1863 -745 1863
rect -791 -1875 -745 -1863
rect -695 1863 -649 1875
rect -695 -1863 -689 1863
rect -655 -1863 -649 1863
rect -695 -1875 -649 -1863
rect -599 1863 -553 1875
rect -599 -1863 -593 1863
rect -559 -1863 -553 1863
rect -599 -1875 -553 -1863
rect -503 1863 -457 1875
rect -503 -1863 -497 1863
rect -463 -1863 -457 1863
rect -503 -1875 -457 -1863
rect -407 1863 -361 1875
rect -407 -1863 -401 1863
rect -367 -1863 -361 1863
rect -407 -1875 -361 -1863
rect -311 1863 -265 1875
rect -311 -1863 -305 1863
rect -271 -1863 -265 1863
rect -311 -1875 -265 -1863
rect -215 1863 -169 1875
rect -215 -1863 -209 1863
rect -175 -1863 -169 1863
rect -215 -1875 -169 -1863
rect -119 1863 -73 1875
rect -119 -1863 -113 1863
rect -79 -1863 -73 1863
rect -119 -1875 -73 -1863
rect -23 1863 23 1875
rect -23 -1863 -17 1863
rect 17 -1863 23 1863
rect -23 -1875 23 -1863
rect 73 1863 119 1875
rect 73 -1863 79 1863
rect 113 -1863 119 1863
rect 73 -1875 119 -1863
rect 169 1863 215 1875
rect 169 -1863 175 1863
rect 209 -1863 215 1863
rect 169 -1875 215 -1863
rect 265 1863 311 1875
rect 265 -1863 271 1863
rect 305 -1863 311 1863
rect 265 -1875 311 -1863
rect 361 1863 407 1875
rect 361 -1863 367 1863
rect 401 -1863 407 1863
rect 361 -1875 407 -1863
rect 457 1863 503 1875
rect 457 -1863 463 1863
rect 497 -1863 503 1863
rect 457 -1875 503 -1863
rect 553 1863 599 1875
rect 553 -1863 559 1863
rect 593 -1863 599 1863
rect 553 -1875 599 -1863
rect 649 1863 695 1875
rect 649 -1863 655 1863
rect 689 -1863 695 1863
rect 649 -1875 695 -1863
rect 745 1863 791 1875
rect 745 -1863 751 1863
rect 785 -1863 791 1863
rect 745 -1875 791 -1863
rect 841 1863 887 1875
rect 841 -1863 847 1863
rect 881 -1863 887 1863
rect 841 -1875 887 -1863
rect 937 1863 983 1875
rect 937 -1863 943 1863
rect 977 -1863 983 1863
rect 937 -1875 983 -1863
rect -941 -1913 -883 -1907
rect -941 -1947 -929 -1913
rect -895 -1947 -883 -1913
rect -941 -1953 -883 -1947
rect -749 -1913 -691 -1907
rect -749 -1947 -737 -1913
rect -703 -1947 -691 -1913
rect -749 -1953 -691 -1947
rect -557 -1913 -499 -1907
rect -557 -1947 -545 -1913
rect -511 -1947 -499 -1913
rect -557 -1953 -499 -1947
rect -365 -1913 -307 -1907
rect -365 -1947 -353 -1913
rect -319 -1947 -307 -1913
rect -365 -1953 -307 -1947
rect -173 -1913 -115 -1907
rect -173 -1947 -161 -1913
rect -127 -1947 -115 -1913
rect -173 -1953 -115 -1947
rect 19 -1913 77 -1907
rect 19 -1947 31 -1913
rect 65 -1947 77 -1913
rect 19 -1953 77 -1947
rect 211 -1913 269 -1907
rect 211 -1947 223 -1913
rect 257 -1947 269 -1913
rect 211 -1953 269 -1947
rect 403 -1913 461 -1907
rect 403 -1947 415 -1913
rect 449 -1947 461 -1913
rect 403 -1953 461 -1947
rect 595 -1913 653 -1907
rect 595 -1947 607 -1913
rect 641 -1947 653 -1913
rect 595 -1953 653 -1947
rect 787 -1913 845 -1907
rect 787 -1947 799 -1913
rect 833 -1947 845 -1913
rect 787 -1953 845 -1947
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -2032 1074 2032
string parameters w 18.75 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
