magic
tech sky130A
magscale 1 2
timestamp 1616191617
<< nwell >>
rect -866 998 1812 1462
rect -472 654 -142 998
rect -472 636 -160 654
rect 210 636 464 998
rect 862 636 1812 998
rect 258 634 442 636
rect 1450 632 1812 636
rect 722 -14 1302 96
rect 1608 -14 1810 632
rect -172 -288 452 -268
rect -172 -650 456 -288
rect 722 -300 1810 -14
rect 1280 -310 1810 -300
rect 1608 -314 1810 -310
rect -172 -652 242 -650
<< pwell >>
rect -858 520 -484 800
rect -860 518 -444 520
rect 184 518 880 520
rect -860 498 166 518
rect 184 498 1500 518
rect -860 196 1478 498
rect -858 194 1478 196
rect -858 192 166 194
rect 866 192 1478 194
rect -858 -754 -380 192
rect -858 -756 1668 -754
rect -866 -1090 1814 -756
<< nmos >>
rect 334 314 364 404
rect 1176 -622 1206 -532
rect 56 -984 86 -894
<< pmos >>
rect 334 710 364 890
rect 56 -588 86 -408
rect 1176 -226 1206 -46
<< ndiff >>
rect 276 392 334 404
rect 276 326 288 392
rect 322 326 334 392
rect 276 314 334 326
rect 364 392 422 404
rect 364 326 376 392
rect 410 326 422 392
rect 364 314 422 326
rect 1118 -544 1176 -532
rect 1118 -610 1130 -544
rect 1164 -610 1176 -544
rect 1118 -622 1176 -610
rect 1206 -544 1264 -532
rect 1206 -610 1218 -544
rect 1252 -610 1264 -544
rect 1206 -622 1264 -610
rect -2 -906 56 -894
rect -2 -972 10 -906
rect 44 -972 56 -906
rect -2 -984 56 -972
rect 86 -906 144 -894
rect 86 -972 98 -906
rect 132 -972 144 -906
rect 86 -984 144 -972
<< pdiff >>
rect 276 878 334 890
rect 276 722 288 878
rect 322 722 334 878
rect 276 710 334 722
rect 364 878 422 890
rect 364 722 376 878
rect 410 722 422 878
rect 364 710 422 722
rect -2 -420 56 -408
rect -2 -576 10 -420
rect 44 -576 56 -420
rect -2 -588 56 -576
rect 86 -420 144 -408
rect 86 -576 98 -420
rect 132 -576 144 -420
rect 86 -588 144 -576
rect 1118 -58 1176 -46
rect 1118 -214 1130 -58
rect 1164 -214 1176 -58
rect 1118 -226 1176 -214
rect 1206 -58 1264 -46
rect 1206 -214 1218 -58
rect 1252 -214 1264 -58
rect 1206 -226 1264 -214
<< ndiffc >>
rect 288 326 322 392
rect 376 326 410 392
rect 1130 -610 1164 -544
rect 1218 -610 1252 -544
rect 10 -972 44 -906
rect 98 -972 132 -906
<< pdiffc >>
rect 288 722 322 878
rect 376 722 410 878
rect 10 -576 44 -420
rect 98 -576 132 -420
rect 1130 -214 1164 -58
rect 1218 -214 1252 -58
<< poly >>
rect 404 1392 960 1462
rect 404 1144 444 1392
rect -436 1102 348 1138
rect 404 1106 586 1144
rect -866 918 -786 946
rect -436 918 -398 1102
rect 316 987 348 1102
rect 554 1078 584 1106
rect 316 971 382 987
rect 316 937 332 971
rect 366 937 382 971
rect 316 921 382 937
rect -866 888 -398 918
rect 334 890 364 921
rect -866 886 -402 888
rect -434 542 -402 886
rect 334 684 364 710
rect -178 610 -112 618
rect -178 558 46 610
rect -178 550 -112 558
rect -434 500 -288 542
rect -318 422 -288 500
rect 334 404 364 436
rect -318 36 -288 308
rect 334 178 364 314
rect -70 142 364 178
rect 34 36 100 51
rect -318 -2 100 36
rect 34 -16 100 -2
rect 56 -311 86 -16
rect 38 -327 104 -311
rect 38 -361 54 -327
rect 88 -361 104 -327
rect 38 -377 104 -361
rect 56 -408 86 -377
rect 56 -614 86 -588
rect 170 -788 204 142
rect 272 -156 338 -136
rect 272 -200 572 -156
rect 272 -204 338 -200
rect 914 -654 960 1392
rect 1200 566 1320 616
rect 1176 51 1206 98
rect 1158 35 1224 51
rect 1158 1 1174 35
rect 1208 1 1224 35
rect 1158 -15 1224 1
rect 1176 -46 1206 -15
rect 1176 -252 1206 -226
rect 1176 -532 1206 -468
rect 648 -686 960 -654
rect 1176 -660 1206 -622
rect 56 -830 204 -788
rect 56 -894 86 -830
rect 56 -1022 86 -984
<< polycont >>
rect 332 937 366 971
rect 54 -361 88 -327
rect 1174 1 1208 35
<< locali >>
rect 316 937 332 971
rect 366 937 382 971
rect 288 878 322 894
rect 288 706 322 722
rect 376 878 410 894
rect 376 706 410 722
rect 288 392 322 408
rect 288 310 322 326
rect 376 392 410 408
rect 376 310 410 326
rect 1158 1 1174 35
rect 1208 1 1224 35
rect 1130 -58 1164 -42
rect 1130 -230 1164 -214
rect 1218 -58 1252 -42
rect 1218 -230 1252 -214
rect 38 -361 54 -327
rect 88 -361 104 -327
rect 10 -420 44 -404
rect 10 -592 44 -576
rect 98 -420 132 -404
rect 98 -592 132 -576
rect 1130 -544 1164 -528
rect 1130 -626 1164 -610
rect 1218 -544 1252 -528
rect 1218 -626 1252 -610
rect 10 -906 44 -890
rect 10 -988 44 -972
rect 98 -906 132 -890
rect 98 -988 132 -972
<< viali >>
rect 332 937 366 971
rect 288 722 322 878
rect 376 722 410 878
rect 1014 518 1072 600
rect -676 424 -618 508
rect 288 326 322 392
rect 376 326 410 392
rect 1174 1 1208 35
rect 1130 -214 1164 -58
rect 1218 -214 1252 -58
rect 54 -361 88 -327
rect 10 -576 44 -420
rect 98 -576 132 -420
rect 1130 -610 1164 -544
rect 1218 -610 1252 -544
rect 10 -972 44 -906
rect 98 -972 132 -906
<< metal1 >>
rect -486 1320 -76 1462
rect -486 1296 796 1320
rect -250 1214 796 1296
rect -342 986 -332 988
rect -362 984 -332 986
rect -620 930 -332 984
rect -342 928 -332 930
rect -274 928 -264 988
rect -130 954 -70 1214
rect 836 1184 1470 1302
rect 1128 1066 1468 1184
rect 318 971 378 986
rect 318 937 332 971
rect 366 937 380 971
rect 318 922 380 937
rect 282 878 328 890
rect -682 508 -612 520
rect -682 424 -676 508
rect -618 490 -612 508
rect -364 490 -330 778
rect -276 608 -242 778
rect 282 722 288 878
rect 322 722 328 878
rect 282 710 328 722
rect 370 878 416 890
rect 370 722 376 878
rect 410 722 416 878
rect 370 710 416 722
rect -276 560 -114 608
rect 288 604 322 710
rect 56 572 322 604
rect -618 452 -328 490
rect -618 424 -612 452
rect -682 412 -612 424
rect -364 362 -330 452
rect -276 362 -242 560
rect 288 404 322 572
rect 376 626 410 710
rect 376 592 696 626
rect 1008 600 1258 622
rect 376 404 410 592
rect 1008 580 1014 600
rect 834 536 1014 580
rect 1008 518 1014 536
rect 1072 570 1258 600
rect 1072 518 1078 570
rect 1196 562 1258 570
rect 1448 546 1458 620
rect 1518 546 1528 620
rect 1008 506 1078 518
rect 282 392 328 404
rect -276 -650 -240 362
rect 282 326 288 392
rect 322 326 328 392
rect 282 314 328 326
rect 370 392 416 404
rect 370 326 376 392
rect 410 326 416 392
rect 1608 360 1666 364
rect 370 314 416 326
rect -106 126 -96 193
rect -30 126 -20 193
rect 288 156 322 314
rect 376 162 410 314
rect 1412 280 1670 360
rect 24 -16 34 51
rect 100 -16 110 51
rect 288 -150 320 156
rect 374 130 1022 162
rect 992 -288 1022 130
rect 1150 122 1160 202
rect 1226 122 1236 202
rect 1162 48 1222 122
rect 1160 35 1222 48
rect 1160 1 1174 35
rect 1208 1 1222 35
rect 1160 -14 1222 1
rect 1124 -58 1170 -46
rect 1124 -214 1130 -58
rect 1164 -214 1170 -58
rect 1124 -226 1170 -214
rect 1212 -58 1258 -46
rect 1212 -214 1218 -58
rect 1252 -214 1258 -58
rect 1212 -226 1258 -214
rect 1130 -288 1164 -226
rect 40 -327 102 -314
rect 40 -361 54 -327
rect 88 -361 102 -327
rect 992 -330 1164 -288
rect 40 -376 102 -361
rect 4 -420 50 -408
rect 4 -576 10 -420
rect 44 -576 50 -420
rect 4 -588 50 -576
rect 92 -420 138 -408
rect 92 -576 98 -420
rect 132 -576 138 -420
rect 1130 -532 1164 -330
rect 1218 -364 1252 -226
rect 1416 -364 1426 -336
rect 1218 -400 1426 -364
rect 1218 -532 1252 -400
rect 1416 -424 1426 -400
rect 1496 -424 1506 -336
rect 92 -588 138 -576
rect 1124 -544 1170 -532
rect 10 -650 44 -588
rect -276 -692 44 -650
rect 10 -894 44 -692
rect 98 -728 132 -588
rect 1124 -610 1130 -544
rect 1164 -610 1170 -544
rect 1124 -622 1170 -610
rect 1212 -544 1258 -532
rect 1212 -610 1218 -544
rect 1252 -610 1258 -544
rect 1212 -622 1258 -610
rect 1148 -724 1158 -657
rect 1224 -724 1234 -657
rect 98 -762 808 -728
rect 98 -894 132 -762
rect 4 -906 50 -894
rect 4 -972 10 -906
rect 44 -972 50 -906
rect 4 -984 50 -972
rect 92 -906 138 -894
rect 92 -972 98 -906
rect 132 -972 138 -906
rect 1608 -966 1666 280
rect 92 -984 138 -972
rect 768 -1072 1666 -966
rect 768 -1074 1664 -1072
<< via1 >>
rect -332 928 -274 988
rect 1458 546 1518 620
rect -96 126 -30 193
rect 34 -16 100 51
rect 1160 122 1226 202
rect 1426 -424 1496 -336
rect 1158 -724 1224 -657
<< metal2 >>
rect -322 998 -172 1004
rect -332 988 -172 998
rect -274 932 -172 988
rect -332 918 -274 928
rect -210 184 -172 932
rect 1458 620 1518 630
rect 1458 536 1518 546
rect -96 193 -30 203
rect -210 132 -96 184
rect 1160 202 1226 212
rect -30 138 1160 184
rect -96 116 -30 126
rect 1160 112 1226 122
rect 34 51 100 61
rect -146 -16 34 46
rect -146 -26 100 -16
rect -144 -660 -108 -26
rect 1472 -326 1504 536
rect 1426 -336 1504 -326
rect 1496 -424 1504 -336
rect 1426 -432 1504 -424
rect 1426 -434 1496 -432
rect 1158 -657 1224 -647
rect -144 -724 1158 -660
rect 1158 -734 1224 -724
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_5
timestamp 1616001657
transform 1 0 67 0 1 -52
box -33 36 33 103
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_2
timestamp 1616001657
transform 1 0 305 0 1 -240
box -33 36 33 103
use nor  nor_1
timestamp 1616102052
transform 1 0 510 0 1 -344
box -62 -746 356 438
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_6
timestamp 1616001657
transform 1 0 1191 0 1 -760
box -33 36 33 103
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615953154
transform 1 0 -303 0 1 361
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_A663FE  sky130_fd_pr__pfet_01v8_A663FE_0
timestamp 1616013451
transform 1 0 -303 0 1 838
box -109 -188 109 154
use inverter2  inverter2_1
timestamp 1616102052
transform 1 0 -774 0 1 1000
box -84 -364 296 458
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_3
timestamp 1616001657
transform 1 0 -63 0 1 90
box -33 36 33 103
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_0
timestamp 1616001657
transform 1 0 -145 0 1 514
box -33 36 33 103
use inverter2  inverter2_0
timestamp 1616102052
transform 1 0 -78 0 1 638
box -84 -364 296 458
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_1
timestamp 1616001657
transform 1 0 677 0 1 540
box -33 36 33 103
use nor  nor_0
timestamp 1616102052
transform 1 0 522 0 1 940
box -62 -746 356 438
use sky130_fd_pr__pfet_01v8_ACP95B  sky130_fd_pr__pfet_01v8_ACP95B_4
timestamp 1616001657
transform 1 0 1227 0 1 520
box -33 36 33 103
use inverter2  inverter2_2
timestamp 1616102052
transform 1 0 1210 0 1 642
box -84 -364 296 458
<< end >>
