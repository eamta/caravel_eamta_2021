magic
tech sky130A
magscale 1 2
timestamp 1623263513
<< nwell >>
rect -186 12450 270 14480
rect 278 12450 9021 14561
rect -186 12322 9021 12450
rect -186 10943 270 12322
rect 278 10943 9021 12322
<< metal1 >>
rect -3925 14353 -3915 14525
rect -133 14353 -123 14525
<< via1 >>
rect -3915 14353 -133 14525
<< metal2 >>
rect -3915 14525 -133 14535
rect -133 14353 13227 14515
rect -3915 14343 13227 14353
rect -771 10896 -197 10906
rect -771 10593 -197 10603
rect 2989 10456 3270 10466
rect 2989 10231 3270 10241
rect 7456 10456 7737 10466
rect 7456 10231 7737 10241
rect 11923 10456 12204 10466
rect 11923 10231 12204 10241
rect 2367 9406 2622 9416
rect 2367 8911 2622 8921
rect 6834 9406 7089 9416
rect 3148 8905 4074 8915
rect 6834 8911 7089 8921
rect 11301 9406 11556 9416
rect 3148 8399 4074 8409
rect 7615 8905 8541 8915
rect 11301 8911 11556 8921
rect 7615 8399 8541 8409
rect 12082 8905 13008 8915
rect 12082 8399 13008 8409
rect -1639 7762 -1307 7772
rect -1639 7058 -1307 7068
rect 159 6 13266 198
<< via2 >>
rect -771 10603 -197 10896
rect 2989 10241 3270 10456
rect 7456 10241 7737 10456
rect 11923 10241 12204 10456
rect 2367 8921 2622 9406
rect 6834 8921 7089 9406
rect 11301 8921 11556 9406
rect 3148 8409 4074 8905
rect 7615 8409 8541 8905
rect 12082 8409 13008 8905
rect -1639 7068 -1307 7762
<< metal3 >>
rect -781 10896 -187 10901
rect -781 10603 -771 10896
rect -197 10603 12214 10896
rect -781 10598 -187 10603
rect 2979 10456 3280 10603
rect 2979 10241 2989 10456
rect 3270 10241 3280 10456
rect 2979 10236 3280 10241
rect 7446 10456 7747 10603
rect 7446 10241 7456 10456
rect 7737 10241 7747 10456
rect 7446 10236 7747 10241
rect 11913 10456 12214 10603
rect 11913 10241 11923 10456
rect 12204 10241 12214 10456
rect 11913 10236 12214 10241
rect -1649 9406 11566 9496
rect -1649 9144 2367 9406
rect -1649 7762 -1297 9144
rect 2357 8921 2367 9144
rect 2622 9144 6834 9406
rect 2622 8921 2632 9144
rect 2357 8916 2632 8921
rect 6824 8921 6834 9144
rect 7089 9144 11301 9406
rect 7089 8921 7099 9144
rect 6824 8916 7099 8921
rect 11291 8921 11301 9144
rect 11556 8921 11566 9406
rect 11291 8916 11566 8921
rect 3138 8905 4084 8910
rect 3138 8409 3148 8905
rect 4074 8409 4084 8905
rect 3138 8404 4084 8409
rect 7605 8905 8551 8910
rect 7605 8409 7615 8905
rect 8541 8409 8551 8905
rect 7605 8404 8551 8409
rect 12072 8905 13018 8910
rect 12072 8409 12082 8905
rect 13008 8409 13018 8905
rect 12072 8404 13018 8409
rect -1649 7068 -1639 7762
rect -1307 7068 -1297 7762
rect -1649 6636 -1297 7068
rect -2387 6051 -1297 6636
use bias_reference  bias_reference_0
timestamp 1623262251
transform 1 0 -3993 0 1 11016
box -54 -3958 3993 3545
use bias  bias_2
timestamp 1623250946
transform 1 0 8360 0 1 852
box 574 -852 5041 13709
use bias  bias_1
timestamp 1623250946
transform 1 0 3893 0 1 852
box 574 -852 5041 13709
use bias  bias_0
timestamp 1623250946
transform 1 0 -574 0 1 852
box 574 -852 5041 13709
<< labels >>
rlabel metal2 -3915 14343 13227 14515 1 vdd
rlabel metal2 159 6 13266 198 1 vss
rlabel metal3 -2387 6051 -1297 6636 1 vref
rlabel via2 3148 8409 4074 8905 1 ibias_1
rlabel via2 7615 8409 8541 8905 1 ibias_2
rlabel via2 12082 8409 13008 8905 1 ibias_3
<< end >>
