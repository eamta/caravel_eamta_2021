magic
tech sky130A
magscale 1 2
timestamp 1623255091
<< error_p >>
rect -927 1581 -865 1587
rect -799 1581 -737 1587
rect -671 1581 -609 1587
rect -543 1581 -481 1587
rect -415 1581 -353 1587
rect -287 1581 -225 1587
rect -159 1581 -97 1587
rect -31 1581 31 1587
rect 97 1581 159 1587
rect 225 1581 287 1587
rect 353 1581 415 1587
rect 481 1581 543 1587
rect 609 1581 671 1587
rect 737 1581 799 1587
rect 865 1581 927 1587
rect -927 1547 -915 1581
rect -799 1547 -787 1581
rect -671 1547 -659 1581
rect -543 1547 -531 1581
rect -415 1547 -403 1581
rect -287 1547 -275 1581
rect -159 1547 -147 1581
rect -31 1547 -19 1581
rect 97 1547 109 1581
rect 225 1547 237 1581
rect 353 1547 365 1581
rect 481 1547 493 1581
rect 609 1547 621 1581
rect 737 1547 749 1581
rect 865 1547 877 1581
rect -927 1541 -865 1547
rect -799 1541 -737 1547
rect -671 1541 -609 1547
rect -543 1541 -481 1547
rect -415 1541 -353 1547
rect -287 1541 -225 1547
rect -159 1541 -97 1547
rect -31 1541 31 1547
rect 97 1541 159 1547
rect 225 1541 287 1547
rect 353 1541 415 1547
rect 481 1541 543 1547
rect 609 1541 671 1547
rect 737 1541 799 1547
rect 865 1541 927 1547
rect -927 -1547 -865 -1541
rect -799 -1547 -737 -1541
rect -671 -1547 -609 -1541
rect -543 -1547 -481 -1541
rect -415 -1547 -353 -1541
rect -287 -1547 -225 -1541
rect -159 -1547 -97 -1541
rect -31 -1547 31 -1541
rect 97 -1547 159 -1541
rect 225 -1547 287 -1541
rect 353 -1547 415 -1541
rect 481 -1547 543 -1541
rect 609 -1547 671 -1541
rect 737 -1547 799 -1541
rect 865 -1547 927 -1541
rect -927 -1581 -915 -1547
rect -799 -1581 -787 -1547
rect -671 -1581 -659 -1547
rect -543 -1581 -531 -1547
rect -415 -1581 -403 -1547
rect -287 -1581 -275 -1547
rect -159 -1581 -147 -1547
rect -31 -1581 -19 -1547
rect 97 -1581 109 -1547
rect 225 -1581 237 -1547
rect 353 -1581 365 -1547
rect 481 -1581 493 -1547
rect 609 -1581 621 -1547
rect 737 -1581 749 -1547
rect 865 -1581 877 -1547
rect -927 -1587 -865 -1581
rect -799 -1587 -737 -1581
rect -671 -1587 -609 -1581
rect -543 -1587 -481 -1581
rect -415 -1587 -353 -1581
rect -287 -1587 -225 -1581
rect -159 -1587 -97 -1581
rect -31 -1587 31 -1581
rect 97 -1587 159 -1581
rect 225 -1587 287 -1581
rect 353 -1587 415 -1581
rect 481 -1587 543 -1581
rect 609 -1587 671 -1581
rect 737 -1587 799 -1581
rect 865 -1587 927 -1581
<< nwell >>
rect -1127 -1719 1127 1719
<< pmoslvt >>
rect -931 -1500 -861 1500
rect -803 -1500 -733 1500
rect -675 -1500 -605 1500
rect -547 -1500 -477 1500
rect -419 -1500 -349 1500
rect -291 -1500 -221 1500
rect -163 -1500 -93 1500
rect -35 -1500 35 1500
rect 93 -1500 163 1500
rect 221 -1500 291 1500
rect 349 -1500 419 1500
rect 477 -1500 547 1500
rect 605 -1500 675 1500
rect 733 -1500 803 1500
rect 861 -1500 931 1500
<< pdiff >>
rect -989 1488 -931 1500
rect -989 -1488 -977 1488
rect -943 -1488 -931 1488
rect -989 -1500 -931 -1488
rect -861 1488 -803 1500
rect -861 -1488 -849 1488
rect -815 -1488 -803 1488
rect -861 -1500 -803 -1488
rect -733 1488 -675 1500
rect -733 -1488 -721 1488
rect -687 -1488 -675 1488
rect -733 -1500 -675 -1488
rect -605 1488 -547 1500
rect -605 -1488 -593 1488
rect -559 -1488 -547 1488
rect -605 -1500 -547 -1488
rect -477 1488 -419 1500
rect -477 -1488 -465 1488
rect -431 -1488 -419 1488
rect -477 -1500 -419 -1488
rect -349 1488 -291 1500
rect -349 -1488 -337 1488
rect -303 -1488 -291 1488
rect -349 -1500 -291 -1488
rect -221 1488 -163 1500
rect -221 -1488 -209 1488
rect -175 -1488 -163 1488
rect -221 -1500 -163 -1488
rect -93 1488 -35 1500
rect -93 -1488 -81 1488
rect -47 -1488 -35 1488
rect -93 -1500 -35 -1488
rect 35 1488 93 1500
rect 35 -1488 47 1488
rect 81 -1488 93 1488
rect 35 -1500 93 -1488
rect 163 1488 221 1500
rect 163 -1488 175 1488
rect 209 -1488 221 1488
rect 163 -1500 221 -1488
rect 291 1488 349 1500
rect 291 -1488 303 1488
rect 337 -1488 349 1488
rect 291 -1500 349 -1488
rect 419 1488 477 1500
rect 419 -1488 431 1488
rect 465 -1488 477 1488
rect 419 -1500 477 -1488
rect 547 1488 605 1500
rect 547 -1488 559 1488
rect 593 -1488 605 1488
rect 547 -1500 605 -1488
rect 675 1488 733 1500
rect 675 -1488 687 1488
rect 721 -1488 733 1488
rect 675 -1500 733 -1488
rect 803 1488 861 1500
rect 803 -1488 815 1488
rect 849 -1488 861 1488
rect 803 -1500 861 -1488
rect 931 1488 989 1500
rect 931 -1488 943 1488
rect 977 -1488 989 1488
rect 931 -1500 989 -1488
<< pdiffc >>
rect -977 -1488 -943 1488
rect -849 -1488 -815 1488
rect -721 -1488 -687 1488
rect -593 -1488 -559 1488
rect -465 -1488 -431 1488
rect -337 -1488 -303 1488
rect -209 -1488 -175 1488
rect -81 -1488 -47 1488
rect 47 -1488 81 1488
rect 175 -1488 209 1488
rect 303 -1488 337 1488
rect 431 -1488 465 1488
rect 559 -1488 593 1488
rect 687 -1488 721 1488
rect 815 -1488 849 1488
rect 943 -1488 977 1488
<< nsubdiff >>
rect -1091 1649 -995 1683
rect 995 1649 1091 1683
rect -1091 1587 -1057 1649
rect 1057 1587 1091 1649
rect -1091 -1649 -1057 -1587
rect 1057 -1649 1091 -1587
rect -1091 -1683 -995 -1649
rect 995 -1683 1091 -1649
<< nsubdiffcont >>
rect -995 1649 995 1683
rect -1091 -1587 -1057 1587
rect 1057 -1587 1091 1587
rect -995 -1683 995 -1649
<< poly >>
rect -931 1581 -861 1597
rect -931 1547 -915 1581
rect -877 1547 -861 1581
rect -931 1500 -861 1547
rect -803 1581 -733 1597
rect -803 1547 -787 1581
rect -749 1547 -733 1581
rect -803 1500 -733 1547
rect -675 1581 -605 1597
rect -675 1547 -659 1581
rect -621 1547 -605 1581
rect -675 1500 -605 1547
rect -547 1581 -477 1597
rect -547 1547 -531 1581
rect -493 1547 -477 1581
rect -547 1500 -477 1547
rect -419 1581 -349 1597
rect -419 1547 -403 1581
rect -365 1547 -349 1581
rect -419 1500 -349 1547
rect -291 1581 -221 1597
rect -291 1547 -275 1581
rect -237 1547 -221 1581
rect -291 1500 -221 1547
rect -163 1581 -93 1597
rect -163 1547 -147 1581
rect -109 1547 -93 1581
rect -163 1500 -93 1547
rect -35 1581 35 1597
rect -35 1547 -19 1581
rect 19 1547 35 1581
rect -35 1500 35 1547
rect 93 1581 163 1597
rect 93 1547 109 1581
rect 147 1547 163 1581
rect 93 1500 163 1547
rect 221 1581 291 1597
rect 221 1547 237 1581
rect 275 1547 291 1581
rect 221 1500 291 1547
rect 349 1581 419 1597
rect 349 1547 365 1581
rect 403 1547 419 1581
rect 349 1500 419 1547
rect 477 1581 547 1597
rect 477 1547 493 1581
rect 531 1547 547 1581
rect 477 1500 547 1547
rect 605 1581 675 1597
rect 605 1547 621 1581
rect 659 1547 675 1581
rect 605 1500 675 1547
rect 733 1581 803 1597
rect 733 1547 749 1581
rect 787 1547 803 1581
rect 733 1500 803 1547
rect 861 1581 931 1597
rect 861 1547 877 1581
rect 915 1547 931 1581
rect 861 1500 931 1547
rect -931 -1547 -861 -1500
rect -931 -1581 -915 -1547
rect -877 -1581 -861 -1547
rect -931 -1597 -861 -1581
rect -803 -1547 -733 -1500
rect -803 -1581 -787 -1547
rect -749 -1581 -733 -1547
rect -803 -1597 -733 -1581
rect -675 -1547 -605 -1500
rect -675 -1581 -659 -1547
rect -621 -1581 -605 -1547
rect -675 -1597 -605 -1581
rect -547 -1547 -477 -1500
rect -547 -1581 -531 -1547
rect -493 -1581 -477 -1547
rect -547 -1597 -477 -1581
rect -419 -1547 -349 -1500
rect -419 -1581 -403 -1547
rect -365 -1581 -349 -1547
rect -419 -1597 -349 -1581
rect -291 -1547 -221 -1500
rect -291 -1581 -275 -1547
rect -237 -1581 -221 -1547
rect -291 -1597 -221 -1581
rect -163 -1547 -93 -1500
rect -163 -1581 -147 -1547
rect -109 -1581 -93 -1547
rect -163 -1597 -93 -1581
rect -35 -1547 35 -1500
rect -35 -1581 -19 -1547
rect 19 -1581 35 -1547
rect -35 -1597 35 -1581
rect 93 -1547 163 -1500
rect 93 -1581 109 -1547
rect 147 -1581 163 -1547
rect 93 -1597 163 -1581
rect 221 -1547 291 -1500
rect 221 -1581 237 -1547
rect 275 -1581 291 -1547
rect 221 -1597 291 -1581
rect 349 -1547 419 -1500
rect 349 -1581 365 -1547
rect 403 -1581 419 -1547
rect 349 -1597 419 -1581
rect 477 -1547 547 -1500
rect 477 -1581 493 -1547
rect 531 -1581 547 -1547
rect 477 -1597 547 -1581
rect 605 -1547 675 -1500
rect 605 -1581 621 -1547
rect 659 -1581 675 -1547
rect 605 -1597 675 -1581
rect 733 -1547 803 -1500
rect 733 -1581 749 -1547
rect 787 -1581 803 -1547
rect 733 -1597 803 -1581
rect 861 -1547 931 -1500
rect 861 -1581 877 -1547
rect 915 -1581 931 -1547
rect 861 -1597 931 -1581
<< polycont >>
rect -915 1547 -877 1581
rect -787 1547 -749 1581
rect -659 1547 -621 1581
rect -531 1547 -493 1581
rect -403 1547 -365 1581
rect -275 1547 -237 1581
rect -147 1547 -109 1581
rect -19 1547 19 1581
rect 109 1547 147 1581
rect 237 1547 275 1581
rect 365 1547 403 1581
rect 493 1547 531 1581
rect 621 1547 659 1581
rect 749 1547 787 1581
rect 877 1547 915 1581
rect -915 -1581 -877 -1547
rect -787 -1581 -749 -1547
rect -659 -1581 -621 -1547
rect -531 -1581 -493 -1547
rect -403 -1581 -365 -1547
rect -275 -1581 -237 -1547
rect -147 -1581 -109 -1547
rect -19 -1581 19 -1547
rect 109 -1581 147 -1547
rect 237 -1581 275 -1547
rect 365 -1581 403 -1547
rect 493 -1581 531 -1547
rect 621 -1581 659 -1547
rect 749 -1581 787 -1547
rect 877 -1581 915 -1547
<< locali >>
rect -1091 1649 -995 1683
rect 995 1649 1091 1683
rect -1091 1587 -1057 1649
rect 1057 1587 1091 1649
rect -931 1547 -915 1581
rect -877 1547 -861 1581
rect -803 1547 -787 1581
rect -749 1547 -733 1581
rect -675 1547 -659 1581
rect -621 1547 -605 1581
rect -547 1547 -531 1581
rect -493 1547 -477 1581
rect -419 1547 -403 1581
rect -365 1547 -349 1581
rect -291 1547 -275 1581
rect -237 1547 -221 1581
rect -163 1547 -147 1581
rect -109 1547 -93 1581
rect -35 1547 -19 1581
rect 19 1547 35 1581
rect 93 1547 109 1581
rect 147 1547 163 1581
rect 221 1547 237 1581
rect 275 1547 291 1581
rect 349 1547 365 1581
rect 403 1547 419 1581
rect 477 1547 493 1581
rect 531 1547 547 1581
rect 605 1547 621 1581
rect 659 1547 675 1581
rect 733 1547 749 1581
rect 787 1547 803 1581
rect 861 1547 877 1581
rect 915 1547 931 1581
rect -977 1488 -943 1504
rect -977 -1504 -943 -1488
rect -849 1488 -815 1504
rect -849 -1504 -815 -1488
rect -721 1488 -687 1504
rect -721 -1504 -687 -1488
rect -593 1488 -559 1504
rect -593 -1504 -559 -1488
rect -465 1488 -431 1504
rect -465 -1504 -431 -1488
rect -337 1488 -303 1504
rect -337 -1504 -303 -1488
rect -209 1488 -175 1504
rect -209 -1504 -175 -1488
rect -81 1488 -47 1504
rect -81 -1504 -47 -1488
rect 47 1488 81 1504
rect 47 -1504 81 -1488
rect 175 1488 209 1504
rect 175 -1504 209 -1488
rect 303 1488 337 1504
rect 303 -1504 337 -1488
rect 431 1488 465 1504
rect 431 -1504 465 -1488
rect 559 1488 593 1504
rect 559 -1504 593 -1488
rect 687 1488 721 1504
rect 687 -1504 721 -1488
rect 815 1488 849 1504
rect 815 -1504 849 -1488
rect 943 1488 977 1504
rect 943 -1504 977 -1488
rect -931 -1581 -915 -1547
rect -877 -1581 -861 -1547
rect -803 -1581 -787 -1547
rect -749 -1581 -733 -1547
rect -675 -1581 -659 -1547
rect -621 -1581 -605 -1547
rect -547 -1581 -531 -1547
rect -493 -1581 -477 -1547
rect -419 -1581 -403 -1547
rect -365 -1581 -349 -1547
rect -291 -1581 -275 -1547
rect -237 -1581 -221 -1547
rect -163 -1581 -147 -1547
rect -109 -1581 -93 -1547
rect -35 -1581 -19 -1547
rect 19 -1581 35 -1547
rect 93 -1581 109 -1547
rect 147 -1581 163 -1547
rect 221 -1581 237 -1547
rect 275 -1581 291 -1547
rect 349 -1581 365 -1547
rect 403 -1581 419 -1547
rect 477 -1581 493 -1547
rect 531 -1581 547 -1547
rect 605 -1581 621 -1547
rect 659 -1581 675 -1547
rect 733 -1581 749 -1547
rect 787 -1581 803 -1547
rect 861 -1581 877 -1547
rect 915 -1581 931 -1547
rect -1091 -1649 -1057 -1587
rect 1057 -1649 1091 -1587
rect -1091 -1683 -995 -1649
rect 995 -1683 1091 -1649
<< viali >>
rect -915 1547 -877 1581
rect -787 1547 -749 1581
rect -659 1547 -621 1581
rect -531 1547 -493 1581
rect -403 1547 -365 1581
rect -275 1547 -237 1581
rect -147 1547 -109 1581
rect -19 1547 19 1581
rect 109 1547 147 1581
rect 237 1547 275 1581
rect 365 1547 403 1581
rect 493 1547 531 1581
rect 621 1547 659 1581
rect 749 1547 787 1581
rect 877 1547 915 1581
rect -977 -1488 -943 1488
rect -849 -1488 -815 1488
rect -721 -1488 -687 1488
rect -593 -1488 -559 1488
rect -465 -1488 -431 1488
rect -337 -1488 -303 1488
rect -209 -1488 -175 1488
rect -81 -1488 -47 1488
rect 47 -1488 81 1488
rect 175 -1488 209 1488
rect 303 -1488 337 1488
rect 431 -1488 465 1488
rect 559 -1488 593 1488
rect 687 -1488 721 1488
rect 815 -1488 849 1488
rect 943 -1488 977 1488
rect -915 -1581 -877 -1547
rect -787 -1581 -749 -1547
rect -659 -1581 -621 -1547
rect -531 -1581 -493 -1547
rect -403 -1581 -365 -1547
rect -275 -1581 -237 -1547
rect -147 -1581 -109 -1547
rect -19 -1581 19 -1547
rect 109 -1581 147 -1547
rect 237 -1581 275 -1547
rect 365 -1581 403 -1547
rect 493 -1581 531 -1547
rect 621 -1581 659 -1547
rect 749 -1581 787 -1547
rect 877 -1581 915 -1547
<< metal1 >>
rect -927 1581 -865 1587
rect -927 1547 -915 1581
rect -877 1547 -865 1581
rect -927 1541 -865 1547
rect -799 1581 -737 1587
rect -799 1547 -787 1581
rect -749 1547 -737 1581
rect -799 1541 -737 1547
rect -671 1581 -609 1587
rect -671 1547 -659 1581
rect -621 1547 -609 1581
rect -671 1541 -609 1547
rect -543 1581 -481 1587
rect -543 1547 -531 1581
rect -493 1547 -481 1581
rect -543 1541 -481 1547
rect -415 1581 -353 1587
rect -415 1547 -403 1581
rect -365 1547 -353 1581
rect -415 1541 -353 1547
rect -287 1581 -225 1587
rect -287 1547 -275 1581
rect -237 1547 -225 1581
rect -287 1541 -225 1547
rect -159 1581 -97 1587
rect -159 1547 -147 1581
rect -109 1547 -97 1581
rect -159 1541 -97 1547
rect -31 1581 31 1587
rect -31 1547 -19 1581
rect 19 1547 31 1581
rect -31 1541 31 1547
rect 97 1581 159 1587
rect 97 1547 109 1581
rect 147 1547 159 1581
rect 97 1541 159 1547
rect 225 1581 287 1587
rect 225 1547 237 1581
rect 275 1547 287 1581
rect 225 1541 287 1547
rect 353 1581 415 1587
rect 353 1547 365 1581
rect 403 1547 415 1581
rect 353 1541 415 1547
rect 481 1581 543 1587
rect 481 1547 493 1581
rect 531 1547 543 1581
rect 481 1541 543 1547
rect 609 1581 671 1587
rect 609 1547 621 1581
rect 659 1547 671 1581
rect 609 1541 671 1547
rect 737 1581 799 1587
rect 737 1547 749 1581
rect 787 1547 799 1581
rect 737 1541 799 1547
rect 865 1581 927 1587
rect 865 1547 877 1581
rect 915 1547 927 1581
rect 865 1541 927 1547
rect -983 1488 -937 1500
rect -983 -1488 -977 1488
rect -943 -1488 -937 1488
rect -983 -1500 -937 -1488
rect -855 1488 -809 1500
rect -855 -1488 -849 1488
rect -815 -1488 -809 1488
rect -855 -1500 -809 -1488
rect -727 1488 -681 1500
rect -727 -1488 -721 1488
rect -687 -1488 -681 1488
rect -727 -1500 -681 -1488
rect -599 1488 -553 1500
rect -599 -1488 -593 1488
rect -559 -1488 -553 1488
rect -599 -1500 -553 -1488
rect -471 1488 -425 1500
rect -471 -1488 -465 1488
rect -431 -1488 -425 1488
rect -471 -1500 -425 -1488
rect -343 1488 -297 1500
rect -343 -1488 -337 1488
rect -303 -1488 -297 1488
rect -343 -1500 -297 -1488
rect -215 1488 -169 1500
rect -215 -1488 -209 1488
rect -175 -1488 -169 1488
rect -215 -1500 -169 -1488
rect -87 1488 -41 1500
rect -87 -1488 -81 1488
rect -47 -1488 -41 1488
rect -87 -1500 -41 -1488
rect 41 1488 87 1500
rect 41 -1488 47 1488
rect 81 -1488 87 1488
rect 41 -1500 87 -1488
rect 169 1488 215 1500
rect 169 -1488 175 1488
rect 209 -1488 215 1488
rect 169 -1500 215 -1488
rect 297 1488 343 1500
rect 297 -1488 303 1488
rect 337 -1488 343 1488
rect 297 -1500 343 -1488
rect 425 1488 471 1500
rect 425 -1488 431 1488
rect 465 -1488 471 1488
rect 425 -1500 471 -1488
rect 553 1488 599 1500
rect 553 -1488 559 1488
rect 593 -1488 599 1488
rect 553 -1500 599 -1488
rect 681 1488 727 1500
rect 681 -1488 687 1488
rect 721 -1488 727 1488
rect 681 -1500 727 -1488
rect 809 1488 855 1500
rect 809 -1488 815 1488
rect 849 -1488 855 1488
rect 809 -1500 855 -1488
rect 937 1488 983 1500
rect 937 -1488 943 1488
rect 977 -1488 983 1488
rect 937 -1500 983 -1488
rect -927 -1547 -865 -1541
rect -927 -1581 -915 -1547
rect -877 -1581 -865 -1547
rect -927 -1587 -865 -1581
rect -799 -1547 -737 -1541
rect -799 -1581 -787 -1547
rect -749 -1581 -737 -1547
rect -799 -1587 -737 -1581
rect -671 -1547 -609 -1541
rect -671 -1581 -659 -1547
rect -621 -1581 -609 -1547
rect -671 -1587 -609 -1581
rect -543 -1547 -481 -1541
rect -543 -1581 -531 -1547
rect -493 -1581 -481 -1547
rect -543 -1587 -481 -1581
rect -415 -1547 -353 -1541
rect -415 -1581 -403 -1547
rect -365 -1581 -353 -1547
rect -415 -1587 -353 -1581
rect -287 -1547 -225 -1541
rect -287 -1581 -275 -1547
rect -237 -1581 -225 -1547
rect -287 -1587 -225 -1581
rect -159 -1547 -97 -1541
rect -159 -1581 -147 -1547
rect -109 -1581 -97 -1547
rect -159 -1587 -97 -1581
rect -31 -1547 31 -1541
rect -31 -1581 -19 -1547
rect 19 -1581 31 -1547
rect -31 -1587 31 -1581
rect 97 -1547 159 -1541
rect 97 -1581 109 -1547
rect 147 -1581 159 -1547
rect 97 -1587 159 -1581
rect 225 -1547 287 -1541
rect 225 -1581 237 -1547
rect 275 -1581 287 -1547
rect 225 -1587 287 -1581
rect 353 -1547 415 -1541
rect 353 -1581 365 -1547
rect 403 -1581 415 -1547
rect 353 -1587 415 -1581
rect 481 -1547 543 -1541
rect 481 -1581 493 -1547
rect 531 -1581 543 -1547
rect 481 -1587 543 -1581
rect 609 -1547 671 -1541
rect 609 -1581 621 -1547
rect 659 -1581 671 -1547
rect 609 -1587 671 -1581
rect 737 -1547 799 -1541
rect 737 -1581 749 -1547
rect 787 -1581 799 -1547
rect 737 -1587 799 -1581
rect 865 -1547 927 -1541
rect 865 -1581 877 -1547
rect 915 -1581 927 -1547
rect 865 -1587 927 -1581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -1074 -1666 1074 1666
string parameters w 15 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
