magic
tech sky130A
magscale 1 2
timestamp 1623887338
<< metal3 >>
rect -4969 4872 -1670 4900
rect -4969 1728 -1754 4872
rect -1690 1728 -1670 4872
rect -4969 1700 -1670 1728
rect -1430 4872 1869 4900
rect -1430 1728 1785 4872
rect 1849 1728 1869 4872
rect -1430 1700 1869 1728
rect 2109 4872 5408 4900
rect 2109 1728 5324 4872
rect 5388 1728 5408 4872
rect 2109 1700 5408 1728
rect -4969 1432 -1670 1460
rect -4969 -1712 -1754 1432
rect -1690 -1712 -1670 1432
rect -4969 -1740 -1670 -1712
rect -1430 1432 1869 1460
rect -1430 -1712 1785 1432
rect 1849 -1712 1869 1432
rect -1430 -1740 1869 -1712
rect 2109 1432 5408 1460
rect 2109 -1712 5324 1432
rect 5388 -1712 5408 1432
rect 2109 -1740 5408 -1712
rect -4969 -2008 -1670 -1980
rect -4969 -5152 -1754 -2008
rect -1690 -5152 -1670 -2008
rect -4969 -5180 -1670 -5152
rect -1430 -2008 1869 -1980
rect -1430 -5152 1785 -2008
rect 1849 -5152 1869 -2008
rect -1430 -5180 1869 -5152
rect 2109 -2008 5408 -1980
rect 2109 -5152 5324 -2008
rect 5388 -5152 5408 -2008
rect 2109 -5180 5408 -5152
<< via3 >>
rect -1754 1728 -1690 4872
rect 1785 1728 1849 4872
rect 5324 1728 5388 4872
rect -1754 -1712 -1690 1432
rect 1785 -1712 1849 1432
rect 5324 -1712 5388 1432
rect -1754 -5152 -1690 -2008
rect 1785 -5152 1849 -2008
rect 5324 -5152 5388 -2008
<< mimcap >>
rect -4869 4760 -1869 4800
rect -4869 1840 -4829 4760
rect -1909 1840 -1869 4760
rect -4869 1800 -1869 1840
rect -1330 4760 1670 4800
rect -1330 1840 -1290 4760
rect 1630 1840 1670 4760
rect -1330 1800 1670 1840
rect 2209 4760 5209 4800
rect 2209 1840 2249 4760
rect 5169 1840 5209 4760
rect 2209 1800 5209 1840
rect -4869 1320 -1869 1360
rect -4869 -1600 -4829 1320
rect -1909 -1600 -1869 1320
rect -4869 -1640 -1869 -1600
rect -1330 1320 1670 1360
rect -1330 -1600 -1290 1320
rect 1630 -1600 1670 1320
rect -1330 -1640 1670 -1600
rect 2209 1320 5209 1360
rect 2209 -1600 2249 1320
rect 5169 -1600 5209 1320
rect 2209 -1640 5209 -1600
rect -4869 -2120 -1869 -2080
rect -4869 -5040 -4829 -2120
rect -1909 -5040 -1869 -2120
rect -4869 -5080 -1869 -5040
rect -1330 -2120 1670 -2080
rect -1330 -5040 -1290 -2120
rect 1630 -5040 1670 -2120
rect -1330 -5080 1670 -5040
rect 2209 -2120 5209 -2080
rect 2209 -5040 2249 -2120
rect 5169 -5040 5209 -2120
rect 2209 -5080 5209 -5040
<< mimcapcontact >>
rect -4829 1840 -1909 4760
rect -1290 1840 1630 4760
rect 2249 1840 5169 4760
rect -4829 -1600 -1909 1320
rect -1290 -1600 1630 1320
rect 2249 -1600 5169 1320
rect -4829 -5040 -1909 -2120
rect -1290 -5040 1630 -2120
rect 2249 -5040 5169 -2120
<< metal4 >>
rect -3421 4761 -3317 4950
rect -1801 4888 -1697 4950
rect -1801 4872 -1674 4888
rect -4830 4760 -1908 4761
rect -4830 1840 -4829 4760
rect -1909 1840 -1908 4760
rect -4830 1839 -1908 1840
rect -3421 1321 -3317 1839
rect -1801 1728 -1754 4872
rect -1690 1728 -1674 4872
rect 118 4761 222 4950
rect 1738 4888 1842 4950
rect 1738 4872 1865 4888
rect -1291 4760 1631 4761
rect -1291 1840 -1290 4760
rect 1630 1840 1631 4760
rect -1291 1839 1631 1840
rect -1801 1712 -1674 1728
rect -1801 1448 -1697 1712
rect -1801 1432 -1674 1448
rect -4830 1320 -1908 1321
rect -4830 -1600 -4829 1320
rect -1909 -1600 -1908 1320
rect -4830 -1601 -1908 -1600
rect -3421 -2119 -3317 -1601
rect -1801 -1712 -1754 1432
rect -1690 -1712 -1674 1432
rect 118 1321 222 1839
rect 1738 1728 1785 4872
rect 1849 1728 1865 4872
rect 3657 4761 3761 4950
rect 5277 4888 5381 4950
rect 5277 4872 5404 4888
rect 2248 4760 5170 4761
rect 2248 1840 2249 4760
rect 5169 1840 5170 4760
rect 2248 1839 5170 1840
rect 1738 1712 1865 1728
rect 1738 1448 1842 1712
rect 1738 1432 1865 1448
rect -1291 1320 1631 1321
rect -1291 -1600 -1290 1320
rect 1630 -1600 1631 1320
rect -1291 -1601 1631 -1600
rect -1801 -1728 -1674 -1712
rect -1801 -1992 -1697 -1728
rect -1801 -2008 -1674 -1992
rect -4830 -2120 -1908 -2119
rect -4830 -5040 -4829 -2120
rect -1909 -5040 -1908 -2120
rect -4830 -5041 -1908 -5040
rect -3421 -5230 -3317 -5041
rect -1801 -5152 -1754 -2008
rect -1690 -5152 -1674 -2008
rect 118 -2119 222 -1601
rect 1738 -1712 1785 1432
rect 1849 -1712 1865 1432
rect 3657 1321 3761 1839
rect 5277 1728 5324 4872
rect 5388 1728 5404 4872
rect 5277 1712 5404 1728
rect 5277 1448 5381 1712
rect 5277 1432 5404 1448
rect 2248 1320 5170 1321
rect 2248 -1600 2249 1320
rect 5169 -1600 5170 1320
rect 2248 -1601 5170 -1600
rect 1738 -1728 1865 -1712
rect 1738 -1992 1842 -1728
rect 1738 -2008 1865 -1992
rect -1291 -2120 1631 -2119
rect -1291 -5040 -1290 -2120
rect 1630 -5040 1631 -2120
rect -1291 -5041 1631 -5040
rect -1801 -5168 -1674 -5152
rect -1801 -5230 -1697 -5168
rect 118 -5230 222 -5041
rect 1738 -5152 1785 -2008
rect 1849 -5152 1865 -2008
rect 3657 -2119 3761 -1601
rect 5277 -1712 5324 1432
rect 5388 -1712 5404 1432
rect 5277 -1728 5404 -1712
rect 5277 -1992 5381 -1728
rect 5277 -2008 5404 -1992
rect 2248 -2120 5170 -2119
rect 2248 -5040 2249 -2120
rect 5169 -5040 5170 -2120
rect 2248 -5041 5170 -5040
rect 1738 -5168 1865 -5152
rect 1738 -5230 1842 -5168
rect 3657 -5230 3761 -5041
rect 5277 -5152 5324 -2008
rect 5388 -5152 5404 -2008
rect 5277 -5168 5404 -5152
rect 5277 -5230 5381 -5168
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1669 1700 4869 4900
string parameters w 15 l 15 val 235.2 carea 1.00 cperi 0.17 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
