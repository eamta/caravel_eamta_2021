magic
tech sky130A
magscale 1 2
timestamp 1614978561
<< nmos >>
rect -15 -90 15 90
<< ndiff >>
rect -73 78 -15 90
rect -73 -78 -61 78
rect -27 -78 -15 78
rect -73 -90 -15 -78
rect 15 78 73 90
rect 15 -78 27 78
rect 61 -78 73 78
rect 15 -90 73 -78
<< ndiffc >>
rect -61 -78 -27 78
rect 27 -78 61 78
<< poly >>
rect -15 90 15 116
rect -15 -116 15 -90
<< locali >>
rect -61 78 -27 94
rect -61 -94 -27 -78
rect 27 78 61 94
rect 27 -94 61 -78
<< viali >>
rect -61 -78 -27 78
rect 27 -78 61 78
<< metal1 >>
rect -67 78 -21 90
rect -67 -78 -61 78
rect -27 -78 -21 78
rect -67 -90 -21 -78
rect 21 78 67 90
rect 21 -78 27 78
rect 61 -78 67 78
rect 21 -90 67 -78
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.9 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
