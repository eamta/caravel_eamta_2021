magic
tech sky130A
magscale 1 2
timestamp 1615311859
<< nmos >>
rect -15 -49 15 49
<< ndiff >>
rect -73 37 -15 49
rect -73 -37 -61 37
rect -27 -37 -15 37
rect -73 -49 -15 -37
rect 15 37 73 49
rect 15 -37 27 37
rect 61 -37 73 37
rect 15 -49 73 -37
<< ndiffc >>
rect -61 -37 -27 37
rect 27 -37 61 37
<< poly >>
rect -15 49 15 75
rect -15 -75 15 -49
<< locali >>
rect -61 37 -27 53
rect -61 -53 -27 -37
rect 27 37 61 53
rect 27 -53 61 -37
<< viali >>
rect -61 -37 -27 37
rect 27 -37 61 37
<< metal1 >>
rect -67 37 -21 49
rect -67 -37 -61 37
rect -27 -37 -21 37
rect -67 -49 -21 -37
rect 21 37 67 49
rect 21 -37 27 37
rect 61 -37 67 37
rect 21 -49 67 -37
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.49 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
