magic
tech sky130A
magscale 1 2
timestamp 1623092848
<< pwell >>
rect -1127 -2085 1127 2085
<< nmos >>
rect -927 -1875 -897 1875
rect -831 -1875 -801 1875
rect -735 -1875 -705 1875
rect -639 -1875 -609 1875
rect -543 -1875 -513 1875
rect -447 -1875 -417 1875
rect -351 -1875 -321 1875
rect -255 -1875 -225 1875
rect -159 -1875 -129 1875
rect -63 -1875 -33 1875
rect 33 -1875 63 1875
rect 129 -1875 159 1875
rect 225 -1875 255 1875
rect 321 -1875 351 1875
rect 417 -1875 447 1875
rect 513 -1875 543 1875
rect 609 -1875 639 1875
rect 705 -1875 735 1875
rect 801 -1875 831 1875
rect 897 -1875 927 1875
<< ndiff >>
rect -989 1863 -927 1875
rect -989 -1863 -977 1863
rect -943 -1863 -927 1863
rect -989 -1875 -927 -1863
rect -897 1863 -831 1875
rect -897 -1863 -881 1863
rect -847 -1863 -831 1863
rect -897 -1875 -831 -1863
rect -801 1863 -735 1875
rect -801 -1863 -785 1863
rect -751 -1863 -735 1863
rect -801 -1875 -735 -1863
rect -705 1863 -639 1875
rect -705 -1863 -689 1863
rect -655 -1863 -639 1863
rect -705 -1875 -639 -1863
rect -609 1863 -543 1875
rect -609 -1863 -593 1863
rect -559 -1863 -543 1863
rect -609 -1875 -543 -1863
rect -513 1863 -447 1875
rect -513 -1863 -497 1863
rect -463 -1863 -447 1863
rect -513 -1875 -447 -1863
rect -417 1863 -351 1875
rect -417 -1863 -401 1863
rect -367 -1863 -351 1863
rect -417 -1875 -351 -1863
rect -321 1863 -255 1875
rect -321 -1863 -305 1863
rect -271 -1863 -255 1863
rect -321 -1875 -255 -1863
rect -225 1863 -159 1875
rect -225 -1863 -209 1863
rect -175 -1863 -159 1863
rect -225 -1875 -159 -1863
rect -129 1863 -63 1875
rect -129 -1863 -113 1863
rect -79 -1863 -63 1863
rect -129 -1875 -63 -1863
rect -33 1863 33 1875
rect -33 -1863 -17 1863
rect 17 -1863 33 1863
rect -33 -1875 33 -1863
rect 63 1863 129 1875
rect 63 -1863 79 1863
rect 113 -1863 129 1863
rect 63 -1875 129 -1863
rect 159 1863 225 1875
rect 159 -1863 175 1863
rect 209 -1863 225 1863
rect 159 -1875 225 -1863
rect 255 1863 321 1875
rect 255 -1863 271 1863
rect 305 -1863 321 1863
rect 255 -1875 321 -1863
rect 351 1863 417 1875
rect 351 -1863 367 1863
rect 401 -1863 417 1863
rect 351 -1875 417 -1863
rect 447 1863 513 1875
rect 447 -1863 463 1863
rect 497 -1863 513 1863
rect 447 -1875 513 -1863
rect 543 1863 609 1875
rect 543 -1863 559 1863
rect 593 -1863 609 1863
rect 543 -1875 609 -1863
rect 639 1863 705 1875
rect 639 -1863 655 1863
rect 689 -1863 705 1863
rect 639 -1875 705 -1863
rect 735 1863 801 1875
rect 735 -1863 751 1863
rect 785 -1863 801 1863
rect 735 -1875 801 -1863
rect 831 1863 897 1875
rect 831 -1863 847 1863
rect 881 -1863 897 1863
rect 831 -1875 897 -1863
rect 927 1863 989 1875
rect 927 -1863 943 1863
rect 977 -1863 989 1863
rect 927 -1875 989 -1863
<< ndiffc >>
rect -977 -1863 -943 1863
rect -881 -1863 -847 1863
rect -785 -1863 -751 1863
rect -689 -1863 -655 1863
rect -593 -1863 -559 1863
rect -497 -1863 -463 1863
rect -401 -1863 -367 1863
rect -305 -1863 -271 1863
rect -209 -1863 -175 1863
rect -113 -1863 -79 1863
rect -17 -1863 17 1863
rect 79 -1863 113 1863
rect 175 -1863 209 1863
rect 271 -1863 305 1863
rect 367 -1863 401 1863
rect 463 -1863 497 1863
rect 559 -1863 593 1863
rect 655 -1863 689 1863
rect 751 -1863 785 1863
rect 847 -1863 881 1863
rect 943 -1863 977 1863
<< psubdiff >>
rect -1091 1953 -1057 2049
rect -1091 -2015 -1057 -1953
rect 1057 -2015 1091 2049
rect -1091 -2049 -995 -2015
rect 995 -2049 1091 -2015
<< psubdiffcont >>
rect -1091 -1953 -1057 1953
rect -995 -2049 995 -2015
<< poly >>
rect -927 1981 945 2017
rect -927 1947 -911 1981
rect 925 1947 945 1981
rect -927 1914 945 1947
rect -927 1875 -897 1914
rect -831 1875 -801 1914
rect -735 1875 -705 1914
rect -639 1875 -609 1914
rect -543 1875 -513 1914
rect -447 1875 -417 1914
rect -351 1875 -321 1914
rect -255 1875 -225 1914
rect -159 1875 -129 1914
rect -63 1875 -33 1914
rect 33 1875 63 1914
rect 129 1875 159 1914
rect 225 1875 255 1914
rect 321 1875 351 1914
rect 417 1875 447 1914
rect 513 1875 543 1914
rect 609 1875 639 1914
rect 705 1875 735 1914
rect 801 1875 831 1914
rect 897 1875 927 1914
rect -927 -1901 -897 -1875
rect -831 -1901 -801 -1875
rect -735 -1901 -705 -1875
rect -639 -1901 -609 -1875
rect -543 -1901 -513 -1875
rect -447 -1901 -417 -1875
rect -351 -1901 -321 -1875
rect -255 -1901 -225 -1875
rect -159 -1901 -129 -1875
rect -63 -1901 -33 -1875
rect 33 -1901 63 -1875
rect 129 -1901 159 -1875
rect 225 -1901 255 -1875
rect 321 -1901 351 -1875
rect 417 -1901 447 -1875
rect 513 -1901 543 -1875
rect 609 -1901 639 -1875
rect 705 -1901 735 -1875
rect 801 -1901 831 -1875
rect 897 -1901 927 -1875
<< polycont >>
rect -911 1947 925 1981
<< locali >>
rect -1091 1953 -1057 2049
rect -927 1983 941 1997
rect -927 1947 -911 1983
rect 925 1947 941 1983
rect -927 1931 941 1947
rect -977 1863 -943 1879
rect -977 -1879 -943 -1863
rect -881 1863 -847 1879
rect -881 -1879 -847 -1863
rect -785 1863 -751 1879
rect -785 -1879 -751 -1863
rect -689 1863 -655 1879
rect -689 -1879 -655 -1863
rect -593 1863 -559 1879
rect -593 -1879 -559 -1863
rect -497 1863 -463 1879
rect -497 -1879 -463 -1863
rect -401 1863 -367 1879
rect -401 -1879 -367 -1863
rect -305 1863 -271 1879
rect -305 -1879 -271 -1863
rect -209 1863 -175 1879
rect -209 -1879 -175 -1863
rect -113 1863 -79 1879
rect -113 -1879 -79 -1863
rect -17 1863 17 1879
rect -17 -1879 17 -1863
rect 79 1863 113 1879
rect 79 -1879 113 -1863
rect 175 1863 209 1879
rect 175 -1879 209 -1863
rect 271 1863 305 1879
rect 271 -1879 305 -1863
rect 367 1863 401 1879
rect 367 -1879 401 -1863
rect 463 1863 497 1879
rect 463 -1879 497 -1863
rect 559 1863 593 1879
rect 559 -1879 593 -1863
rect 655 1863 689 1879
rect 655 -1879 689 -1863
rect 751 1863 785 1879
rect 751 -1879 785 -1863
rect 847 1863 881 1879
rect 847 -1879 881 -1863
rect 943 1863 977 1879
rect 943 -1879 977 -1863
rect -1091 -2015 -1057 -1953
rect 1057 -2015 1091 2049
rect -1091 -2049 -995 -2015
rect 995 -2049 1091 -2015
<< viali >>
rect -911 1981 925 1983
rect -911 1947 925 1981
rect -977 -1863 -943 1863
rect -881 -1863 -847 1863
rect -785 -1863 -751 1863
rect -689 -1863 -655 1863
rect -593 -1863 -559 1863
rect -497 -1863 -463 1863
rect -401 -1863 -367 1863
rect -305 -1863 -271 1863
rect -209 -1863 -175 1863
rect -113 -1863 -79 1863
rect -17 -1863 17 1863
rect 79 -1863 113 1863
rect 175 -1863 209 1863
rect 271 -1863 305 1863
rect 367 -1863 401 1863
rect 463 -1863 497 1863
rect 559 -1863 593 1863
rect 655 -1863 689 1863
rect 751 -1863 785 1863
rect 847 -1863 881 1863
rect 943 -1863 977 1863
<< metal1 >>
rect -927 1983 941 1997
rect -927 1947 -911 1983
rect 925 1947 941 1983
rect -927 1931 941 1947
rect -983 1863 -937 1875
rect -983 -1863 -977 1863
rect -943 -1863 -937 1863
rect -983 -1875 -937 -1863
rect -887 1863 -841 1931
rect -887 -1863 -881 1863
rect -847 -1863 -841 1863
rect -887 -1875 -841 -1863
rect -791 1863 -745 1875
rect -791 -1863 -785 1863
rect -751 -1863 -745 1863
rect -791 -1875 -745 -1863
rect -695 1863 -649 1931
rect -695 -1863 -689 1863
rect -655 -1863 -649 1863
rect -695 -1875 -649 -1863
rect -599 1863 -553 1875
rect -599 -1863 -593 1863
rect -559 -1863 -553 1863
rect -599 -1875 -553 -1863
rect -503 1863 -457 1931
rect -503 -1863 -497 1863
rect -463 -1863 -457 1863
rect -503 -1875 -457 -1863
rect -407 1863 -361 1875
rect -407 -1863 -401 1863
rect -367 -1863 -361 1863
rect -407 -1875 -361 -1863
rect -311 1863 -265 1931
rect -311 -1863 -305 1863
rect -271 -1863 -265 1863
rect -311 -1875 -265 -1863
rect -215 1863 -169 1875
rect -215 -1863 -209 1863
rect -175 -1863 -169 1863
rect -215 -1875 -169 -1863
rect -119 1863 -73 1931
rect -119 -1863 -113 1863
rect -79 -1863 -73 1863
rect -119 -1875 -73 -1863
rect -23 1863 23 1875
rect -23 -1863 -17 1863
rect 17 -1863 23 1863
rect -23 -1875 23 -1863
rect 73 1863 119 1931
rect 73 -1863 79 1863
rect 113 -1863 119 1863
rect 73 -1875 119 -1863
rect 169 1863 215 1875
rect 169 -1863 175 1863
rect 209 -1863 215 1863
rect 169 -1875 215 -1863
rect 265 1863 311 1931
rect 265 -1863 271 1863
rect 305 -1863 311 1863
rect 265 -1875 311 -1863
rect 361 1863 407 1875
rect 361 -1863 367 1863
rect 401 -1863 407 1863
rect 361 -1875 407 -1863
rect 457 1863 503 1931
rect 457 -1863 463 1863
rect 497 -1863 503 1863
rect 457 -1875 503 -1863
rect 553 1863 599 1875
rect 553 -1863 559 1863
rect 593 -1863 599 1863
rect 553 -1875 599 -1863
rect 649 1863 695 1931
rect 649 -1863 655 1863
rect 689 -1863 695 1863
rect 649 -1875 695 -1863
rect 745 1863 791 1875
rect 745 -1863 751 1863
rect 785 -1863 791 1863
rect 745 -1875 791 -1863
rect 841 1863 887 1931
rect 841 -1863 847 1863
rect 881 -1863 887 1863
rect 841 -1875 887 -1863
rect 937 1863 983 1875
rect 937 -1863 943 1863
rect 977 -1863 983 1863
rect 937 -1875 983 -1863
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -2032 1074 2032
string parameters w 18.75 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
