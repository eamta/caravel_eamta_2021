magic
tech sky130A
magscale 1 2
timestamp 1615944125
<< error_p >>
rect -1445 341 -1387 347
rect -1327 341 -1269 347
rect -1209 341 -1151 347
rect -1091 341 -1033 347
rect -973 341 -915 347
rect -855 341 -797 347
rect -737 341 -679 347
rect -619 341 -561 347
rect -501 341 -443 347
rect -383 341 -325 347
rect -265 341 -207 347
rect -147 341 -89 347
rect -29 341 29 347
rect 89 341 147 347
rect 207 341 265 347
rect 325 341 383 347
rect 443 341 501 347
rect 561 341 619 347
rect 679 341 737 347
rect 797 341 855 347
rect 915 341 973 347
rect 1033 341 1091 347
rect 1151 341 1209 347
rect 1269 341 1327 347
rect 1387 341 1445 347
rect -1445 307 -1433 341
rect -1327 307 -1315 341
rect -1209 307 -1197 341
rect -1091 307 -1079 341
rect -973 307 -961 341
rect -855 307 -843 341
rect -737 307 -725 341
rect -619 307 -607 341
rect -501 307 -489 341
rect -383 307 -371 341
rect -265 307 -253 341
rect -147 307 -135 341
rect -29 307 -17 341
rect 89 307 101 341
rect 207 307 219 341
rect 325 307 337 341
rect 443 307 455 341
rect 561 307 573 341
rect 679 307 691 341
rect 797 307 809 341
rect 915 307 927 341
rect 1033 307 1045 341
rect 1151 307 1163 341
rect 1269 307 1281 341
rect 1387 307 1399 341
rect -1445 301 -1387 307
rect -1327 301 -1269 307
rect -1209 301 -1151 307
rect -1091 301 -1033 307
rect -973 301 -915 307
rect -855 301 -797 307
rect -737 301 -679 307
rect -619 301 -561 307
rect -501 301 -443 307
rect -383 301 -325 307
rect -265 301 -207 307
rect -147 301 -89 307
rect -29 301 29 307
rect 89 301 147 307
rect 207 301 265 307
rect 325 301 383 307
rect 443 301 501 307
rect 561 301 619 307
rect 679 301 737 307
rect 797 301 855 307
rect 915 301 973 307
rect 1033 301 1091 307
rect 1151 301 1209 307
rect 1269 301 1327 307
rect 1387 301 1445 307
<< pwell >>
rect -1642 -479 1642 479
<< nmos >>
rect -1446 -331 -1386 269
rect -1328 -331 -1268 269
rect -1210 -331 -1150 269
rect -1092 -331 -1032 269
rect -974 -331 -914 269
rect -856 -331 -796 269
rect -738 -331 -678 269
rect -620 -331 -560 269
rect -502 -331 -442 269
rect -384 -331 -324 269
rect -266 -331 -206 269
rect -148 -331 -88 269
rect -30 -331 30 269
rect 88 -331 148 269
rect 206 -331 266 269
rect 324 -331 384 269
rect 442 -331 502 269
rect 560 -331 620 269
rect 678 -331 738 269
rect 796 -331 856 269
rect 914 -331 974 269
rect 1032 -331 1092 269
rect 1150 -331 1210 269
rect 1268 -331 1328 269
rect 1386 -331 1446 269
<< ndiff >>
rect -1504 257 -1446 269
rect -1504 -319 -1492 257
rect -1458 -319 -1446 257
rect -1504 -331 -1446 -319
rect -1386 257 -1328 269
rect -1386 -319 -1374 257
rect -1340 -319 -1328 257
rect -1386 -331 -1328 -319
rect -1268 257 -1210 269
rect -1268 -319 -1256 257
rect -1222 -319 -1210 257
rect -1268 -331 -1210 -319
rect -1150 257 -1092 269
rect -1150 -319 -1138 257
rect -1104 -319 -1092 257
rect -1150 -331 -1092 -319
rect -1032 257 -974 269
rect -1032 -319 -1020 257
rect -986 -319 -974 257
rect -1032 -331 -974 -319
rect -914 257 -856 269
rect -914 -319 -902 257
rect -868 -319 -856 257
rect -914 -331 -856 -319
rect -796 257 -738 269
rect -796 -319 -784 257
rect -750 -319 -738 257
rect -796 -331 -738 -319
rect -678 257 -620 269
rect -678 -319 -666 257
rect -632 -319 -620 257
rect -678 -331 -620 -319
rect -560 257 -502 269
rect -560 -319 -548 257
rect -514 -319 -502 257
rect -560 -331 -502 -319
rect -442 257 -384 269
rect -442 -319 -430 257
rect -396 -319 -384 257
rect -442 -331 -384 -319
rect -324 257 -266 269
rect -324 -319 -312 257
rect -278 -319 -266 257
rect -324 -331 -266 -319
rect -206 257 -148 269
rect -206 -319 -194 257
rect -160 -319 -148 257
rect -206 -331 -148 -319
rect -88 257 -30 269
rect -88 -319 -76 257
rect -42 -319 -30 257
rect -88 -331 -30 -319
rect 30 257 88 269
rect 30 -319 42 257
rect 76 -319 88 257
rect 30 -331 88 -319
rect 148 257 206 269
rect 148 -319 160 257
rect 194 -319 206 257
rect 148 -331 206 -319
rect 266 257 324 269
rect 266 -319 278 257
rect 312 -319 324 257
rect 266 -331 324 -319
rect 384 257 442 269
rect 384 -319 396 257
rect 430 -319 442 257
rect 384 -331 442 -319
rect 502 257 560 269
rect 502 -319 514 257
rect 548 -319 560 257
rect 502 -331 560 -319
rect 620 257 678 269
rect 620 -319 632 257
rect 666 -319 678 257
rect 620 -331 678 -319
rect 738 257 796 269
rect 738 -319 750 257
rect 784 -319 796 257
rect 738 -331 796 -319
rect 856 257 914 269
rect 856 -319 868 257
rect 902 -319 914 257
rect 856 -331 914 -319
rect 974 257 1032 269
rect 974 -319 986 257
rect 1020 -319 1032 257
rect 974 -331 1032 -319
rect 1092 257 1150 269
rect 1092 -319 1104 257
rect 1138 -319 1150 257
rect 1092 -331 1150 -319
rect 1210 257 1268 269
rect 1210 -319 1222 257
rect 1256 -319 1268 257
rect 1210 -331 1268 -319
rect 1328 257 1386 269
rect 1328 -319 1340 257
rect 1374 -319 1386 257
rect 1328 -331 1386 -319
rect 1446 257 1504 269
rect 1446 -319 1458 257
rect 1492 -319 1504 257
rect 1446 -331 1504 -319
<< ndiffc >>
rect -1492 -319 -1458 257
rect -1374 -319 -1340 257
rect -1256 -319 -1222 257
rect -1138 -319 -1104 257
rect -1020 -319 -986 257
rect -902 -319 -868 257
rect -784 -319 -750 257
rect -666 -319 -632 257
rect -548 -319 -514 257
rect -430 -319 -396 257
rect -312 -319 -278 257
rect -194 -319 -160 257
rect -76 -319 -42 257
rect 42 -319 76 257
rect 160 -319 194 257
rect 278 -319 312 257
rect 396 -319 430 257
rect 514 -319 548 257
rect 632 -319 666 257
rect 750 -319 784 257
rect 868 -319 902 257
rect 986 -319 1020 257
rect 1104 -319 1138 257
rect 1222 -319 1256 257
rect 1340 -319 1374 257
rect 1458 -319 1492 257
<< psubdiff >>
rect -1606 409 -1510 443
rect 1510 409 1606 443
rect -1606 347 -1572 409
rect 1572 347 1606 409
rect -1606 -409 -1572 -347
rect 1572 -409 1606 -347
rect -1606 -443 -1510 -409
rect 1510 -443 1606 -409
<< psubdiffcont >>
rect -1510 409 1510 443
rect -1606 -347 -1572 347
rect 1572 -347 1606 347
rect -1510 -443 1510 -409
<< poly >>
rect -1449 341 -1383 357
rect -1449 307 -1433 341
rect -1399 307 -1383 341
rect -1449 291 -1383 307
rect -1331 341 -1265 357
rect -1331 307 -1315 341
rect -1281 307 -1265 341
rect -1331 291 -1265 307
rect -1213 341 -1147 357
rect -1213 307 -1197 341
rect -1163 307 -1147 341
rect -1213 291 -1147 307
rect -1095 341 -1029 357
rect -1095 307 -1079 341
rect -1045 307 -1029 341
rect -1095 291 -1029 307
rect -977 341 -911 357
rect -977 307 -961 341
rect -927 307 -911 341
rect -977 291 -911 307
rect -859 341 -793 357
rect -859 307 -843 341
rect -809 307 -793 341
rect -859 291 -793 307
rect -741 341 -675 357
rect -741 307 -725 341
rect -691 307 -675 341
rect -741 291 -675 307
rect -623 341 -557 357
rect -623 307 -607 341
rect -573 307 -557 341
rect -623 291 -557 307
rect -505 341 -439 357
rect -505 307 -489 341
rect -455 307 -439 341
rect -505 291 -439 307
rect -387 341 -321 357
rect -387 307 -371 341
rect -337 307 -321 341
rect -387 291 -321 307
rect -269 341 -203 357
rect -269 307 -253 341
rect -219 307 -203 341
rect -269 291 -203 307
rect -151 341 -85 357
rect -151 307 -135 341
rect -101 307 -85 341
rect -151 291 -85 307
rect -33 341 33 357
rect -33 307 -17 341
rect 17 307 33 341
rect -33 291 33 307
rect 85 341 151 357
rect 85 307 101 341
rect 135 307 151 341
rect 85 291 151 307
rect 203 341 269 357
rect 203 307 219 341
rect 253 307 269 341
rect 203 291 269 307
rect 321 341 387 357
rect 321 307 337 341
rect 371 307 387 341
rect 321 291 387 307
rect 439 341 505 357
rect 439 307 455 341
rect 489 307 505 341
rect 439 291 505 307
rect 557 341 623 357
rect 557 307 573 341
rect 607 307 623 341
rect 557 291 623 307
rect 675 341 741 357
rect 675 307 691 341
rect 725 307 741 341
rect 675 291 741 307
rect 793 341 859 357
rect 793 307 809 341
rect 843 307 859 341
rect 793 291 859 307
rect 911 341 977 357
rect 911 307 927 341
rect 961 307 977 341
rect 911 291 977 307
rect 1029 341 1095 357
rect 1029 307 1045 341
rect 1079 307 1095 341
rect 1029 291 1095 307
rect 1147 341 1213 357
rect 1147 307 1163 341
rect 1197 307 1213 341
rect 1147 291 1213 307
rect 1265 341 1331 357
rect 1265 307 1281 341
rect 1315 307 1331 341
rect 1265 291 1331 307
rect 1383 341 1449 357
rect 1383 307 1399 341
rect 1433 307 1449 341
rect 1383 291 1449 307
rect -1446 269 -1386 291
rect -1328 269 -1268 291
rect -1210 269 -1150 291
rect -1092 269 -1032 291
rect -974 269 -914 291
rect -856 269 -796 291
rect -738 269 -678 291
rect -620 269 -560 291
rect -502 269 -442 291
rect -384 269 -324 291
rect -266 269 -206 291
rect -148 269 -88 291
rect -30 269 30 291
rect 88 269 148 291
rect 206 269 266 291
rect 324 269 384 291
rect 442 269 502 291
rect 560 269 620 291
rect 678 269 738 291
rect 796 269 856 291
rect 914 269 974 291
rect 1032 269 1092 291
rect 1150 269 1210 291
rect 1268 269 1328 291
rect 1386 269 1446 291
rect -1446 -357 -1386 -331
rect -1328 -357 -1268 -331
rect -1210 -357 -1150 -331
rect -1092 -357 -1032 -331
rect -974 -357 -914 -331
rect -856 -357 -796 -331
rect -738 -357 -678 -331
rect -620 -357 -560 -331
rect -502 -357 -442 -331
rect -384 -357 -324 -331
rect -266 -357 -206 -331
rect -148 -357 -88 -331
rect -30 -357 30 -331
rect 88 -357 148 -331
rect 206 -357 266 -331
rect 324 -357 384 -331
rect 442 -357 502 -331
rect 560 -357 620 -331
rect 678 -357 738 -331
rect 796 -357 856 -331
rect 914 -357 974 -331
rect 1032 -357 1092 -331
rect 1150 -357 1210 -331
rect 1268 -357 1328 -331
rect 1386 -357 1446 -331
<< polycont >>
rect -1433 307 -1399 341
rect -1315 307 -1281 341
rect -1197 307 -1163 341
rect -1079 307 -1045 341
rect -961 307 -927 341
rect -843 307 -809 341
rect -725 307 -691 341
rect -607 307 -573 341
rect -489 307 -455 341
rect -371 307 -337 341
rect -253 307 -219 341
rect -135 307 -101 341
rect -17 307 17 341
rect 101 307 135 341
rect 219 307 253 341
rect 337 307 371 341
rect 455 307 489 341
rect 573 307 607 341
rect 691 307 725 341
rect 809 307 843 341
rect 927 307 961 341
rect 1045 307 1079 341
rect 1163 307 1197 341
rect 1281 307 1315 341
rect 1399 307 1433 341
<< locali >>
rect -1606 409 -1510 443
rect 1510 409 1606 443
rect -1606 347 -1572 409
rect 1572 347 1606 409
rect -1449 307 -1433 341
rect -1399 307 -1383 341
rect -1331 307 -1315 341
rect -1281 307 -1265 341
rect -1213 307 -1197 341
rect -1163 307 -1147 341
rect -1095 307 -1079 341
rect -1045 307 -1029 341
rect -977 307 -961 341
rect -927 307 -911 341
rect -859 307 -843 341
rect -809 307 -793 341
rect -741 307 -725 341
rect -691 307 -675 341
rect -623 307 -607 341
rect -573 307 -557 341
rect -505 307 -489 341
rect -455 307 -439 341
rect -387 307 -371 341
rect -337 307 -321 341
rect -269 307 -253 341
rect -219 307 -203 341
rect -151 307 -135 341
rect -101 307 -85 341
rect -33 307 -17 341
rect 17 307 33 341
rect 85 307 101 341
rect 135 307 151 341
rect 203 307 219 341
rect 253 307 269 341
rect 321 307 337 341
rect 371 307 387 341
rect 439 307 455 341
rect 489 307 505 341
rect 557 307 573 341
rect 607 307 623 341
rect 675 307 691 341
rect 725 307 741 341
rect 793 307 809 341
rect 843 307 859 341
rect 911 307 927 341
rect 961 307 977 341
rect 1029 307 1045 341
rect 1079 307 1095 341
rect 1147 307 1163 341
rect 1197 307 1213 341
rect 1265 307 1281 341
rect 1315 307 1331 341
rect 1383 307 1399 341
rect 1433 307 1449 341
rect -1492 257 -1458 273
rect -1492 -335 -1458 -319
rect -1374 257 -1340 273
rect -1374 -335 -1340 -319
rect -1256 257 -1222 273
rect -1256 -335 -1222 -319
rect -1138 257 -1104 273
rect -1138 -335 -1104 -319
rect -1020 257 -986 273
rect -1020 -335 -986 -319
rect -902 257 -868 273
rect -902 -335 -868 -319
rect -784 257 -750 273
rect -784 -335 -750 -319
rect -666 257 -632 273
rect -666 -335 -632 -319
rect -548 257 -514 273
rect -548 -335 -514 -319
rect -430 257 -396 273
rect -430 -335 -396 -319
rect -312 257 -278 273
rect -312 -335 -278 -319
rect -194 257 -160 273
rect -194 -335 -160 -319
rect -76 257 -42 273
rect -76 -335 -42 -319
rect 42 257 76 273
rect 42 -335 76 -319
rect 160 257 194 273
rect 160 -335 194 -319
rect 278 257 312 273
rect 278 -335 312 -319
rect 396 257 430 273
rect 396 -335 430 -319
rect 514 257 548 273
rect 514 -335 548 -319
rect 632 257 666 273
rect 632 -335 666 -319
rect 750 257 784 273
rect 750 -335 784 -319
rect 868 257 902 273
rect 868 -335 902 -319
rect 986 257 1020 273
rect 986 -335 1020 -319
rect 1104 257 1138 273
rect 1104 -335 1138 -319
rect 1222 257 1256 273
rect 1222 -335 1256 -319
rect 1340 257 1374 273
rect 1340 -335 1374 -319
rect 1458 257 1492 273
rect 1458 -335 1492 -319
rect -1606 -409 -1572 -347
rect 1572 -409 1606 -347
rect -1606 -443 -1510 -409
rect 1510 -443 1606 -409
<< viali >>
rect -1433 307 -1399 341
rect -1315 307 -1281 341
rect -1197 307 -1163 341
rect -1079 307 -1045 341
rect -961 307 -927 341
rect -843 307 -809 341
rect -725 307 -691 341
rect -607 307 -573 341
rect -489 307 -455 341
rect -371 307 -337 341
rect -253 307 -219 341
rect -135 307 -101 341
rect -17 307 17 341
rect 101 307 135 341
rect 219 307 253 341
rect 337 307 371 341
rect 455 307 489 341
rect 573 307 607 341
rect 691 307 725 341
rect 809 307 843 341
rect 927 307 961 341
rect 1045 307 1079 341
rect 1163 307 1197 341
rect 1281 307 1315 341
rect 1399 307 1433 341
rect -1492 -319 -1458 257
rect -1374 -319 -1340 257
rect -1256 -319 -1222 257
rect -1138 -319 -1104 257
rect -1020 -319 -986 257
rect -902 -319 -868 257
rect -784 -319 -750 257
rect -666 -319 -632 257
rect -548 -319 -514 257
rect -430 -319 -396 257
rect -312 -319 -278 257
rect -194 -319 -160 257
rect -76 -319 -42 257
rect 42 -319 76 257
rect 160 -319 194 257
rect 278 -319 312 257
rect 396 -319 430 257
rect 514 -319 548 257
rect 632 -319 666 257
rect 750 -319 784 257
rect 868 -319 902 257
rect 986 -319 1020 257
rect 1104 -319 1138 257
rect 1222 -319 1256 257
rect 1340 -319 1374 257
rect 1458 -319 1492 257
<< metal1 >>
rect -1445 341 -1387 347
rect -1445 307 -1433 341
rect -1399 307 -1387 341
rect -1445 301 -1387 307
rect -1327 341 -1269 347
rect -1327 307 -1315 341
rect -1281 307 -1269 341
rect -1327 301 -1269 307
rect -1209 341 -1151 347
rect -1209 307 -1197 341
rect -1163 307 -1151 341
rect -1209 301 -1151 307
rect -1091 341 -1033 347
rect -1091 307 -1079 341
rect -1045 307 -1033 341
rect -1091 301 -1033 307
rect -973 341 -915 347
rect -973 307 -961 341
rect -927 307 -915 341
rect -973 301 -915 307
rect -855 341 -797 347
rect -855 307 -843 341
rect -809 307 -797 341
rect -855 301 -797 307
rect -737 341 -679 347
rect -737 307 -725 341
rect -691 307 -679 341
rect -737 301 -679 307
rect -619 341 -561 347
rect -619 307 -607 341
rect -573 307 -561 341
rect -619 301 -561 307
rect -501 341 -443 347
rect -501 307 -489 341
rect -455 307 -443 341
rect -501 301 -443 307
rect -383 341 -325 347
rect -383 307 -371 341
rect -337 307 -325 341
rect -383 301 -325 307
rect -265 341 -207 347
rect -265 307 -253 341
rect -219 307 -207 341
rect -265 301 -207 307
rect -147 341 -89 347
rect -147 307 -135 341
rect -101 307 -89 341
rect -147 301 -89 307
rect -29 341 29 347
rect -29 307 -17 341
rect 17 307 29 341
rect -29 301 29 307
rect 89 341 147 347
rect 89 307 101 341
rect 135 307 147 341
rect 89 301 147 307
rect 207 341 265 347
rect 207 307 219 341
rect 253 307 265 341
rect 207 301 265 307
rect 325 341 383 347
rect 325 307 337 341
rect 371 307 383 341
rect 325 301 383 307
rect 443 341 501 347
rect 443 307 455 341
rect 489 307 501 341
rect 443 301 501 307
rect 561 341 619 347
rect 561 307 573 341
rect 607 307 619 341
rect 561 301 619 307
rect 679 341 737 347
rect 679 307 691 341
rect 725 307 737 341
rect 679 301 737 307
rect 797 341 855 347
rect 797 307 809 341
rect 843 307 855 341
rect 797 301 855 307
rect 915 341 973 347
rect 915 307 927 341
rect 961 307 973 341
rect 915 301 973 307
rect 1033 341 1091 347
rect 1033 307 1045 341
rect 1079 307 1091 341
rect 1033 301 1091 307
rect 1151 341 1209 347
rect 1151 307 1163 341
rect 1197 307 1209 341
rect 1151 301 1209 307
rect 1269 341 1327 347
rect 1269 307 1281 341
rect 1315 307 1327 341
rect 1269 301 1327 307
rect 1387 341 1445 347
rect 1387 307 1399 341
rect 1433 307 1445 341
rect 1387 301 1445 307
rect -1498 257 -1452 269
rect -1498 -319 -1492 257
rect -1458 -319 -1452 257
rect -1498 -331 -1452 -319
rect -1380 257 -1334 269
rect -1380 -319 -1374 257
rect -1340 -319 -1334 257
rect -1380 -331 -1334 -319
rect -1262 257 -1216 269
rect -1262 -319 -1256 257
rect -1222 -319 -1216 257
rect -1262 -331 -1216 -319
rect -1144 257 -1098 269
rect -1144 -319 -1138 257
rect -1104 -319 -1098 257
rect -1144 -331 -1098 -319
rect -1026 257 -980 269
rect -1026 -319 -1020 257
rect -986 -319 -980 257
rect -1026 -331 -980 -319
rect -908 257 -862 269
rect -908 -319 -902 257
rect -868 -319 -862 257
rect -908 -331 -862 -319
rect -790 257 -744 269
rect -790 -319 -784 257
rect -750 -319 -744 257
rect -790 -331 -744 -319
rect -672 257 -626 269
rect -672 -319 -666 257
rect -632 -319 -626 257
rect -672 -331 -626 -319
rect -554 257 -508 269
rect -554 -319 -548 257
rect -514 -319 -508 257
rect -554 -331 -508 -319
rect -436 257 -390 269
rect -436 -319 -430 257
rect -396 -319 -390 257
rect -436 -331 -390 -319
rect -318 257 -272 269
rect -318 -319 -312 257
rect -278 -319 -272 257
rect -318 -331 -272 -319
rect -200 257 -154 269
rect -200 -319 -194 257
rect -160 -319 -154 257
rect -200 -331 -154 -319
rect -82 257 -36 269
rect -82 -319 -76 257
rect -42 -319 -36 257
rect -82 -331 -36 -319
rect 36 257 82 269
rect 36 -319 42 257
rect 76 -319 82 257
rect 36 -331 82 -319
rect 154 257 200 269
rect 154 -319 160 257
rect 194 -319 200 257
rect 154 -331 200 -319
rect 272 257 318 269
rect 272 -319 278 257
rect 312 -319 318 257
rect 272 -331 318 -319
rect 390 257 436 269
rect 390 -319 396 257
rect 430 -319 436 257
rect 390 -331 436 -319
rect 508 257 554 269
rect 508 -319 514 257
rect 548 -319 554 257
rect 508 -331 554 -319
rect 626 257 672 269
rect 626 -319 632 257
rect 666 -319 672 257
rect 626 -331 672 -319
rect 744 257 790 269
rect 744 -319 750 257
rect 784 -319 790 257
rect 744 -331 790 -319
rect 862 257 908 269
rect 862 -319 868 257
rect 902 -319 908 257
rect 862 -331 908 -319
rect 980 257 1026 269
rect 980 -319 986 257
rect 1020 -319 1026 257
rect 980 -331 1026 -319
rect 1098 257 1144 269
rect 1098 -319 1104 257
rect 1138 -319 1144 257
rect 1098 -331 1144 -319
rect 1216 257 1262 269
rect 1216 -319 1222 257
rect 1256 -319 1262 257
rect 1216 -331 1262 -319
rect 1334 257 1380 269
rect 1334 -319 1340 257
rect 1374 -319 1380 257
rect 1334 -331 1380 -319
rect 1452 257 1498 269
rect 1452 -319 1458 257
rect 1492 -319 1498 257
rect 1452 -331 1498 -319
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1589 -426 1589 426
string parameters w 3 l 0.3 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
