magic
tech sky130A
magscale 1 2
timestamp 1619042384
<< pwell >>
rect -839 -360 839 360
<< nmos >>
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
<< ndiff >>
rect -701 138 -639 150
rect -701 -138 -689 138
rect -655 -138 -639 138
rect -701 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 701 150
rect 639 -138 655 138
rect 689 -138 701 138
rect 639 -150 701 -138
<< ndiffc >>
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
<< psubdiff >>
rect -803 290 -707 324
rect 707 290 803 324
rect -803 228 -769 290
rect 769 228 803 290
rect -803 -290 -769 -228
rect 769 -290 803 -228
rect -803 -324 -707 -290
rect 707 -324 803 -290
<< psubdiffcont >>
rect -707 290 707 324
rect -803 -228 -769 228
rect 769 -228 803 228
rect -707 -324 707 -290
<< poly >>
rect -639 225 639 238
rect -639 191 -593 225
rect 582 191 639 225
rect -639 172 639 191
rect -639 150 -609 172
rect -543 150 -513 172
rect -447 150 -417 172
rect -351 150 -321 172
rect -255 150 -225 172
rect -159 150 -129 172
rect -63 150 -33 172
rect 33 150 63 172
rect 129 150 159 172
rect 225 150 255 172
rect 321 150 351 172
rect 417 150 447 172
rect 513 150 543 172
rect 609 150 639 172
rect -639 -178 -609 -150
rect -543 -176 -513 -150
rect -447 -178 -417 -150
rect -351 -176 -321 -150
rect -255 -178 -225 -150
rect -159 -176 -129 -150
rect -63 -178 -33 -150
rect 33 -176 63 -150
rect 129 -178 159 -150
rect 225 -176 255 -150
rect 321 -178 351 -150
rect 417 -176 447 -150
rect 513 -178 543 -150
rect 609 -176 639 -150
<< polycont >>
rect -593 191 582 225
<< locali >>
rect -803 290 -707 324
rect 707 290 803 324
rect -803 228 -769 290
rect 769 228 803 290
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect -803 -290 -769 -228
rect 769 -290 803 -228
rect -803 -324 -707 -290
rect 707 -324 803 -290
<< viali >>
rect -621 225 612 226
rect -621 191 -593 225
rect -593 191 582 225
rect 582 191 612 225
rect -621 190 612 191
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
<< metal1 >>
rect -633 226 624 232
rect -633 190 -621 226
rect 612 190 624 226
rect -633 184 624 190
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -786 -307 786 307
string parameters w 1.5 l 0.150 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
