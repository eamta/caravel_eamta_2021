magic
tech sky130A
magscale 1 2
timestamp 1623019696
<< error_p >>
rect -845 972 -787 978
rect -653 972 -595 978
rect -461 972 -403 978
rect -269 972 -211 978
rect -77 972 -19 978
rect 115 972 173 978
rect 307 972 365 978
rect 499 972 557 978
rect 691 972 749 978
rect 883 972 941 978
rect -845 938 -833 972
rect -653 938 -641 972
rect -461 938 -449 972
rect -269 938 -257 972
rect -77 938 -65 972
rect 115 938 127 972
rect 307 938 319 972
rect 499 938 511 972
rect 691 938 703 972
rect 883 938 895 972
rect -845 932 -787 938
rect -653 932 -595 938
rect -461 932 -403 938
rect -269 932 -211 938
rect -77 932 -19 938
rect 115 932 173 938
rect 307 932 365 938
rect 499 932 557 938
rect 691 932 749 938
rect 883 932 941 938
rect -941 -938 -883 -932
rect -749 -938 -691 -932
rect -557 -938 -499 -932
rect -365 -938 -307 -932
rect -173 -938 -115 -932
rect 19 -938 77 -932
rect 211 -938 269 -932
rect 403 -938 461 -932
rect 595 -938 653 -932
rect 787 -938 845 -932
rect -941 -972 -929 -938
rect -749 -972 -737 -938
rect -557 -972 -545 -938
rect -365 -972 -353 -938
rect -173 -972 -161 -938
rect 19 -972 31 -938
rect 211 -972 223 -938
rect 403 -972 415 -938
rect 595 -972 607 -938
rect 787 -972 799 -938
rect -941 -978 -883 -972
rect -749 -978 -691 -972
rect -557 -978 -499 -972
rect -365 -978 -307 -972
rect -173 -978 -115 -972
rect 19 -978 77 -972
rect 211 -978 269 -972
rect 403 -978 461 -972
rect 595 -978 653 -972
rect 787 -978 845 -972
<< pwell >>
rect -1127 -1110 1127 1110
<< nmos >>
rect -927 -900 -897 900
rect -831 -900 -801 900
rect -735 -900 -705 900
rect -639 -900 -609 900
rect -543 -900 -513 900
rect -447 -900 -417 900
rect -351 -900 -321 900
rect -255 -900 -225 900
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
rect 225 -900 255 900
rect 321 -900 351 900
rect 417 -900 447 900
rect 513 -900 543 900
rect 609 -900 639 900
rect 705 -900 735 900
rect 801 -900 831 900
rect 897 -900 927 900
<< ndiff >>
rect -989 888 -927 900
rect -989 -888 -977 888
rect -943 -888 -927 888
rect -989 -900 -927 -888
rect -897 888 -831 900
rect -897 -888 -881 888
rect -847 -888 -831 888
rect -897 -900 -831 -888
rect -801 888 -735 900
rect -801 -888 -785 888
rect -751 -888 -735 888
rect -801 -900 -735 -888
rect -705 888 -639 900
rect -705 -888 -689 888
rect -655 -888 -639 888
rect -705 -900 -639 -888
rect -609 888 -543 900
rect -609 -888 -593 888
rect -559 -888 -543 888
rect -609 -900 -543 -888
rect -513 888 -447 900
rect -513 -888 -497 888
rect -463 -888 -447 888
rect -513 -900 -447 -888
rect -417 888 -351 900
rect -417 -888 -401 888
rect -367 -888 -351 888
rect -417 -900 -351 -888
rect -321 888 -255 900
rect -321 -888 -305 888
rect -271 -888 -255 888
rect -321 -900 -255 -888
rect -225 888 -159 900
rect -225 -888 -209 888
rect -175 -888 -159 888
rect -225 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 225 900
rect 159 -888 175 888
rect 209 -888 225 888
rect 159 -900 225 -888
rect 255 888 321 900
rect 255 -888 271 888
rect 305 -888 321 888
rect 255 -900 321 -888
rect 351 888 417 900
rect 351 -888 367 888
rect 401 -888 417 888
rect 351 -900 417 -888
rect 447 888 513 900
rect 447 -888 463 888
rect 497 -888 513 888
rect 447 -900 513 -888
rect 543 888 609 900
rect 543 -888 559 888
rect 593 -888 609 888
rect 543 -900 609 -888
rect 639 888 705 900
rect 639 -888 655 888
rect 689 -888 705 888
rect 639 -900 705 -888
rect 735 888 801 900
rect 735 -888 751 888
rect 785 -888 801 888
rect 735 -900 801 -888
rect 831 888 897 900
rect 831 -888 847 888
rect 881 -888 897 888
rect 831 -900 897 -888
rect 927 888 989 900
rect 927 -888 943 888
rect 977 -888 989 888
rect 927 -900 989 -888
<< ndiffc >>
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
<< psubdiff >>
rect -1091 1040 -995 1074
rect 995 1040 1091 1074
rect -1091 978 -1057 1040
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1040
rect -1091 -1074 1091 -1040
<< psubdiffcont >>
rect -995 1040 995 1074
rect -1091 -978 -1057 978
<< poly >>
rect -849 972 -783 988
rect -849 938 -833 972
rect -799 938 -783 972
rect -927 900 -897 926
rect -849 922 -783 938
rect -657 972 -591 988
rect -657 938 -641 972
rect -607 938 -591 972
rect -831 900 -801 922
rect -735 900 -705 926
rect -657 922 -591 938
rect -465 972 -399 988
rect -465 938 -449 972
rect -415 938 -399 972
rect -639 900 -609 922
rect -543 900 -513 926
rect -465 922 -399 938
rect -273 972 -207 988
rect -273 938 -257 972
rect -223 938 -207 972
rect -447 900 -417 922
rect -351 900 -321 926
rect -273 922 -207 938
rect -81 972 -15 988
rect -81 938 -65 972
rect -31 938 -15 972
rect -255 900 -225 922
rect -159 900 -129 926
rect -81 922 -15 938
rect 111 972 177 988
rect 111 938 127 972
rect 161 938 177 972
rect -63 900 -33 922
rect 33 900 63 926
rect 111 922 177 938
rect 303 972 369 988
rect 303 938 319 972
rect 353 938 369 972
rect 129 900 159 922
rect 225 900 255 926
rect 303 922 369 938
rect 495 972 561 988
rect 495 938 511 972
rect 545 938 561 972
rect 321 900 351 922
rect 417 900 447 926
rect 495 922 561 938
rect 687 972 753 988
rect 687 938 703 972
rect 737 938 753 972
rect 513 900 543 922
rect 609 900 639 926
rect 687 922 753 938
rect 879 972 945 988
rect 879 938 895 972
rect 929 938 945 972
rect 705 900 735 922
rect 801 900 831 926
rect 879 922 945 938
rect 897 900 927 922
rect -927 -922 -897 -900
rect -945 -938 -879 -922
rect -831 -926 -801 -900
rect -735 -922 -705 -900
rect -945 -972 -929 -938
rect -895 -972 -879 -938
rect -945 -988 -879 -972
rect -753 -938 -687 -922
rect -639 -926 -609 -900
rect -543 -922 -513 -900
rect -753 -972 -737 -938
rect -703 -972 -687 -938
rect -753 -988 -687 -972
rect -561 -938 -495 -922
rect -447 -926 -417 -900
rect -351 -922 -321 -900
rect -561 -972 -545 -938
rect -511 -972 -495 -938
rect -561 -988 -495 -972
rect -369 -938 -303 -922
rect -255 -926 -225 -900
rect -159 -922 -129 -900
rect -369 -972 -353 -938
rect -319 -972 -303 -938
rect -369 -988 -303 -972
rect -177 -938 -111 -922
rect -63 -926 -33 -900
rect 33 -922 63 -900
rect -177 -972 -161 -938
rect -127 -972 -111 -938
rect -177 -988 -111 -972
rect 15 -938 81 -922
rect 129 -926 159 -900
rect 225 -922 255 -900
rect 15 -972 31 -938
rect 65 -972 81 -938
rect 15 -988 81 -972
rect 207 -938 273 -922
rect 321 -926 351 -900
rect 417 -922 447 -900
rect 207 -972 223 -938
rect 257 -972 273 -938
rect 207 -988 273 -972
rect 399 -938 465 -922
rect 513 -926 543 -900
rect 609 -922 639 -900
rect 399 -972 415 -938
rect 449 -972 465 -938
rect 399 -988 465 -972
rect 591 -938 657 -922
rect 705 -926 735 -900
rect 801 -922 831 -900
rect 591 -972 607 -938
rect 641 -972 657 -938
rect 591 -988 657 -972
rect 783 -938 849 -922
rect 897 -926 927 -900
rect 783 -972 799 -938
rect 833 -972 849 -938
rect 783 -988 849 -972
<< polycont >>
rect -833 938 -799 972
rect -641 938 -607 972
rect -449 938 -415 972
rect -257 938 -223 972
rect -65 938 -31 972
rect 127 938 161 972
rect 319 938 353 972
rect 511 938 545 972
rect 703 938 737 972
rect 895 938 929 972
rect -929 -972 -895 -938
rect -737 -972 -703 -938
rect -545 -972 -511 -938
rect -353 -972 -319 -938
rect -161 -972 -127 -938
rect 31 -972 65 -938
rect 223 -972 257 -938
rect 415 -972 449 -938
rect 607 -972 641 -938
rect 799 -972 833 -938
<< locali >>
rect -1091 1040 -995 1074
rect 995 1040 1091 1074
rect -1091 978 -1057 1040
rect -849 938 -833 972
rect -799 938 -783 972
rect -657 938 -641 972
rect -607 938 -591 972
rect -465 938 -449 972
rect -415 938 -399 972
rect -273 938 -257 972
rect -223 938 -207 972
rect -81 938 -65 972
rect -31 938 -15 972
rect 111 938 127 972
rect 161 938 177 972
rect 303 938 319 972
rect 353 938 369 972
rect 495 938 511 972
rect 545 938 561 972
rect 687 938 703 972
rect 737 938 753 972
rect 879 938 895 972
rect 929 938 945 972
rect -977 888 -943 904
rect -977 -904 -943 -888
rect -881 888 -847 904
rect -881 -904 -847 -888
rect -785 888 -751 904
rect -785 -904 -751 -888
rect -689 888 -655 904
rect -689 -904 -655 -888
rect -593 888 -559 904
rect -593 -904 -559 -888
rect -497 888 -463 904
rect -497 -904 -463 -888
rect -401 888 -367 904
rect -401 -904 -367 -888
rect -305 888 -271 904
rect -305 -904 -271 -888
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect 271 888 305 904
rect 271 -904 305 -888
rect 367 888 401 904
rect 367 -904 401 -888
rect 463 888 497 904
rect 463 -904 497 -888
rect 559 888 593 904
rect 559 -904 593 -888
rect 655 888 689 904
rect 655 -904 689 -888
rect 751 888 785 904
rect 751 -904 785 -888
rect 847 888 881 904
rect 847 -904 881 -888
rect 943 888 977 904
rect 943 -904 977 -888
rect -945 -972 -929 -938
rect -895 -972 -879 -938
rect -753 -972 -737 -938
rect -703 -972 -687 -938
rect -561 -972 -545 -938
rect -511 -972 -495 -938
rect -369 -972 -353 -938
rect -319 -972 -303 -938
rect -177 -972 -161 -938
rect -127 -972 -111 -938
rect 15 -972 31 -938
rect 65 -972 81 -938
rect 207 -972 223 -938
rect 257 -972 273 -938
rect 399 -972 415 -938
rect 449 -972 465 -938
rect 591 -972 607 -938
rect 641 -972 657 -938
rect 783 -972 799 -938
rect 833 -972 849 -938
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1040
rect -1091 -1074 1091 -1040
<< viali >>
rect -833 938 -799 972
rect -641 938 -607 972
rect -449 938 -415 972
rect -257 938 -223 972
rect -65 938 -31 972
rect 127 938 161 972
rect 319 938 353 972
rect 511 938 545 972
rect 703 938 737 972
rect 895 938 929 972
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
rect -929 -972 -895 -938
rect -737 -972 -703 -938
rect -545 -972 -511 -938
rect -353 -972 -319 -938
rect -161 -972 -127 -938
rect 31 -972 65 -938
rect 223 -972 257 -938
rect 415 -972 449 -938
rect 607 -972 641 -938
rect 799 -972 833 -938
<< metal1 >>
rect -845 972 -787 978
rect -845 938 -833 972
rect -799 938 -787 972
rect -845 932 -787 938
rect -653 972 -595 978
rect -653 938 -641 972
rect -607 938 -595 972
rect -653 932 -595 938
rect -461 972 -403 978
rect -461 938 -449 972
rect -415 938 -403 972
rect -461 932 -403 938
rect -269 972 -211 978
rect -269 938 -257 972
rect -223 938 -211 972
rect -269 932 -211 938
rect -77 972 -19 978
rect -77 938 -65 972
rect -31 938 -19 972
rect -77 932 -19 938
rect 115 972 173 978
rect 115 938 127 972
rect 161 938 173 972
rect 115 932 173 938
rect 307 972 365 978
rect 307 938 319 972
rect 353 938 365 972
rect 307 932 365 938
rect 499 972 557 978
rect 499 938 511 972
rect 545 938 557 972
rect 499 932 557 938
rect 691 972 749 978
rect 691 938 703 972
rect 737 938 749 972
rect 691 932 749 938
rect 883 972 941 978
rect 883 938 895 972
rect 929 938 941 972
rect 883 932 941 938
rect -983 888 -937 900
rect -983 -888 -977 888
rect -943 -888 -937 888
rect -983 -900 -937 -888
rect -887 888 -841 900
rect -887 -888 -881 888
rect -847 -888 -841 888
rect -887 -900 -841 -888
rect -791 888 -745 900
rect -791 -888 -785 888
rect -751 -888 -745 888
rect -791 -900 -745 -888
rect -695 888 -649 900
rect -695 -888 -689 888
rect -655 -888 -649 888
rect -695 -900 -649 -888
rect -599 888 -553 900
rect -599 -888 -593 888
rect -559 -888 -553 888
rect -599 -900 -553 -888
rect -503 888 -457 900
rect -503 -888 -497 888
rect -463 -888 -457 888
rect -503 -900 -457 -888
rect -407 888 -361 900
rect -407 -888 -401 888
rect -367 -888 -361 888
rect -407 -900 -361 -888
rect -311 888 -265 900
rect -311 -888 -305 888
rect -271 -888 -265 888
rect -311 -900 -265 -888
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect 265 888 311 900
rect 265 -888 271 888
rect 305 -888 311 888
rect 265 -900 311 -888
rect 361 888 407 900
rect 361 -888 367 888
rect 401 -888 407 888
rect 361 -900 407 -888
rect 457 888 503 900
rect 457 -888 463 888
rect 497 -888 503 888
rect 457 -900 503 -888
rect 553 888 599 900
rect 553 -888 559 888
rect 593 -888 599 888
rect 553 -900 599 -888
rect 649 888 695 900
rect 649 -888 655 888
rect 689 -888 695 888
rect 649 -900 695 -888
rect 745 888 791 900
rect 745 -888 751 888
rect 785 -888 791 888
rect 745 -900 791 -888
rect 841 888 887 900
rect 841 -888 847 888
rect 881 -888 887 888
rect 841 -900 887 -888
rect 937 888 983 900
rect 937 -888 943 888
rect 977 -888 983 888
rect 937 -900 983 -888
rect -941 -938 -883 -932
rect -941 -972 -929 -938
rect -895 -972 -883 -938
rect -941 -978 -883 -972
rect -749 -938 -691 -932
rect -749 -972 -737 -938
rect -703 -972 -691 -938
rect -749 -978 -691 -972
rect -557 -938 -499 -932
rect -557 -972 -545 -938
rect -511 -972 -499 -938
rect -557 -978 -499 -972
rect -365 -938 -307 -932
rect -365 -972 -353 -938
rect -319 -972 -307 -938
rect -365 -978 -307 -972
rect -173 -938 -115 -932
rect -173 -972 -161 -938
rect -127 -972 -115 -938
rect -173 -978 -115 -972
rect 19 -938 77 -932
rect 19 -972 31 -938
rect 65 -972 77 -938
rect 19 -978 77 -972
rect 211 -938 269 -932
rect 211 -972 223 -938
rect 257 -972 269 -938
rect 211 -978 269 -972
rect 403 -938 461 -932
rect 403 -972 415 -938
rect 449 -972 461 -938
rect 403 -978 461 -972
rect 595 -938 653 -932
rect 595 -972 607 -938
rect 641 -972 653 -938
rect 595 -978 653 -972
rect 787 -938 845 -932
rect 787 -972 799 -938
rect 833 -972 845 -938
rect 787 -978 845 -972
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -1057 1074 1057
string parameters w 9 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
