magic
tech sky130A
magscale 1 2
timestamp 1615222810
<< error_p >>
rect -77 171 -19 177
rect 115 171 173 177
rect -77 137 -65 171
rect 115 137 127 171
rect -77 131 -19 137
rect 115 131 173 137
rect -173 -137 -115 -131
rect 19 -137 77 -131
rect -173 -171 -161 -137
rect 19 -171 31 -137
rect -173 -177 -115 -171
rect 19 -177 77 -171
<< nwell >>
rect -161 152 257 190
rect -257 -152 257 152
rect -257 -190 161 -152
<< pmos >>
rect -159 -90 -129 90
rect -63 -90 -33 90
rect 33 -90 63 90
rect 129 -90 159 90
<< pdiff >>
rect -221 78 -159 90
rect -221 -78 -209 78
rect -175 -78 -159 78
rect -221 -90 -159 -78
rect -129 78 -63 90
rect -129 -78 -113 78
rect -79 -78 -63 78
rect -129 -90 -63 -78
rect -33 78 33 90
rect -33 -78 -17 78
rect 17 -78 33 78
rect -33 -90 33 -78
rect 63 78 129 90
rect 63 -78 79 78
rect 113 -78 129 78
rect 63 -90 129 -78
rect 159 78 221 90
rect 159 -78 175 78
rect 209 -78 221 78
rect 159 -90 221 -78
<< pdiffc >>
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
<< poly >>
rect -81 171 -15 187
rect -81 137 -65 171
rect -31 137 -15 171
rect -81 121 -15 137
rect 111 171 177 187
rect 111 137 127 171
rect 161 137 177 171
rect 111 121 177 137
rect -159 90 -129 116
rect -63 90 -33 121
rect 33 90 63 116
rect 129 90 159 121
rect -159 -121 -129 -90
rect -63 -116 -33 -90
rect 33 -121 63 -90
rect 129 -116 159 -90
rect -177 -137 -111 -121
rect -177 -171 -161 -137
rect -127 -171 -111 -137
rect -177 -187 -111 -171
rect 15 -137 81 -121
rect 15 -171 31 -137
rect 65 -171 81 -137
rect 15 -187 81 -171
<< polycont >>
rect -65 137 -31 171
rect 127 137 161 171
rect -161 -171 -127 -137
rect 31 -171 65 -137
<< locali >>
rect -81 137 -65 171
rect -31 137 -15 171
rect 111 137 127 171
rect 161 137 177 171
rect -209 78 -175 94
rect -209 -94 -175 -78
rect -113 78 -79 94
rect -113 -94 -79 -78
rect -17 78 17 94
rect -17 -94 17 -78
rect 79 78 113 94
rect 79 -94 113 -78
rect 175 78 209 94
rect 175 -94 209 -78
rect -177 -171 -161 -137
rect -127 -171 -111 -137
rect 15 -171 31 -137
rect 65 -171 81 -137
<< viali >>
rect -65 137 -31 171
rect 127 137 161 171
rect -209 -78 -175 78
rect -113 -78 -79 78
rect -17 -78 17 78
rect 79 -78 113 78
rect 175 -78 209 78
rect -161 -171 -127 -137
rect 31 -171 65 -137
<< metal1 >>
rect -77 171 -19 177
rect -77 137 -65 171
rect -31 137 -19 171
rect -77 131 -19 137
rect 115 171 173 177
rect 115 137 127 171
rect 161 137 173 171
rect 115 131 173 137
rect -215 78 -169 90
rect -215 -78 -209 78
rect -175 -78 -169 78
rect -215 -90 -169 -78
rect -119 78 -73 90
rect -119 -78 -113 78
rect -79 -78 -73 78
rect -119 -90 -73 -78
rect -23 78 23 90
rect -23 -78 -17 78
rect 17 -78 23 78
rect -23 -90 23 -78
rect 73 78 119 90
rect 73 -78 79 78
rect 113 -78 119 78
rect 73 -90 119 -78
rect 169 78 215 90
rect 169 -78 175 78
rect 209 -78 215 78
rect 169 -90 215 -78
rect -173 -137 -115 -131
rect -173 -171 -161 -137
rect -127 -171 -115 -137
rect -173 -177 -115 -171
rect 19 -137 77 -131
rect 19 -171 31 -137
rect 65 -171 77 -137
rect 19 -177 77 -171
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.9 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
