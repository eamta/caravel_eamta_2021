magic
tech sky130A
magscale 1 2
timestamp 1616024728
<< nwell >>
rect -104 -76 10001 2080
<< pmos >>
rect 3447 167 3587 1567
rect 3645 167 3785 1567
rect 3843 167 3983 1567
rect 4041 167 4181 1567
rect 4239 167 4379 1567
rect 4437 167 4577 1567
rect 4635 167 4775 1567
rect 4833 167 4973 1567
rect 5031 167 5171 1567
rect 5229 167 5369 1567
rect 5427 167 5567 1567
rect 5625 167 5765 1567
rect 5823 167 5963 1567
rect 6021 167 6161 1567
rect 6219 167 6359 1567
rect 6751 167 6891 1567
rect 6949 167 7089 1567
rect 7147 167 7287 1567
rect 7345 167 7485 1567
rect 7543 167 7683 1567
rect 7741 167 7881 1567
rect 7939 167 8079 1567
rect 8137 167 8277 1567
rect 8335 167 8475 1567
rect 8533 167 8673 1567
rect 8731 167 8871 1567
rect 8929 167 9069 1567
rect 9127 167 9267 1567
rect 9325 167 9465 1567
rect 9523 167 9663 1567
<< pdiff >>
rect 3389 1555 3447 1567
rect 3389 179 3401 1555
rect 3435 179 3447 1555
rect 3389 167 3447 179
rect 3587 1555 3645 1567
rect 3587 179 3599 1555
rect 3633 179 3645 1555
rect 3587 167 3645 179
rect 3785 1555 3843 1567
rect 3785 179 3797 1555
rect 3831 179 3843 1555
rect 3785 167 3843 179
rect 3983 1555 4041 1567
rect 3983 179 3995 1555
rect 4029 179 4041 1555
rect 3983 167 4041 179
rect 4181 1555 4239 1567
rect 4181 179 4193 1555
rect 4227 179 4239 1555
rect 4181 167 4239 179
rect 4379 1555 4437 1567
rect 4379 179 4391 1555
rect 4425 179 4437 1555
rect 4379 167 4437 179
rect 4577 1555 4635 1567
rect 4577 179 4589 1555
rect 4623 179 4635 1555
rect 4577 167 4635 179
rect 4775 1555 4833 1567
rect 4775 179 4787 1555
rect 4821 179 4833 1555
rect 4775 167 4833 179
rect 4973 1555 5031 1567
rect 4973 179 4985 1555
rect 5019 179 5031 1555
rect 4973 167 5031 179
rect 5171 1555 5229 1567
rect 5171 179 5183 1555
rect 5217 179 5229 1555
rect 5171 167 5229 179
rect 5369 1555 5427 1567
rect 5369 179 5381 1555
rect 5415 179 5427 1555
rect 5369 167 5427 179
rect 5567 1555 5625 1567
rect 5567 179 5579 1555
rect 5613 179 5625 1555
rect 5567 167 5625 179
rect 5765 1555 5823 1567
rect 5765 179 5777 1555
rect 5811 179 5823 1555
rect 5765 167 5823 179
rect 5963 1555 6021 1567
rect 5963 179 5975 1555
rect 6009 179 6021 1555
rect 5963 167 6021 179
rect 6161 1555 6219 1567
rect 6161 179 6173 1555
rect 6207 179 6219 1555
rect 6161 167 6219 179
rect 6359 1555 6417 1567
rect 6359 179 6371 1555
rect 6405 179 6417 1555
rect 6359 167 6417 179
rect 6693 1555 6751 1567
rect 6693 179 6705 1555
rect 6739 179 6751 1555
rect 6693 167 6751 179
rect 6891 1555 6949 1567
rect 6891 179 6903 1555
rect 6937 179 6949 1555
rect 6891 167 6949 179
rect 7089 1555 7147 1567
rect 7089 179 7101 1555
rect 7135 179 7147 1555
rect 7089 167 7147 179
rect 7287 1555 7345 1567
rect 7287 179 7299 1555
rect 7333 179 7345 1555
rect 7287 167 7345 179
rect 7485 1555 7543 1567
rect 7485 179 7497 1555
rect 7531 179 7543 1555
rect 7485 167 7543 179
rect 7683 1555 7741 1567
rect 7683 179 7695 1555
rect 7729 179 7741 1555
rect 7683 167 7741 179
rect 7881 1555 7939 1567
rect 7881 179 7893 1555
rect 7927 179 7939 1555
rect 7881 167 7939 179
rect 8079 1555 8137 1567
rect 8079 179 8091 1555
rect 8125 179 8137 1555
rect 8079 167 8137 179
rect 8277 1555 8335 1567
rect 8277 179 8289 1555
rect 8323 179 8335 1555
rect 8277 167 8335 179
rect 8475 1555 8533 1567
rect 8475 179 8487 1555
rect 8521 179 8533 1555
rect 8475 167 8533 179
rect 8673 1555 8731 1567
rect 8673 179 8685 1555
rect 8719 179 8731 1555
rect 8673 167 8731 179
rect 8871 1555 8929 1567
rect 8871 179 8883 1555
rect 8917 179 8929 1555
rect 8871 167 8929 179
rect 9069 1555 9127 1567
rect 9069 179 9081 1555
rect 9115 179 9127 1555
rect 9069 167 9127 179
rect 9267 1555 9325 1567
rect 9267 179 9279 1555
rect 9313 179 9325 1555
rect 9267 167 9325 179
rect 9465 1555 9523 1567
rect 9465 179 9477 1555
rect 9511 179 9523 1555
rect 9465 167 9523 179
rect 9663 1555 9721 1567
rect 9663 179 9675 1555
rect 9709 179 9721 1555
rect 9663 167 9721 179
<< pdiffc >>
rect 3401 179 3435 1555
rect 3599 179 3633 1555
rect 3797 179 3831 1555
rect 3995 179 4029 1555
rect 4193 179 4227 1555
rect 4391 179 4425 1555
rect 4589 179 4623 1555
rect 4787 179 4821 1555
rect 4985 179 5019 1555
rect 5183 179 5217 1555
rect 5381 179 5415 1555
rect 5579 179 5613 1555
rect 5777 179 5811 1555
rect 5975 179 6009 1555
rect 6173 179 6207 1555
rect 6371 179 6405 1555
rect 6705 179 6739 1555
rect 6903 179 6937 1555
rect 7101 179 7135 1555
rect 7299 179 7333 1555
rect 7497 179 7531 1555
rect 7695 179 7729 1555
rect 7893 179 7927 1555
rect 8091 179 8125 1555
rect 8289 179 8323 1555
rect 8487 179 8521 1555
rect 8685 179 8719 1555
rect 8883 179 8917 1555
rect 9081 179 9115 1555
rect 9279 179 9313 1555
rect 9477 179 9511 1555
rect 9675 179 9709 1555
<< nsubdiff >>
rect 3287 1645 3383 1679
rect 6423 1645 6519 1679
rect 3287 1582 3321 1645
rect 6485 1582 6519 1645
rect 3287 17 3321 80
rect 6485 17 6519 80
rect 3287 -17 3383 17
rect 6423 -17 6519 17
rect 6591 1645 6687 1679
rect 9727 1645 9823 1679
rect 6591 1582 6625 1645
rect 9789 1582 9823 1645
rect 6591 17 6625 80
rect 9789 17 9823 80
rect 6591 -17 6687 17
rect 9727 -17 9823 17
<< nsubdiffcont >>
rect 3383 1645 6423 1679
rect 3287 80 3321 1582
rect 6485 80 6519 1582
rect 3383 -17 6423 17
rect 6687 1645 9727 1679
rect 6591 80 6625 1582
rect 9789 80 9823 1582
rect 6687 -17 9727 17
<< poly >>
rect 3447 1567 3587 1593
rect 3645 1567 3785 1593
rect 3843 1567 3983 1593
rect 4041 1567 4181 1593
rect 4239 1567 4379 1593
rect 4437 1567 4577 1593
rect 4635 1567 4775 1593
rect 4833 1567 4973 1593
rect 5031 1567 5171 1593
rect 5229 1567 5369 1593
rect 5427 1567 5567 1593
rect 5625 1567 5765 1593
rect 5823 1567 5963 1593
rect 6021 1567 6161 1593
rect 6219 1567 6359 1593
rect 3447 120 3587 167
rect 3447 86 3463 120
rect 3571 86 3587 120
rect 3447 70 3587 86
rect 3645 120 3785 167
rect 3645 86 3661 120
rect 3769 86 3785 120
rect 3645 70 3785 86
rect 3843 120 3983 167
rect 3843 86 3859 120
rect 3967 86 3983 120
rect 3843 70 3983 86
rect 4041 120 4181 167
rect 4041 86 4057 120
rect 4165 86 4181 120
rect 4041 70 4181 86
rect 4239 120 4379 167
rect 4239 86 4255 120
rect 4363 86 4379 120
rect 4239 70 4379 86
rect 4437 120 4577 167
rect 4437 86 4453 120
rect 4561 86 4577 120
rect 4437 70 4577 86
rect 4635 120 4775 167
rect 4635 86 4651 120
rect 4759 86 4775 120
rect 4635 70 4775 86
rect 4833 120 4973 167
rect 4833 86 4849 120
rect 4957 86 4973 120
rect 4833 70 4973 86
rect 5031 120 5171 167
rect 5031 86 5047 120
rect 5155 86 5171 120
rect 5031 70 5171 86
rect 5229 120 5369 167
rect 5229 86 5245 120
rect 5353 86 5369 120
rect 5229 70 5369 86
rect 5427 120 5567 167
rect 5427 86 5443 120
rect 5551 86 5567 120
rect 5427 70 5567 86
rect 5625 120 5765 167
rect 5625 86 5641 120
rect 5749 86 5765 120
rect 5625 70 5765 86
rect 5823 120 5963 167
rect 5823 86 5839 120
rect 5947 86 5963 120
rect 5823 70 5963 86
rect 6021 120 6161 167
rect 6021 86 6037 120
rect 6145 86 6161 120
rect 6021 70 6161 86
rect 6219 120 6359 167
rect 6219 86 6235 120
rect 6343 86 6359 120
rect 6219 70 6359 86
rect 6751 1567 6891 1593
rect 6949 1567 7089 1593
rect 7147 1567 7287 1593
rect 7345 1567 7485 1593
rect 7543 1567 7683 1593
rect 7741 1567 7881 1593
rect 7939 1567 8079 1593
rect 8137 1567 8277 1593
rect 8335 1567 8475 1593
rect 8533 1567 8673 1593
rect 8731 1567 8871 1593
rect 8929 1567 9069 1593
rect 9127 1567 9267 1593
rect 9325 1567 9465 1593
rect 9523 1567 9663 1593
rect 6751 120 6891 167
rect 6751 86 6767 120
rect 6875 86 6891 120
rect 6751 70 6891 86
rect 6949 120 7089 167
rect 6949 86 6965 120
rect 7073 86 7089 120
rect 6949 70 7089 86
rect 7147 120 7287 167
rect 7147 86 7163 120
rect 7271 86 7287 120
rect 7147 70 7287 86
rect 7345 120 7485 167
rect 7345 86 7361 120
rect 7469 86 7485 120
rect 7345 70 7485 86
rect 7543 120 7683 167
rect 7543 86 7559 120
rect 7667 86 7683 120
rect 7543 70 7683 86
rect 7741 120 7881 167
rect 7741 86 7757 120
rect 7865 86 7881 120
rect 7741 70 7881 86
rect 7939 120 8079 167
rect 7939 86 7955 120
rect 8063 86 8079 120
rect 7939 70 8079 86
rect 8137 120 8277 167
rect 8137 86 8153 120
rect 8261 86 8277 120
rect 8137 70 8277 86
rect 8335 120 8475 167
rect 8335 86 8351 120
rect 8459 86 8475 120
rect 8335 70 8475 86
rect 8533 120 8673 167
rect 8533 86 8549 120
rect 8657 86 8673 120
rect 8533 70 8673 86
rect 8731 120 8871 167
rect 8731 86 8747 120
rect 8855 86 8871 120
rect 8731 70 8871 86
rect 8929 120 9069 167
rect 8929 86 8945 120
rect 9053 86 9069 120
rect 8929 70 9069 86
rect 9127 120 9267 167
rect 9127 86 9143 120
rect 9251 86 9267 120
rect 9127 70 9267 86
rect 9325 120 9465 167
rect 9325 86 9341 120
rect 9449 86 9465 120
rect 9325 70 9465 86
rect 9523 120 9663 167
rect 9523 86 9539 120
rect 9647 86 9663 120
rect 9523 70 9663 86
<< polycont >>
rect 3463 86 3571 120
rect 3661 86 3769 120
rect 3859 86 3967 120
rect 4057 86 4165 120
rect 4255 86 4363 120
rect 4453 86 4561 120
rect 4651 86 4759 120
rect 4849 86 4957 120
rect 5047 86 5155 120
rect 5245 86 5353 120
rect 5443 86 5551 120
rect 5641 86 5749 120
rect 5839 86 5947 120
rect 6037 86 6145 120
rect 6235 86 6343 120
rect 6767 86 6875 120
rect 6965 86 7073 120
rect 7163 86 7271 120
rect 7361 86 7469 120
rect 7559 86 7667 120
rect 7757 86 7865 120
rect 7955 86 8063 120
rect 8153 86 8261 120
rect 8351 86 8459 120
rect 8549 86 8657 120
rect 8747 86 8855 120
rect 8945 86 9053 120
rect 9143 86 9251 120
rect 9341 86 9449 120
rect 9539 86 9647 120
<< locali >>
rect 3287 1645 3383 1679
rect 6423 1645 6519 1679
rect 3287 1582 3321 1645
rect 6485 1582 6519 1645
rect 3401 1555 3435 1571
rect 3401 163 3435 179
rect 3599 1555 3633 1571
rect 3599 163 3633 179
rect 3797 1555 3831 1571
rect 3797 163 3831 179
rect 3995 1555 4029 1571
rect 3995 163 4029 179
rect 4193 1555 4227 1571
rect 4193 163 4227 179
rect 4391 1555 4425 1571
rect 4391 163 4425 179
rect 4589 1555 4623 1571
rect 4589 163 4623 179
rect 4787 1555 4821 1571
rect 4787 163 4821 179
rect 4985 1555 5019 1571
rect 4985 163 5019 179
rect 5183 1555 5217 1571
rect 5183 163 5217 179
rect 5381 1555 5415 1571
rect 5381 163 5415 179
rect 5579 1555 5613 1571
rect 5579 163 5613 179
rect 5777 1555 5811 1571
rect 5777 163 5811 179
rect 5975 1555 6009 1571
rect 5975 163 6009 179
rect 6173 1555 6207 1571
rect 6173 163 6207 179
rect 6371 1555 6405 1571
rect 6371 163 6405 179
rect 3447 86 3463 120
rect 3571 86 3587 120
rect 3645 86 3661 120
rect 3769 86 3785 120
rect 3843 86 3859 120
rect 3967 86 3983 120
rect 4041 86 4057 120
rect 4165 86 4181 120
rect 4239 86 4255 120
rect 4363 86 4379 120
rect 4437 86 4453 120
rect 4561 86 4577 120
rect 4635 86 4651 120
rect 4759 86 4775 120
rect 4833 86 4849 120
rect 4957 86 4973 120
rect 5031 86 5047 120
rect 5155 86 5171 120
rect 5229 86 5245 120
rect 5353 86 5369 120
rect 5427 86 5443 120
rect 5551 86 5567 120
rect 5625 86 5641 120
rect 5749 86 5765 120
rect 5823 86 5839 120
rect 5947 86 5963 120
rect 6021 86 6037 120
rect 6145 86 6161 120
rect 6219 86 6235 120
rect 6343 86 6359 120
rect 3287 17 3321 80
rect 6485 17 6519 80
rect 3287 -17 3383 17
rect 6423 -17 6519 17
rect 6591 1645 6687 1679
rect 9727 1645 9823 1679
rect 6591 1582 6625 1645
rect 9789 1582 9823 1645
rect 6705 1555 6739 1571
rect 6705 163 6739 179
rect 6903 1555 6937 1571
rect 6903 163 6937 179
rect 7101 1555 7135 1571
rect 7101 163 7135 179
rect 7299 1555 7333 1571
rect 7299 163 7333 179
rect 7497 1555 7531 1571
rect 7497 163 7531 179
rect 7695 1555 7729 1571
rect 7695 163 7729 179
rect 7893 1555 7927 1571
rect 7893 163 7927 179
rect 8091 1555 8125 1571
rect 8091 163 8125 179
rect 8289 1555 8323 1571
rect 8289 163 8323 179
rect 8487 1555 8521 1571
rect 8487 163 8521 179
rect 8685 1555 8719 1571
rect 8685 163 8719 179
rect 8883 1555 8917 1571
rect 8883 163 8917 179
rect 9081 1555 9115 1571
rect 9081 163 9115 179
rect 9279 1555 9313 1571
rect 9279 163 9313 179
rect 9477 1555 9511 1571
rect 9477 163 9511 179
rect 9675 1555 9709 1571
rect 9675 163 9709 179
rect 6751 86 6767 120
rect 6875 86 6891 120
rect 6949 86 6965 120
rect 7073 86 7089 120
rect 7147 86 7163 120
rect 7271 86 7287 120
rect 7345 86 7361 120
rect 7469 86 7485 120
rect 7543 86 7559 120
rect 7667 86 7683 120
rect 7741 86 7757 120
rect 7865 86 7881 120
rect 7939 86 7955 120
rect 8063 86 8079 120
rect 8137 86 8153 120
rect 8261 86 8277 120
rect 8335 86 8351 120
rect 8459 86 8475 120
rect 8533 86 8549 120
rect 8657 86 8673 120
rect 8731 86 8747 120
rect 8855 86 8871 120
rect 8929 86 8945 120
rect 9053 86 9069 120
rect 9127 86 9143 120
rect 9251 86 9267 120
rect 9325 86 9341 120
rect 9449 86 9465 120
rect 9523 86 9539 120
rect 9647 86 9663 120
rect 6591 17 6625 80
rect 9789 17 9823 80
rect 6591 -17 6687 17
rect 9727 -17 9823 17
<< viali >>
rect 3401 179 3435 1555
rect 3599 179 3633 1555
rect 3797 179 3831 1555
rect 3995 179 4029 1555
rect 4193 179 4227 1555
rect 4391 179 4425 1555
rect 4589 179 4623 1555
rect 4787 179 4821 1555
rect 4985 179 5019 1555
rect 5183 179 5217 1555
rect 5381 179 5415 1555
rect 5579 179 5613 1555
rect 5777 179 5811 1555
rect 5975 179 6009 1555
rect 6173 179 6207 1555
rect 6371 179 6405 1555
rect 3463 86 3571 120
rect 3661 86 3769 120
rect 3859 86 3967 120
rect 4057 86 4165 120
rect 4255 86 4363 120
rect 4453 86 4561 120
rect 4651 86 4759 120
rect 4849 86 4957 120
rect 5047 86 5155 120
rect 5245 86 5353 120
rect 5443 86 5551 120
rect 5641 86 5749 120
rect 5839 86 5947 120
rect 6037 86 6145 120
rect 6235 86 6343 120
rect 6705 179 6739 1555
rect 6903 179 6937 1555
rect 7101 179 7135 1555
rect 7299 179 7333 1555
rect 7497 179 7531 1555
rect 7695 179 7729 1555
rect 7893 179 7927 1555
rect 8091 179 8125 1555
rect 8289 179 8323 1555
rect 8487 179 8521 1555
rect 8685 179 8719 1555
rect 8883 179 8917 1555
rect 9081 179 9115 1555
rect 9279 179 9313 1555
rect 9477 179 9511 1555
rect 9675 179 9709 1555
rect 6767 86 6875 120
rect 6965 86 7073 120
rect 7163 86 7271 120
rect 7361 86 7469 120
rect 7559 86 7667 120
rect 7757 86 7865 120
rect 7955 86 8063 120
rect 8153 86 8261 120
rect 8351 86 8459 120
rect 8549 86 8657 120
rect 8747 86 8855 120
rect 8945 86 9053 120
rect 9143 86 9251 120
rect 9341 86 9449 120
rect 9539 86 9647 120
<< metal1 >>
rect 91 167 137 1743
rect 276 179 286 1555
rect 338 179 348 1555
rect 487 167 533 1743
rect 672 179 682 1555
rect 734 179 744 1555
rect 883 167 929 1743
rect 1068 179 1078 1555
rect 1130 179 1140 1555
rect 1279 167 1325 1743
rect 1464 179 1474 1555
rect 1526 179 1536 1555
rect 1675 167 1721 1743
rect 1860 179 1870 1555
rect 1922 179 1932 1555
rect 2071 167 2117 1743
rect 2256 179 2266 1555
rect 2318 179 2328 1555
rect 2467 167 2513 1743
rect 2652 179 2662 1555
rect 2714 179 2724 1555
rect 2863 167 2909 1743
rect 3395 1555 3441 1743
rect 3593 1555 3639 1567
rect 3791 1555 3837 1743
rect 3989 1555 4035 1567
rect 4187 1555 4233 1743
rect 4385 1555 4431 1567
rect 4583 1555 4629 1743
rect 4781 1555 4827 1567
rect 4979 1555 5025 1743
rect 5177 1555 5223 1567
rect 5375 1555 5421 1743
rect 5573 1555 5619 1567
rect 5771 1555 5817 1743
rect 5969 1555 6015 1567
rect 6167 1555 6213 1743
rect 6365 1555 6411 1567
rect 6699 1555 6745 1743
rect 6897 1555 6943 1567
rect 7095 1555 7141 1743
rect 7293 1555 7339 1567
rect 7491 1555 7537 1743
rect 7689 1555 7735 1567
rect 7887 1555 7933 1743
rect 8085 1555 8131 1567
rect 8283 1555 8329 1743
rect 8481 1555 8527 1567
rect 8679 1555 8725 1743
rect 8877 1555 8923 1567
rect 9075 1555 9121 1743
rect 9273 1555 9319 1567
rect 9471 1555 9517 1743
rect 9669 1555 9715 1567
rect 3048 179 3058 1555
rect 3110 179 3120 1555
rect 3395 179 3401 1555
rect 3435 179 3441 1555
rect 3580 179 3590 1555
rect 3642 179 3652 1555
rect 3791 179 3797 1555
rect 3831 179 3837 1555
rect 3976 179 3986 1555
rect 4038 179 4048 1555
rect 4187 179 4193 1555
rect 4227 179 4233 1555
rect 4372 179 4382 1555
rect 4434 179 4444 1555
rect 4583 179 4589 1555
rect 4623 179 4629 1555
rect 4768 179 4778 1555
rect 4830 179 4840 1555
rect 4979 179 4985 1555
rect 5019 179 5025 1555
rect 5164 179 5174 1555
rect 5226 179 5236 1555
rect 5375 179 5381 1555
rect 5415 179 5421 1555
rect 5560 179 5570 1555
rect 5622 179 5632 1555
rect 5771 179 5777 1555
rect 5811 179 5817 1555
rect 5956 179 5966 1555
rect 6018 179 6028 1555
rect 6167 179 6173 1555
rect 6207 179 6213 1555
rect 6352 179 6362 1555
rect 6414 179 6424 1555
rect 6699 179 6705 1555
rect 6739 179 6745 1555
rect 6884 179 6894 1555
rect 6946 179 6956 1555
rect 7095 179 7101 1555
rect 7135 179 7141 1555
rect 7280 179 7290 1555
rect 7342 179 7352 1555
rect 7491 179 7497 1555
rect 7531 179 7537 1555
rect 7676 179 7686 1555
rect 7738 179 7748 1555
rect 7887 179 7893 1555
rect 7927 179 7933 1555
rect 8072 179 8082 1555
rect 8134 179 8144 1555
rect 8283 179 8289 1555
rect 8323 179 8329 1555
rect 8468 179 8478 1555
rect 8530 179 8540 1555
rect 8679 179 8685 1555
rect 8719 179 8725 1555
rect 8864 179 8874 1555
rect 8926 179 8936 1555
rect 9075 179 9081 1555
rect 9115 179 9121 1555
rect 9260 179 9270 1555
rect 9322 179 9332 1555
rect 9471 179 9477 1555
rect 9511 179 9517 1555
rect 9656 179 9666 1555
rect 9718 179 9728 1555
rect 3395 167 3441 179
rect 3593 167 3639 179
rect 3791 167 3837 179
rect 3989 167 4035 179
rect 4187 167 4233 179
rect 4385 167 4431 179
rect 4583 167 4629 179
rect 4781 167 4827 179
rect 4979 167 5025 179
rect 5177 167 5223 179
rect 5375 167 5421 179
rect 5573 167 5619 179
rect 5771 167 5817 179
rect 5969 167 6015 179
rect 6167 167 6213 179
rect 6365 167 6411 179
rect 6699 167 6745 179
rect 6897 167 6943 179
rect 7095 167 7141 179
rect 7293 167 7339 179
rect 7491 167 7537 179
rect 7689 167 7735 179
rect 7887 167 7933 179
rect 8085 167 8131 179
rect 8283 167 8329 179
rect 8481 167 8527 179
rect 8679 167 8725 179
rect 8877 167 8923 179
rect 9075 167 9121 179
rect 9273 167 9319 179
rect 9471 167 9517 179
rect 9669 167 9715 179
rect 147 80 3051 126
rect 3451 120 6355 126
rect 3451 86 3463 120
rect 3571 86 3661 120
rect 3769 86 3859 120
rect 3967 86 4057 120
rect 4165 86 4255 120
rect 4363 86 4453 120
rect 4561 86 4651 120
rect 4759 86 4849 120
rect 4957 86 5047 120
rect 5155 86 5245 120
rect 5353 86 5443 120
rect 5551 86 5641 120
rect 5749 86 5839 120
rect 5947 86 6037 120
rect 6145 86 6235 120
rect 6343 86 6355 120
rect 3451 80 6355 86
rect 6755 120 9659 126
rect 6755 86 6767 120
rect 6875 86 6965 120
rect 7073 86 7163 120
rect 7271 86 7361 120
rect 7469 86 7559 120
rect 7667 86 7757 120
rect 7865 86 7955 120
rect 8063 86 8153 120
rect 8261 86 8351 120
rect 8459 86 8549 120
rect 8657 86 8747 120
rect 8855 86 8945 120
rect 9053 86 9143 120
rect 9251 86 9341 120
rect 9449 86 9539 120
rect 9647 86 9659 120
rect 6755 80 9659 86
rect 1545 -100 1653 80
rect 1545 -188 1555 -100
rect 1642 -188 1653 -100
rect 1545 -198 1653 -188
rect 4849 -100 4957 80
rect 4849 -188 4859 -100
rect 4946 -188 4957 -100
rect 4849 -198 4957 -188
rect 8153 -100 8261 80
rect 8153 -188 8163 -100
rect 8250 -188 8261 -100
rect 8153 -198 8261 -188
<< via1 >>
rect 286 179 338 1555
rect 682 179 734 1555
rect 1078 179 1130 1555
rect 1474 179 1526 1555
rect 1870 179 1922 1555
rect 2266 179 2318 1555
rect 2662 179 2714 1555
rect 3058 179 3110 1555
rect 3590 179 3599 1555
rect 3599 179 3633 1555
rect 3633 179 3642 1555
rect 3986 179 3995 1555
rect 3995 179 4029 1555
rect 4029 179 4038 1555
rect 4382 179 4391 1555
rect 4391 179 4425 1555
rect 4425 179 4434 1555
rect 4778 179 4787 1555
rect 4787 179 4821 1555
rect 4821 179 4830 1555
rect 5174 179 5183 1555
rect 5183 179 5217 1555
rect 5217 179 5226 1555
rect 5570 179 5579 1555
rect 5579 179 5613 1555
rect 5613 179 5622 1555
rect 5966 179 5975 1555
rect 5975 179 6009 1555
rect 6009 179 6018 1555
rect 6362 179 6371 1555
rect 6371 179 6405 1555
rect 6405 179 6414 1555
rect 6894 179 6903 1555
rect 6903 179 6937 1555
rect 6937 179 6946 1555
rect 7290 179 7299 1555
rect 7299 179 7333 1555
rect 7333 179 7342 1555
rect 7686 179 7695 1555
rect 7695 179 7729 1555
rect 7729 179 7738 1555
rect 8082 179 8091 1555
rect 8091 179 8125 1555
rect 8125 179 8134 1555
rect 8478 179 8487 1555
rect 8487 179 8521 1555
rect 8521 179 8530 1555
rect 8874 179 8883 1555
rect 8883 179 8917 1555
rect 8917 179 8926 1555
rect 9270 179 9279 1555
rect 9279 179 9313 1555
rect 9313 179 9322 1555
rect 9666 179 9675 1555
rect 9675 179 9709 1555
rect 9709 179 9718 1555
rect 1555 -188 1642 -100
rect 4859 -188 4946 -100
rect 8163 -188 8250 -100
<< metal2 >>
rect 286 1555 338 1565
rect 286 -305 338 179
rect 682 1555 734 1565
rect 682 -305 734 179
rect 1078 1555 1130 1565
rect 1078 -305 1130 179
rect 1474 1555 1526 1565
rect 1474 -305 1526 179
rect 1870 1555 1922 1565
rect 1555 -100 1642 -90
rect 1555 -198 1642 -188
rect 1870 -305 1922 179
rect 2266 1555 2318 1565
rect 2266 -305 2318 179
rect 2662 1555 2714 1565
rect 2662 -305 2714 179
rect 3058 1555 3110 1565
rect 3058 -305 3110 179
rect 3590 1555 3642 1565
rect 3590 -305 3642 179
rect 3986 1555 4038 1565
rect 3986 -305 4038 179
rect 4382 1555 4434 1565
rect 4382 -305 4434 179
rect 4778 1555 4830 1565
rect 4778 -305 4830 179
rect 5174 1555 5226 1565
rect 4859 -100 4946 -90
rect 4859 -198 4946 -188
rect 5174 -305 5226 179
rect 5570 1555 5622 1565
rect 5570 -305 5622 179
rect 5966 1555 6018 1565
rect 5966 -305 6018 179
rect 6362 1555 6414 1565
rect 6362 -305 6414 179
rect 6894 1555 6946 1565
rect 6894 -305 6946 179
rect 7290 1555 7342 1565
rect 7290 -305 7342 179
rect 7686 1555 7738 1565
rect 7686 -305 7738 179
rect 8082 1555 8134 1565
rect 8082 -305 8134 179
rect 8478 1555 8530 1565
rect 8163 -100 8250 -90
rect 8163 -198 8250 -188
rect 8478 -305 8530 179
rect 8874 1555 8926 1565
rect 8874 -305 8926 179
rect 9270 1555 9322 1565
rect 9270 -305 9322 179
rect 9666 1555 9718 1565
rect 9666 -305 9718 179
rect 271 -315 351 -305
rect 271 -375 281 -315
rect 341 -375 351 -315
rect 271 -385 351 -375
rect 667 -315 747 -305
rect 667 -375 677 -315
rect 737 -375 747 -315
rect 667 -385 747 -375
rect 1063 -315 1143 -305
rect 1063 -375 1073 -315
rect 1133 -375 1143 -315
rect 1063 -385 1143 -375
rect 1459 -315 1539 -305
rect 1459 -375 1469 -315
rect 1529 -375 1539 -315
rect 1459 -385 1539 -375
rect 1855 -315 1935 -305
rect 1855 -375 1865 -315
rect 1925 -375 1935 -315
rect 1855 -385 1935 -375
rect 2251 -315 2331 -305
rect 2251 -375 2261 -315
rect 2321 -375 2331 -315
rect 2251 -385 2331 -375
rect 2647 -315 2727 -305
rect 2647 -375 2657 -315
rect 2717 -375 2727 -315
rect 2647 -385 2727 -375
rect 3043 -315 3123 -305
rect 3043 -375 3053 -315
rect 3113 -375 3123 -315
rect 3043 -385 3123 -375
rect 3575 -315 3655 -305
rect 3575 -375 3585 -315
rect 3645 -375 3655 -315
rect 3575 -385 3655 -375
rect 3971 -315 4051 -305
rect 3971 -375 3981 -315
rect 4041 -375 4051 -315
rect 3971 -385 4051 -375
rect 4367 -315 4447 -305
rect 4367 -375 4377 -315
rect 4437 -375 4447 -315
rect 4367 -385 4447 -375
rect 4763 -315 4843 -305
rect 4763 -375 4773 -315
rect 4833 -375 4843 -315
rect 4763 -385 4843 -375
rect 5159 -315 5239 -305
rect 5159 -375 5169 -315
rect 5229 -375 5239 -315
rect 5159 -385 5239 -375
rect 5555 -315 5635 -305
rect 5555 -375 5565 -315
rect 5625 -375 5635 -315
rect 5555 -385 5635 -375
rect 5951 -315 6031 -305
rect 5951 -375 5961 -315
rect 6021 -375 6031 -315
rect 5951 -385 6031 -375
rect 6347 -315 6427 -305
rect 6347 -375 6357 -315
rect 6417 -375 6427 -315
rect 6347 -385 6427 -375
rect 6879 -315 6959 -305
rect 6879 -375 6889 -315
rect 6949 -375 6959 -315
rect 6879 -385 6959 -375
rect 7275 -315 7355 -305
rect 7275 -375 7285 -315
rect 7345 -375 7355 -315
rect 7275 -385 7355 -375
rect 7671 -315 7751 -305
rect 7671 -375 7681 -315
rect 7741 -375 7751 -315
rect 7671 -385 7751 -375
rect 8067 -315 8147 -305
rect 8067 -375 8077 -315
rect 8137 -375 8147 -315
rect 8067 -385 8147 -375
rect 8463 -315 8543 -305
rect 8463 -375 8473 -315
rect 8533 -375 8543 -315
rect 8463 -385 8543 -375
rect 8859 -315 8939 -305
rect 8859 -375 8869 -315
rect 8929 -375 8939 -315
rect 8859 -385 8939 -375
rect 9255 -315 9335 -305
rect 9255 -375 9265 -315
rect 9325 -375 9335 -315
rect 9255 -385 9335 -375
rect 9651 -315 9731 -305
rect 9651 -375 9661 -315
rect 9721 -375 9731 -315
rect 9651 -385 9731 -375
<< via2 >>
rect 1555 -188 1642 -100
rect 4859 -188 4946 -100
rect 8163 -188 8250 -100
rect 281 -375 341 -315
rect 677 -375 737 -315
rect 1073 -375 1133 -315
rect 1469 -375 1529 -315
rect 1865 -375 1925 -315
rect 2261 -375 2321 -315
rect 2657 -375 2717 -315
rect 3053 -375 3113 -315
rect 3585 -375 3645 -315
rect 3981 -375 4041 -315
rect 4377 -375 4437 -315
rect 4773 -375 4833 -315
rect 5169 -375 5229 -315
rect 5565 -375 5625 -315
rect 5961 -375 6021 -315
rect 6357 -375 6417 -315
rect 6889 -375 6949 -315
rect 7285 -375 7345 -315
rect 7681 -375 7741 -315
rect 8077 -375 8137 -315
rect 8473 -375 8533 -315
rect 8869 -375 8929 -315
rect 9265 -375 9325 -315
rect 9661 -375 9721 -315
<< metal3 >>
rect 1545 -100 8261 -90
rect 1545 -188 1555 -100
rect 1642 -188 4859 -100
rect 4946 -188 8163 -100
rect 8250 -188 8261 -100
rect 1545 -198 8261 -188
rect 271 -315 9735 -305
rect 271 -375 281 -315
rect 341 -375 677 -315
rect 737 -375 1073 -315
rect 1133 -375 1469 -315
rect 1529 -375 1865 -315
rect 1925 -375 2261 -315
rect 2321 -375 2657 -315
rect 2717 -375 3053 -315
rect 3113 -375 3585 -315
rect 3645 -375 3981 -315
rect 4041 -375 4377 -315
rect 4437 -375 4773 -315
rect 4833 -375 5169 -315
rect 5229 -375 5565 -315
rect 5625 -375 5961 -315
rect 6021 -375 6357 -315
rect 6417 -375 6889 -315
rect 6949 -375 7285 -315
rect 7345 -375 7681 -315
rect 7741 -375 8077 -315
rect 8137 -375 8473 -315
rect 8533 -375 8869 -315
rect 8929 -375 9265 -315
rect 9325 -375 9661 -315
rect 9721 -375 9735 -315
rect 271 -385 9735 -375
use sky130_fd_pr__pfet_01v8_DDZS4V  sky130_fd_pr__pfet_01v8_DDZS4V_0
timestamp 1616017086
transform 1 0 1599 0 1 831
box -1652 -884 1652 884
<< end >>
