magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect 667 1042 702 1076
rect 129 919 187 925
rect 129 885 141 919
rect 129 879 187 885
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1042
rect 668 1023 702 1042
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 687 530 702 1023
rect 721 989 756 1023
rect 721 530 755 989
rect 2512 957 2547 991
rect 2513 938 2547 957
rect 867 921 925 927
rect 867 887 879 921
rect 1037 898 1071 916
rect 867 881 925 887
rect 1037 862 1107 898
rect 1054 828 1125 862
rect 1405 828 1440 862
rect 1828 845 1863 863
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1054 477 1124 828
rect 1406 809 1440 828
rect 1792 830 1863 845
rect 1236 760 1294 766
rect 1236 726 1248 760
rect 1236 720 1294 726
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1425 424 1440 809
rect 1459 775 1494 809
rect 1459 424 1493 775
rect 1605 707 1663 713
rect 1605 673 1617 707
rect 1605 667 1663 673
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2163 318 2178 864
rect 2197 318 2231 918
rect 2343 889 2401 895
rect 2343 855 2355 889
rect 2343 849 2401 855
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2532 265 2547 938
rect 2566 904 2601 938
rect 2566 265 2600 904
rect 2712 836 2770 842
rect 2712 802 2724 836
rect 2712 796 2770 802
rect 2882 633 2916 651
rect 4726 639 4761 673
rect 2882 597 2952 633
rect 4727 620 4761 639
rect 2899 563 2970 597
rect 3250 563 3285 597
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 2899 212 2969 563
rect 3251 544 3285 563
rect 3081 495 3139 501
rect 3081 461 3093 495
rect 3081 455 3139 461
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2899 176 2952 212
rect 3270 159 3285 544
rect 3304 510 3339 544
rect 3619 510 3654 544
rect 4042 527 4077 545
rect 3304 159 3338 510
rect 3620 491 3654 510
rect 4006 512 4077 527
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 491
rect 3673 457 3708 491
rect 3673 106 3707 457
rect 3819 389 3877 395
rect 3819 355 3831 389
rect 3819 349 3877 355
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4006 53 4076 512
rect 4188 444 4246 450
rect 4188 410 4200 444
rect 4188 404 4246 410
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4006 17 4059 53
rect 4377 0 4392 546
rect 4411 0 4445 600
rect 4557 571 4615 577
rect 4557 537 4569 571
rect 4557 531 4615 537
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 620
rect 4780 586 4815 620
rect 4780 -53 4814 586
rect 4926 518 4984 524
rect 4926 484 4938 518
rect 4926 478 4984 484
rect 5096 315 5130 333
rect 5096 279 5166 315
rect 5113 245 5184 279
rect 5464 245 5499 279
rect 5887 262 5922 280
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5113 -106 5183 245
rect 5465 226 5499 245
rect 5851 247 5922 262
rect 5295 177 5353 183
rect 5295 143 5307 177
rect 5295 137 5353 143
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5113 -142 5166 -106
rect 5484 -159 5499 226
rect 5518 192 5553 226
rect 5518 -159 5552 192
rect 5664 124 5722 130
rect 5664 90 5676 124
rect 5664 84 5722 90
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5518 -193 5533 -159
rect 5851 -212 5921 247
rect 6033 179 6091 185
rect 6033 145 6045 179
rect 6203 156 6237 174
rect 6033 139 6091 145
rect 6203 120 6273 156
rect 6220 86 6291 120
rect 6571 86 6606 120
rect 6994 103 7029 121
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5851 -248 5904 -212
rect 6220 -265 6290 86
rect 6572 67 6606 86
rect 6958 88 7029 103
rect 7309 88 7344 122
rect 6402 18 6460 24
rect 6402 -16 6414 18
rect 6402 -22 6460 -16
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6220 -301 6273 -265
rect 6591 -318 6606 67
rect 6625 33 6660 67
rect 6625 -318 6659 33
rect 6771 -35 6829 -29
rect 6771 -69 6783 -35
rect 6771 -75 6829 -69
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6625 -352 6640 -318
rect 6958 -371 7028 88
rect 7310 69 7344 88
rect 7140 20 7198 26
rect 7140 -14 7152 20
rect 7140 -20 7198 -14
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6958 -407 7011 -371
rect 7329 -424 7344 69
rect 7363 35 7398 69
rect 7363 -424 7397 35
rect 7509 -33 7567 -27
rect 7509 -67 7521 -33
rect 7679 -56 7713 -38
rect 7509 -73 7567 -67
rect 7679 -92 7749 -56
rect 7696 -126 7767 -92
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7363 -458 7378 -424
rect 7696 -477 7766 -126
rect 7878 -194 7936 -188
rect 7878 -228 7890 -194
rect 7878 -234 7936 -228
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7696 -513 7749 -477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use sky130_fd_pr__pfet_01v8_XYCVAL  XM6
timestamp 1624053917
transform 1 0 2372 0 1 628
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM7
timestamp 1624053917
transform 1 0 2741 0 1 575
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM8
timestamp 1624053917
transform 1 0 3110 0 1 378
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM10
timestamp 1624053917
transform 1 0 3848 0 1 272
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM14
timestamp 1624053917
transform 1 0 5324 0 1 60
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM13
timestamp 1624053917
transform 1 0 4955 0 1 257
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM12
timestamp 1624053917
transform 1 0 4586 0 1 310
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XSLFBL  XM11
timestamp 1624053917
transform 1 0 4217 0 1 273
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM18
timestamp 1624053917
transform 1 0 6800 0 1 -152
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM17
timestamp 1624053917
transform 1 0 6431 0 1 -99
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM16
timestamp 1624053917
transform 1 0 6062 0 1 8
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM15
timestamp 1624053917
transform 1 0 5693 0 1 7
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM21
timestamp 1624053917
transform 1 0 7907 0 1 -311
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM20
timestamp 1624053917
transform 1 0 7538 0 1 -204
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM19
timestamp 1624053917
transform 1 0 7169 0 1 -151
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM0
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM3
timestamp 1624053917
transform 1 0 1265 0 1 643
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1624053917
transform 1 0 1634 0 1 590
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Q
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 D
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 CLK
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 CLR
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Qb
port 7 nsew
<< end >>
