magic
tech sky130A
magscale 1 2
timestamp 1623095677
<< nwell >>
rect -1127 -1234 1161 1234
<< pmos >>
rect -931 -1014 -861 1086
rect -803 -1014 -733 1086
rect -675 -1014 -605 1086
rect -547 -1014 -477 1086
rect -419 -1014 -349 1086
rect -291 -1014 -221 1086
rect -163 -1014 -93 1086
rect -35 -1014 35 1086
rect 93 -1014 163 1086
rect 221 -1014 291 1086
rect 349 -1014 419 1086
rect 477 -1014 547 1086
rect 605 -1014 675 1086
rect 733 -1014 803 1086
rect 861 -1014 931 1086
<< pdiff >>
rect -989 1074 -931 1086
rect -989 -1002 -977 1074
rect -943 -1002 -931 1074
rect -989 -1014 -931 -1002
rect -861 1074 -803 1086
rect -861 -1002 -849 1074
rect -815 -1002 -803 1074
rect -861 -1014 -803 -1002
rect -733 1074 -675 1086
rect -733 -1002 -721 1074
rect -687 -1002 -675 1074
rect -733 -1014 -675 -1002
rect -605 1074 -547 1086
rect -605 -1002 -593 1074
rect -559 -1002 -547 1074
rect -605 -1014 -547 -1002
rect -477 1074 -419 1086
rect -477 -1002 -465 1074
rect -431 -1002 -419 1074
rect -477 -1014 -419 -1002
rect -349 1074 -291 1086
rect -349 -1002 -337 1074
rect -303 -1002 -291 1074
rect -349 -1014 -291 -1002
rect -221 1074 -163 1086
rect -221 -1002 -209 1074
rect -175 -1002 -163 1074
rect -221 -1014 -163 -1002
rect -93 1074 -35 1086
rect -93 -1002 -81 1074
rect -47 -1002 -35 1074
rect -93 -1014 -35 -1002
rect 35 1074 93 1086
rect 35 -1002 47 1074
rect 81 -1002 93 1074
rect 35 -1014 93 -1002
rect 163 1074 221 1086
rect 163 -1002 175 1074
rect 209 -1002 221 1074
rect 163 -1014 221 -1002
rect 291 1074 349 1086
rect 291 -1002 303 1074
rect 337 -1002 349 1074
rect 291 -1014 349 -1002
rect 419 1074 477 1086
rect 419 -1002 431 1074
rect 465 -1002 477 1074
rect 419 -1014 477 -1002
rect 547 1074 605 1086
rect 547 -1002 559 1074
rect 593 -1002 605 1074
rect 547 -1014 605 -1002
rect 675 1074 733 1086
rect 675 -1002 687 1074
rect 721 -1002 733 1074
rect 675 -1014 733 -1002
rect 803 1074 861 1086
rect 803 -1002 815 1074
rect 849 -1002 861 1074
rect 803 -1014 861 -1002
rect 931 1074 989 1086
rect 931 -1002 943 1074
rect 977 -1002 989 1074
rect 931 -1014 989 -1002
<< pdiffc >>
rect -977 -1002 -943 1074
rect -849 -1002 -815 1074
rect -721 -1002 -687 1074
rect -593 -1002 -559 1074
rect -465 -1002 -431 1074
rect -337 -1002 -303 1074
rect -209 -1002 -175 1074
rect -81 -1002 -47 1074
rect 47 -1002 81 1074
rect 175 -1002 209 1074
rect 303 -1002 337 1074
rect 431 -1002 465 1074
rect 559 -1002 593 1074
rect 687 -1002 721 1074
rect 815 -1002 849 1074
rect 943 -1002 977 1074
<< nsubdiff >>
rect -1091 1164 -995 1198
rect 995 1164 1125 1198
rect -1091 1101 -1057 1164
rect 1057 1101 1125 1164
rect -1091 -1164 -1057 -1101
rect 1057 -1039 1125 -1014
rect -1091 -1198 -995 -1164
rect 995 -1198 1125 -1164
<< nsubdiffcont >>
rect -995 1164 995 1198
rect -1091 -1101 -1057 1101
rect 1057 -1014 1125 1101
rect -995 -1198 995 -1164
<< poly >>
rect -931 1086 -861 1112
rect -803 1086 -733 1112
rect -675 1086 -605 1112
rect -547 1086 -477 1112
rect -419 1086 -349 1112
rect -291 1086 -221 1112
rect -163 1086 -93 1112
rect -35 1086 35 1112
rect 93 1086 163 1112
rect 221 1086 291 1112
rect 349 1086 419 1112
rect 477 1086 547 1112
rect 605 1086 675 1112
rect 733 1086 803 1112
rect 861 1086 931 1112
rect -931 -1061 -861 -1014
rect -931 -1095 -915 -1061
rect -877 -1095 -861 -1061
rect -931 -1111 -861 -1095
rect -803 -1061 -733 -1014
rect -803 -1095 -787 -1061
rect -749 -1095 -733 -1061
rect -803 -1111 -733 -1095
rect -675 -1061 -605 -1014
rect -675 -1095 -659 -1061
rect -621 -1095 -605 -1061
rect -675 -1111 -605 -1095
rect -547 -1061 -477 -1014
rect -547 -1095 -531 -1061
rect -493 -1095 -477 -1061
rect -547 -1111 -477 -1095
rect -419 -1061 -349 -1014
rect -419 -1095 -403 -1061
rect -365 -1095 -349 -1061
rect -419 -1111 -349 -1095
rect -291 -1061 -221 -1014
rect -291 -1095 -275 -1061
rect -237 -1095 -221 -1061
rect -291 -1111 -221 -1095
rect -163 -1061 -93 -1014
rect -163 -1095 -147 -1061
rect -109 -1095 -93 -1061
rect -163 -1111 -93 -1095
rect -35 -1061 35 -1014
rect -35 -1095 -19 -1061
rect 19 -1095 35 -1061
rect -35 -1111 35 -1095
rect 93 -1061 163 -1014
rect 93 -1095 109 -1061
rect 147 -1095 163 -1061
rect 93 -1111 163 -1095
rect 221 -1061 291 -1014
rect 221 -1095 237 -1061
rect 275 -1095 291 -1061
rect 221 -1111 291 -1095
rect 349 -1061 419 -1014
rect 349 -1095 365 -1061
rect 403 -1095 419 -1061
rect 349 -1111 419 -1095
rect 477 -1061 547 -1014
rect 477 -1095 493 -1061
rect 531 -1095 547 -1061
rect 477 -1111 547 -1095
rect 605 -1061 675 -1014
rect 605 -1095 621 -1061
rect 659 -1095 675 -1061
rect 605 -1111 675 -1095
rect 733 -1061 803 -1014
rect 733 -1095 749 -1061
rect 787 -1095 803 -1061
rect 733 -1111 803 -1095
rect 861 -1061 931 -1014
rect 861 -1095 877 -1061
rect 915 -1095 931 -1061
rect 861 -1111 931 -1095
<< polycont >>
rect -915 -1095 -877 -1061
rect -787 -1095 -749 -1061
rect -659 -1095 -621 -1061
rect -531 -1095 -493 -1061
rect -403 -1095 -365 -1061
rect -275 -1095 -237 -1061
rect -147 -1095 -109 -1061
rect -19 -1095 19 -1061
rect 109 -1095 147 -1061
rect 237 -1095 275 -1061
rect 365 -1095 403 -1061
rect 493 -1095 531 -1061
rect 621 -1095 659 -1061
rect 749 -1095 787 -1061
rect 877 -1095 915 -1061
<< locali >>
rect -1091 1164 -995 1198
rect 995 1164 1125 1198
rect -1091 1101 -1057 1164
rect 1057 1101 1125 1164
rect -977 1074 -943 1090
rect -977 -1018 -943 -1002
rect -849 1074 -815 1090
rect -849 -1018 -815 -1002
rect -721 1074 -687 1090
rect -721 -1018 -687 -1002
rect -593 1074 -559 1090
rect -593 -1018 -559 -1002
rect -465 1074 -431 1090
rect -465 -1018 -431 -1002
rect -337 1074 -303 1090
rect -337 -1018 -303 -1002
rect -209 1074 -175 1090
rect -209 -1018 -175 -1002
rect -81 1074 -47 1090
rect -81 -1018 -47 -1002
rect 47 1074 81 1090
rect 47 -1018 81 -1002
rect 175 1074 209 1090
rect 175 -1018 209 -1002
rect 303 1074 337 1090
rect 303 -1018 337 -1002
rect 431 1074 465 1090
rect 431 -1018 465 -1002
rect 559 1074 593 1090
rect 559 -1018 593 -1002
rect 687 1074 721 1090
rect 687 -1018 721 -1002
rect 815 1074 849 1090
rect 815 -1018 849 -1002
rect 943 1074 977 1090
rect 943 -1018 977 -1002
rect 1057 -1039 1125 -1014
rect -931 -1095 -915 -1061
rect -877 -1095 -861 -1061
rect -803 -1095 -787 -1061
rect -749 -1095 -733 -1061
rect -675 -1095 -659 -1061
rect -621 -1095 -605 -1061
rect -547 -1095 -531 -1061
rect -493 -1095 -477 -1061
rect -419 -1095 -403 -1061
rect -365 -1095 -349 -1061
rect -291 -1095 -275 -1061
rect -237 -1095 -221 -1061
rect -163 -1095 -147 -1061
rect -109 -1095 -93 -1061
rect -35 -1095 -19 -1061
rect 19 -1095 35 -1061
rect 93 -1095 109 -1061
rect 147 -1095 163 -1061
rect 221 -1095 237 -1061
rect 275 -1095 291 -1061
rect 349 -1095 365 -1061
rect 403 -1095 419 -1061
rect 477 -1095 493 -1061
rect 531 -1095 547 -1061
rect 605 -1095 621 -1061
rect 659 -1095 675 -1061
rect 733 -1095 749 -1061
rect 787 -1095 803 -1061
rect 861 -1095 877 -1061
rect 915 -1095 931 -1061
rect -1091 -1164 -1057 -1101
rect -1091 -1198 -995 -1164
rect 995 -1198 1125 -1164
<< viali >>
rect -977 -1002 -943 1074
rect -849 -1002 -815 1074
rect -721 -1002 -687 1074
rect -593 -1002 -559 1074
rect -465 -1002 -431 1074
rect -337 -1002 -303 1074
rect -209 -1002 -175 1074
rect -81 -1002 -47 1074
rect 47 -1002 81 1074
rect 175 -1002 209 1074
rect 303 -1002 337 1074
rect 431 -1002 465 1074
rect 559 -1002 593 1074
rect 687 -1002 721 1074
rect 815 -1002 849 1074
rect 943 -1002 977 1074
rect -915 -1095 -877 -1061
rect -787 -1095 -749 -1061
rect -659 -1095 -621 -1061
rect -531 -1095 -493 -1061
rect -403 -1095 -365 -1061
rect -275 -1095 -237 -1061
rect -147 -1095 -109 -1061
rect -19 -1095 19 -1061
rect 109 -1095 147 -1061
rect 237 -1095 275 -1061
rect 365 -1095 403 -1061
rect 493 -1095 531 -1061
rect 621 -1095 659 -1061
rect 749 -1095 787 -1061
rect 877 -1095 915 -1061
<< metal1 >>
rect -983 1074 -937 1086
rect -983 -1002 -977 1074
rect -943 -1002 -937 1074
rect -983 -1014 -937 -1002
rect -855 1074 -809 1086
rect -855 -1002 -849 1074
rect -815 -1002 -809 1074
rect -855 -1014 -809 -1002
rect -727 1074 -681 1086
rect -727 -1002 -721 1074
rect -687 -1002 -681 1074
rect -727 -1014 -681 -1002
rect -599 1074 -553 1086
rect -599 -1002 -593 1074
rect -559 -1002 -553 1074
rect -599 -1014 -553 -1002
rect -471 1074 -425 1086
rect -471 -1002 -465 1074
rect -431 -1002 -425 1074
rect -471 -1014 -425 -1002
rect -343 1074 -297 1086
rect -343 -1002 -337 1074
rect -303 -1002 -297 1074
rect -343 -1014 -297 -1002
rect -215 1074 -169 1086
rect -215 -1002 -209 1074
rect -175 -1002 -169 1074
rect -215 -1014 -169 -1002
rect -87 1074 -41 1086
rect -87 -1002 -81 1074
rect -47 -1002 -41 1074
rect -87 -1014 -41 -1002
rect 41 1074 87 1086
rect 41 -1002 47 1074
rect 81 -1002 87 1074
rect 41 -1014 87 -1002
rect 169 1074 215 1086
rect 169 -1002 175 1074
rect 209 -1002 215 1074
rect 169 -1014 215 -1002
rect 297 1074 343 1086
rect 297 -1002 303 1074
rect 337 -1002 343 1074
rect 297 -1014 343 -1002
rect 425 1074 471 1086
rect 425 -1002 431 1074
rect 465 -1002 471 1074
rect 425 -1014 471 -1002
rect 553 1074 599 1086
rect 553 -1002 559 1074
rect 593 -1002 599 1074
rect 553 -1014 599 -1002
rect 681 1074 727 1086
rect 681 -1002 687 1074
rect 721 -1002 727 1074
rect 681 -1014 727 -1002
rect 809 1074 855 1086
rect 809 -1002 815 1074
rect 849 -1002 855 1074
rect 809 -1014 855 -1002
rect 937 1074 983 1086
rect 937 -1002 943 1074
rect 977 -1002 983 1074
rect 937 -1014 983 -1002
rect -931 -1061 931 -1055
rect -931 -1095 -915 -1061
rect -877 -1095 -787 -1061
rect -749 -1095 -659 -1061
rect -621 -1095 -531 -1061
rect -493 -1095 -403 -1061
rect -365 -1095 -275 -1061
rect -237 -1095 -147 -1061
rect -109 -1095 -19 -1061
rect 19 -1095 109 -1061
rect 147 -1095 237 -1061
rect 275 -1095 365 -1061
rect 403 -1095 493 -1061
rect 531 -1095 621 -1061
rect 659 -1095 749 -1061
rect 787 -1095 877 -1061
rect 915 -1095 931 -1061
rect -931 -1101 931 -1095
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1074 -1181 1074 1181
string parameters w 10.5 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
