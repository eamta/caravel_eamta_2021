magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< nwell >>
rect -17 306 296 869
<< pwell >>
rect -17 -20 296 306
<< psubdiff >>
rect 180 -3 204 31
rect 239 -3 263 31
<< nsubdiff >>
rect 148 794 172 828
rect 206 794 231 828
<< psubdiffcont >>
rect 204 -3 239 31
<< nsubdiffcont >>
rect 172 794 206 828
<< poly >>
rect 80 340 110 375
rect 168 340 198 385
rect 44 324 110 340
rect 44 290 60 324
rect 94 290 110 324
rect 44 274 110 290
rect 152 324 218 340
rect 152 290 168 324
rect 202 290 218 324
rect 152 274 218 290
rect 80 202 110 274
rect 168 202 198 274
<< polycont >>
rect 60 290 94 324
rect 168 290 202 324
<< locali >>
rect 44 324 109 340
rect 44 290 60 324
rect 94 290 109 324
rect 44 274 109 290
rect 152 324 218 340
rect 152 290 168 324
rect 202 290 218 324
rect 152 274 218 290
<< viali >>
rect 148 794 172 828
rect 172 794 206 828
rect 206 794 231 828
rect 60 290 94 324
rect 168 290 202 324
rect 180 -3 204 31
rect 204 -3 239 31
rect 239 -3 263 31
<< metal1 >>
rect -14 828 292 835
rect -14 794 148 828
rect 231 794 292 828
rect -14 789 292 794
rect 34 368 68 789
rect 136 788 243 789
rect 204 378 290 738
rect 44 324 109 340
rect 44 290 60 324
rect 94 290 109 324
rect 44 274 109 290
rect 152 324 218 340
rect 152 290 168 324
rect 202 290 218 324
rect 152 274 218 290
rect 256 243 290 378
rect 122 209 290 243
rect 34 35 68 181
rect 122 87 156 209
rect 210 37 244 181
rect 168 35 275 37
rect -17 31 296 35
rect -17 -3 180 31
rect 263 -3 296 31
rect -17 -11 296 -3
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_0
timestamp 1615302329
transform 1 0 95 0 1 558
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_1
timestamp 1615302329
transform 1 0 183 0 1 558
box -109 -242 109 242
use sky130_fd_pr__nfet_01v8_NNQ2PV  sky130_fd_pr__nfet_01v8_NNQ2PV_0
timestamp 1615600491
transform 1 0 95 0 1 136
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_NNQ2PV  sky130_fd_pr__nfet_01v8_NNQ2PV_1
timestamp 1615600491
transform 1 0 183 0 1 136
box -73 -71 73 71
<< labels >>
rlabel nwell 172 794 206 828 1 vdd!
rlabel pwell 180 -3 263 31 1 vss!
<< end >>
