magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 2619 4771 4272 4806
rect 2971 4695 3068 4716
rect 3098 4695 3175 4716
rect 3716 4695 3793 4716
rect 3823 4695 3920 4716
rect 2999 4667 3068 4688
rect 3098 4667 3175 4688
rect 3716 4667 3793 4688
rect 3823 4667 3892 4688
rect 7734 4654 7769 4688
rect 3414 4633 3432 4645
rect 3460 4633 3462 4644
rect 3383 4630 3432 4633
rect -491 4161 -438 4618
rect 3383 4570 3420 4630
rect 3429 4570 3432 4630
rect 3383 4567 3432 4570
rect 3471 4567 3508 4633
rect 7365 4618 7400 4635
rect 7329 4601 7400 4618
rect 3414 4555 3432 4567
rect 6996 4548 7031 4582
rect 229 4495 264 4529
rect 230 4476 264 4495
rect 6627 4495 6662 4529
rect 60 4427 118 4433
rect 60 4393 72 4427
rect 60 4387 118 4393
rect 60 4119 118 4125
rect 60 4085 72 4119
rect 60 4079 118 4085
rect 249 3983 264 4476
rect 283 4442 318 4476
rect 598 4442 633 4476
rect 283 3983 317 4442
rect 599 4423 633 4442
rect 6258 4442 6293 4476
rect 429 4374 487 4380
rect 429 4340 441 4374
rect 429 4334 487 4340
rect 429 4066 487 4072
rect 429 4032 441 4066
rect 429 4026 487 4032
rect 283 3949 298 3983
rect 618 3930 633 4423
rect 652 4389 687 4423
rect 967 4389 1002 4423
rect 652 3930 686 4389
rect 968 4370 1002 4389
rect 5889 4389 5924 4423
rect 798 4321 856 4327
rect 798 4287 810 4321
rect 798 4281 856 4287
rect 798 4013 856 4019
rect 798 3979 810 4013
rect 798 3973 856 3979
rect 652 3896 667 3930
rect 987 3877 1002 4370
rect 1021 4336 1056 4370
rect 1336 4336 1371 4370
rect 1021 3877 1055 4336
rect 1337 4317 1371 4336
rect 3412 4332 3441 4354
rect 3397 4320 3441 4332
rect 3450 4332 3479 4354
rect 5520 4336 5555 4370
rect 3450 4320 3494 4332
rect 1167 4268 1225 4274
rect 1167 4234 1179 4268
rect 1167 4228 1225 4234
rect 1167 3960 1225 3966
rect 1167 3926 1179 3960
rect 1167 3920 1225 3926
rect 1021 3843 1036 3877
rect 1356 3824 1371 4317
rect 1390 4283 1425 4317
rect 1705 4300 1740 4317
rect 3397 4304 3429 4320
rect 3462 4304 3494 4320
rect 5151 4300 5186 4317
rect 1705 4283 1776 4300
rect 1390 3824 1424 4283
rect 1706 4264 1776 4283
rect 5115 4283 5186 4300
rect 1723 4230 1794 4264
rect 2074 4230 2109 4264
rect 1536 4215 1594 4221
rect 1536 4181 1548 4215
rect 1536 4175 1594 4181
rect 1536 3907 1594 3913
rect 1536 3873 1548 3907
rect 1536 3867 1594 3873
rect 1390 3790 1405 3824
rect 1723 3771 1793 4230
rect 2075 4211 2109 4230
rect 1905 4162 1963 4168
rect 1905 4128 1917 4162
rect 1905 4122 1963 4128
rect 1905 3872 1963 3878
rect 1905 3838 1917 3872
rect 1905 3832 1963 3838
rect 1723 3735 1776 3771
rect 2094 3736 2109 4211
rect 2128 4177 2163 4211
rect 2443 4177 2478 4211
rect 2128 3736 2162 4177
rect 2444 4158 2478 4177
rect 2274 4109 2332 4115
rect 2274 4075 2286 4109
rect 2274 4069 2332 4075
rect 2274 3819 2332 3825
rect 2274 3785 2286 3819
rect 2325 3785 2332 3819
rect 2274 3779 2332 3785
rect 2353 3751 2360 3811
rect 2128 3702 2143 3736
rect 2463 3683 2478 4158
rect 2497 4124 2532 4158
rect 2552 4141 2883 4194
rect 3309 4184 3311 4245
rect 3337 4212 3339 4273
rect 3414 4233 3432 4245
rect 3460 4233 3462 4244
rect 3383 4230 3432 4233
rect 2497 3683 2531 4124
rect 2552 3937 3252 4141
rect 3383 4080 3420 4230
rect 3429 4080 3432 4230
rect 3383 4077 3432 4080
rect 3471 4077 3508 4233
rect 3552 4212 3554 4273
rect 3580 4184 3582 4245
rect 4782 4230 4817 4264
rect 4008 4141 4339 4194
rect 4413 4177 4448 4211
rect 3414 4065 3432 4077
rect 3639 3937 4339 4141
rect 2552 3903 4339 3937
rect 2552 3867 3252 3903
rect 3639 3867 4339 3903
rect 2611 3816 2645 3867
rect 2699 3816 2733 3867
rect 2643 3766 2701 3772
rect 2643 3732 2655 3766
rect 2643 3726 2701 3732
rect 2497 3649 2512 3683
rect 2832 3630 2847 3867
rect 2866 3630 2900 3867
rect 2866 3596 2881 3630
rect 4010 3596 4025 3867
rect 4044 3664 4078 3867
rect 4158 3816 4192 3867
rect 4246 3816 4280 3867
rect 4190 3766 4248 3772
rect 4190 3732 4202 3766
rect 4190 3726 4248 3732
rect 4044 3630 4079 3664
rect 4379 3649 4394 4158
rect 4413 3717 4447 4177
rect 4559 4109 4617 4115
rect 4559 4075 4571 4109
rect 4559 4069 4617 4075
rect 4559 3819 4617 3825
rect 4531 3751 4538 3811
rect 4559 3785 4571 3819
rect 4559 3779 4617 3785
rect 4413 3683 4448 3717
rect 4748 3702 4763 4211
rect 4782 3770 4816 4230
rect 4928 4162 4986 4168
rect 4928 4128 4940 4162
rect 4928 4122 4986 4128
rect 4928 3872 4986 3878
rect 4928 3838 4940 3872
rect 4928 3832 4986 3838
rect 5115 3805 5185 4283
rect 5297 4215 5355 4221
rect 5297 4181 5309 4215
rect 5297 4175 5355 4181
rect 5297 3907 5355 3913
rect 5297 3873 5309 3907
rect 5297 3867 5355 3873
rect 5115 3771 5186 3805
rect 5486 3790 5501 4317
rect 5520 3858 5554 4336
rect 5666 4268 5724 4274
rect 5666 4234 5678 4268
rect 5666 4228 5724 4234
rect 5666 3960 5724 3966
rect 5666 3926 5678 3960
rect 5666 3920 5724 3926
rect 5520 3824 5555 3858
rect 5855 3843 5870 4370
rect 5889 3911 5923 4389
rect 6035 4321 6093 4327
rect 6035 4287 6047 4321
rect 6035 4281 6093 4287
rect 6035 4013 6093 4019
rect 6035 3979 6047 4013
rect 6035 3973 6093 3979
rect 5889 3877 5924 3911
rect 6224 3896 6239 4423
rect 6258 3964 6292 4442
rect 6404 4374 6462 4380
rect 6404 4340 6416 4374
rect 6404 4334 6462 4340
rect 6404 4066 6462 4072
rect 6404 4032 6416 4066
rect 6404 4026 6462 4032
rect 6258 3930 6293 3964
rect 6593 3949 6608 4476
rect 6627 4017 6661 4495
rect 6773 4427 6831 4433
rect 6773 4393 6785 4427
rect 6773 4387 6831 4393
rect 6773 4119 6831 4125
rect 6773 4085 6785 4119
rect 6773 4079 6831 4085
rect 6627 3983 6662 4017
rect 6962 4002 6977 4529
rect 6996 4070 7030 4548
rect 7142 4480 7200 4486
rect 7142 4446 7154 4480
rect 7142 4440 7200 4446
rect 7329 4231 7399 4601
rect 7511 4533 7569 4539
rect 7511 4499 7523 4533
rect 7511 4493 7569 4499
rect 7511 4333 7569 4339
rect 7511 4299 7523 4333
rect 7511 4293 7569 4299
rect 7329 4197 7400 4231
rect 7700 4216 7715 4635
rect 7734 4284 7768 4654
rect 7880 4586 7938 4592
rect 7880 4552 7892 4586
rect 7880 4546 7938 4552
rect 7880 4386 7938 4392
rect 7880 4352 7892 4386
rect 7880 4346 7938 4352
rect 7734 4250 7769 4284
rect 7142 4172 7200 4178
rect 7142 4138 7154 4172
rect 7329 4161 7382 4197
rect 7142 4132 7200 4138
rect 6996 4036 7031 4070
rect 4782 3736 4817 3770
rect 5115 3735 5168 3771
rect 194 2281 229 2315
rect 3608 2281 3643 2315
rect 7022 2281 7057 2315
rect 10436 2281 10471 2315
rect 195 2262 229 2281
rect 3609 2262 3643 2281
rect 7023 2262 7057 2281
rect 10437 2262 10471 2281
rect 25 2213 83 2219
rect 25 2179 37 2213
rect 25 2173 83 2179
rect 87 1968 127 1986
rect 214 1968 229 2262
rect 248 2228 283 2262
rect 248 1968 282 2228
rect 394 2160 452 2166
rect 394 2126 406 2160
rect 394 2120 452 2126
rect 362 1974 396 2008
rect 450 1974 484 2008
rect 564 1974 598 2173
rect 986 2155 1021 2173
rect 950 2140 1021 2155
rect 1301 2140 1336 2174
rect 617 2085 652 2119
rect 617 1974 651 2085
rect 950 2023 1020 2140
rect 1302 2121 1336 2140
rect 1132 2072 1190 2078
rect 1132 2038 1144 2072
rect 1132 2032 1190 2038
rect 775 2008 809 2012
rect 759 1983 825 2008
rect 933 2000 1020 2023
rect 933 1974 1088 2000
rect 1100 1974 1134 2008
rect 1188 1974 1222 2008
rect 1321 2000 1336 2121
rect 1355 2087 1390 2121
rect 1670 2087 1705 2121
rect 1355 2000 1389 2087
rect 1671 2068 1705 2087
rect 1234 1974 1302 2000
rect 1321 1974 1389 2000
rect 291 1968 1020 1974
rect -140 1941 1020 1968
rect 1066 1941 1234 1974
rect 1302 1941 1389 1974
rect -140 1940 1389 1941
rect -140 1929 366 1940
rect 481 1929 496 1940
rect -140 1879 408 1929
rect 416 1880 426 1921
rect 438 1908 496 1929
rect 438 1899 498 1908
rect 438 1879 488 1899
rect -1524 1777 -1489 1811
rect -1523 1758 -1489 1777
rect -140 1792 366 1879
rect 393 1836 394 1879
rect 406 1836 440 1839
rect -140 1768 391 1792
rect 439 1768 469 1785
rect 564 1768 598 1940
rect -140 1759 502 1768
rect 516 1759 568 1768
rect 583 1763 598 1768
rect 583 1759 603 1763
rect -1693 1709 -1635 1715
rect -1693 1675 -1681 1709
rect -1693 1669 -1635 1675
rect -1737 1581 -1679 1599
rect -1649 1581 -1591 1599
rect -1504 1581 -1489 1758
rect -1470 1724 -1435 1758
rect -1155 1741 -1120 1758
rect -1155 1724 -1084 1741
rect -1470 1581 -1436 1724
rect -1154 1705 -1084 1724
rect -140 1734 615 1759
rect -1137 1671 -1066 1705
rect -1024 1671 -751 1705
rect -1324 1656 -1266 1662
rect -1324 1636 -1312 1656
rect -1324 1634 -1310 1636
rect -1280 1634 -1278 1636
rect -1137 1634 -1067 1671
rect -785 1652 -751 1671
rect -766 1651 -751 1652
rect -732 1651 -697 1652
rect -1375 1581 -1067 1634
rect -970 1643 -785 1651
rect -417 1650 -382 1652
rect -970 1637 -717 1643
rect -970 1617 -859 1637
rect -819 1617 -717 1637
rect -655 1632 -382 1650
rect -140 1635 366 1734
rect 419 1672 427 1734
rect 381 1669 439 1672
rect 453 1669 487 1734
rect 583 1681 615 1734
rect 617 1715 651 1940
rect 719 1933 734 1940
rect 719 1929 765 1933
rect 719 1899 777 1929
rect 819 1902 853 1933
rect 933 1916 1020 1940
rect 1135 1916 1140 1921
rect 1163 1916 1168 1921
rect 1211 1916 1234 1925
rect 1321 1916 1336 1940
rect 719 1884 734 1899
rect 725 1873 731 1875
rect 719 1867 731 1873
rect 757 1870 777 1899
rect 853 1880 878 1885
rect 742 1867 777 1870
rect 719 1855 777 1867
rect 844 1865 865 1880
rect 813 1864 865 1865
rect 933 1864 1234 1916
rect 1246 1878 1256 1890
rect 731 1851 749 1855
rect 697 1837 711 1847
rect 757 1837 777 1855
rect 807 1863 1234 1864
rect 1242 1863 1256 1878
rect 1258 1874 1281 1878
rect 1258 1863 1292 1874
rect 1302 1863 1336 1916
rect 1355 1863 1389 1940
rect 1540 1880 1557 1914
rect 1589 1905 1603 1908
rect 1588 1890 1603 1905
rect 1558 1863 1603 1890
rect 1671 1893 1682 1904
rect 1690 1893 1705 2068
rect 1608 1863 1625 1880
rect 1671 1863 1705 1893
rect 1724 2034 1759 2068
rect 1724 1863 1758 2034
rect 3293 1968 3327 2219
rect 3395 1973 3441 1983
rect 3395 1968 3452 1973
rect 3501 1968 3541 1986
rect 3628 1968 3643 2262
rect 3662 2228 3697 2262
rect 3662 1968 3696 2228
rect 6853 2213 6911 2219
rect 6853 2179 6865 2213
rect 3978 2119 4012 2173
rect 4400 2155 4435 2173
rect 4364 2140 4435 2155
rect 4715 2140 4750 2174
rect 6853 2173 6911 2179
rect 3747 2099 3932 2116
rect 3770 2071 3816 2088
rect 3858 2071 3904 2088
rect 3274 1963 3780 1968
rect 1948 1928 2040 1954
rect 2074 1928 2110 1954
rect 3274 1929 3810 1963
rect 3864 1929 3898 1963
rect 1974 1923 2026 1928
rect 1906 1889 1957 1913
rect 1973 1895 2026 1923
rect 2040 1895 2074 1928
rect 2110 1895 2136 1928
rect 2986 1920 3932 1929
rect 2986 1895 3930 1920
rect 1973 1894 2136 1895
rect 3274 1894 3930 1895
rect 3978 1895 3983 1983
rect 3997 1895 4012 2119
rect 1906 1887 1960 1889
rect 1939 1885 1960 1887
rect 1826 1863 1828 1885
rect 807 1849 1828 1863
rect 1920 1859 1960 1885
rect 1935 1856 1960 1859
rect 807 1846 1866 1849
rect 2040 1848 2074 1894
rect 807 1837 878 1846
rect 697 1835 887 1837
rect 699 1827 887 1835
rect 699 1817 715 1827
rect 807 1814 859 1827
rect 867 1823 878 1827
rect 752 1770 759 1791
rect 810 1783 825 1814
rect 844 1798 859 1814
rect 933 1821 1866 1846
rect 1972 1834 2110 1848
rect 3274 1844 3780 1894
rect 3822 1886 3843 1894
rect 933 1810 1739 1821
rect 1758 1817 1866 1821
rect 1758 1810 1892 1817
rect 1947 1810 2110 1834
rect 2325 1818 2422 1839
rect 2452 1818 2529 1839
rect 867 1798 878 1803
rect 794 1744 828 1748
rect 694 1715 705 1744
rect 794 1715 840 1744
rect 844 1715 878 1798
rect 933 1780 2110 1810
rect 2353 1790 2422 1811
rect 2452 1790 2529 1811
rect 3259 1793 3780 1844
rect 3804 1870 3843 1886
rect 3804 1860 3870 1870
rect 3804 1841 3859 1860
rect 3867 1841 3870 1860
rect 3801 1836 3892 1841
rect 3801 1826 3859 1836
rect 3804 1820 3859 1826
rect 2155 1780 2189 1784
rect 933 1768 1972 1780
rect 933 1762 1994 1768
rect 933 1751 944 1762
rect 950 1757 1994 1762
rect 2040 1757 2074 1780
rect 2089 1757 2110 1780
rect 2143 1757 2189 1780
rect 933 1715 946 1728
rect 617 1681 669 1715
rect 694 1712 946 1715
rect 950 1712 2110 1757
rect 2155 1721 2189 1757
rect 2331 1722 2335 1755
rect 2337 1722 2465 1780
rect 2519 1722 2665 1762
rect 2725 1755 2774 1768
rect 2284 1721 2337 1722
rect 694 1681 2110 1712
rect 2143 1687 2337 1721
rect 419 1665 427 1669
rect -268 1632 366 1635
rect -655 1617 366 1632
rect -970 1609 -936 1617
rect -970 1603 -897 1609
rect -1744 1337 -1067 1581
rect -1506 1284 -1067 1337
rect -1562 1135 -1504 1141
rect -1562 1101 -1550 1135
rect -1373 1111 -1358 1284
rect -1339 1111 -1305 1284
rect -1135 1231 -1103 1284
rect -1101 1255 -1067 1284
rect -1023 1560 -1013 1564
rect -1004 1560 -989 1598
rect -1101 1197 -1069 1255
rect -1193 1188 -1135 1194
rect -1193 1154 -1181 1188
rect -1135 1154 -1131 1188
rect -1101 1159 -1097 1197
rect -1023 1193 -989 1560
rect -970 1583 -893 1603
rect -766 1587 -751 1617
rect -785 1583 -751 1587
rect -970 1569 -936 1583
rect -970 1563 -897 1569
rect -970 1526 -936 1563
rect -785 1555 -744 1583
rect -987 1338 -936 1526
rect -824 1549 -744 1555
rect -824 1515 -806 1549
rect -785 1515 -744 1549
rect -824 1509 -751 1515
rect -890 1494 -865 1506
rect -894 1354 -865 1494
rect -785 1499 -751 1509
rect -785 1490 -780 1499
rect -766 1490 -751 1499
rect -802 1472 -751 1490
rect -890 1342 -865 1354
rect -856 1456 -831 1472
rect -802 1456 -734 1472
rect -732 1468 -698 1617
rect -654 1601 366 1617
rect 453 1601 469 1669
rect 583 1665 603 1681
rect 794 1658 840 1681
rect 694 1654 840 1658
rect 794 1650 828 1654
rect 844 1618 878 1681
rect 950 1678 2110 1681
rect 930 1674 2110 1678
rect 918 1656 2110 1674
rect 2267 1686 2337 1687
rect 2465 1686 2533 1722
rect 2665 1687 2706 1722
rect 2725 1716 2780 1755
rect 3128 1739 3178 1793
rect 3232 1792 3780 1793
rect 3813 1798 3847 1820
rect 3901 1802 3904 1845
rect 3813 1792 3839 1798
rect 3232 1768 3901 1792
rect 3978 1768 4012 1895
rect 4031 2085 4066 2119
rect 4031 1768 4065 2085
rect 4364 2023 4434 2140
rect 4716 2121 4750 2140
rect 4068 1928 4099 1929
rect 4145 1928 4179 1962
rect 4233 1928 4267 1962
rect 4347 1954 4434 2023
rect 4518 2019 4538 2106
rect 4546 2072 4604 2078
rect 4546 2038 4566 2072
rect 4546 2032 4604 2038
rect 4480 2011 4538 2019
rect 4508 1983 4554 1991
rect 4347 1928 4502 1954
rect 4514 1928 4548 1979
rect 4602 1928 4636 1979
rect 4735 1954 4750 2121
rect 4769 2087 4804 2121
rect 5084 2087 5119 2121
rect 4769 1954 4803 2087
rect 5085 2068 5119 2087
rect 4849 1954 4893 1960
rect 4648 1928 4716 1954
rect 4735 1929 4893 1954
rect 4750 1928 4893 1929
rect 4068 1916 4434 1928
rect 4480 1916 4648 1928
rect 4068 1895 4648 1916
rect 4716 1895 4750 1928
rect 4769 1895 4803 1928
rect 4849 1926 4917 1928
rect 4849 1895 4927 1926
rect 4068 1894 4927 1895
rect 4133 1880 4148 1894
rect 4267 1880 4292 1885
rect 4347 1880 4644 1894
rect 4133 1855 4191 1880
rect 4131 1850 4191 1855
rect 4141 1833 4191 1850
rect 4173 1830 4191 1833
rect 4221 1863 4644 1880
rect 4716 1863 4750 1894
rect 4769 1863 4803 1894
rect 4883 1863 4917 1894
rect 5085 1893 5096 1904
rect 5104 1893 5119 2068
rect 5085 1863 5119 1893
rect 5138 2034 5173 2068
rect 5138 1863 5172 2034
rect 6915 1968 6955 1986
rect 7042 1968 7057 2262
rect 7076 2228 7111 2262
rect 7076 1968 7110 2228
rect 10267 2213 10325 2219
rect 10267 2179 10279 2213
rect 7222 2160 7280 2166
rect 7222 2126 7234 2160
rect 7222 2120 7280 2126
rect 7392 2119 7426 2173
rect 7814 2155 7849 2173
rect 7778 2140 7849 2155
rect 8129 2140 8164 2174
rect 10267 2173 10325 2179
rect 5280 1916 5298 1935
rect 5328 1916 5346 1932
rect 5279 1892 5320 1907
rect 5279 1886 5325 1892
rect 5340 1886 5363 1889
rect 5248 1885 5325 1886
rect 5328 1885 5378 1886
rect 5240 1863 5363 1885
rect 4221 1850 5255 1863
rect 4221 1846 4271 1850
rect 4347 1848 5255 1850
rect 4221 1833 4273 1846
rect 4221 1830 4239 1833
rect 4173 1783 4188 1806
rect 4189 1800 4204 1806
rect 4224 1800 4239 1817
rect 4189 1783 4239 1800
rect 4177 1777 4188 1783
rect 4204 1777 4235 1783
rect 4139 1768 4154 1772
rect 3232 1750 3947 1768
rect 3244 1746 3947 1750
rect 3274 1739 3947 1746
rect 2725 1687 2871 1716
rect 2665 1686 2871 1687
rect 930 1634 2110 1656
rect 2143 1652 2181 1657
rect 2267 1652 2665 1686
rect 2725 1678 2871 1686
rect 2737 1674 2771 1678
rect 2780 1674 2859 1678
rect 2143 1634 2201 1652
rect 2231 1634 2377 1652
rect 930 1618 2377 1634
rect 2407 1651 2453 1652
rect 2465 1651 2533 1652
rect 2636 1651 2665 1652
rect 2780 1669 2830 1674
rect 2956 1673 2990 1696
rect 3044 1673 3078 1696
rect 2780 1662 3075 1669
rect 3148 1662 3178 1739
rect 2780 1661 3178 1662
rect 3182 1734 3947 1739
rect 3995 1734 4012 1768
rect 4020 1734 4066 1768
rect 4139 1752 4166 1768
rect 4258 1766 4273 1833
rect 4347 1810 5251 1848
rect 5263 1846 5363 1863
rect 5263 1836 5298 1846
rect 5306 1834 5325 1846
rect 5328 1836 5329 1846
rect 5252 1821 5277 1833
rect 5252 1810 5281 1821
rect 5334 1812 5363 1846
rect 6660 1820 6666 1921
rect 5334 1810 5353 1812
rect 4347 1807 5382 1810
rect 4281 1788 4292 1799
rect 4238 1762 4273 1766
rect 4284 1762 4292 1788
rect 4226 1752 4292 1762
rect 4139 1749 4160 1752
rect 4232 1749 4235 1752
rect 4238 1745 4292 1752
rect 3182 1712 3780 1734
rect 3182 1681 3232 1712
rect 3274 1711 3780 1712
rect 2780 1654 3075 1661
rect 3090 1654 3120 1661
rect 3148 1654 3166 1661
rect 2780 1651 3166 1654
rect 2407 1630 2665 1651
rect 2703 1640 3166 1651
rect 2391 1624 2665 1630
rect 2759 1628 3166 1640
rect 2391 1618 2698 1624
rect 492 1601 569 1618
rect 802 1617 924 1618
rect -654 1600 569 1601
rect -654 1596 523 1600
rect -654 1507 -644 1596
rect -637 1590 523 1596
rect 844 1590 878 1617
rect 918 1615 924 1617
rect 930 1617 2698 1618
rect 930 1611 2562 1617
rect 930 1608 2377 1611
rect 918 1601 2377 1608
rect 2391 1601 2478 1611
rect 918 1600 2478 1601
rect 918 1596 2343 1600
rect 2391 1598 2419 1600
rect 918 1590 946 1596
rect 950 1594 2343 1596
rect 2366 1596 2418 1598
rect 2425 1596 2478 1600
rect 950 1592 2337 1594
rect 958 1590 998 1592
rect 1012 1590 1026 1592
rect 1046 1590 1086 1592
rect 1092 1590 1152 1592
rect 1160 1590 1240 1592
rect 1319 1590 2337 1592
rect 2366 1590 2425 1596
rect 2444 1590 2478 1596
rect 2519 1608 2562 1611
rect 2519 1590 2577 1608
rect 2619 1594 2670 1617
rect -637 1572 569 1590
rect 774 1589 2354 1590
rect -637 1507 523 1572
rect 808 1554 2354 1589
rect 2366 1587 2577 1590
rect 2636 1588 2670 1594
rect 2371 1583 2577 1587
rect 2619 1583 2670 1588
rect 2377 1574 2491 1583
rect 2493 1582 2670 1583
rect 2377 1572 2487 1574
rect 2377 1554 2407 1572
rect 2410 1555 2428 1572
rect 2444 1555 2478 1572
rect 2493 1556 2528 1582
rect 2531 1578 2565 1582
rect 2568 1562 2670 1582
rect 2497 1555 2528 1556
rect 2541 1555 2670 1562
rect 2689 1608 2724 1617
rect 2759 1616 3075 1628
rect 3132 1616 3166 1628
rect 3182 1616 3219 1681
rect 3274 1662 3781 1711
rect 3833 1696 3847 1734
rect 3813 1673 3847 1696
rect 3833 1662 3847 1673
rect 3867 1696 3901 1734
rect 4031 1716 4065 1734
rect 4020 1715 4108 1716
rect 4258 1715 4292 1745
rect 4347 1757 5386 1807
rect 5454 1792 5465 1803
rect 5477 1792 5488 1803
rect 5454 1757 5488 1792
rect 6688 1792 7194 1968
rect 7222 1870 7280 1876
rect 7222 1839 7234 1870
rect 7222 1836 7268 1839
rect 7222 1830 7280 1836
rect 6688 1768 7219 1792
rect 4347 1732 5524 1757
rect 4334 1721 5524 1732
rect 6051 1722 6197 1744
rect 4334 1716 5532 1721
rect 5597 1716 5681 1721
rect 4334 1715 5681 1716
rect 3867 1673 3935 1696
rect 4020 1681 4166 1715
rect 4226 1687 5681 1715
rect 4226 1681 5524 1687
rect 4020 1678 4129 1681
rect 4032 1674 4066 1678
rect 3867 1662 3901 1673
rect 3274 1661 4075 1662
rect 3274 1656 3801 1661
rect 3821 1656 4075 1661
rect 3274 1640 4075 1656
rect 3274 1628 4016 1640
rect 3274 1616 3821 1628
rect 2759 1608 3821 1616
rect 2689 1599 3821 1608
rect 2689 1555 2723 1599
rect 2760 1594 3821 1599
rect 2760 1564 3799 1594
rect 3801 1573 3821 1594
rect 3867 1618 3901 1628
rect 3916 1618 3982 1623
rect 3867 1594 3982 1618
rect 3867 1590 3975 1594
rect 4067 1590 4075 1640
rect 4258 1608 4292 1681
rect 4334 1608 4360 1681
rect 4226 1590 4292 1608
rect 4314 1590 4360 1608
rect 4364 1650 5524 1681
rect 5663 1674 5681 1678
rect 5698 1674 5751 1722
rect 6051 1686 6052 1722
rect 6084 1686 6109 1705
rect 6120 1687 6197 1722
rect 6276 1737 6312 1747
rect 6688 1739 7330 1768
rect 5786 1675 5838 1686
rect 5874 1685 5926 1686
rect 5973 1685 6050 1686
rect 5797 1674 5827 1675
rect 5873 1674 5927 1685
rect 5961 1674 6050 1685
rect 5651 1662 6050 1674
rect 5533 1654 5571 1657
rect 5533 1653 5579 1654
rect 5663 1653 6050 1662
rect 6051 1655 6109 1686
rect 6139 1669 6244 1687
rect 6276 1669 6510 1737
rect 6596 1734 7330 1739
rect 7411 1734 7426 2119
rect 7445 2085 7480 2119
rect 7445 1734 7479 2085
rect 7778 2023 7848 2140
rect 8130 2121 8164 2140
rect 7960 2072 8018 2078
rect 7960 2038 7972 2072
rect 7960 2032 8018 2038
rect 7591 2017 7649 2023
rect 7591 1983 7603 2017
rect 7591 1977 7649 1983
rect 7761 1916 7848 2023
rect 7681 1880 7706 1885
rect 7672 1855 7693 1880
rect 7761 1863 8058 1916
rect 8149 1863 8164 2121
rect 8183 2087 8218 2121
rect 8498 2087 8533 2121
rect 8183 1863 8217 2087
rect 8499 2068 8533 2087
rect 8329 2019 8387 2025
rect 8329 1985 8341 2019
rect 8329 1979 8387 1985
rect 7672 1846 7684 1855
rect 7761 1847 8427 1863
rect 8518 1847 8533 2068
rect 8552 2034 8587 2068
rect 8552 1847 8586 2034
rect 8698 1966 8756 1972
rect 10329 1968 10369 1986
rect 10456 1968 10471 2262
rect 10490 2228 10525 2262
rect 10490 1968 10524 2228
rect 10636 2160 10694 2166
rect 10636 2126 10648 2160
rect 10636 2120 10694 2126
rect 10806 2119 10840 2173
rect 11228 2155 11263 2173
rect 11192 2140 11263 2155
rect 11543 2140 11578 2174
rect 8698 1932 8710 1966
rect 8698 1926 8756 1932
rect 7591 1817 7649 1823
rect 7591 1783 7603 1817
rect 7638 1783 7653 1817
rect 7672 1784 7687 1846
rect 7761 1810 8766 1847
rect 7591 1777 7649 1783
rect 7672 1741 7706 1784
rect 7761 1777 8796 1810
rect 7778 1757 8796 1777
rect 10102 1792 10608 1968
rect 10636 1870 10694 1876
rect 10636 1839 10648 1870
rect 10636 1836 10682 1839
rect 10636 1830 10694 1836
rect 10102 1768 10633 1792
rect 7778 1741 8938 1757
rect 6596 1705 7194 1734
rect 6139 1655 6265 1669
rect 6288 1665 6322 1667
rect 6376 1665 6410 1667
rect 6464 1665 6487 1667
rect 6051 1654 6265 1655
rect 5533 1650 5591 1653
rect 4364 1634 5591 1650
rect 5681 1652 6050 1653
rect 5681 1634 5768 1652
rect 5973 1651 6041 1652
rect 4364 1632 5768 1634
rect 4364 1624 5777 1632
rect 5858 1624 6050 1651
rect 6098 1640 6150 1651
rect 6109 1624 6139 1640
rect 4364 1608 5785 1624
rect 5858 1622 6139 1624
rect 5854 1617 6139 1622
rect 5805 1608 5839 1614
rect 5854 1608 5892 1617
rect 5926 1614 5964 1617
rect 5967 1615 6041 1617
rect 4364 1594 5892 1608
rect 5908 1608 5964 1614
rect 5973 1608 6041 1615
rect 5908 1594 6041 1608
rect 4364 1592 6041 1594
rect 4372 1590 4398 1592
rect 4399 1590 4412 1592
rect 4427 1590 6041 1592
rect 6069 1590 6084 1617
rect 6103 1610 6139 1617
rect 6173 1633 6208 1650
rect 6173 1632 6453 1633
rect 6173 1616 6489 1632
rect 6596 1616 6630 1705
rect 6633 1665 6664 1705
rect 6688 1635 7194 1705
rect 7445 1706 7460 1734
rect 7606 1715 8938 1741
rect 10102 1734 10744 1768
rect 10825 1734 10840 2119
rect 10859 2085 10894 2119
rect 10859 1734 10893 2085
rect 11192 2023 11262 2140
rect 11544 2121 11578 2140
rect 11374 2072 11432 2078
rect 11374 2038 11386 2072
rect 11374 2032 11432 2038
rect 11005 2017 11063 2023
rect 11005 1983 11017 2017
rect 11005 1977 11063 1983
rect 11175 1916 11262 2023
rect 11095 1880 11120 1885
rect 11086 1855 11107 1880
rect 11175 1863 11472 1916
rect 11563 1863 11578 2121
rect 11597 2087 11632 2121
rect 11912 2087 11947 2121
rect 11597 1863 11631 2087
rect 11913 2068 11947 2087
rect 11743 2019 11801 2025
rect 11743 1985 11755 2019
rect 11743 1979 11801 1985
rect 11086 1846 11098 1855
rect 11005 1817 11063 1823
rect 11005 1783 11017 1817
rect 11052 1783 11067 1817
rect 11086 1784 11101 1846
rect 11175 1810 11841 1863
rect 11932 1810 11947 2068
rect 11966 2034 12001 2068
rect 11966 1810 12000 2034
rect 12112 1966 12170 1972
rect 12112 1932 12124 1966
rect 12112 1926 12170 1932
rect 11005 1777 11063 1783
rect 9112 1721 9165 1722
rect 7541 1706 8938 1715
rect 7445 1688 8938 1706
rect 7237 1635 7351 1688
rect 7409 1645 8938 1688
rect 9094 1687 9165 1721
rect 9095 1686 9165 1687
rect 6688 1616 7351 1635
rect 6103 1608 6150 1610
rect 6173 1608 7351 1616
rect 6103 1599 7351 1608
rect 6103 1590 6137 1599
rect 6174 1596 7351 1599
rect 3867 1577 4111 1590
rect 2760 1563 3444 1564
rect 3498 1563 3585 1564
rect 3638 1563 3799 1564
rect 2760 1555 3813 1563
rect 2410 1554 3813 1555
rect -654 1493 523 1507
rect 569 1539 3813 1554
rect 3867 1560 3901 1577
rect 3920 1560 4111 1577
rect 3867 1555 4111 1560
rect 4222 1589 6137 1590
rect 4222 1584 6041 1589
rect 4222 1580 5827 1584
rect 5839 1580 5965 1584
rect 6050 1583 6084 1589
rect 4222 1564 5839 1580
rect 4222 1555 5768 1564
rect 3867 1551 3917 1555
rect 3920 1554 5768 1555
rect 5805 1558 5839 1564
rect 5805 1554 5822 1558
rect 5824 1554 5839 1558
rect 5858 1558 5965 1580
rect 5858 1554 5892 1558
rect 5915 1554 5965 1558
rect 5982 1554 6084 1583
rect 6103 1554 6137 1589
rect 3867 1539 3901 1551
rect 3920 1547 6150 1554
rect 3920 1539 6174 1547
rect 569 1538 6174 1539
rect 569 1531 782 1538
rect 808 1531 6174 1538
rect 6191 1531 7351 1596
rect 7608 1554 7623 1645
rect 7636 1634 8938 1645
rect 9112 1652 9183 1686
rect 9218 1652 9464 1686
rect 9112 1634 9182 1652
rect 7636 1598 9182 1634
rect 9272 1624 9464 1651
rect 9587 1633 9622 1650
rect 9587 1632 9833 1633
rect 9272 1618 9526 1624
rect 9272 1617 9368 1618
rect 9430 1617 9526 1618
rect 7636 1592 9219 1598
rect 7636 1590 8075 1592
rect 8147 1590 9219 1592
rect 7636 1564 9219 1590
rect 7636 1554 9182 1564
rect 9219 1554 9236 1564
rect 9238 1554 9253 1598
rect 9272 1588 9306 1617
rect 9483 1590 9498 1617
rect 9272 1584 9340 1588
rect 9272 1583 9356 1584
rect 9464 1583 9498 1590
rect 9272 1554 9306 1583
rect 9396 1554 9498 1583
rect 9517 1608 9552 1617
rect 9587 1616 9903 1632
rect 10010 1616 10044 1650
rect 10102 1616 10608 1734
rect 10859 1700 10874 1734
rect 11086 1715 11120 1784
rect 11175 1777 12210 1810
rect 10955 1681 11120 1715
rect 11192 1757 12210 1777
rect 11192 1706 12352 1757
rect 12526 1721 12579 1722
rect 11188 1681 12352 1706
rect 12508 1687 12579 1721
rect 12509 1686 12579 1687
rect 9587 1608 10608 1616
rect 9517 1599 10608 1608
rect 9517 1554 9551 1599
rect 9588 1564 10608 1599
rect 11086 1590 11120 1681
rect 11192 1619 12352 1681
rect 12526 1652 12597 1686
rect 12877 1652 12912 1686
rect 11192 1592 12354 1619
rect 11402 1590 11436 1592
rect 11455 1590 11489 1592
rect 11561 1590 12354 1592
rect 12526 1590 12596 1652
rect 12878 1633 12912 1652
rect 12897 1590 12912 1633
rect 10749 1589 10765 1590
rect 9588 1563 10272 1564
rect 10326 1563 10413 1564
rect 10481 1563 10514 1564
rect 9588 1554 10641 1563
rect 569 1527 793 1531
rect 808 1527 7351 1531
rect 569 1520 7351 1527
rect 7416 1531 9551 1554
rect 9605 1531 10641 1554
rect 7416 1520 10641 1531
rect 569 1493 603 1520
rect -654 1486 725 1493
rect -732 1456 -700 1468
rect -890 1338 -862 1342
rect -970 1301 -936 1338
rect -970 1295 -897 1301
rect -970 1261 -936 1295
rect -868 1288 -862 1338
rect -856 1316 -827 1456
rect -856 1304 -831 1316
rect -785 1300 -700 1456
rect -785 1288 -734 1300
rect -785 1279 -780 1288
rect -766 1284 -734 1288
rect -732 1288 -700 1300
rect -654 1459 615 1486
rect 629 1459 637 1486
rect 667 1484 725 1486
rect 667 1472 751 1484
rect 689 1470 751 1472
rect 678 1459 751 1470
rect -654 1414 523 1459
rect 569 1438 603 1459
rect 691 1440 751 1459
rect 752 1440 779 1512
rect 808 1494 5768 1520
rect 808 1440 2354 1494
rect 2361 1473 5768 1494
rect 5805 1503 5839 1520
rect 5844 1509 5916 1520
rect 6000 1515 6004 1520
rect 6016 1515 6029 1520
rect 5844 1503 5894 1509
rect 5936 1503 5970 1507
rect 5805 1487 5894 1503
rect 5921 1496 5982 1503
rect 5921 1495 5993 1496
rect 5921 1487 5930 1495
rect 5936 1487 5993 1495
rect 6050 1490 6084 1520
rect 5805 1486 5993 1487
rect 5805 1481 5982 1486
rect 2361 1452 5778 1473
rect 2361 1448 2388 1452
rect 2391 1445 5778 1452
rect 5805 1445 5839 1481
rect 555 1433 614 1438
rect 555 1414 615 1433
rect -654 1357 615 1414
rect 691 1426 2354 1440
rect 691 1413 725 1426
rect 672 1396 725 1413
rect -654 1341 527 1357
rect -654 1310 523 1341
rect 555 1338 615 1357
rect 657 1395 725 1396
rect 744 1424 2354 1426
rect 2374 1424 5778 1445
rect 744 1406 2370 1424
rect 744 1398 779 1406
rect 744 1396 778 1398
rect 801 1396 2370 1406
rect 2391 1423 5778 1424
rect 5788 1440 5839 1445
rect 5848 1474 5982 1481
rect 5848 1468 6006 1474
rect 6026 1472 6084 1490
rect 6103 1512 6137 1520
rect 6191 1512 7351 1520
rect 7431 1516 7465 1520
rect 6103 1509 7351 1512
rect 5848 1440 6018 1468
rect 6026 1467 6094 1472
rect 6103 1467 6137 1509
rect 6166 1484 6177 1493
rect 6191 1488 7351 1509
rect 6183 1484 7351 1488
rect 6026 1456 6137 1467
rect 6048 1440 6137 1456
rect 6140 1481 7351 1484
rect 6140 1440 6148 1481
rect 5788 1423 5827 1440
rect 2391 1422 5827 1423
rect 5836 1426 6148 1440
rect 6166 1446 7351 1481
rect 7422 1469 7474 1474
rect 7375 1446 7521 1469
rect 7525 1446 7560 1474
rect 6166 1440 7560 1446
rect 5836 1422 6147 1426
rect 2391 1417 6147 1422
rect 2391 1416 5827 1417
rect 5836 1416 6147 1417
rect 2391 1406 6147 1416
rect 2391 1398 5839 1406
rect 5842 1398 5844 1406
rect 5848 1398 5894 1406
rect 5936 1398 5970 1406
rect 2391 1396 5894 1398
rect 657 1391 740 1395
rect 744 1392 789 1396
rect 801 1395 2371 1396
rect 794 1392 2371 1395
rect 743 1391 2371 1392
rect 657 1379 2371 1391
rect 643 1338 645 1348
rect 549 1310 615 1338
rect 637 1336 645 1338
rect -654 1309 529 1310
rect -766 1279 -751 1284
rect -970 1255 -897 1261
rect -970 1193 -936 1255
rect -785 1247 -751 1279
rect -824 1241 -751 1247
rect -824 1227 -812 1241
rect -785 1227 -751 1241
rect -828 1207 -751 1227
rect -824 1201 -751 1207
rect -785 1193 -751 1201
rect -1023 1164 -751 1193
rect -732 1164 -698 1288
rect -654 1251 534 1309
rect -654 1164 -644 1251
rect -637 1228 534 1251
rect -637 1227 176 1228
rect 190 1227 204 1228
rect -637 1209 170 1227
rect 208 1209 282 1228
rect 322 1209 464 1228
rect -637 1191 464 1209
rect -637 1174 409 1191
rect -637 1164 -30 1174
rect -1193 1148 -1135 1154
rect -1023 1148 -30 1164
rect -1022 1111 -30 1148
rect -1562 1095 -1504 1101
rect -1391 1070 -30 1111
rect -1391 1069 -584 1070
rect -1391 1016 -953 1069
rect -399 1017 -30 1070
rect -28 1053 -13 1174
rect 6 1103 41 1174
rect 6 1053 40 1103
rect 48 1099 74 1174
rect 166 1170 182 1174
rect 196 1170 212 1174
rect 236 1170 245 1174
rect 130 1162 136 1170
rect 166 1168 245 1170
rect 166 1162 182 1168
rect 117 1149 182 1162
rect 196 1153 212 1168
rect 117 1142 198 1149
rect 117 1136 210 1142
rect 117 1115 182 1136
rect 148 1111 182 1115
rect 124 1103 182 1111
rect 195 1103 210 1136
rect 124 1096 210 1103
rect 223 1126 245 1168
rect 266 1145 409 1174
rect 223 1111 251 1126
rect 273 1111 288 1145
rect 301 1111 409 1145
rect 424 1179 464 1191
rect 475 1184 534 1228
rect 549 1224 623 1310
rect 549 1212 557 1224
rect 555 1208 557 1212
rect 569 1191 623 1224
rect 637 1224 649 1336
rect 637 1212 645 1224
rect 643 1208 645 1212
rect 657 1212 689 1379
rect 691 1366 2371 1379
rect 2374 1394 5894 1396
rect 5927 1394 5970 1398
rect 2374 1366 5892 1394
rect 5921 1393 5970 1394
rect 5916 1382 5970 1393
rect 691 1358 2370 1366
rect 2385 1365 5892 1366
rect 5893 1366 5898 1370
rect 5893 1365 5904 1366
rect 691 1356 2354 1358
rect 691 1354 2365 1356
rect 2377 1354 5904 1365
rect 691 1316 5904 1354
rect 5914 1354 5970 1382
rect 5972 1385 6006 1406
rect 6050 1395 6147 1406
rect 6166 1395 7351 1440
rect 7387 1419 7421 1440
rect 7383 1418 7421 1419
rect 7383 1403 7433 1418
rect 6048 1391 6147 1395
rect 6151 1391 7351 1395
rect 7375 1392 7433 1403
rect 5972 1373 6018 1385
rect 6048 1379 7351 1391
rect 6048 1373 6097 1379
rect 6103 1373 7351 1379
rect 5972 1369 6034 1373
rect 6048 1372 7351 1373
rect 6048 1369 6097 1372
rect 5972 1354 6040 1369
rect 5914 1345 6040 1354
rect 6050 1357 6097 1369
rect 6103 1357 7351 1372
rect 5914 1335 6034 1345
rect 5921 1323 6034 1335
rect 691 1226 834 1316
rect 837 1288 877 1316
rect 886 1304 915 1316
rect 886 1288 889 1304
rect 837 1273 889 1288
rect 837 1258 877 1273
rect 837 1226 892 1258
rect 918 1257 1001 1316
rect 691 1212 892 1226
rect 896 1212 898 1252
rect 924 1214 926 1252
rect 930 1226 1001 1257
rect 1007 1282 5904 1316
rect 5915 1317 6034 1323
rect 5915 1288 6040 1317
rect 6050 1295 7351 1357
rect 7356 1332 7362 1378
rect 7371 1338 7433 1392
rect 7460 1380 7463 1391
rect 7475 1380 7521 1440
rect 7371 1301 7421 1338
rect 6050 1291 7358 1295
rect 7371 1291 7417 1301
rect 5915 1284 6046 1288
rect 1007 1279 5898 1282
rect 5915 1279 5973 1284
rect 1007 1263 5973 1279
rect 5988 1275 6046 1284
rect 5982 1263 6046 1275
rect 1007 1260 6046 1263
rect 1007 1245 5973 1260
rect 1007 1242 5961 1245
rect 1007 1235 5898 1242
rect 5911 1235 5961 1242
rect 5982 1241 6046 1260
rect 6050 1241 7364 1291
rect 1007 1227 5904 1235
rect 946 1214 1001 1226
rect 1006 1226 5904 1227
rect 1006 1214 1037 1226
rect 1049 1224 5844 1226
rect 1060 1214 5844 1224
rect 5852 1214 5904 1226
rect 5905 1226 5961 1235
rect 5905 1214 5945 1226
rect 5965 1214 5967 1235
rect 657 1208 677 1212
rect 577 1187 623 1191
rect 569 1184 623 1187
rect 672 1185 677 1208
rect 691 1211 840 1212
rect 691 1207 740 1211
rect 744 1208 789 1211
rect 691 1185 737 1207
rect 744 1185 778 1208
rect 794 1207 828 1211
rect 843 1208 898 1212
rect 801 1197 824 1207
rect 852 1185 898 1208
rect 946 1212 1007 1214
rect 1012 1212 1040 1214
rect 946 1208 995 1212
rect 946 1198 992 1208
rect 475 1179 523 1184
rect 424 1118 469 1179
rect 477 1145 524 1179
rect 527 1145 623 1184
rect 631 1167 831 1185
rect 477 1137 623 1145
rect 477 1130 535 1137
rect 489 1126 492 1130
rect 424 1111 470 1118
rect 527 1113 535 1130
rect 565 1130 623 1137
rect 565 1117 615 1130
rect 223 1103 294 1111
rect 124 1093 174 1096
rect 223 1093 238 1103
rect 244 1093 294 1103
rect 301 1103 316 1111
rect 322 1103 409 1111
rect 301 1099 409 1103
rect 313 1095 316 1099
rect 124 1081 294 1093
rect 124 1075 174 1081
rect 223 1075 238 1081
rect 124 1068 238 1075
rect 244 1075 294 1081
rect 322 1082 409 1099
rect 322 1081 356 1082
rect 322 1075 324 1081
rect 244 1071 325 1075
rect 341 1071 356 1081
rect 375 1071 409 1082
rect 124 1061 174 1068
rect 6 1034 21 1053
rect 182 1035 216 1068
rect 244 1061 294 1071
rect 322 1045 324 1071
rect 341 1054 409 1071
rect 412 1103 470 1111
rect 412 1061 462 1103
rect 565 1099 617 1117
rect 520 1087 521 1099
rect 565 1093 620 1099
rect 566 1087 620 1093
rect 493 1071 520 1087
rect 521 1083 548 1087
rect 521 1071 589 1083
rect 601 1071 625 1087
rect 691 1077 725 1167
rect 744 1143 778 1167
rect 850 1163 898 1185
rect 918 1184 992 1198
rect 1007 1188 1040 1212
rect 1012 1184 1040 1188
rect 1043 1184 5839 1214
rect 5852 1188 5945 1214
rect 5993 1198 5995 1235
rect 5999 1228 7364 1241
rect 5999 1227 7009 1228
rect 7018 1227 7032 1228
rect 5999 1221 7018 1227
rect 7043 1221 7110 1228
rect 7157 1227 7198 1228
rect 5999 1209 7110 1221
rect 7116 1209 7198 1227
rect 5999 1207 7198 1209
rect 5999 1198 6046 1207
rect 5852 1186 5904 1188
rect 5905 1186 5945 1188
rect 5988 1191 6046 1198
rect 5988 1189 6034 1191
rect 6045 1189 6046 1191
rect 6050 1201 6156 1207
rect 6050 1189 6147 1201
rect 917 1173 992 1184
rect 1060 1174 5839 1184
rect 5858 1182 5898 1186
rect 5858 1174 5896 1182
rect 5899 1174 5946 1186
rect 5988 1174 6045 1189
rect 6050 1174 6084 1189
rect 6088 1185 6147 1189
rect 6103 1176 6147 1185
rect 6154 1182 6156 1201
rect 6154 1176 6163 1182
rect 6103 1174 6163 1176
rect 917 1163 980 1173
rect 850 1161 892 1163
rect 850 1158 904 1161
rect 846 1151 904 1158
rect 918 1156 992 1163
rect 918 1151 1040 1156
rect 846 1143 861 1151
rect 868 1143 1040 1151
rect 744 1135 1040 1143
rect 1060 1153 6163 1174
rect 6166 1175 7198 1207
rect 6166 1170 6616 1175
rect 6618 1170 6638 1175
rect 6646 1170 6704 1175
rect 6727 1174 7198 1175
rect 6727 1170 6822 1174
rect 6166 1168 6822 1170
rect 6166 1153 6704 1168
rect 1060 1142 6157 1153
rect 1060 1140 6084 1142
rect 744 1117 992 1135
rect 744 1113 904 1117
rect 744 1086 778 1113
rect 846 1107 904 1113
rect 846 1102 892 1107
rect 795 1094 812 1102
rect 824 1099 892 1102
rect 946 1099 992 1117
rect 824 1094 917 1099
rect 795 1086 917 1094
rect 945 1086 992 1099
rect 999 1128 1014 1132
rect 1026 1128 1053 1132
rect 999 1086 1053 1128
rect 1060 1086 5839 1140
rect 5858 1139 5892 1140
rect 5899 1139 6045 1140
rect 6103 1139 6157 1142
rect 6166 1152 6692 1153
rect 6695 1152 6704 1153
rect 6166 1142 6704 1152
rect 6727 1142 6822 1168
rect 6166 1140 6822 1142
rect 6166 1139 6704 1140
rect 5858 1136 6704 1139
rect 6712 1136 6822 1140
rect 5858 1122 6617 1136
rect 6618 1130 6638 1136
rect 5858 1121 6208 1122
rect 6213 1121 6271 1122
rect 6301 1121 6389 1122
rect 6401 1121 6453 1122
rect 5858 1105 6453 1121
rect 5877 1094 5896 1105
rect 5905 1094 5957 1105
rect 5999 1099 6045 1105
rect 6103 1099 6453 1105
rect 5911 1089 5957 1094
rect 5930 1086 5957 1089
rect 5993 1086 6045 1099
rect 6077 1096 6453 1099
rect 6103 1087 6453 1096
rect 6113 1086 6147 1087
rect 520 1067 521 1071
rect 532 1067 648 1071
rect 341 1045 356 1054
rect 322 1034 356 1045
rect -1391 963 -1322 1016
rect 6 1000 356 1034
rect 375 1033 409 1054
rect 517 1060 648 1067
rect 691 1060 741 1077
rect 744 1066 779 1086
rect 784 1075 6147 1086
rect 6154 1077 6163 1087
rect 6166 1077 6200 1087
rect 795 1071 998 1075
rect 999 1071 1053 1075
rect 795 1066 1053 1071
rect 1060 1071 6147 1075
rect 6150 1071 6200 1077
rect 744 1060 1037 1066
rect 1060 1064 5852 1071
rect 5893 1068 6200 1071
rect 5893 1064 6147 1068
rect 1060 1060 6147 1064
rect 6150 1060 6200 1068
rect 6213 1060 6259 1087
rect 6308 1083 6447 1087
rect 6307 1071 6447 1083
rect 6467 1071 6469 1122
rect 6472 1113 6527 1122
rect 6302 1060 6447 1071
rect 517 1049 6447 1060
rect 517 1035 583 1049
rect 601 1035 631 1049
rect 691 1045 6200 1049
rect 691 1043 2606 1045
rect 707 1042 2606 1043
rect 2632 1042 2715 1045
rect 2799 1043 6200 1045
rect 2799 1042 6184 1043
rect 707 1041 6184 1042
rect 6213 1041 6359 1049
rect 6389 1041 6447 1049
rect 6472 1043 6516 1113
rect 6532 1111 6617 1122
rect 6532 1099 6616 1111
rect 6535 1081 6616 1099
rect 6535 1068 6604 1081
rect 6608 1071 6610 1081
rect 6636 1071 6638 1130
rect 6646 1120 6822 1136
rect 6658 1111 6822 1120
rect 6646 1102 6822 1111
rect 6646 1099 6704 1102
rect 6712 1099 6822 1102
rect 6646 1096 6822 1099
rect 6646 1081 6704 1096
rect 6734 1081 6822 1096
rect 6658 1068 6692 1081
rect 6740 1071 6780 1081
rect 6698 1068 6780 1071
rect 6788 1068 6822 1081
rect 6472 1041 6501 1043
rect 6558 1041 6792 1068
rect 517 1033 691 1035
rect 375 1029 423 1033
rect 483 1029 691 1033
rect 375 999 691 1029
rect 707 1026 2826 1041
rect 2840 1026 6184 1041
rect 6271 1035 6301 1041
rect 6308 1035 6359 1041
rect 6401 1037 6435 1041
rect 6200 1033 6359 1035
rect 6472 1034 6482 1041
rect 6568 1034 6734 1041
rect 6807 1034 6822 1068
rect 6841 1168 6944 1174
rect 6955 1168 6972 1174
rect 6841 1115 6948 1168
rect 6949 1164 6976 1168
rect 7001 1164 7009 1174
rect 7031 1164 7130 1174
rect 6955 1160 6976 1164
rect 6958 1155 6976 1160
rect 6984 1155 7010 1164
rect 6958 1141 7010 1155
rect 6841 1034 6885 1115
rect 6501 1033 6516 1034
rect 6200 1026 6516 1033
rect 375 987 409 999
rect 437 991 489 999
rect 437 987 505 991
rect 168 980 322 987
rect 356 981 538 987
rect 356 980 691 981
rect 6 970 691 980
rect 710 970 725 1026
rect 744 1024 917 1026
rect 744 1022 921 1024
rect 744 1020 936 1022
rect 727 1018 936 1020
rect 952 1018 2606 1026
rect 727 998 2606 1018
rect 2621 1017 2726 1026
rect 2840 1017 4069 1026
rect 4095 1022 5978 1026
rect 4095 1018 5989 1022
rect 727 992 795 998
rect 849 996 2606 998
rect 849 992 895 996
rect 727 988 779 992
rect 852 988 895 992
rect 727 986 795 988
rect 744 970 812 986
rect 6 966 812 970
rect 6 946 41 966
rect 94 957 124 966
rect 83 946 135 957
rect 168 956 340 966
rect -363 893 -328 927
rect -732 840 -697 874
rect -955 719 -897 725
rect -1101 696 -1067 714
rect -1470 626 -1435 660
rect -1693 505 -1635 511
rect -1693 471 -1681 505
rect -1693 465 -1635 471
rect -1693 305 -1635 311
rect -1693 271 -1681 305
rect -1693 265 -1635 271
rect -1504 188 -1489 607
rect -1470 256 -1436 626
rect -1324 558 -1266 564
rect -1324 524 -1312 558
rect -1324 518 -1266 524
rect -1324 358 -1266 364
rect -1324 324 -1312 358
rect -1324 318 -1266 324
rect -1137 309 -1067 696
rect -955 685 -943 719
rect -955 679 -897 685
rect -955 411 -897 417
rect -955 377 -943 411
rect -955 371 -897 377
rect -1137 275 -1066 309
rect -766 294 -751 821
rect -732 362 -698 840
rect -586 772 -528 778
rect -586 738 -574 772
rect -586 732 -528 738
rect -586 464 -528 470
rect -586 430 -574 464
rect -586 424 -528 430
rect -732 328 -697 362
rect -397 347 -382 874
rect -363 415 -329 893
rect -217 825 -159 831
rect -217 791 -205 825
rect -217 785 -159 791
rect -140 757 -131 768
rect -132 564 -121 568
rect -104 536 -93 568
rect -217 517 -159 523
rect -217 483 -205 517
rect -217 477 -159 483
rect -363 381 -328 415
rect -28 400 -13 927
rect 6 898 40 946
rect 168 919 324 956
rect 341 954 812 966
rect 849 984 895 988
rect 902 984 936 988
rect 952 984 2606 996
rect 849 983 2606 984
rect 849 954 883 983
rect 886 980 2606 983
rect 886 958 995 980
rect 1060 968 2606 980
rect 2840 979 4068 1017
rect 4095 998 6005 1018
rect 886 954 921 958
rect 923 954 995 958
rect 1049 954 2606 968
rect 2621 954 2726 963
rect 2731 954 2823 979
rect 2840 965 2911 979
rect 2945 970 4068 979
rect 4112 970 4122 998
rect 4131 986 4209 998
rect 4263 996 6005 998
rect 4131 970 4146 986
rect 4163 971 4233 986
rect 4163 970 4209 971
rect 2945 965 4209 970
rect 2840 962 2927 965
rect 2945 963 4221 965
rect 4263 963 5844 996
rect 2945 962 5844 963
rect 341 953 2826 954
rect 2840 953 2910 962
rect 341 920 2910 953
rect 341 919 567 920
rect 236 914 237 919
rect 248 914 282 919
rect 236 912 282 914
rect 124 909 166 912
rect 236 899 251 912
rect 322 909 370 919
rect 375 909 409 919
rect 322 907 409 909
rect 275 899 409 907
rect 424 913 458 919
rect 424 904 443 913
rect 470 904 567 919
rect 579 909 2910 920
rect 583 904 2910 909
rect 424 902 567 904
rect 579 902 2910 904
rect 424 899 605 902
rect 6 869 148 898
rect 152 881 166 884
rect 236 873 409 899
rect 195 869 210 873
rect 223 869 409 873
rect 412 897 605 899
rect 412 869 538 897
rect 6 868 166 869
rect 195 868 214 869
rect 6 838 214 868
rect 6 834 166 838
rect 6 830 170 834
rect 6 801 41 830
rect 48 823 74 830
rect 48 801 82 823
rect 86 804 96 825
rect 130 810 182 830
rect 196 828 214 838
rect 223 855 251 869
rect 223 823 266 855
rect 275 823 282 869
rect 223 819 282 823
rect 313 835 370 869
rect 313 819 316 835
rect 322 823 370 835
rect 375 823 409 869
rect 423 850 538 869
rect 223 810 292 819
rect 86 801 88 804
rect 136 801 182 810
rect 6 740 182 801
rect 202 796 204 797
rect 197 785 212 796
rect 236 789 292 810
rect 224 785 292 789
rect 6 685 41 740
rect 48 685 82 740
rect 86 704 88 740
rect 114 704 116 740
rect 120 686 170 740
rect 174 704 176 740
rect 202 704 204 785
rect 208 751 292 785
rect 322 801 409 823
rect 424 801 538 850
rect 543 887 598 897
rect 543 881 595 887
rect 637 882 683 902
rect 689 899 2910 902
rect 2927 933 2961 962
rect 3047 954 5844 962
rect 5864 992 5898 996
rect 5864 988 5865 992
rect 5910 988 5978 996
rect 5864 954 5898 988
rect 5910 984 5989 988
rect 5910 962 6005 984
rect 5910 958 5989 962
rect 5910 954 5978 958
rect 6046 954 6047 1026
rect 6113 979 6147 1026
rect 6166 999 6516 1026
rect 6535 1015 6885 1034
rect 6892 1087 6948 1115
rect 6952 1138 7010 1141
rect 7046 1155 7130 1164
rect 7046 1141 7112 1155
rect 7157 1141 7198 1174
rect 7210 1202 7364 1228
rect 7377 1279 7417 1291
rect 7429 1290 7433 1338
rect 7471 1319 7521 1380
rect 7437 1291 7446 1295
rect 7437 1290 7452 1291
rect 7429 1289 7452 1290
rect 7465 1289 7521 1319
rect 7429 1279 7458 1289
rect 7377 1242 7458 1279
rect 7459 1258 7463 1289
rect 7465 1258 7517 1289
rect 7459 1242 7517 1258
rect 7377 1224 7517 1242
rect 7377 1212 7392 1224
rect 7383 1208 7392 1212
rect 7412 1212 7517 1224
rect 7412 1208 7480 1212
rect 7492 1208 7505 1212
rect 7210 1141 7307 1202
rect 7046 1139 7122 1141
rect 6952 1133 6998 1138
rect 7001 1133 7010 1138
rect 6952 1121 7017 1133
rect 7022 1121 7045 1123
rect 6952 1103 7033 1121
rect 7042 1117 7045 1121
rect 7042 1103 7049 1117
rect 7064 1103 7122 1139
rect 7152 1140 7307 1141
rect 7312 1184 7364 1202
rect 7412 1192 7458 1208
rect 7429 1184 7458 1192
rect 7312 1140 7361 1184
rect 7365 1140 7458 1184
rect 7477 1140 7480 1202
rect 7526 1140 7560 1440
rect 7589 1421 7623 1520
rect 7579 1414 7614 1421
rect 7636 1418 9182 1520
rect 7629 1414 9182 1418
rect 7579 1392 9182 1414
rect 7571 1316 9182 1392
rect 9219 1509 9418 1520
rect 9430 1515 9443 1520
rect 9219 1503 9253 1509
rect 9272 1507 9306 1509
rect 9262 1503 9306 1507
rect 9350 1503 9384 1507
rect 9219 1495 9308 1503
rect 9338 1495 9396 1503
rect 9219 1392 9253 1495
rect 9256 1481 9306 1495
rect 9344 1487 9396 1495
rect 9464 1490 9498 1520
rect 9440 1487 9498 1490
rect 9344 1481 9432 1487
rect 9256 1392 9258 1417
rect 9262 1392 9306 1481
rect 9312 1463 9330 1475
rect 9350 1473 9432 1481
rect 9338 1468 9432 1473
rect 9440 1468 9512 1487
rect 9338 1467 9418 1468
rect 9440 1467 9508 1468
rect 9517 1467 9551 1520
rect 9338 1463 9432 1467
rect 9308 1437 9432 1463
rect 9440 1456 9551 1467
rect 9462 1437 9551 1456
rect 9308 1429 9420 1437
rect 9338 1419 9384 1429
rect 7571 1266 7717 1316
rect 7721 1311 7832 1316
rect 7834 1311 7945 1316
rect 7721 1296 7945 1311
rect 7958 1296 9182 1316
rect 7721 1295 9182 1296
rect 7721 1285 7771 1295
rect 7777 1266 9182 1295
rect 7571 1263 9182 1266
rect 7571 1261 8334 1263
rect 8374 1261 9182 1263
rect 7571 1252 7835 1261
rect 7843 1255 7846 1261
rect 7571 1238 7727 1252
rect 7777 1245 7835 1252
rect 7871 1247 7874 1261
rect 7877 1247 8334 1261
rect 7777 1238 7823 1245
rect 7571 1224 7739 1238
rect 7775 1224 7823 1238
rect 7571 1212 7623 1224
rect 7152 1115 7298 1140
rect 7152 1111 7254 1115
rect 7124 1103 7254 1111
rect 7273 1106 7298 1115
rect 7312 1111 7560 1140
rect 7359 1106 7560 1111
rect 7290 1103 7292 1106
rect 6964 1099 7049 1103
rect 7076 1099 7110 1103
rect 7124 1099 7198 1103
rect 6966 1087 7049 1099
rect 7124 1087 7191 1099
rect 7210 1087 7245 1103
rect 7400 1098 7459 1106
rect 7328 1087 7459 1098
rect 6892 1077 7244 1087
rect 6892 1065 7158 1077
rect 7191 1065 7244 1077
rect 6892 1064 6952 1065
rect 6960 1064 7158 1065
rect 6892 1053 7163 1064
rect 6892 1015 6916 1053
rect 6920 1015 6944 1053
rect 6996 1051 7073 1053
rect 6994 1049 7073 1051
rect 7010 1035 7044 1049
rect 7157 1045 7163 1053
rect 7176 1045 7191 1053
rect 6994 1019 7060 1035
rect 7157 1015 7191 1045
rect 6535 1004 7071 1015
rect 7080 1007 7191 1015
rect 7091 1004 7191 1007
rect 6535 1001 7060 1004
rect 6535 1000 6952 1001
rect 6166 981 6200 999
rect 6482 981 6516 999
rect 6841 992 6952 1000
rect 6841 981 6963 992
rect 6994 984 7060 1001
rect 7102 992 7191 1004
rect 7091 981 7191 992
rect 6166 980 6516 981
rect 6166 979 6482 980
rect 6501 979 6516 980
rect 6113 954 6516 979
rect 3047 949 6516 954
rect 3041 947 6516 949
rect 3041 939 6358 947
rect 3035 933 6358 939
rect 6359 933 6516 947
rect 6535 941 6885 980
rect 7210 962 7244 1065
rect 7328 1026 7348 1087
rect 7356 1064 7414 1070
rect 7356 1053 7418 1064
rect 7356 1045 7376 1053
rect 7352 1030 7376 1045
rect 7352 1024 7414 1030
rect 7352 1014 7376 1024
rect 7429 1014 7459 1087
rect 7477 1085 7480 1106
rect 7526 1066 7560 1106
rect 7579 1106 7623 1212
rect 7642 1216 7739 1224
rect 7642 1212 7727 1216
rect 7732 1212 7739 1216
rect 7642 1208 7739 1212
rect 7642 1193 7676 1208
rect 7681 1193 7739 1208
rect 7781 1212 7823 1224
rect 7827 1212 7835 1245
rect 7865 1243 8334 1247
rect 8372 1243 9182 1261
rect 7865 1228 9182 1243
rect 9190 1228 9216 1370
rect 9219 1366 9306 1392
rect 9219 1228 9253 1366
rect 9256 1323 9258 1366
rect 9262 1354 9312 1366
rect 9262 1323 9306 1354
rect 9308 1323 9312 1354
rect 9316 1323 9318 1366
rect 9344 1323 9346 1394
rect 9350 1335 9384 1419
rect 9352 1323 9384 1335
rect 9386 1357 9420 1429
rect 9464 1395 9551 1437
rect 9462 1391 9551 1395
rect 9588 1510 10641 1520
rect 10748 1510 10765 1589
rect 11050 1554 12596 1590
rect 12720 1584 12754 1588
rect 12878 1554 12912 1590
rect 12931 1608 12966 1633
rect 12931 1599 13155 1608
rect 13246 1599 13281 1633
rect 12931 1554 12965 1599
rect 13247 1580 13281 1599
rect 10830 1531 12965 1554
rect 13051 1531 13123 1554
rect 10830 1520 13123 1531
rect 9588 1446 10765 1510
rect 10939 1446 10974 1474
rect 9588 1440 10974 1446
rect 9430 1369 9448 1373
rect 9462 1369 9570 1391
rect 9430 1357 9454 1369
rect 9386 1323 9454 1357
rect 9262 1319 9324 1323
rect 9352 1319 9454 1323
rect 9272 1297 9324 1319
rect 9272 1292 9306 1297
rect 9308 1292 9324 1297
rect 9272 1228 9324 1292
rect 9374 1288 9454 1319
rect 9464 1300 9570 1369
rect 9386 1285 9460 1288
rect 9386 1284 9390 1285
rect 9340 1242 9346 1276
rect 9352 1263 9356 1276
rect 9414 1275 9460 1285
rect 9396 1263 9460 1275
rect 9352 1260 9460 1263
rect 9352 1250 9356 1260
rect 9396 1241 9460 1260
rect 9464 1275 9498 1300
rect 9502 1275 9570 1300
rect 9464 1241 9570 1275
rect 9414 1228 9570 1241
rect 7865 1212 9253 1228
rect 7781 1208 7827 1212
rect 7877 1208 9253 1212
rect 7781 1193 7815 1208
rect 7820 1193 7827 1208
rect 7895 1198 9253 1208
rect 7895 1193 8716 1198
rect 8736 1194 9253 1198
rect 7642 1167 7659 1193
rect 7676 1186 8716 1193
rect 7676 1174 8703 1186
rect 8708 1182 8716 1186
rect 8739 1186 9253 1194
rect 9266 1186 9324 1228
rect 9402 1207 9570 1228
rect 9402 1189 9460 1207
rect 9464 1201 9570 1207
rect 9588 1295 10765 1440
rect 10797 1392 10850 1406
rect 10770 1332 10776 1378
rect 10785 1338 10850 1392
rect 10906 1392 10919 1396
rect 10785 1322 10832 1338
rect 9588 1291 10772 1295
rect 10785 1291 10831 1322
rect 10885 1319 10894 1329
rect 10879 1317 10894 1319
rect 10851 1291 10860 1295
rect 9588 1228 10778 1291
rect 9588 1227 10423 1228
rect 10432 1227 10446 1228
rect 9588 1209 10412 1227
rect 10415 1209 10423 1227
rect 10457 1209 10524 1228
rect 10571 1209 10612 1228
rect 9464 1189 9548 1201
rect 8739 1182 9182 1186
rect 9190 1182 9253 1186
rect 9272 1182 9287 1186
rect 9306 1182 9312 1186
rect 9414 1185 9448 1189
rect 7681 1167 8703 1174
rect 7642 1159 8703 1167
rect 7693 1133 7739 1159
rect 7681 1124 7739 1133
rect 7745 1156 7761 1159
rect 7790 1156 7827 1159
rect 7745 1124 7773 1156
rect 7775 1132 7827 1156
rect 7895 1150 8703 1159
rect 8711 1154 8716 1182
rect 8743 1174 9182 1182
rect 9219 1174 9287 1182
rect 9464 1174 9498 1189
rect 9502 1185 9551 1189
rect 9517 1174 9551 1185
rect 8743 1157 9551 1174
rect 7775 1125 7881 1132
rect 7775 1124 7849 1125
rect 7579 1066 7613 1106
rect 7623 1086 7657 1102
rect 7659 1086 7677 1102
rect 7623 1072 7677 1086
rect 7623 1066 7651 1072
rect 7655 1066 7677 1072
rect 7681 1087 7727 1124
rect 7732 1087 7739 1124
rect 7790 1116 7849 1124
rect 7861 1116 7881 1125
rect 7681 1066 7739 1087
rect 7793 1082 7881 1116
rect 7793 1072 7849 1082
rect 7509 1057 7739 1066
rect 7509 1011 7721 1057
rect 7745 1038 7773 1072
rect 7775 1066 7849 1072
rect 7861 1066 7881 1082
rect 7895 1123 8028 1150
rect 8094 1124 8106 1150
rect 8137 1124 8152 1150
rect 7775 1058 7827 1066
rect 7793 1054 7815 1058
rect 7895 1048 7982 1123
rect 8094 1118 8152 1124
rect 8165 1096 8180 1150
rect 8066 1090 8180 1096
rect 8283 1076 8298 1150
rect 8264 1063 8298 1076
rect 7787 1038 7982 1048
rect 7745 1030 7982 1038
rect 8235 1045 8298 1063
rect 8317 1135 8703 1150
rect 8754 1146 8784 1157
rect 8798 1154 8804 1157
rect 8317 1116 8714 1135
rect 8317 1101 8742 1116
rect 8317 1095 8711 1101
rect 8317 1077 8703 1095
rect 8712 1085 8742 1101
rect 8317 1067 8711 1077
rect 8317 1065 8703 1067
rect 7725 1011 7745 1017
rect 7787 1011 7982 1030
rect 7509 998 7749 1011
rect 7755 1006 7982 1011
rect 7336 996 7398 998
rect 7272 991 7317 996
rect 7267 987 7283 991
rect 7254 970 7366 987
rect 7545 986 7614 998
rect 7687 997 7749 998
rect 7751 997 7982 1006
rect 7545 970 7560 986
rect 7577 971 7647 986
rect 7687 983 7982 997
rect 8050 1008 8150 1034
rect 8235 1029 8313 1045
rect 8317 1029 8351 1065
rect 8459 1055 8472 1065
rect 8498 1055 8703 1065
rect 8485 1044 8703 1055
rect 8850 1044 8884 1157
rect 8903 1086 8937 1157
rect 9148 1148 9551 1157
rect 9588 1175 10612 1209
rect 9588 1152 10027 1175
rect 9148 1140 9189 1148
rect 9236 1142 9551 1148
rect 9236 1141 9498 1142
rect 9244 1140 9498 1141
rect 8939 1124 8975 1140
rect 9148 1138 9153 1140
rect 8939 1120 8989 1124
rect 8939 1106 9005 1120
rect 9219 1099 9230 1110
rect 9238 1099 9253 1140
rect 9272 1139 9306 1140
rect 9517 1139 9551 1142
rect 9272 1108 9575 1139
rect 9602 1122 10027 1152
rect 10028 1170 10030 1175
rect 10032 1170 10052 1175
rect 10060 1170 10106 1175
rect 10155 1174 10612 1175
rect 10028 1136 10106 1170
rect 9602 1121 9622 1122
rect 9627 1121 9676 1122
rect 9727 1121 9761 1122
rect 9833 1121 9867 1122
rect 9272 1106 9553 1108
rect 9272 1105 9307 1106
rect 9339 1105 9391 1106
rect 9449 1105 9553 1106
rect 9219 1086 9253 1099
rect 9517 1098 9553 1105
rect 9517 1087 9528 1098
rect 9613 1087 9867 1121
rect 9886 1087 9920 1122
rect 8903 1072 9039 1086
rect 9049 1075 9101 1086
rect 9137 1075 9253 1086
rect 8903 1064 8938 1072
rect 9060 1064 9090 1075
rect 9148 1069 9253 1075
rect 9236 1064 9253 1069
rect 8903 1052 9289 1064
rect 8934 1044 9289 1052
rect 9481 1051 9543 1065
rect 9727 1053 9761 1087
rect 8431 1033 8464 1037
rect 8419 1031 8464 1033
rect 8050 996 8153 1008
rect 8062 992 8096 996
rect 8264 995 8351 1029
rect 8364 997 8464 1031
rect 8485 1021 9289 1044
rect 9886 1041 9915 1087
rect 9972 1068 9974 1122
rect 9984 1102 10024 1122
rect 10028 1120 10030 1136
rect 10032 1130 10052 1136
rect 10060 1120 10106 1136
rect 9984 1068 10018 1102
rect 10072 1068 10106 1120
rect 10160 1068 10194 1174
rect 10202 1068 10236 1174
rect 9972 1041 10206 1068
rect 10019 1034 10071 1041
rect 10107 1034 10159 1041
rect 10221 1034 10236 1068
rect 10255 1103 10323 1174
rect 10415 1164 10423 1174
rect 10398 1155 10424 1164
rect 10378 1138 10424 1155
rect 10378 1133 10412 1138
rect 10415 1133 10424 1138
rect 10478 1151 10494 1164
rect 10378 1117 10431 1133
rect 10456 1117 10459 1123
rect 10378 1115 10447 1117
rect 10382 1103 10447 1115
rect 10456 1103 10463 1117
rect 10478 1103 10497 1151
rect 10255 1034 10289 1103
rect 10290 1099 10323 1103
rect 10397 1075 10463 1103
rect 10490 1099 10497 1103
rect 10571 1103 10612 1174
rect 10397 1067 10487 1075
rect 10410 1051 10487 1067
rect 10408 1049 10487 1051
rect 10424 1035 10458 1049
rect 10571 1045 10577 1103
rect 10590 1099 10612 1103
rect 10590 1045 10605 1099
rect 7577 970 7614 971
rect 7254 962 7614 970
rect 2927 899 2967 933
rect 689 894 2967 899
rect 689 882 812 894
rect 824 891 895 894
rect 637 881 649 882
rect 543 867 589 881
rect 643 878 645 881
rect 637 876 645 878
rect 637 867 649 876
rect 657 867 812 882
rect 846 867 917 891
rect 543 858 601 867
rect 543 850 611 858
rect 543 813 623 850
rect 631 837 689 867
rect 691 837 725 867
rect 726 837 737 867
rect 744 837 812 867
rect 837 863 917 867
rect 918 863 1014 894
rect 837 837 1014 863
rect 637 824 649 837
rect 657 830 824 837
rect 637 813 645 824
rect 657 823 779 830
rect 807 823 824 830
rect 846 834 1014 837
rect 1049 846 2967 894
rect 2987 880 2995 915
rect 3007 911 3021 915
rect 3035 911 6516 933
rect 6520 929 6885 941
rect 3007 910 3027 911
rect 3035 910 6156 911
rect 3007 906 6156 910
rect 3007 905 5852 906
rect 3007 899 5863 905
rect 2996 894 5863 899
rect 5893 894 6156 906
rect 2996 892 5831 894
rect 2996 880 3891 892
rect 2987 860 3891 880
rect 2987 846 3873 860
rect 3930 846 3964 892
rect 3969 864 5831 892
rect 5905 878 5957 894
rect 3969 846 5827 864
rect 1049 834 5827 846
rect 5911 863 5957 878
rect 5961 863 5979 875
rect 5988 873 6067 894
rect 5987 863 6067 873
rect 6088 867 6156 894
rect 5911 848 6067 863
rect 6076 848 6156 867
rect 5911 837 6046 848
rect 6076 837 6147 848
rect 5911 836 6147 837
rect 846 829 1037 834
rect 846 823 904 829
rect 657 822 904 823
rect 657 813 677 822
rect 680 813 683 822
rect 689 819 904 822
rect 946 820 1037 829
rect 1049 820 5831 834
rect 5911 833 6046 836
rect 689 818 895 819
rect 689 817 824 818
rect 837 817 894 818
rect 689 813 778 817
rect 543 812 778 813
rect 551 808 623 812
rect 643 808 645 812
rect 657 808 677 812
rect 322 789 470 801
rect 208 740 270 751
rect 322 740 370 789
rect 375 740 470 789
rect 208 739 470 740
rect 208 704 264 739
rect 270 711 292 739
rect 322 719 324 739
rect 341 735 370 739
rect 341 719 356 735
rect 322 711 356 719
rect 375 711 443 739
rect 120 685 181 686
rect 208 685 258 704
rect 270 686 443 711
rect 447 704 470 739
rect 475 704 534 801
rect 481 693 534 704
rect 551 693 557 808
rect 577 805 623 808
rect 558 789 565 800
rect 569 712 623 805
rect 691 791 725 812
rect 672 773 725 791
rect 727 790 737 812
rect 730 773 737 790
rect 672 769 740 773
rect 744 769 778 812
rect 807 792 824 817
rect 672 757 778 769
rect 691 712 778 757
rect 794 730 812 773
rect 824 769 828 773
rect 824 757 834 769
rect 820 745 834 757
rect 820 730 840 745
rect 270 685 453 686
rect 6 652 270 685
rect 288 652 461 685
rect 6 651 461 652
rect 481 682 523 693
rect 527 682 534 693
rect 569 686 778 712
rect 782 712 840 730
rect 846 730 894 817
rect 946 800 5831 820
rect 5899 829 6046 833
rect 5899 818 5957 829
rect 5987 819 6046 829
rect 5879 817 5994 818
rect 896 769 940 794
rect 946 790 992 800
rect 1007 790 1037 800
rect 1049 796 5831 800
rect 1060 794 5831 796
rect 946 774 1037 790
rect 946 769 1012 774
rect 1040 770 5831 794
rect 5877 790 5879 817
rect 5899 790 5957 817
rect 5879 789 5966 790
rect 5899 788 5957 789
rect 1018 769 5831 770
rect 896 762 898 769
rect 930 766 992 769
rect 1012 766 1052 769
rect 924 765 980 766
rect 919 762 980 765
rect 984 762 992 766
rect 1006 762 1058 766
rect 1060 762 5831 769
rect 898 741 980 762
rect 992 759 5831 762
rect 992 741 1012 759
rect 1026 746 5831 759
rect 5839 746 5865 770
rect 5899 769 5945 788
rect 5965 771 5966 789
rect 5993 771 5994 817
rect 5997 817 6046 819
rect 6067 817 6147 836
rect 5997 769 6045 817
rect 6067 810 6076 817
rect 6113 813 6147 817
rect 6095 791 6147 813
rect 6154 808 6156 848
rect 6166 909 6259 911
rect 6166 897 6200 909
rect 6213 897 6259 909
rect 6166 881 6259 897
rect 6301 909 6396 911
rect 6301 897 6398 909
rect 6301 896 6359 897
rect 6308 881 6359 896
rect 6367 891 6370 897
rect 6166 791 6200 881
rect 6213 878 6259 881
rect 6213 867 6265 878
rect 6313 867 6356 881
rect 6395 867 6398 897
rect 6401 872 6408 911
rect 6432 903 6516 911
rect 6535 927 6885 929
rect 7042 927 7144 941
rect 7210 928 7614 962
rect 7687 969 7717 983
rect 7721 980 7982 983
rect 8053 980 8087 984
rect 7721 977 7821 980
rect 7721 969 7723 977
rect 7725 971 7821 977
rect 7777 969 7821 971
rect 7687 965 7821 969
rect 7895 968 7982 980
rect 8047 968 8099 980
rect 7687 961 7787 965
rect 7789 961 7821 965
rect 7687 943 7821 961
rect 7254 927 7613 928
rect 6535 911 6860 927
rect 6535 907 6569 911
rect 6570 907 6603 911
rect 6698 909 6724 911
rect 6608 907 6610 909
rect 6535 903 6610 907
rect 6432 899 6612 903
rect 6422 872 6447 899
rect 6401 867 6447 872
rect 6213 850 6271 867
rect 6280 850 6359 867
rect 6368 850 6447 867
rect 6213 837 6447 850
rect 6213 822 6265 837
rect 6268 822 6447 837
rect 6213 821 6447 822
rect 6221 817 6435 821
rect 6095 779 6163 791
rect 6166 779 6219 791
rect 6063 769 6067 773
rect 6079 769 6097 773
rect 6113 769 6147 779
rect 6163 769 6219 779
rect 5899 766 5961 769
rect 5877 746 5879 762
rect 1026 741 5885 746
rect 930 735 980 741
rect 896 730 898 734
rect 846 723 904 730
rect 924 723 926 734
rect 930 730 964 735
rect 930 723 976 730
rect 984 723 986 734
rect 1012 730 1014 734
rect 1026 730 1052 741
rect 1060 730 5885 741
rect 844 712 904 723
rect 782 710 904 712
rect 918 720 976 723
rect 918 719 980 720
rect 918 710 976 719
rect 782 700 976 710
rect 1006 716 5885 730
rect 5905 723 5907 762
rect 5911 735 5961 766
rect 6025 761 6033 769
rect 6025 746 6045 761
rect 5915 723 5961 735
rect 5965 723 5967 743
rect 5987 723 6045 746
rect 6051 746 6099 769
rect 5915 716 5973 723
rect 1006 700 5831 716
rect 794 686 964 700
rect 1012 695 1014 700
rect 1018 686 1052 700
rect 1060 686 5831 700
rect 6 468 41 651
rect 48 468 74 651
rect 86 604 88 645
rect 114 629 116 645
rect 120 629 170 651
rect 114 617 124 629
rect 136 617 170 629
rect 174 617 176 645
rect 202 617 204 645
rect 208 629 258 651
rect 224 617 258 629
rect 86 589 96 604
rect 136 570 182 617
rect 198 576 258 617
rect 190 570 258 576
rect 136 536 258 570
rect 136 520 182 536
rect 190 530 210 536
rect 212 520 214 536
rect 136 468 170 520
rect 218 509 258 536
rect 218 502 264 509
rect 224 468 264 502
rect 270 468 292 481
rect 322 468 324 651
rect 6 441 292 468
rect 341 453 356 651
rect 375 583 443 651
rect 375 521 410 583
rect 481 521 515 682
rect 569 670 5831 686
rect 557 639 565 670
rect 567 664 5831 670
rect 567 663 2237 664
rect 567 651 1868 663
rect 1877 659 1945 663
rect 567 639 614 651
rect 517 623 527 639
rect 557 623 614 639
rect 517 589 614 623
rect 691 601 778 651
rect 794 628 828 651
rect 902 642 977 651
rect 918 628 952 642
rect 1018 628 1052 651
rect 1060 642 1868 651
rect 1883 654 1945 659
rect 1883 642 1917 654
rect 1921 642 1945 654
rect 1060 628 1870 642
rect 1871 641 1945 642
rect 1871 628 1948 641
rect 517 573 527 589
rect 557 573 603 589
rect 569 521 603 573
rect 691 585 740 601
rect 691 574 725 585
rect 744 574 778 601
rect 782 589 840 628
rect 794 585 828 589
rect 918 586 976 628
rect 1006 610 1948 628
rect 1006 598 1546 610
rect 1006 586 1499 598
rect 1531 586 1546 598
rect 930 582 964 586
rect 1018 582 1052 586
rect 1060 574 1499 586
rect 691 571 862 574
rect 896 571 1499 574
rect 691 557 1499 571
rect 1656 568 1661 610
rect 1675 568 1690 610
rect 691 551 1094 557
rect 691 542 793 551
rect 691 521 725 542
rect 744 540 793 542
rect 851 548 1094 551
rect 851 541 1006 548
rect 851 540 903 541
rect 1053 540 1094 548
rect 1340 546 1374 557
rect 1656 546 1690 568
rect 375 487 615 521
rect 629 487 637 521
rect 678 510 725 521
rect 1340 535 1411 546
rect 1447 535 1560 546
rect 1340 523 1400 535
rect 1458 523 1560 535
rect 1574 530 1690 546
rect 1602 523 1690 530
rect 1340 512 1411 523
rect 1458 516 1571 523
rect 1519 512 1571 516
rect 1591 512 1690 523
rect 689 498 725 510
rect 714 487 725 498
rect 1709 493 1743 610
rect 1769 557 1803 610
rect 1851 601 1854 610
rect 1867 595 1948 610
rect 1955 608 2017 663
rect 1851 583 1948 595
rect 1971 594 2017 608
rect 1871 582 1948 583
rect 1986 582 2017 594
rect 2025 640 2226 663
rect 2238 659 2320 664
rect 2325 659 2374 664
rect 2238 647 2314 659
rect 2238 640 2277 647
rect 2280 640 2314 647
rect 2331 640 2374 659
rect 2377 640 2386 664
rect 2394 663 5831 664
rect 2394 652 4866 663
rect 2394 640 4497 652
rect 2025 624 4497 640
rect 2025 612 2059 624
rect 1929 575 1959 582
rect 1991 578 2019 582
rect 1889 569 1901 573
rect 1917 569 1959 575
rect 1877 561 1959 569
rect 1769 527 1797 557
rect 1887 555 1913 561
rect 1917 551 1959 561
rect 1915 535 1973 541
rect 1911 527 1951 535
rect 1769 495 1803 527
rect 1911 501 1977 527
rect 1915 495 1973 501
rect 1769 493 1797 495
rect 2001 493 2019 578
rect 2025 544 2039 612
rect 2041 572 2059 608
rect 2075 606 4497 624
rect 2044 544 2059 572
rect 2025 514 2059 544
rect 2025 493 2031 514
rect 381 441 410 487
rect 6 434 41 441
rect 83 434 135 441
rect 171 434 223 441
rect 270 413 292 441
rect 447 413 470 481
rect 475 453 515 487
rect 569 453 603 487
rect 1709 470 1740 493
rect 1812 487 1864 493
rect 1803 482 1864 487
rect 1877 487 2031 493
rect 2044 487 2059 514
rect 1803 470 1812 482
rect 1823 470 1853 482
rect 1709 466 1751 470
rect 1803 469 1864 470
rect 1877 469 2059 487
rect 1709 462 1762 466
rect 1709 459 1774 462
rect 475 441 498 453
rect 1690 425 1740 428
rect -32 345 23 379
rect 464 339 470 408
rect 1735 394 1740 425
rect 1769 399 1774 459
rect 1790 459 2059 469
rect 2078 459 2119 606
rect 1790 433 1803 459
rect 1905 433 2007 459
rect 2078 448 2093 459
rect 2104 448 2119 459
rect 2138 486 2172 606
rect 2180 604 2231 606
rect 2180 589 2238 604
rect 2249 600 2370 606
rect 2371 600 4497 606
rect 4503 624 4514 646
rect 4517 635 4560 652
rect 4563 635 4571 652
rect 4577 651 4653 652
rect 4577 647 4648 651
rect 4577 635 4611 647
rect 4614 635 4648 647
rect 4517 631 4648 635
rect 4526 624 4648 631
rect 4503 617 4648 624
rect 4660 617 4699 652
rect 4503 612 4654 617
rect 4659 612 4699 617
rect 4702 651 4748 652
rect 4702 612 4753 651
rect 4503 604 4514 612
rect 2249 594 2326 600
rect 2249 589 2342 594
rect 2192 586 2231 589
rect 2238 586 2268 589
rect 2280 588 2310 589
rect 2315 588 2342 589
rect 2343 588 2370 600
rect 2192 585 2206 586
rect 2280 556 2370 588
rect 2377 584 2388 600
rect 2394 584 2407 600
rect 2411 584 4497 600
rect 2371 572 4497 584
rect 2280 554 2346 556
rect 2284 548 2310 554
rect 2315 548 2346 554
rect 2224 542 2282 548
rect 2224 524 2236 542
rect 2246 524 2286 542
rect 2319 538 2346 548
rect 2377 538 2388 572
rect 2394 532 2407 572
rect 2411 550 4497 572
rect 4521 602 4562 612
rect 4565 608 4648 612
rect 4659 608 4753 612
rect 4521 594 4556 602
rect 4565 594 4642 608
rect 4659 604 4711 608
rect 4521 589 4642 594
rect 4653 589 4711 604
rect 4521 556 4611 589
rect 4623 558 4653 589
rect 4660 586 4699 589
rect 4665 585 4699 586
rect 2411 532 2893 550
rect 2908 539 3983 550
rect 2908 534 3995 539
rect 2224 520 2286 524
rect 2361 520 2380 532
rect 2394 520 2893 532
rect 2220 508 2286 520
rect 2371 516 2893 520
rect 2224 502 2282 508
rect 2196 486 2310 496
rect 2394 486 2893 516
rect 2138 469 2893 486
rect 2138 466 2630 469
rect 2138 452 2407 466
rect 2394 448 2407 452
rect 2411 461 2630 466
rect 2772 461 2797 469
rect 2411 448 2524 461
rect 2075 433 2524 448
rect 1790 431 2524 433
rect 1801 425 2524 431
rect 1801 422 1900 425
rect 1812 410 1900 422
rect 1801 399 1900 410
rect 1901 422 2042 425
rect 1901 410 2031 422
rect 2075 416 2524 425
rect 2816 427 2831 469
rect 2896 464 3995 534
rect 3998 528 4497 550
rect 4545 554 4611 556
rect 4545 548 4576 554
rect 4581 548 4607 554
rect 4545 538 4572 548
rect 4609 542 4667 548
rect 3998 486 4503 528
rect 4511 520 4530 532
rect 4605 524 4645 542
rect 4605 520 4667 524
rect 4605 508 4671 520
rect 4719 514 4753 608
rect 4609 502 4667 508
rect 4719 503 4730 514
rect 4581 486 4695 496
rect 4738 494 4753 514
rect 4719 486 4753 494
rect 3998 469 4753 486
rect 2908 441 3983 464
rect 1901 399 2042 410
rect 890 391 924 393
rect -1470 222 -1435 256
rect -1137 239 -1084 275
rect 242 253 264 311
rect 270 281 292 339
rect 447 281 470 339
rect 492 311 498 380
rect 861 369 924 391
rect 2075 380 2464 416
rect 918 363 924 365
rect 2143 363 2144 380
rect 2155 372 2189 380
rect 2243 372 2277 380
rect 2331 372 2365 380
rect 2419 372 2453 380
rect 2464 370 2465 380
rect 2519 370 2532 398
rect 2155 363 2223 370
rect 833 341 924 363
rect 2816 356 2824 427
rect 2958 426 3002 441
rect 2958 425 3005 426
rect 2958 420 3008 425
rect 2958 414 3005 420
rect 2958 404 3002 414
rect 2934 391 2977 398
rect 2925 386 2977 391
rect 3120 386 3124 399
rect 3132 386 3166 441
rect 3185 435 3219 441
rect 3287 439 3335 441
rect 3356 439 3390 441
rect 3458 439 3487 441
rect 3290 435 3320 439
rect 3322 435 3333 439
rect 3345 435 3390 439
rect 3182 401 3219 435
rect 3285 417 3320 435
rect 3345 417 3411 435
rect 2909 357 2975 386
rect 3074 373 3166 386
rect 3132 356 3140 373
rect 3148 367 3166 373
rect 2816 352 2850 356
rect 3132 352 3143 356
rect 2816 345 3143 352
rect 2816 339 3132 345
rect 2816 319 3070 339
rect 3090 319 3120 339
rect 3151 319 3166 367
rect 2816 318 3178 319
rect 475 253 498 311
rect 2825 302 2859 306
rect 2816 293 2871 302
rect 2825 284 2859 293
rect 3151 265 3178 318
rect 3185 299 3219 401
rect 3185 284 3232 299
rect 3246 284 3248 384
rect 3274 284 3276 368
rect 3327 367 3411 417
rect 3327 351 3390 367
rect 3356 340 3367 351
rect 3379 340 3390 351
rect 3501 351 3535 441
rect 3556 439 3604 441
rect 3558 435 3569 439
rect 3571 435 3601 439
rect 3672 435 3706 441
rect 3571 401 3606 435
rect 3643 401 3659 435
rect 3672 401 3709 435
rect 3725 407 3759 441
rect 3889 426 3933 441
rect 4060 427 4075 469
rect 4094 461 4129 469
rect 4261 466 4753 469
rect 4261 461 4480 466
rect 3886 425 3933 426
rect 3883 420 3933 425
rect 3886 414 3933 420
rect 3571 351 3601 401
rect 3672 384 3706 401
rect 3672 373 3683 384
rect 3691 373 3706 384
rect 3501 340 3512 351
rect 3524 340 3535 351
rect 3672 319 3706 373
rect 3725 384 3743 407
rect 3751 386 3759 407
rect 3889 404 3933 414
rect 3767 386 3771 399
rect 3914 391 3957 398
rect 3914 386 3966 391
rect 3751 384 3817 386
rect 3725 373 3817 384
rect 3725 352 3759 373
rect 3916 357 3982 386
rect 4067 356 4075 427
rect 4367 448 4480 461
rect 4484 452 4753 466
rect 4772 452 4813 652
rect 4814 608 4866 652
rect 4880 612 4882 617
rect 4886 612 4936 663
rect 4946 659 5014 663
rect 4946 654 5008 659
rect 4946 641 4970 654
rect 4974 642 5008 654
rect 5023 642 5831 663
rect 4974 641 5020 642
rect 4832 493 4866 608
rect 4874 608 4936 612
rect 4943 628 5020 641
rect 5021 640 5831 642
rect 5839 674 5865 716
rect 5877 695 5879 716
rect 5927 710 5973 716
rect 5921 676 5973 710
rect 5987 716 6047 723
rect 5987 696 6037 716
rect 5939 674 5995 676
rect 5839 640 5873 674
rect 5927 666 6005 674
rect 6041 666 6047 716
rect 6051 681 6071 746
rect 6079 743 6097 746
rect 6079 705 6103 743
rect 6113 735 6219 769
rect 6079 681 6097 705
rect 6113 681 6147 735
rect 6151 681 6219 735
rect 6051 666 6109 681
rect 5927 651 6109 666
rect 6113 666 6219 681
rect 6246 666 6259 817
rect 6271 805 6314 817
rect 6356 805 6402 817
rect 6407 805 6414 817
rect 6271 801 6322 805
rect 6356 801 6414 805
rect 6271 800 6328 801
rect 6271 795 6333 800
rect 6274 793 6333 795
rect 6362 793 6410 801
rect 6274 768 6322 793
rect 6268 753 6322 768
rect 6326 753 6333 793
rect 6368 753 6410 793
rect 6268 723 6326 753
rect 6364 723 6422 753
rect 6268 708 6322 723
rect 6274 696 6322 708
rect 6268 682 6322 696
rect 6268 681 6287 682
rect 6288 681 6322 682
rect 6326 681 6333 723
rect 6368 687 6410 723
rect 6362 682 6410 687
rect 6362 681 6370 682
rect 6376 681 6410 682
rect 6268 670 6326 681
rect 6362 670 6422 681
rect 6276 666 6334 670
rect 6113 659 6334 666
rect 6364 659 6422 670
rect 6430 659 6435 817
rect 6467 805 6469 899
rect 6464 801 6469 805
rect 6458 793 6469 801
rect 6458 753 6463 793
rect 6464 789 6469 793
rect 6482 869 6616 899
rect 6482 823 6516 869
rect 6534 835 6612 869
rect 6534 833 6603 835
rect 6534 829 6604 833
rect 6608 829 6610 835
rect 6482 753 6532 823
rect 6534 822 6610 829
rect 6636 822 6638 909
rect 6696 899 6698 909
rect 6646 884 6704 899
rect 6724 884 6726 909
rect 6727 899 6860 911
rect 6646 881 6724 884
rect 6646 878 6704 881
rect 6727 878 6792 899
rect 6646 869 6792 878
rect 6658 855 6792 869
rect 6646 829 6792 855
rect 6870 898 6885 927
rect 6904 916 6963 927
rect 7042 919 7110 927
rect 7111 919 7163 927
rect 7176 919 7613 927
rect 6904 904 6952 916
rect 6904 898 6963 904
rect 7042 898 7286 919
rect 6870 894 7286 898
rect 7298 909 7613 919
rect 7677 909 7711 943
rect 7723 909 7823 943
rect 7877 909 7999 968
rect 8053 958 8099 968
rect 7298 902 7723 909
rect 6870 893 7254 894
rect 6870 863 7078 893
rect 6870 859 7114 863
rect 6870 852 7130 859
rect 6842 830 7130 852
rect 6842 829 6885 830
rect 6646 822 6885 829
rect 6534 821 6885 822
rect 6534 819 6569 821
rect 6599 819 6604 821
rect 6616 819 6630 821
rect 6452 723 6532 753
rect 6458 681 6463 723
rect 6482 681 6532 723
rect 6452 674 6532 681
rect 6535 783 6569 819
rect 6570 817 6604 819
rect 6535 723 6550 783
rect 6535 674 6569 723
rect 6113 651 6422 659
rect 6452 651 6569 674
rect 6599 659 6603 817
rect 6636 805 6638 821
rect 6658 817 6692 821
rect 6633 801 6667 805
rect 6679 801 6692 817
rect 6724 818 6885 821
rect 6904 818 6948 830
rect 6724 805 6948 818
rect 6721 804 6948 805
rect 6721 801 6779 804
rect 6809 801 6814 804
rect 6817 801 6843 804
rect 6621 780 6683 801
rect 6621 696 6623 780
rect 6627 777 6631 780
rect 6633 777 6683 780
rect 6626 743 6683 777
rect 6687 768 6692 801
rect 6709 797 6771 801
rect 6710 790 6771 797
rect 6694 743 6771 790
rect 6775 768 6779 801
rect 6803 776 6849 801
rect 6803 768 6807 776
rect 6817 768 6849 776
rect 6627 696 6631 743
rect 6633 709 6771 743
rect 6817 724 6843 768
rect 6633 696 6683 709
rect 5927 642 6097 651
rect 5927 640 5973 642
rect 6005 640 6097 642
rect 6113 640 6147 651
rect 6151 640 6410 651
rect 6464 640 6569 651
rect 5021 628 6219 640
rect 6246 632 6550 640
rect 4943 610 6219 628
rect 4874 594 4920 608
rect 4943 595 5024 610
rect 5079 601 5082 610
rect 4943 594 5042 595
rect 4874 582 4905 594
rect 4962 583 5040 594
rect 4962 582 5020 583
rect 4872 578 4900 582
rect 4872 551 4890 578
rect 4974 575 5004 582
rect 4962 569 5004 575
rect 4962 561 5014 569
rect 5088 568 5109 610
rect 4962 551 5004 561
rect 5088 557 5099 568
rect 4914 541 4932 551
rect 4914 535 4976 541
rect 4914 527 4932 535
rect 4940 527 4980 535
rect 5114 527 5122 610
rect 4914 501 4980 527
rect 4914 495 4976 501
rect 5088 495 5122 527
rect 4914 493 4932 495
rect 5114 493 5122 495
rect 5148 493 5182 610
rect 5201 568 5216 610
rect 5230 568 5235 610
rect 5345 607 6219 610
rect 6254 607 6550 632
rect 6621 636 6683 696
rect 5345 606 6550 607
rect 5345 598 5885 606
rect 5345 586 5360 598
rect 5392 586 5885 598
rect 5915 586 5973 606
rect 6051 589 6109 606
rect 5201 546 5235 568
rect 5392 574 5831 586
rect 5839 582 5873 586
rect 5927 582 5961 586
rect 6063 585 6097 589
rect 6113 574 6147 606
rect 6151 601 6219 606
rect 6151 589 6197 601
rect 6288 589 6410 606
rect 6151 585 6200 589
rect 6166 574 6200 585
rect 5392 572 6200 574
rect 5392 571 5995 572
rect 6029 571 6200 572
rect 5392 557 6200 571
rect 5517 546 5521 557
rect 5201 512 5317 546
rect 5331 535 5444 546
rect 5480 535 5521 546
rect 5797 551 6200 557
rect 5797 548 6040 551
rect 5797 540 5838 548
rect 5885 541 6040 548
rect 5988 540 6040 541
rect 6098 542 6200 551
rect 6098 540 6147 542
rect 5331 523 5433 535
rect 5491 523 5521 535
rect 5320 516 5433 523
rect 5320 512 5372 516
rect 5480 512 5532 523
rect 6166 521 6200 542
rect 6288 573 6334 589
rect 6364 573 6374 589
rect 6288 521 6322 573
rect 6376 521 6410 589
rect 6482 600 6569 606
rect 6575 600 6618 613
rect 6482 583 6532 600
rect 6482 521 6516 583
rect 4832 469 5014 493
rect 5027 487 5079 493
rect 5027 482 5088 487
rect 5038 470 5068 482
rect 5079 470 5088 482
rect 5151 478 5182 493
rect 6166 508 6224 521
rect 6166 498 6202 508
rect 6166 487 6177 498
rect 6262 487 6516 521
rect 6535 487 6569 600
rect 6575 572 6590 585
rect 5151 470 5181 478
rect 5027 469 5088 470
rect 4832 459 5101 469
rect 5140 466 5182 470
rect 5129 462 5182 466
rect 4484 448 4497 452
rect 4772 448 4787 452
rect 4798 448 4813 452
rect 4367 433 4816 448
rect 4908 433 4962 445
rect 5088 433 5101 459
rect 4367 425 5101 433
rect 4367 416 4816 425
rect 4849 422 4973 425
rect 5002 422 5101 425
rect 4427 380 4816 416
rect 4860 410 4962 422
rect 5013 410 5101 422
rect 4849 399 4973 410
rect 5002 399 5101 410
rect 5117 459 5182 462
rect 5117 399 5122 459
rect 6376 453 6410 487
rect 6535 441 6564 487
rect 6621 468 6623 636
rect 6633 629 6683 636
rect 6721 629 6771 709
rect 6809 719 6843 724
rect 6851 752 6948 804
rect 6851 741 6885 752
rect 6892 741 6948 752
rect 6958 741 6976 830
rect 7010 791 7130 830
rect 6984 772 6998 782
rect 7010 775 7112 791
rect 6984 770 7004 772
rect 6980 752 7004 770
rect 6984 741 7004 752
rect 7010 770 7094 775
rect 7164 770 7174 782
rect 7010 769 7110 770
rect 7010 751 7140 769
rect 7010 744 7094 751
rect 7110 748 7140 751
rect 7130 744 7140 748
rect 7164 751 7178 770
rect 7006 741 7010 744
rect 6851 740 7010 741
rect 6851 736 6877 740
rect 6851 719 6885 736
rect 6809 711 6885 719
rect 6904 711 6948 740
rect 6958 711 6976 740
rect 6984 711 7004 740
rect 7012 732 7032 744
rect 7042 732 7058 744
rect 7064 740 7152 744
rect 7164 740 7174 751
rect 7186 740 7198 893
rect 7220 865 7254 893
rect 7298 874 7366 902
rect 7371 874 7372 902
rect 7383 874 7417 902
rect 7471 874 7505 902
rect 7517 875 7723 902
rect 7755 875 7999 909
rect 8056 908 8087 958
rect 8090 928 8125 958
rect 8137 951 8152 964
rect 8134 928 8152 951
rect 8090 924 8156 928
rect 8090 908 8099 924
rect 8134 918 8152 924
rect 8165 923 8180 992
rect 8264 979 8313 995
rect 8264 968 8275 979
rect 8283 944 8298 979
rect 8056 893 8099 908
rect 8162 894 8180 923
rect 8056 890 8087 893
rect 8162 890 8190 894
rect 8264 890 8298 944
rect 7517 874 7585 875
rect 7273 865 7298 874
rect 7220 778 7298 865
rect 7369 840 7517 874
rect 7527 840 7539 874
rect 7545 841 7623 874
rect 7723 855 7791 875
rect 7577 840 7623 841
rect 7371 813 7372 840
rect 7517 819 7585 840
rect 7589 819 7623 840
rect 7704 830 7711 855
rect 7723 821 7823 855
rect 7877 821 7911 875
rect 7912 857 7999 875
rect 7912 856 8028 857
rect 8053 856 8087 890
rect 8165 856 8199 890
rect 8264 856 8299 890
rect 7912 822 8099 856
rect 8131 822 8299 856
rect 7912 821 8028 822
rect 7642 819 7723 821
rect 7517 818 7723 819
rect 7517 813 7585 818
rect 7371 812 7585 813
rect 7220 751 7320 778
rect 7220 740 7254 751
rect 7273 740 7298 751
rect 7064 739 7298 740
rect 7076 735 7086 739
rect 7122 732 7152 739
rect 7164 735 7174 739
rect 7186 735 7198 739
rect 7220 735 7240 739
rect 7012 711 7058 732
rect 7106 713 7152 732
rect 6809 685 7006 711
rect 7012 704 7052 711
rect 7018 685 7052 704
rect 7106 685 7140 713
rect 7220 711 7254 735
rect 7273 711 7307 739
rect 7152 685 7307 711
rect 7391 704 7410 806
rect 7419 772 7477 778
rect 7419 738 7438 772
rect 7419 732 7477 738
rect 7589 730 7600 741
rect 7608 730 7623 818
rect 7441 712 7543 713
rect 7589 712 7623 730
rect 7642 787 7677 818
rect 7777 800 8028 821
rect 7835 798 7865 800
rect 7824 790 7876 798
rect 7642 712 7676 787
rect 7713 769 7790 790
rect 7820 769 7889 790
rect 7912 786 8028 800
rect 8283 796 8287 822
rect 8292 800 8299 822
rect 8317 803 8351 995
rect 8419 987 8430 997
rect 8431 987 8464 997
rect 8419 963 8464 987
rect 8498 1016 9289 1021
rect 8498 976 8920 1016
rect 10255 1000 10270 1034
rect 10571 1015 10605 1045
rect 10325 1004 10485 1015
rect 10494 1007 10605 1015
rect 10505 1004 10605 1007
rect 10336 1001 10474 1004
rect 10336 992 10366 1001
rect 10325 981 10377 992
rect 10408 987 10474 1001
rect 10516 992 10605 1004
rect 10505 987 10605 992
rect 10624 987 10658 1228
rect 10666 1099 10692 1228
rect 10704 1103 10706 1228
rect 10726 1184 10778 1228
rect 10791 1279 10831 1291
rect 10843 1279 10872 1291
rect 10791 1224 10872 1279
rect 10791 1212 10806 1224
rect 10797 1208 10806 1212
rect 10826 1184 10872 1224
rect 10879 1224 10898 1317
rect 10879 1212 10894 1224
rect 10885 1208 10894 1212
rect 10906 1212 10931 1392
rect 10940 1212 10974 1440
rect 11050 1421 12596 1520
rect 12642 1509 12832 1520
rect 12676 1503 12710 1507
rect 12764 1503 12798 1507
rect 12664 1495 12722 1503
rect 12752 1495 12810 1503
rect 12670 1481 12716 1495
rect 12758 1481 12810 1495
rect 10993 1392 12596 1421
rect 12676 1445 12716 1481
rect 12726 1463 12744 1475
rect 12764 1473 12810 1481
rect 12752 1463 12810 1473
rect 10985 1387 12596 1392
rect 10985 1359 11028 1387
rect 11050 1359 12596 1387
rect 10985 1316 12596 1359
rect 10985 1224 11061 1316
rect 11085 1258 11119 1316
rect 11120 1266 11131 1316
rect 11135 1285 11237 1316
rect 11191 1269 11201 1285
rect 11203 1269 11237 1285
rect 11191 1266 11237 1269
rect 11120 1258 11237 1266
rect 11085 1252 11237 1258
rect 11085 1238 11141 1252
rect 11191 1238 11237 1252
rect 11085 1224 11153 1238
rect 11189 1224 11237 1238
rect 11291 1296 11359 1316
rect 11419 1296 12596 1316
rect 11291 1263 12596 1296
rect 11291 1243 11748 1263
rect 11788 1261 12596 1263
rect 11786 1243 12596 1261
rect 11291 1228 12596 1243
rect 12604 1228 12630 1370
rect 12642 1295 12644 1417
rect 12670 1407 12672 1417
rect 12676 1407 12710 1445
rect 12722 1429 12810 1463
rect 12752 1423 12788 1429
rect 12795 1423 12810 1429
rect 12752 1419 12810 1423
rect 12664 1369 12710 1407
rect 12664 1366 12726 1369
rect 12670 1323 12672 1366
rect 12676 1335 12726 1366
rect 12692 1323 12726 1335
rect 12730 1323 12732 1366
rect 12758 1323 12760 1394
rect 12762 1369 12810 1419
rect 12828 1369 12832 1373
rect 12844 1369 12862 1373
rect 12790 1335 12804 1369
rect 12794 1323 12804 1335
rect 12816 1323 12864 1369
rect 12692 1310 12738 1323
rect 12794 1319 12798 1323
rect 12686 1276 12738 1310
rect 12822 1297 12836 1323
rect 12822 1295 12832 1297
rect 12828 1285 12832 1295
rect 12704 1228 12738 1276
rect 12754 1242 12760 1276
rect 12844 1228 12862 1323
rect 11291 1224 12650 1228
rect 10985 1212 11028 1224
rect 11107 1216 11153 1224
rect 11107 1212 11141 1216
rect 11146 1212 11153 1216
rect 10906 1208 10919 1212
rect 10726 1174 10872 1184
rect 10726 1111 10766 1174
rect 10771 1171 10872 1174
rect 10771 1137 10886 1171
rect 10814 1123 10886 1137
rect 10814 1111 10872 1123
rect 10814 1098 10873 1111
rect 10742 1087 10873 1098
rect 10742 1026 10762 1087
rect 10770 1064 10828 1070
rect 10770 1053 10832 1064
rect 10770 1045 10790 1053
rect 10766 1030 10790 1045
rect 10766 1024 10828 1030
rect 10766 1014 10790 1024
rect 10843 1014 10873 1087
rect 10891 1085 10894 1208
rect 10940 1197 10953 1212
rect 10959 1197 10974 1212
rect 10940 1167 10974 1197
rect 10940 1156 10951 1167
rect 10959 1066 10974 1167
rect 10993 1066 11027 1212
rect 11107 1133 11153 1212
rect 11095 1124 11153 1133
rect 11159 1156 11175 1184
rect 11195 1163 11229 1224
rect 11309 1212 12650 1224
rect 11234 1163 11241 1212
rect 11326 1210 12650 1212
rect 11326 1186 12135 1210
rect 12157 1186 12650 1210
rect 12680 1186 12738 1228
rect 12816 1189 12874 1228
rect 11326 1166 12117 1186
rect 11195 1156 11241 1163
rect 11159 1124 11187 1156
rect 11189 1132 11241 1156
rect 11309 1150 12117 1166
rect 12157 1174 12596 1186
rect 12604 1182 12638 1186
rect 12692 1182 12726 1186
rect 12828 1185 12862 1189
rect 12878 1174 12912 1520
rect 12931 1391 12965 1520
rect 13089 1509 13123 1520
rect 13073 1497 13139 1509
rect 13073 1487 13091 1497
rect 13041 1450 13091 1487
rect 13121 1481 13139 1497
rect 13247 1499 13258 1510
rect 13266 1503 13281 1580
rect 13300 1546 13335 1580
rect 13300 1503 13334 1546
rect 13266 1499 13334 1503
rect 13247 1469 13334 1499
rect 13247 1458 13258 1469
rect 13266 1455 13281 1469
rect 13033 1437 13091 1450
rect 13121 1438 13144 1450
rect 13033 1422 13079 1437
rect 12931 1373 12984 1391
rect 12916 1201 12984 1373
rect 13045 1389 13079 1422
rect 13121 1435 13167 1438
rect 13121 1401 13129 1435
rect 13045 1282 13087 1389
rect 13053 1239 13087 1282
rect 13091 1270 13098 1400
rect 13133 1389 13167 1435
rect 13172 1401 13179 1450
rect 13247 1423 13281 1455
rect 13133 1282 13175 1389
rect 13141 1270 13175 1282
rect 13091 1239 13099 1270
rect 13053 1223 13099 1239
rect 13123 1223 13175 1270
rect 12916 1189 12962 1201
rect 13053 1189 13175 1223
rect 12916 1185 12965 1189
rect 12931 1174 12965 1185
rect 12157 1171 12760 1174
rect 12794 1171 12965 1174
rect 12157 1157 12965 1171
rect 11309 1144 11379 1150
rect 11385 1144 11396 1150
rect 11189 1124 11263 1132
rect 11037 1086 11061 1102
rect 11073 1086 11091 1102
rect 11037 1066 11065 1086
rect 11069 1066 11091 1086
rect 11095 1087 11141 1124
rect 11146 1087 11153 1124
rect 11095 1066 11153 1087
rect 11195 1116 11263 1124
rect 11275 1116 11295 1132
rect 11195 1082 11295 1116
rect 11195 1072 11263 1082
rect 10923 1057 11153 1066
rect 10923 1011 11135 1057
rect 11159 1038 11187 1072
rect 11189 1066 11263 1072
rect 11275 1066 11295 1082
rect 11189 1058 11241 1066
rect 11207 1054 11229 1058
rect 11309 1048 11396 1144
rect 11508 1124 11520 1150
rect 11551 1124 11566 1150
rect 11508 1118 11566 1124
rect 11579 1096 11594 1150
rect 11480 1090 11594 1096
rect 11697 1076 11712 1150
rect 11678 1063 11712 1076
rect 11201 1038 11396 1048
rect 11159 1032 11396 1038
rect 11649 1045 11712 1063
rect 11731 1065 12117 1150
rect 12562 1151 12965 1157
rect 12562 1148 12805 1151
rect 12562 1140 12603 1148
rect 12650 1141 12805 1148
rect 12753 1140 12805 1141
rect 12863 1142 12965 1151
rect 12863 1140 12912 1142
rect 12931 1121 12965 1142
rect 13053 1173 13099 1189
rect 13129 1173 13139 1189
rect 13053 1121 13087 1173
rect 13141 1121 13175 1189
rect 13247 1183 13297 1423
rect 13247 1121 13281 1183
rect 12931 1108 12989 1121
rect 12931 1098 12967 1108
rect 12931 1087 12942 1098
rect 13027 1087 13281 1121
rect 13300 1087 13334 1469
rect 13343 1435 13368 1469
rect 13474 1397 13490 1401
rect 13444 1229 13448 1385
rect 13486 1217 13490 1389
rect 13532 1229 13536 1385
rect 13474 1186 13490 1217
rect 13442 1120 13444 1186
rect 13474 1170 13508 1186
rect 13458 1136 13508 1170
rect 13474 1120 13508 1136
rect 11159 1030 11309 1032
rect 11139 1011 11159 1017
rect 11201 1011 11309 1030
rect 10923 998 11163 1011
rect 11169 1006 11309 1011
rect 10750 996 10812 998
rect 10686 991 10731 996
rect 10681 987 10697 991
rect 10408 984 10780 987
rect 8498 963 8703 976
rect 8708 965 8742 976
rect 8796 965 8830 976
rect 8884 965 8918 976
rect 8920 963 8930 976
rect 8417 959 8452 963
rect 8417 943 8434 959
rect 8507 958 8533 963
rect 8544 958 8559 963
rect 8507 947 8559 958
rect 8507 943 8563 947
rect 8417 921 8419 943
rect 8435 919 8534 939
rect 8572 915 8587 952
rect 8649 929 8667 963
rect 10219 945 10274 979
rect 10410 970 10780 984
rect 10959 986 11028 998
rect 11101 997 11163 998
rect 11165 1002 11309 1006
rect 11326 1002 11396 1032
rect 11165 997 11396 1002
rect 10959 970 10974 986
rect 10991 971 11061 986
rect 11101 983 11396 997
rect 11464 1008 11564 1034
rect 11649 1029 11727 1045
rect 11731 1029 11765 1065
rect 11873 1055 11886 1065
rect 11845 1033 11878 1037
rect 11833 1031 11878 1033
rect 11464 996 11567 1008
rect 11476 992 11510 996
rect 11678 995 11765 1029
rect 11778 997 11878 1031
rect 11899 1033 11966 1055
rect 12047 1049 12078 1065
rect 13141 1053 13175 1087
rect 12047 1046 12081 1049
rect 12047 1038 12058 1046
rect 12070 1038 12081 1046
rect 13300 1041 13329 1087
rect 13616 1068 13620 1401
rect 13386 1041 13620 1068
rect 11899 1021 11979 1033
rect 10991 970 11028 971
rect 10410 945 11028 970
rect 8463 905 8521 911
rect 8460 891 8521 905
rect 8384 875 8385 879
rect 8460 875 8518 891
rect 8372 831 8405 875
rect 8460 871 8547 875
rect 8460 855 8518 871
rect 8372 803 8418 831
rect 8472 803 8506 855
rect 8560 803 8605 837
rect 8633 803 8667 929
rect 10110 821 10112 911
rect 10138 804 10140 939
rect 10588 928 11028 945
rect 11101 969 11131 983
rect 11135 980 11396 983
rect 11467 980 11501 984
rect 11135 977 11235 980
rect 11135 969 11137 977
rect 11139 971 11235 977
rect 11191 969 11235 971
rect 11101 965 11235 969
rect 11101 961 11201 965
rect 11203 961 11235 965
rect 11101 943 11235 961
rect 11309 968 11396 980
rect 11461 968 11513 980
rect 10588 919 11027 928
rect 10590 894 10612 919
rect 10666 894 10700 919
rect 10712 909 11027 919
rect 11091 909 11125 943
rect 11137 909 11237 943
rect 11309 909 11413 968
rect 11467 958 11513 968
rect 10712 902 11137 909
rect 10712 892 10780 902
rect 10785 892 10786 902
rect 10797 894 10831 902
rect 10885 894 10919 902
rect 10931 892 11137 902
rect 10957 875 11137 892
rect 11169 875 11413 909
rect 11470 908 11501 958
rect 11504 928 11539 958
rect 11551 951 11566 964
rect 11548 928 11566 951
rect 11504 924 11570 928
rect 11504 908 11513 924
rect 11548 918 11566 924
rect 11579 923 11594 992
rect 11678 979 11727 995
rect 11678 968 11689 979
rect 11697 944 11712 979
rect 11470 893 11513 908
rect 11576 894 11594 923
rect 11470 890 11501 893
rect 11576 890 11604 894
rect 11678 890 11712 944
rect 10957 839 10999 875
rect 11137 839 11205 875
rect 11326 856 11413 875
rect 11467 856 11501 890
rect 11579 856 11613 890
rect 11678 856 11713 890
rect 11326 839 11513 856
rect 11362 822 11513 839
rect 11545 822 11713 856
rect 11379 812 11413 822
rect 8317 800 8353 803
rect 8317 788 8332 800
rect 7713 753 7790 762
rect 7820 753 7917 762
rect 7713 741 7917 753
rect 7760 734 7874 741
rect 7414 686 7433 691
rect 7441 686 7784 712
rect 7788 706 7846 725
rect 7958 720 7964 786
rect 8317 769 8321 788
rect 8372 785 8606 803
rect 8649 788 8667 803
rect 11697 796 11701 822
rect 11706 800 11713 822
rect 11731 803 11765 995
rect 11833 987 11844 997
rect 11845 987 11878 997
rect 11833 963 11878 987
rect 11921 994 12000 1021
rect 12047 997 12081 1038
rect 13444 1034 13474 1041
rect 13532 1034 13562 1041
rect 11921 984 11979 994
rect 11831 959 11866 963
rect 11831 943 11848 959
rect 11921 958 11947 984
rect 11964 980 11979 984
rect 11958 969 11979 980
rect 12056 976 12081 997
rect 11958 958 11973 969
rect 11921 947 11973 958
rect 11921 943 11977 947
rect 11831 921 11833 943
rect 11849 919 11948 939
rect 11986 915 12001 952
rect 12063 929 12081 976
rect 11877 905 11935 911
rect 11874 891 11935 905
rect 11798 875 11799 879
rect 11874 875 11932 891
rect 11786 831 11819 875
rect 11874 871 11961 875
rect 11874 855 11932 871
rect 11786 803 11832 831
rect 11886 803 11920 855
rect 11974 803 12019 837
rect 12047 803 12081 929
rect 11731 800 11767 803
rect 8430 780 8460 785
rect 8518 780 8548 785
rect 8419 769 8471 780
rect 8507 769 8559 780
rect 8656 777 8667 788
rect 11127 769 11204 790
rect 11234 769 11303 790
rect 11731 788 11746 800
rect 11731 769 11735 788
rect 11786 785 12020 803
rect 12063 788 12081 803
rect 11844 780 11874 785
rect 11932 780 11962 785
rect 11833 769 11885 780
rect 11921 769 11973 780
rect 12070 777 12081 788
rect 11127 741 11204 762
rect 11234 741 11331 762
rect 7958 712 7992 720
rect 7850 686 8028 712
rect 6633 604 6667 629
rect 6721 617 6755 629
rect 6633 600 6688 604
rect 6633 502 6673 600
rect 6677 570 6679 586
rect 6688 576 6701 600
rect 6681 570 6701 576
rect 6709 570 6755 617
rect 6809 613 6843 685
rect 6844 652 6938 685
rect 6984 652 7152 685
rect 7186 652 7254 685
rect 7256 652 7290 685
rect 6844 651 7290 652
rect 7387 679 7419 685
rect 7420 679 7543 686
rect 7555 679 8244 686
rect 7387 651 8269 679
rect 6677 536 6755 570
rect 6677 520 6679 536
rect 6681 530 6701 536
rect 6709 520 6755 536
rect 6633 468 6667 502
rect 6721 468 6755 520
rect 6817 502 6843 613
rect 6809 468 6843 502
rect 6851 468 6885 651
rect 6621 441 6855 468
rect 6668 434 6720 441
rect 6756 434 6808 441
rect 6870 434 6885 468
rect 6904 434 6938 651
rect 7108 481 7126 505
rect 5151 425 5201 428
rect 5151 394 5156 425
rect 6904 400 6919 434
rect 7239 381 7254 651
rect 7273 381 7307 651
rect 7387 523 7421 651
rect 7475 523 7509 651
rect 7419 464 7477 470
rect 7419 430 7431 464
rect 7419 424 7477 430
rect 4427 372 4472 380
rect 4526 372 4560 380
rect 4614 372 4648 380
rect 4702 372 4736 380
rect 4427 370 4440 372
rect 4748 363 4816 380
rect 4041 352 4075 356
rect 3725 339 4075 352
rect 6868 345 6923 379
rect 7273 347 7288 381
rect 3725 319 3760 339
rect 3771 319 3801 339
rect 3821 319 4075 339
rect 3279 288 3331 299
rect 3290 284 3320 288
rect 3452 284 3473 299
rect 3560 288 3612 299
rect 3571 284 3601 288
rect 3688 284 3706 319
rect 3185 265 3432 284
rect 3452 265 3706 284
rect 3713 318 4075 319
rect 3713 265 3760 318
rect 3867 281 3884 318
rect 3895 281 3912 318
rect 4032 302 4066 306
rect 4020 293 4075 302
rect 4032 284 4066 293
rect 82 221 88 232
rect 3151 231 3166 265
rect 3274 251 3276 265
rect 3244 231 3278 234
rect 3332 231 3366 234
rect 3525 231 3559 234
rect 3613 231 3647 234
rect 3725 231 3740 265
rect 130 221 136 228
rect 169 221 176 228
rect 218 221 228 228
rect 82 200 96 204
rect 82 193 136 200
rect 169 193 200 200
rect 197 59 200 193
rect 225 59 228 221
rect 6660 221 6673 311
rect 2353 169 2422 190
rect 2452 169 2529 190
rect 3491 168 3510 204
rect 3519 168 3538 204
rect 4475 169 4538 190
rect 2325 141 2422 162
rect 2452 141 2529 162
rect 242 59 258 109
rect 3282 104 3284 168
rect 3310 104 3312 168
rect 4475 141 4566 162
rect 6660 140 6666 221
rect 6688 193 6701 339
rect 7608 328 7623 651
rect 7642 328 7676 651
rect 7756 613 7790 642
rect 7844 613 7878 642
rect 7975 626 8046 651
rect 8107 626 8265 651
rect 8326 626 8361 660
rect 7642 294 7657 328
rect 7975 275 8045 626
rect 8327 607 8361 626
rect 8157 558 8215 564
rect 8157 524 8169 558
rect 8157 518 8215 524
rect 8157 358 8215 364
rect 8157 324 8169 358
rect 8157 318 8215 324
rect 7975 239 8028 275
rect 8346 222 8361 607
rect 8380 573 8415 607
rect 8380 222 8414 573
rect 8526 505 8584 511
rect 8526 471 8538 505
rect 8526 465 8584 471
rect 8526 305 8584 311
rect 8526 271 8538 305
rect 8526 265 8584 271
rect 6688 183 6694 193
rect 8380 188 8395 222
rect 6688 168 6722 183
rect 6711 140 6722 155
rect 270 59 286 81
rect 513 -1031 548 -997
rect 3927 -1031 3962 -997
rect 7341 -1031 7376 -997
rect 10755 -1031 10790 -997
rect 514 -1050 548 -1031
rect 3928 -1050 3962 -1031
rect 7342 -1050 7376 -1031
rect 10756 -1050 10790 -1031
rect 533 -1287 548 -1050
rect 567 -1084 602 -1050
rect 882 -1084 917 -1050
rect 567 -1287 601 -1084
rect 883 -1103 917 -1084
rect 713 -1152 771 -1146
rect 713 -1186 725 -1152
rect 713 -1192 771 -1186
rect 681 -1287 715 -1236
rect 769 -1287 803 -1236
rect 162 -1323 862 -1287
rect 0 -1357 862 -1323
rect 162 -1561 862 -1357
rect 531 -1614 862 -1561
rect 902 -1578 917 -1103
rect 936 -1137 971 -1103
rect 1251 -1137 1286 -1103
rect 936 -1578 970 -1137
rect 1252 -1156 1286 -1137
rect 1638 -1156 1691 -1155
rect 1054 -1231 1061 -1171
rect 1082 -1205 1140 -1199
rect 1082 -1239 1094 -1205
rect 1082 -1245 1140 -1239
rect 1082 -1495 1140 -1489
rect 1082 -1529 1094 -1495
rect 1082 -1535 1140 -1529
rect 936 -1612 951 -1578
rect 362 -1660 862 -1614
rect 1271 -1631 1286 -1156
rect 1305 -1190 1340 -1156
rect 1620 -1190 1691 -1156
rect 1305 -1631 1339 -1190
rect 1621 -1191 1691 -1190
rect 1638 -1225 1709 -1191
rect 1989 -1225 2024 -1191
rect 1451 -1258 1509 -1252
rect 1451 -1292 1463 -1258
rect 1451 -1298 1509 -1292
rect 1451 -1548 1509 -1542
rect 1451 -1582 1463 -1548
rect 1451 -1588 1509 -1582
rect 0 -1713 862 -1660
rect 1305 -1665 1320 -1631
rect -140 -1727 862 -1713
rect 1638 -1684 1708 -1225
rect 1990 -1244 2024 -1225
rect 1820 -1293 1878 -1287
rect 1820 -1327 1832 -1293
rect 1820 -1333 1878 -1327
rect 1820 -1601 1878 -1595
rect 1820 -1635 1832 -1601
rect 1820 -1641 1878 -1635
rect 1638 -1720 1691 -1684
rect 2009 -1702 2024 -1244
rect 1990 -1703 2024 -1702
rect 1705 -1720 2024 -1703
rect 2043 -1278 2078 -1244
rect 2358 -1278 2393 -1244
rect 2043 -1720 2077 -1278
rect 2359 -1297 2393 -1278
rect 3947 -1287 3962 -1050
rect 3981 -1084 4016 -1050
rect 4296 -1084 4331 -1050
rect 3981 -1287 4015 -1084
rect 4297 -1103 4331 -1084
rect 4127 -1152 4185 -1146
rect 4127 -1186 4139 -1152
rect 4127 -1192 4185 -1186
rect 4095 -1287 4129 -1236
rect 4183 -1287 4217 -1236
rect 3275 -1288 3421 -1287
rect 2189 -1346 2247 -1340
rect 2189 -1380 2201 -1346
rect 2189 -1386 2247 -1380
rect 2189 -1654 2247 -1648
rect 2189 -1667 2201 -1654
rect 2378 -1667 2393 -1297
rect 2412 -1331 2447 -1297
rect 2727 -1331 2762 -1297
rect 2412 -1667 2446 -1331
rect 2728 -1350 2762 -1331
rect 3274 -1323 3421 -1288
rect 3576 -1323 4276 -1287
rect 2530 -1431 2553 -1365
rect 2558 -1399 2616 -1393
rect 2558 -1433 2581 -1399
rect 2558 -1439 2616 -1433
rect 2747 -1614 2762 -1350
rect 2781 -1384 2816 -1350
rect 3096 -1384 3131 -1350
rect 3274 -1357 4276 -1323
rect 3274 -1367 3421 -1357
rect 2781 -1614 2815 -1384
rect 3097 -1403 3131 -1384
rect 2944 -1519 3051 -1505
rect 2916 -1545 2935 -1533
rect 2929 -1547 2935 -1545
rect 2977 -1547 3023 -1533
rect 3116 -1561 3131 -1403
rect 3150 -1437 3185 -1403
rect 3465 -1431 3500 -1403
rect 3257 -1437 3500 -1431
rect 3150 -1561 3184 -1437
rect 3323 -1485 3376 -1471
rect 3311 -1539 3376 -1485
rect 3432 -1485 3445 -1481
rect 3311 -1555 3358 -1539
rect 2830 -1586 3252 -1561
rect 3289 -1586 3298 -1582
rect 3311 -1586 3357 -1555
rect 3411 -1560 3420 -1548
rect 3377 -1586 3386 -1582
rect 2830 -1614 3270 -1586
rect 3289 -1598 3304 -1586
rect 2461 -1667 3270 -1614
rect 2092 -1720 3270 -1667
rect 3285 -1632 3304 -1598
rect 3317 -1598 3357 -1586
rect 3369 -1598 3398 -1586
rect 3317 -1632 3398 -1598
rect 3285 -1691 3298 -1632
rect 3323 -1653 3398 -1632
rect 3323 -1669 3332 -1653
rect 3289 -1693 3298 -1691
rect 3352 -1693 3398 -1653
rect 3411 -1653 3424 -1560
rect 3411 -1669 3420 -1653
rect 3432 -1665 3457 -1485
rect 3466 -1665 3500 -1437
rect 3576 -1456 4276 -1357
rect 3519 -1485 4276 -1456
rect 3511 -1490 4276 -1485
rect 3511 -1518 3554 -1490
rect 3576 -1518 4276 -1490
rect 3511 -1561 4276 -1518
rect 3511 -1653 3587 -1561
rect 3611 -1653 4276 -1561
rect 4316 -1578 4331 -1103
rect 4350 -1137 4385 -1103
rect 4665 -1137 4700 -1103
rect 4350 -1578 4384 -1137
rect 4666 -1156 4700 -1137
rect 5052 -1156 5105 -1155
rect 4468 -1231 4475 -1171
rect 4496 -1231 4503 -1199
rect 4518 -1431 4538 -1249
rect 4546 -1457 4566 -1277
rect 4496 -1495 4554 -1489
rect 4496 -1529 4508 -1495
rect 4496 -1535 4554 -1529
rect 4350 -1596 4365 -1578
rect 4350 -1597 4384 -1596
rect 4350 -1616 4446 -1597
rect 4350 -1631 4661 -1616
rect 4685 -1631 4700 -1156
rect 4719 -1190 4754 -1156
rect 5034 -1190 5105 -1156
rect 4719 -1631 4753 -1190
rect 5035 -1191 5105 -1190
rect 5052 -1225 5123 -1191
rect 5403 -1225 5438 -1191
rect 4865 -1258 4923 -1252
rect 4865 -1292 4877 -1258
rect 4865 -1298 4923 -1292
rect 4865 -1548 4923 -1542
rect 4865 -1582 4877 -1548
rect 4865 -1588 4923 -1582
rect 4719 -1649 4734 -1631
rect 4719 -1650 4753 -1649
rect 3511 -1665 3554 -1653
rect 3432 -1669 3445 -1665
rect 3289 -1703 3398 -1693
rect 1705 -1737 3270 -1720
rect 1723 -1766 3270 -1737
rect 3297 -1706 3398 -1703
rect 3466 -1680 3479 -1665
rect 3485 -1680 3500 -1665
rect 3297 -1740 3412 -1706
rect 3466 -1710 3500 -1680
rect 3466 -1721 3477 -1710
rect 3340 -1754 3412 -1740
rect 3340 -1766 3398 -1754
rect 1723 -1773 3252 -1766
rect 1723 -1790 1794 -1773
rect 1390 -1825 1425 -1791
rect 179 -1899 249 -1879
rect 616 -1897 693 -1861
rect 1021 -1878 1056 -1844
rect 103 -1914 249 -1899
rect 303 -1914 616 -1897
rect 103 -1950 317 -1914
rect 403 -1950 437 -1914
rect 491 -1950 525 -1914
rect 625 -1919 693 -1897
rect 726 -1898 850 -1897
rect 726 -1908 767 -1898
rect 839 -1908 850 -1898
rect 737 -1919 767 -1908
rect 625 -1950 794 -1919
rect 103 -1967 247 -1950
rect -122 -1975 111 -1967
rect -103 -2002 -102 -1975
rect -24 -1987 31 -1975
rect -103 -2003 -91 -2002
rect -24 -2003 -3 -1987
rect 43 -2003 111 -1975
rect 115 -2003 149 -1969
rect 249 -1984 633 -1950
rect 249 -2003 318 -1984
rect -103 -2037 44 -2003
rect 81 -2037 264 -2003
rect -125 -2103 -105 -2056
rect -103 -2064 -51 -2037
rect 43 -2058 111 -2037
rect 230 -2058 264 -2037
rect 43 -2059 264 -2058
rect 43 -2064 111 -2059
rect -103 -2065 111 -2064
rect -91 -2069 -52 -2065
rect -309 -2158 -251 -2152
rect -455 -2181 -421 -2163
rect -824 -2251 -789 -2217
rect -1047 -2372 -989 -2366
rect -1047 -2406 -1035 -2372
rect -1047 -2412 -989 -2406
rect -1047 -2572 -989 -2566
rect -1047 -2606 -1035 -2572
rect -1047 -2612 -989 -2606
rect -858 -2689 -843 -2270
rect -824 -2621 -790 -2251
rect -678 -2319 -620 -2313
rect -678 -2353 -666 -2319
rect -678 -2359 -620 -2353
rect -678 -2519 -620 -2513
rect -678 -2553 -666 -2519
rect -678 -2559 -620 -2553
rect -491 -2568 -421 -2181
rect -309 -2192 -297 -2158
rect -309 -2198 -251 -2192
rect -309 -2466 -251 -2460
rect -309 -2500 -297 -2466
rect -309 -2506 -251 -2500
rect -491 -2602 -420 -2568
rect -120 -2583 -105 -2103
rect -86 -2165 -52 -2069
rect 161 -2085 164 -2059
rect 249 -2087 264 -2059
rect 283 -2012 318 -2003
rect 283 -2065 351 -2012
rect 403 -2036 437 -1984
rect 491 -2014 525 -1984
rect 599 -2012 633 -1984
rect 403 -2047 449 -2036
rect 475 -2047 525 -2014
rect 565 -2046 633 -2012
rect 652 -1983 794 -1950
rect 652 -1987 809 -1983
rect 403 -2065 525 -2047
rect 579 -2065 647 -2046
rect 283 -2076 318 -2065
rect 410 -2076 513 -2065
rect 599 -2076 633 -2065
rect 283 -2077 633 -2076
rect 283 -2087 317 -2077
rect 399 -2083 475 -2077
rect 479 -2083 529 -2077
rect 399 -2086 529 -2083
rect 401 -2087 415 -2086
rect 239 -2108 317 -2087
rect 346 -2108 415 -2087
rect 425 -2087 443 -2086
rect 465 -2087 487 -2086
rect 425 -2092 487 -2087
rect 425 -2102 433 -2092
rect 249 -2115 264 -2108
rect 283 -2115 317 -2108
rect 493 -2115 515 -2086
rect 239 -2136 317 -2115
rect 346 -2120 515 -2115
rect 346 -2136 443 -2120
rect 473 -2133 523 -2127
rect 230 -2147 241 -2136
rect 249 -2147 264 -2136
rect -6 -2165 184 -2164
rect 230 -2165 264 -2147
rect 283 -2165 317 -2136
rect 385 -2147 400 -2136
rect 385 -2165 443 -2147
rect -86 -2177 443 -2165
rect 473 -2148 494 -2133
rect 522 -2148 531 -2133
rect 473 -2177 479 -2148
rect -86 -2191 431 -2177
rect 485 -2191 519 -2157
rect 599 -2165 633 -2077
rect 652 -2076 687 -1987
rect 691 -2076 720 -1987
rect 779 -2002 825 -1987
rect 794 -2026 825 -2002
rect 767 -2047 825 -2026
rect 844 -2033 847 -1999
rect 766 -2076 825 -2047
rect 652 -2077 825 -2076
rect 652 -2165 686 -2077
rect 691 -2081 720 -2077
rect 776 -2078 780 -2077
rect 754 -2092 782 -2080
rect 754 -2148 800 -2092
rect 766 -2157 800 -2148
rect 531 -2191 754 -2165
rect 766 -2191 804 -2157
rect -86 -2224 -51 -2191
rect -30 -2224 -18 -2191
rect -6 -2224 804 -2191
rect -86 -2225 804 -2224
rect -86 -2515 -52 -2225
rect 0 -2226 800 -2225
rect 28 -2354 62 -2226
rect 116 -2354 150 -2226
rect 32 -2400 146 -2379
rect 187 -2400 200 -2280
rect 60 -2428 118 -2407
rect 215 -2428 228 -2308
rect 60 -2447 72 -2428
rect 60 -2453 118 -2447
rect -86 -2549 -51 -2515
rect 249 -2530 264 -2226
rect 283 -2462 317 -2226
rect 387 -2308 391 -2285
rect 397 -2301 431 -2226
rect 485 -2301 519 -2226
rect 401 -2428 415 -2326
rect 429 -2360 487 -2354
rect 429 -2394 443 -2360
rect 429 -2400 487 -2394
rect 283 -2496 318 -2462
rect 618 -2477 633 -2226
rect 652 -2409 686 -2226
rect 766 -2248 800 -2226
rect 798 -2307 856 -2301
rect 798 -2341 810 -2307
rect 798 -2347 856 -2341
rect 652 -2443 687 -2409
rect 987 -2424 1002 -1897
rect 1021 -2356 1055 -1878
rect 1167 -1946 1225 -1940
rect 1167 -1980 1179 -1946
rect 1167 -1986 1225 -1980
rect 1167 -2254 1225 -2248
rect 1167 -2288 1179 -2254
rect 1167 -2294 1225 -2288
rect 1021 -2390 1056 -2356
rect 1356 -2371 1371 -1844
rect 1390 -2303 1424 -1825
rect 1536 -1893 1594 -1887
rect 1536 -1927 1548 -1893
rect 1536 -1933 1594 -1927
rect 1536 -2201 1594 -2195
rect 1536 -2235 1548 -2201
rect 1536 -2241 1594 -2235
rect 1723 -2250 1793 -1790
rect 2007 -1826 3252 -1773
rect 3340 -1779 3399 -1766
rect 3334 -1790 3399 -1779
rect 3308 -1824 3358 -1813
rect 1905 -1858 1963 -1852
rect 1905 -1892 1917 -1858
rect 1905 -1898 1963 -1892
rect 1905 -2148 1963 -2142
rect 1905 -2182 1917 -2148
rect 1905 -2188 1963 -2182
rect 1723 -2284 1794 -2250
rect 2094 -2265 2109 -1826
rect 2128 -2197 2162 -1826
rect 2274 -1839 2286 -1826
rect 2325 -1839 2332 -1826
rect 2353 -1831 2360 -1826
rect 2274 -1845 2332 -1839
rect 2376 -1879 3252 -1826
rect 3369 -1863 3399 -1790
rect 3485 -1804 3500 -1710
rect 3519 -1804 3553 -1665
rect 3633 -1684 4276 -1653
rect 4316 -1665 4394 -1650
rect 3633 -1704 4292 -1684
rect 4353 -1703 4543 -1670
rect 4719 -1684 4815 -1650
rect 5052 -1684 5122 -1225
rect 5404 -1244 5438 -1225
rect 5234 -1293 5292 -1287
rect 5234 -1327 5246 -1293
rect 5234 -1333 5292 -1327
rect 5234 -1601 5292 -1595
rect 5234 -1635 5246 -1601
rect 5234 -1641 5292 -1635
rect 5052 -1702 5105 -1684
rect 5052 -1703 5122 -1702
rect 4353 -1704 4667 -1703
rect 3633 -1727 4291 -1704
rect 4379 -1725 4394 -1704
rect 3633 -1744 3922 -1727
rect 3621 -1771 3922 -1744
rect 3991 -1769 4025 -1727
rect 4030 -1753 4120 -1727
rect 4151 -1733 4181 -1727
rect 4144 -1736 4181 -1733
rect 4204 -1736 4215 -1727
rect 4223 -1736 4238 -1727
rect 4034 -1759 4092 -1753
rect 3563 -1791 3587 -1775
rect 3599 -1791 3617 -1775
rect 3563 -1804 3591 -1791
rect 3474 -1811 3591 -1804
rect 3595 -1811 3617 -1791
rect 3621 -1778 3923 -1771
rect 3621 -1811 3922 -1778
rect 3968 -1781 4025 -1769
rect 4044 -1781 4078 -1759
rect 4105 -1781 4120 -1753
rect 3968 -1787 4120 -1781
rect 4186 -1746 4238 -1736
rect 4257 -1736 4291 -1727
rect 4186 -1752 4248 -1746
rect 4186 -1786 4252 -1752
rect 3968 -1803 4036 -1787
rect 4044 -1803 4078 -1787
rect 3449 -1879 3922 -1811
rect 3991 -1843 4078 -1803
rect 4090 -1791 4112 -1787
rect 4090 -1824 4136 -1791
rect 4186 -1792 4248 -1786
rect 4186 -1802 4238 -1792
rect 4204 -1814 4238 -1802
rect 4175 -1820 4238 -1814
rect 4257 -1801 4286 -1736
rect 4368 -1738 4394 -1725
rect 4257 -1802 4290 -1801
rect 4257 -1820 4291 -1802
rect 4365 -1816 4394 -1738
rect 4413 -1725 4448 -1704
rect 4413 -1737 4496 -1725
rect 4509 -1737 4667 -1704
rect 4685 -1718 4763 -1703
rect 4728 -1737 4763 -1718
rect 4413 -1765 4447 -1737
rect 4729 -1756 4763 -1737
rect 5052 -1737 5184 -1703
rect 5423 -1737 5438 -1244
rect 5457 -1278 5492 -1244
rect 5772 -1278 5807 -1244
rect 4413 -1772 4481 -1765
rect 4399 -1806 4447 -1772
rect 4449 -1806 4481 -1772
rect 4413 -1816 4447 -1806
rect 4165 -1824 4238 -1820
rect 4246 -1824 4291 -1820
rect 4338 -1822 4527 -1816
rect 4090 -1843 4112 -1824
rect 3990 -1869 4112 -1843
rect 4120 -1869 4136 -1824
rect 3990 -1875 4136 -1869
rect 2274 -2095 2332 -2089
rect 2274 -2129 2286 -2095
rect 2274 -2135 2332 -2129
rect 2128 -2231 2163 -2197
rect 2463 -2212 2478 -1879
rect 2497 -2144 2531 -1879
rect 2611 -1887 2645 -1879
rect 2699 -1887 2733 -1879
rect 2745 -1887 3252 -1879
rect 2552 -1907 3252 -1887
rect 3485 -1891 3554 -1879
rect 3627 -1887 3922 -1879
rect 3959 -1881 4136 -1875
rect 4146 -1881 4291 -1824
rect 4337 -1831 4527 -1822
rect 4531 -1831 4538 -1772
rect 4573 -1789 4584 -1778
rect 4596 -1789 4607 -1778
rect 4573 -1799 4607 -1789
rect 4559 -1805 4617 -1799
rect 4337 -1840 4394 -1831
rect 4337 -1844 4405 -1840
rect 4337 -1856 4411 -1844
rect 4413 -1856 4447 -1831
rect 4555 -1839 4571 -1805
rect 4573 -1839 4607 -1805
rect 4459 -1844 4481 -1840
rect 3959 -1885 4036 -1881
rect 4044 -1885 4078 -1881
rect 4090 -1885 4112 -1881
rect 3959 -1887 4078 -1885
rect 4124 -1887 4136 -1881
rect 4151 -1887 4291 -1881
rect 3627 -1891 4339 -1887
rect 3485 -1907 3500 -1891
rect 3517 -1906 3587 -1891
rect 3517 -1907 3563 -1906
rect 2552 -1923 3563 -1907
rect 3617 -1923 4339 -1891
rect 2552 -1957 4339 -1923
rect 2552 -1963 3563 -1957
rect 2552 -1968 3569 -1963
rect 3583 -1968 3597 -1963
rect 3617 -1968 4339 -1957
rect 2552 -1975 4339 -1968
rect 2497 -2178 2532 -2144
rect 2552 -2161 3252 -1975
rect 3289 -2032 3308 -1975
rect 3311 -2031 3312 -1975
rect 3317 -1995 3357 -1975
rect 3411 -1995 3445 -1975
rect 3317 -2031 3336 -1995
rect 3457 -2002 4339 -1975
rect 3457 -2031 3525 -2002
rect 3529 -2031 3569 -2002
rect 3583 -2031 3597 -2002
rect 3617 -2031 4339 -2002
rect 3311 -2064 3369 -2031
rect 3399 -2047 3429 -2031
rect 3432 -2047 4339 -2031
rect 3399 -2059 4339 -2047
rect 3399 -2064 3457 -2059
rect 3311 -2065 3457 -2064
rect 3323 -2069 3339 -2065
rect 3349 -2069 3357 -2065
rect 3411 -2069 3445 -2065
rect 3289 -2103 3305 -2081
rect 3383 -2085 3420 -2081
rect 3429 -2085 3441 -2069
rect 3495 -2070 3500 -2059
rect 3371 -2100 3432 -2085
rect 3460 -2097 3462 -2086
rect 3471 -2097 3479 -2081
rect 3495 -2085 3508 -2070
rect 3495 -2097 3514 -2085
rect 2552 -2214 2883 -2161
rect 3306 -2191 3317 -2137
rect 3371 -2147 3420 -2100
rect 3429 -2147 3432 -2100
rect 3471 -2132 3514 -2097
rect 3471 -2147 3520 -2132
rect 3371 -2157 3432 -2147
rect 3350 -2165 3432 -2157
rect 3334 -2177 3432 -2165
rect 3462 -2165 3520 -2147
rect 3526 -2165 3542 -2059
rect 3552 -2165 3566 -2059
rect 3583 -2081 3597 -2059
rect 3617 -2063 4339 -2059
rect 3583 -2085 3620 -2081
rect 3632 -2085 4339 -2063
rect 4360 -1922 4447 -1856
rect 4453 -1859 4505 -1844
rect 4559 -1845 4617 -1839
rect 4360 -1938 4405 -1922
rect 4413 -1938 4447 -1922
rect 4459 -1877 4505 -1859
rect 4539 -1877 4561 -1873
rect 4459 -1938 4481 -1877
rect 4489 -1922 4499 -1877
rect 4493 -1934 4499 -1922
rect 4515 -1934 4561 -1877
rect 4360 -1966 4447 -1938
rect 4521 -1960 4531 -1934
rect 4521 -1962 4527 -1960
rect 4360 -1972 4461 -1966
rect 4360 -2074 4394 -1972
rect 4399 -2006 4447 -1972
rect 4449 -2006 4481 -1972
rect 4403 -2012 4461 -2006
rect 4413 -2074 4447 -2012
rect 4539 -2020 4561 -1934
rect 4573 -2020 4607 -1845
rect 4515 -2057 4607 -2020
rect 4527 -2061 4561 -2057
rect 4573 -2074 4607 -2057
rect 4615 -2061 4641 -1873
rect 3574 -2100 3620 -2085
rect 3639 -2090 4339 -2085
rect 4353 -2089 4607 -2074
rect 4353 -2090 4617 -2089
rect 3639 -2095 4617 -2090
rect 3580 -2132 3594 -2100
rect 3574 -2147 3594 -2132
rect 3639 -2108 4511 -2095
rect 4555 -2097 4607 -2095
rect 4544 -2108 4607 -2097
rect 3574 -2165 3632 -2147
rect 3639 -2161 4339 -2108
rect 3462 -2177 3632 -2165
rect 3662 -2165 3720 -2161
rect 3780 -2165 3838 -2161
rect 3662 -2177 3735 -2165
rect 3334 -2191 3420 -2177
rect 3429 -2191 3432 -2177
rect 3471 -2191 3620 -2177
rect 3674 -2191 3735 -2177
rect 3765 -2177 3838 -2165
rect 3868 -2177 3914 -2161
rect 3962 -2171 3965 -2161
rect 3765 -2191 3826 -2177
rect 3880 -2191 3914 -2177
rect 3968 -2191 4002 -2161
rect 4008 -2191 4339 -2161
rect 4379 -2178 4394 -2108
rect 4413 -2178 4447 -2108
rect 4559 -2129 4571 -2108
rect 4559 -2135 4617 -2129
rect 3360 -2224 3542 -2191
rect 3552 -2214 4339 -2191
rect 4413 -2212 4428 -2178
rect 3552 -2224 4124 -2214
rect 4134 -2224 4218 -2214
rect 3360 -2225 4218 -2224
rect 3309 -2265 3311 -2232
rect 1390 -2337 1425 -2303
rect 1723 -2320 1776 -2284
rect 3337 -2293 3339 -2232
rect 3383 -2250 3420 -2225
rect 3429 -2250 3432 -2225
rect 3383 -2253 3432 -2250
rect 3471 -2253 3508 -2225
rect 3414 -2265 3432 -2253
rect 3355 -2310 3429 -2282
rect 3462 -2310 3536 -2282
rect 3552 -2293 3554 -2232
rect 3580 -2265 3582 -2232
rect 3586 -2253 3620 -2225
rect 3674 -2253 3708 -2225
rect 3792 -2253 3826 -2225
rect 3880 -2253 3914 -2225
rect 3968 -2253 4002 -2225
rect 4056 -2253 4090 -2225
rect 4168 -2253 4202 -2225
rect 4748 -2231 4763 -1756
rect 4782 -1790 4817 -1756
rect 5052 -1773 5168 -1737
rect 5097 -1790 5168 -1773
rect 5457 -1756 5491 -1278
rect 5773 -1297 5807 -1278
rect 7361 -1287 7376 -1050
rect 7395 -1084 7430 -1050
rect 7710 -1084 7745 -1050
rect 7395 -1287 7429 -1084
rect 7711 -1103 7745 -1084
rect 7541 -1152 7599 -1146
rect 7541 -1186 7553 -1152
rect 7541 -1192 7599 -1186
rect 7509 -1287 7543 -1236
rect 7597 -1287 7631 -1236
rect 6689 -1288 6835 -1287
rect 5603 -1346 5661 -1340
rect 5603 -1380 5615 -1346
rect 5603 -1386 5661 -1380
rect 5603 -1654 5661 -1648
rect 5603 -1688 5615 -1654
rect 5603 -1694 5661 -1688
rect 5457 -1790 5555 -1756
rect 5792 -1790 5807 -1297
rect 5826 -1331 5861 -1297
rect 6141 -1331 6176 -1297
rect 4782 -2231 4816 -1790
rect 5098 -1791 5168 -1790
rect 5115 -1825 5186 -1791
rect 5423 -1824 5501 -1791
rect 5466 -1825 5501 -1824
rect 4928 -1858 4986 -1852
rect 4928 -1892 4940 -1858
rect 4928 -1898 4986 -1892
rect 4928 -2148 4986 -2142
rect 4928 -2182 4940 -2148
rect 4928 -2188 4986 -2182
rect 4782 -2265 4797 -2231
rect 5115 -2284 5185 -1825
rect 5467 -1844 5501 -1825
rect 5826 -1809 5860 -1331
rect 6142 -1350 6176 -1331
rect 6688 -1323 6835 -1288
rect 6990 -1323 7690 -1287
rect 5972 -1399 6030 -1393
rect 5972 -1433 5984 -1399
rect 5972 -1439 6030 -1433
rect 5972 -1707 6030 -1701
rect 5972 -1741 5984 -1707
rect 5972 -1747 6030 -1741
rect 5826 -1843 5924 -1809
rect 6161 -1843 6176 -1350
rect 6195 -1384 6230 -1350
rect 6510 -1384 6545 -1350
rect 6688 -1357 7690 -1323
rect 6688 -1367 6835 -1357
rect 5297 -1893 5355 -1887
rect 5297 -1927 5309 -1893
rect 5297 -1933 5355 -1927
rect 5297 -2201 5355 -2195
rect 5297 -2235 5309 -2201
rect 5297 -2241 5355 -2235
rect 5115 -2320 5168 -2284
rect 3412 -2374 3441 -2340
rect 3450 -2374 3479 -2340
rect 3802 -2439 3829 -2321
rect 5486 -2337 5501 -1844
rect 5520 -1878 5555 -1844
rect 5792 -1877 5870 -1844
rect 5835 -1878 5870 -1877
rect 5520 -2337 5554 -1878
rect 5836 -1897 5870 -1878
rect 6195 -1862 6229 -1384
rect 6511 -1403 6545 -1384
rect 6341 -1452 6399 -1446
rect 6341 -1486 6353 -1452
rect 6341 -1492 6399 -1486
rect 6341 -1760 6399 -1754
rect 6341 -1794 6353 -1760
rect 6341 -1800 6399 -1794
rect 6195 -1896 6293 -1862
rect 6530 -1896 6545 -1403
rect 6564 -1437 6599 -1403
rect 6879 -1431 6914 -1403
rect 6671 -1437 6914 -1431
rect 5666 -1946 5724 -1940
rect 5666 -1980 5678 -1946
rect 5666 -1986 5724 -1980
rect 5666 -2254 5724 -2248
rect 5666 -2288 5678 -2254
rect 5666 -2294 5724 -2288
rect 3830 -2411 3857 -2349
rect 5520 -2371 5535 -2337
rect 5855 -2390 5870 -1897
rect 5889 -1931 5924 -1897
rect 6161 -1930 6239 -1897
rect 6204 -1931 6239 -1930
rect 5889 -2390 5923 -1931
rect 6205 -1950 6239 -1931
rect 6564 -1915 6598 -1437
rect 6737 -1485 6790 -1471
rect 6725 -1539 6790 -1485
rect 6846 -1485 6859 -1481
rect 6725 -1555 6772 -1539
rect 6703 -1586 6712 -1582
rect 6725 -1586 6771 -1555
rect 6825 -1558 6834 -1548
rect 6819 -1560 6834 -1558
rect 6791 -1586 6800 -1582
rect 6703 -1598 6718 -1586
rect 6699 -1632 6718 -1598
rect 6731 -1598 6771 -1586
rect 6783 -1598 6812 -1586
rect 6731 -1632 6812 -1598
rect 6819 -1632 6838 -1560
rect 6699 -1691 6712 -1632
rect 6737 -1653 6812 -1632
rect 6737 -1669 6746 -1653
rect 6703 -1693 6712 -1691
rect 6766 -1693 6812 -1653
rect 6825 -1653 6838 -1632
rect 6825 -1669 6834 -1653
rect 6846 -1665 6871 -1485
rect 6880 -1665 6914 -1437
rect 6990 -1456 7690 -1357
rect 6933 -1485 7690 -1456
rect 6925 -1490 7690 -1485
rect 6925 -1518 6968 -1490
rect 6990 -1518 7690 -1490
rect 6925 -1561 7690 -1518
rect 6925 -1653 7001 -1561
rect 7025 -1619 7059 -1561
rect 7060 -1611 7071 -1561
rect 7075 -1592 7177 -1561
rect 7131 -1608 7141 -1592
rect 7143 -1608 7177 -1592
rect 7131 -1611 7177 -1608
rect 7060 -1619 7177 -1611
rect 7025 -1625 7177 -1619
rect 7025 -1639 7081 -1625
rect 7131 -1639 7177 -1625
rect 7025 -1653 7093 -1639
rect 7129 -1653 7177 -1639
rect 7231 -1581 7299 -1561
rect 7359 -1581 7690 -1561
rect 7730 -1578 7745 -1103
rect 7764 -1137 7799 -1103
rect 8079 -1137 8114 -1103
rect 7764 -1578 7798 -1137
rect 8080 -1156 8114 -1137
rect 8466 -1156 8519 -1155
rect 7882 -1231 7889 -1171
rect 7910 -1205 7968 -1199
rect 7910 -1239 7922 -1205
rect 7910 -1245 7968 -1239
rect 7910 -1495 7968 -1489
rect 7910 -1529 7922 -1495
rect 7910 -1535 7968 -1529
rect 7231 -1614 7690 -1581
rect 7764 -1612 7779 -1578
rect 7231 -1634 7688 -1614
rect 7764 -1631 8075 -1616
rect 8099 -1631 8114 -1156
rect 8133 -1190 8168 -1156
rect 8448 -1190 8519 -1156
rect 8133 -1631 8167 -1190
rect 8449 -1191 8519 -1190
rect 8466 -1225 8537 -1191
rect 8817 -1225 8852 -1191
rect 8279 -1258 8337 -1252
rect 8279 -1292 8291 -1258
rect 8279 -1298 8337 -1292
rect 8279 -1548 8337 -1542
rect 8279 -1582 8291 -1548
rect 8279 -1588 8337 -1582
rect 7231 -1653 7690 -1634
rect 6925 -1665 6968 -1653
rect 7047 -1661 7093 -1653
rect 7047 -1665 7081 -1661
rect 7086 -1665 7093 -1661
rect 6846 -1669 6859 -1665
rect 6703 -1703 6812 -1693
rect 6711 -1706 6812 -1703
rect 6880 -1680 6893 -1665
rect 6899 -1680 6914 -1665
rect 6711 -1740 6826 -1706
rect 6880 -1710 6914 -1680
rect 6880 -1721 6891 -1710
rect 6754 -1754 6826 -1740
rect 6754 -1766 6812 -1754
rect 6754 -1779 6813 -1766
rect 6748 -1790 6813 -1779
rect 6722 -1824 6772 -1813
rect 6783 -1863 6813 -1790
rect 6899 -1811 6914 -1710
rect 6933 -1811 6967 -1665
rect 7047 -1744 7093 -1665
rect 7035 -1753 7093 -1744
rect 7099 -1721 7115 -1693
rect 7135 -1714 7169 -1653
rect 7249 -1665 7690 -1653
rect 8133 -1665 8148 -1631
rect 7174 -1714 7181 -1665
rect 7266 -1670 7690 -1665
rect 7266 -1704 7706 -1670
rect 8466 -1684 8536 -1225
rect 8818 -1244 8852 -1225
rect 8648 -1293 8706 -1287
rect 8648 -1327 8660 -1293
rect 8648 -1333 8706 -1327
rect 8648 -1601 8706 -1595
rect 8648 -1635 8660 -1601
rect 8648 -1641 8706 -1635
rect 7266 -1711 7705 -1704
rect 7135 -1721 7181 -1714
rect 7099 -1753 7127 -1721
rect 7129 -1745 7181 -1721
rect 7249 -1727 7705 -1711
rect 8466 -1720 8519 -1684
rect 7249 -1733 7319 -1727
rect 7325 -1733 7336 -1727
rect 7129 -1753 7203 -1745
rect 6977 -1791 7001 -1775
rect 7013 -1791 7031 -1775
rect 6977 -1811 7005 -1791
rect 7009 -1811 7031 -1791
rect 7035 -1790 7081 -1753
rect 7086 -1790 7093 -1753
rect 7035 -1811 7093 -1790
rect 7135 -1761 7203 -1753
rect 7215 -1761 7235 -1745
rect 7135 -1795 7235 -1761
rect 7135 -1805 7203 -1795
rect 6863 -1820 7093 -1811
rect 6863 -1866 7075 -1820
rect 7099 -1839 7127 -1805
rect 7129 -1811 7203 -1805
rect 7215 -1811 7235 -1795
rect 7129 -1819 7181 -1811
rect 7147 -1823 7169 -1819
rect 7249 -1829 7336 -1733
rect 7448 -1753 7460 -1727
rect 7491 -1753 7506 -1727
rect 7448 -1759 7506 -1753
rect 7519 -1781 7534 -1727
rect 7420 -1787 7534 -1781
rect 7637 -1801 7652 -1727
rect 7618 -1814 7652 -1801
rect 7141 -1839 7336 -1829
rect 7099 -1845 7336 -1839
rect 7589 -1832 7652 -1814
rect 7671 -1832 7705 -1727
rect 8837 -1737 8852 -1244
rect 8871 -1278 8906 -1244
rect 9186 -1278 9221 -1244
rect 8871 -1737 8905 -1278
rect 9187 -1297 9221 -1278
rect 10775 -1287 10790 -1050
rect 10809 -1084 10844 -1050
rect 11124 -1084 11159 -1050
rect 10809 -1287 10843 -1084
rect 11125 -1103 11159 -1084
rect 10955 -1152 11013 -1146
rect 10955 -1186 10967 -1152
rect 10955 -1192 11013 -1186
rect 10923 -1287 10957 -1236
rect 11011 -1287 11045 -1236
rect 10103 -1288 10249 -1287
rect 9017 -1346 9075 -1340
rect 9017 -1380 9029 -1346
rect 9017 -1386 9075 -1380
rect 9017 -1654 9075 -1648
rect 9017 -1688 9029 -1654
rect 9017 -1694 9075 -1688
rect 7817 -1772 7875 -1766
rect 8871 -1771 8886 -1737
rect 7817 -1806 7829 -1772
rect 9206 -1790 9221 -1297
rect 9240 -1331 9275 -1297
rect 9555 -1331 9590 -1297
rect 9240 -1790 9274 -1331
rect 9556 -1350 9590 -1331
rect 10102 -1323 10249 -1288
rect 10404 -1323 11104 -1287
rect 9386 -1399 9444 -1393
rect 9386 -1433 9398 -1399
rect 9386 -1439 9444 -1433
rect 9386 -1707 9444 -1701
rect 9386 -1741 9398 -1707
rect 9386 -1747 9444 -1741
rect 7817 -1812 7875 -1806
rect 9240 -1824 9255 -1790
rect 7099 -1847 7249 -1845
rect 7079 -1866 7099 -1860
rect 7141 -1866 7249 -1847
rect 6863 -1879 7103 -1866
rect 7109 -1871 7249 -1866
rect 6899 -1891 6968 -1879
rect 7041 -1880 7103 -1879
rect 7105 -1875 7249 -1871
rect 7266 -1875 7336 -1845
rect 7105 -1880 7336 -1875
rect 6899 -1907 6914 -1891
rect 6931 -1906 7001 -1891
rect 7041 -1894 7336 -1880
rect 7404 -1869 7504 -1843
rect 7589 -1848 7667 -1832
rect 7671 -1848 7704 -1832
rect 9575 -1843 9590 -1350
rect 9609 -1384 9644 -1350
rect 9924 -1384 9959 -1350
rect 10102 -1357 11104 -1323
rect 10102 -1367 10249 -1357
rect 9609 -1843 9643 -1384
rect 9925 -1403 9959 -1384
rect 9755 -1452 9813 -1446
rect 9755 -1486 9767 -1452
rect 9755 -1492 9813 -1486
rect 9755 -1760 9813 -1754
rect 9755 -1794 9767 -1760
rect 9755 -1800 9813 -1794
rect 7404 -1881 7507 -1869
rect 7416 -1885 7450 -1881
rect 7618 -1882 7704 -1848
rect 9609 -1877 9624 -1843
rect 6931 -1907 6968 -1906
rect 6657 -1915 6968 -1907
rect 6564 -1949 6968 -1915
rect 7041 -1908 7071 -1894
rect 7075 -1897 7336 -1894
rect 7407 -1897 7441 -1893
rect 7075 -1900 7175 -1897
rect 7075 -1908 7077 -1900
rect 7079 -1906 7175 -1900
rect 7131 -1908 7175 -1906
rect 7041 -1912 7175 -1908
rect 7249 -1909 7336 -1897
rect 7401 -1909 7453 -1897
rect 7041 -1916 7141 -1912
rect 7143 -1916 7175 -1912
rect 7041 -1934 7175 -1916
rect 6035 -1999 6093 -1993
rect 6035 -2033 6047 -1999
rect 6035 -2039 6093 -2033
rect 6035 -2307 6093 -2301
rect 6035 -2341 6047 -2307
rect 6035 -2347 6093 -2341
rect 5889 -2424 5904 -2390
rect 6224 -2443 6239 -1950
rect 6258 -1984 6293 -1950
rect 6530 -1983 6608 -1950
rect 6657 -1968 6967 -1949
rect 7031 -1968 7065 -1934
rect 7077 -1968 7177 -1934
rect 7231 -1968 7353 -1909
rect 7407 -1919 7453 -1909
rect 6657 -1975 7077 -1968
rect 6573 -1984 6608 -1983
rect 6258 -2443 6292 -1984
rect 6574 -2003 6608 -1984
rect 6725 -2003 6726 -1975
rect 6737 -2003 6771 -1975
rect 6825 -2003 6859 -1975
rect 6871 -2002 7077 -1975
rect 7109 -2002 7353 -1968
rect 7410 -1969 7441 -1919
rect 7444 -1949 7479 -1919
rect 7491 -1926 7506 -1913
rect 7488 -1949 7506 -1926
rect 7444 -1953 7510 -1949
rect 7444 -1969 7453 -1953
rect 7488 -1959 7506 -1953
rect 7519 -1954 7534 -1885
rect 7618 -1898 7667 -1882
rect 7671 -1898 7701 -1882
rect 9944 -1896 9959 -1403
rect 9978 -1437 10013 -1403
rect 10293 -1431 10328 -1403
rect 10085 -1437 10328 -1431
rect 9978 -1896 10012 -1437
rect 10151 -1485 10204 -1471
rect 10139 -1539 10204 -1485
rect 10260 -1485 10273 -1481
rect 10139 -1555 10186 -1539
rect 10117 -1586 10126 -1582
rect 10139 -1586 10185 -1555
rect 10239 -1558 10248 -1548
rect 10233 -1560 10248 -1558
rect 10205 -1586 10214 -1582
rect 10117 -1598 10132 -1586
rect 10113 -1632 10132 -1598
rect 10145 -1598 10185 -1586
rect 10197 -1598 10226 -1586
rect 10145 -1632 10226 -1598
rect 10233 -1632 10252 -1560
rect 10113 -1691 10126 -1632
rect 10151 -1653 10226 -1632
rect 10151 -1669 10160 -1653
rect 10117 -1693 10126 -1691
rect 10180 -1693 10226 -1653
rect 10239 -1653 10252 -1632
rect 10239 -1669 10248 -1653
rect 10260 -1665 10285 -1485
rect 10294 -1665 10328 -1437
rect 10404 -1456 11104 -1357
rect 10347 -1485 11104 -1456
rect 10339 -1490 11104 -1485
rect 10339 -1518 10382 -1490
rect 10404 -1518 11104 -1490
rect 10339 -1561 11104 -1518
rect 10339 -1653 10415 -1561
rect 10439 -1619 10473 -1561
rect 10474 -1611 10485 -1561
rect 10489 -1592 10591 -1561
rect 10545 -1608 10555 -1592
rect 10557 -1608 10591 -1592
rect 10545 -1611 10591 -1608
rect 10474 -1619 10591 -1611
rect 10439 -1625 10591 -1619
rect 10439 -1639 10495 -1625
rect 10545 -1639 10591 -1625
rect 10439 -1653 10507 -1639
rect 10543 -1653 10591 -1639
rect 10645 -1581 10713 -1561
rect 10773 -1581 11104 -1561
rect 11144 -1578 11159 -1103
rect 11178 -1137 11213 -1103
rect 11493 -1137 11528 -1103
rect 11178 -1578 11212 -1137
rect 11494 -1156 11528 -1137
rect 11880 -1156 11933 -1155
rect 11296 -1231 11303 -1171
rect 11324 -1205 11382 -1199
rect 11324 -1239 11336 -1205
rect 11324 -1245 11382 -1239
rect 11324 -1495 11382 -1489
rect 11324 -1529 11336 -1495
rect 11324 -1535 11382 -1529
rect 10645 -1614 11104 -1581
rect 11178 -1612 11193 -1578
rect 10645 -1634 11102 -1614
rect 11178 -1631 11489 -1616
rect 11513 -1631 11528 -1156
rect 11547 -1190 11582 -1156
rect 11862 -1190 11933 -1156
rect 11547 -1631 11581 -1190
rect 11863 -1191 11933 -1190
rect 11880 -1225 11951 -1191
rect 12231 -1225 12266 -1191
rect 11693 -1258 11751 -1252
rect 11693 -1292 11705 -1258
rect 11693 -1298 11751 -1292
rect 11693 -1548 11751 -1542
rect 11693 -1582 11705 -1548
rect 11693 -1588 11751 -1582
rect 10645 -1653 11104 -1634
rect 10339 -1665 10382 -1653
rect 10461 -1661 10507 -1653
rect 10461 -1665 10495 -1661
rect 10500 -1665 10507 -1661
rect 10260 -1669 10273 -1665
rect 10117 -1703 10226 -1693
rect 10125 -1706 10226 -1703
rect 10294 -1680 10307 -1665
rect 10313 -1680 10328 -1665
rect 10125 -1740 10240 -1706
rect 10294 -1710 10328 -1680
rect 10294 -1721 10305 -1710
rect 10168 -1754 10240 -1740
rect 10168 -1766 10226 -1754
rect 10168 -1779 10227 -1766
rect 10162 -1790 10227 -1779
rect 10136 -1824 10186 -1813
rect 10197 -1863 10227 -1790
rect 10313 -1811 10328 -1710
rect 10347 -1811 10381 -1665
rect 10461 -1744 10507 -1665
rect 10449 -1753 10507 -1744
rect 10513 -1721 10529 -1693
rect 10549 -1714 10583 -1653
rect 10663 -1665 11104 -1653
rect 11547 -1665 11562 -1631
rect 10588 -1714 10595 -1665
rect 10680 -1670 11104 -1665
rect 10680 -1704 11120 -1670
rect 11880 -1684 11950 -1225
rect 12232 -1244 12266 -1225
rect 12062 -1293 12120 -1287
rect 12062 -1327 12074 -1293
rect 12062 -1333 12120 -1327
rect 12062 -1601 12120 -1595
rect 12062 -1635 12074 -1601
rect 12062 -1641 12120 -1635
rect 10680 -1711 11119 -1704
rect 10549 -1721 10595 -1714
rect 10513 -1753 10541 -1721
rect 10543 -1745 10595 -1721
rect 10663 -1727 11119 -1711
rect 11880 -1720 11933 -1684
rect 10663 -1733 10733 -1727
rect 10739 -1733 10750 -1727
rect 10543 -1753 10617 -1745
rect 10391 -1791 10415 -1775
rect 10427 -1791 10445 -1775
rect 10391 -1811 10419 -1791
rect 10423 -1811 10445 -1791
rect 10449 -1790 10495 -1753
rect 10500 -1790 10507 -1753
rect 10449 -1811 10507 -1790
rect 10549 -1761 10617 -1753
rect 10629 -1761 10649 -1745
rect 10549 -1795 10649 -1761
rect 10549 -1805 10617 -1795
rect 10277 -1820 10507 -1811
rect 10277 -1866 10489 -1820
rect 10513 -1839 10541 -1805
rect 10543 -1811 10617 -1805
rect 10629 -1811 10649 -1795
rect 10543 -1819 10595 -1811
rect 10561 -1823 10583 -1819
rect 10663 -1829 10750 -1733
rect 10862 -1753 10874 -1727
rect 10905 -1753 10920 -1727
rect 10862 -1759 10920 -1753
rect 10933 -1781 10948 -1727
rect 10834 -1787 10948 -1781
rect 11051 -1801 11066 -1727
rect 11032 -1814 11066 -1801
rect 10555 -1839 10750 -1829
rect 10513 -1845 10750 -1839
rect 11003 -1832 11066 -1814
rect 11085 -1832 11119 -1727
rect 12251 -1737 12266 -1244
rect 12285 -1278 12320 -1244
rect 12600 -1278 12635 -1244
rect 12285 -1737 12319 -1278
rect 12601 -1297 12635 -1278
rect 12431 -1346 12489 -1340
rect 12431 -1380 12443 -1346
rect 12431 -1386 12489 -1380
rect 12431 -1654 12489 -1648
rect 12431 -1688 12443 -1654
rect 12431 -1694 12489 -1688
rect 11231 -1772 11289 -1766
rect 12285 -1771 12300 -1737
rect 11231 -1806 11243 -1772
rect 12620 -1790 12635 -1297
rect 12654 -1331 12689 -1297
rect 12969 -1331 13004 -1297
rect 12654 -1790 12688 -1331
rect 12970 -1350 13004 -1331
rect 12800 -1399 12858 -1393
rect 12800 -1433 12812 -1399
rect 12800 -1439 12858 -1433
rect 12800 -1707 12858 -1701
rect 12800 -1741 12812 -1707
rect 12800 -1747 12858 -1741
rect 11231 -1812 11289 -1806
rect 12654 -1824 12669 -1790
rect 10513 -1847 10663 -1845
rect 10493 -1866 10513 -1860
rect 10555 -1866 10663 -1847
rect 10277 -1879 10517 -1866
rect 10523 -1871 10663 -1866
rect 10313 -1891 10382 -1879
rect 10455 -1880 10517 -1879
rect 10519 -1875 10663 -1871
rect 10680 -1875 10750 -1845
rect 10519 -1880 10750 -1875
rect 7618 -1909 7629 -1898
rect 7637 -1933 7652 -1898
rect 7410 -1984 7453 -1969
rect 7516 -1983 7534 -1954
rect 7410 -1987 7441 -1984
rect 7516 -1987 7544 -1983
rect 7618 -1987 7652 -1933
rect 6871 -2003 6939 -2002
rect 6404 -2052 6462 -2046
rect 6404 -2086 6416 -2052
rect 6404 -2092 6462 -2086
rect 6404 -2360 6462 -2354
rect 6404 -2394 6416 -2360
rect 6404 -2400 6462 -2394
rect 6258 -2477 6273 -2443
rect 6593 -2496 6608 -2003
rect 6627 -2037 6662 -2003
rect 6723 -2037 6871 -2003
rect 6881 -2037 6893 -2003
rect 6899 -2036 6977 -2003
rect 7077 -2022 7145 -2002
rect 6931 -2037 6977 -2036
rect 6627 -2496 6661 -2037
rect 6725 -2064 6726 -2037
rect 6871 -2058 6939 -2037
rect 6943 -2058 6977 -2037
rect 7058 -2047 7065 -2022
rect 7077 -2056 7177 -2022
rect 7231 -2056 7265 -2002
rect 7266 -2020 7353 -2002
rect 7266 -2021 7382 -2020
rect 7407 -2021 7441 -1987
rect 7519 -2021 7553 -1987
rect 7618 -2021 7653 -1987
rect 7266 -2055 7453 -2021
rect 7485 -2055 7653 -2021
rect 7266 -2056 7382 -2055
rect 6996 -2058 7077 -2056
rect 6871 -2059 7077 -2058
rect 6871 -2064 6939 -2059
rect 6725 -2065 6939 -2064
rect 6943 -2147 6954 -2136
rect 6962 -2147 6977 -2059
rect 6795 -2165 6897 -2164
rect 6943 -2165 6977 -2147
rect 6996 -2090 7031 -2059
rect 7131 -2077 7382 -2056
rect 7189 -2079 7219 -2077
rect 7178 -2087 7230 -2079
rect 6996 -2165 7030 -2090
rect 7067 -2108 7144 -2087
rect 7174 -2108 7243 -2087
rect 7266 -2091 7382 -2077
rect 7637 -2081 7641 -2055
rect 7646 -2077 7653 -2055
rect 7671 -2074 7705 -1898
rect 9978 -1930 9993 -1896
rect 10313 -1907 10328 -1891
rect 10345 -1906 10415 -1891
rect 10455 -1894 10750 -1880
rect 10818 -1869 10918 -1843
rect 11003 -1848 11081 -1832
rect 11085 -1848 11118 -1832
rect 12989 -1843 13004 -1350
rect 13023 -1384 13058 -1350
rect 13338 -1384 13373 -1350
rect 13023 -1843 13057 -1384
rect 13339 -1403 13373 -1384
rect 13169 -1452 13227 -1446
rect 13169 -1486 13181 -1452
rect 13169 -1492 13227 -1486
rect 13169 -1760 13227 -1754
rect 13169 -1794 13181 -1760
rect 13169 -1800 13227 -1794
rect 10818 -1881 10921 -1869
rect 10830 -1885 10864 -1881
rect 11032 -1882 11118 -1848
rect 13023 -1877 13038 -1843
rect 10345 -1907 10382 -1906
rect 10071 -1949 10382 -1907
rect 10455 -1908 10485 -1894
rect 10489 -1897 10750 -1894
rect 10821 -1897 10855 -1893
rect 10489 -1900 10589 -1897
rect 10489 -1908 10491 -1900
rect 10493 -1906 10589 -1900
rect 10545 -1908 10589 -1906
rect 10455 -1912 10589 -1908
rect 10455 -1916 10555 -1912
rect 10557 -1916 10589 -1912
rect 10455 -1934 10589 -1916
rect 10663 -1909 10750 -1897
rect 10815 -1909 10867 -1897
rect 7817 -1972 7875 -1966
rect 10071 -1968 10381 -1949
rect 10445 -1968 10479 -1934
rect 10491 -1968 10591 -1934
rect 10663 -1968 10767 -1909
rect 10821 -1919 10867 -1909
rect 7817 -2006 7829 -1972
rect 10071 -1975 10491 -1968
rect 10139 -1985 10140 -1975
rect 10151 -1983 10185 -1975
rect 10239 -1983 10273 -1975
rect 10285 -1985 10491 -1975
rect 10311 -2002 10491 -1985
rect 10523 -2002 10767 -1968
rect 10824 -1969 10855 -1919
rect 10858 -1949 10893 -1919
rect 10905 -1926 10920 -1913
rect 10902 -1949 10920 -1926
rect 10858 -1953 10924 -1949
rect 10858 -1969 10867 -1953
rect 10902 -1959 10920 -1953
rect 10933 -1954 10948 -1885
rect 11032 -1898 11081 -1882
rect 11085 -1898 11115 -1882
rect 13358 -1896 13373 -1403
rect 11032 -1909 11043 -1898
rect 11051 -1933 11066 -1898
rect 10824 -1984 10867 -1969
rect 10930 -1983 10948 -1954
rect 10824 -1987 10855 -1984
rect 10930 -1987 10958 -1983
rect 11032 -1987 11066 -1933
rect 7817 -2012 7875 -2006
rect 10311 -2038 10353 -2002
rect 10491 -2038 10559 -2002
rect 10680 -2021 10767 -2002
rect 10821 -2021 10855 -1987
rect 10933 -2021 10967 -1987
rect 11032 -2021 11067 -1987
rect 10680 -2038 10867 -2021
rect 10716 -2055 10867 -2038
rect 10899 -2055 11067 -2021
rect 10733 -2065 10767 -2055
rect 7671 -2077 7707 -2074
rect 7671 -2089 7686 -2077
rect 11051 -2081 11055 -2055
rect 11060 -2077 11067 -2055
rect 11085 -2074 11119 -1898
rect 11231 -1972 11289 -1966
rect 11231 -2006 11243 -1972
rect 11231 -2012 11289 -2006
rect 14094 -2038 14147 -1581
rect 11085 -2077 11121 -2074
rect 7067 -2124 7144 -2115
rect 7174 -2124 7271 -2115
rect 7067 -2136 7271 -2124
rect 7114 -2143 7228 -2136
rect 6768 -2191 6787 -2186
rect 6795 -2191 7138 -2165
rect 7142 -2171 7200 -2152
rect 7312 -2157 7318 -2091
rect 7671 -2108 7675 -2089
rect 10481 -2108 10558 -2087
rect 10588 -2108 10657 -2087
rect 11085 -2089 11100 -2077
rect 11085 -2108 11089 -2089
rect 10481 -2136 10558 -2115
rect 10588 -2136 10685 -2115
rect 7312 -2165 7346 -2157
rect 7204 -2191 7382 -2165
rect 6741 -2198 6773 -2192
rect 6774 -2198 6897 -2191
rect 6909 -2198 7598 -2191
rect 6741 -2226 7623 -2198
rect 6741 -2354 6775 -2226
rect 6829 -2354 6863 -2226
rect 6773 -2413 6831 -2407
rect 6773 -2447 6785 -2413
rect 6773 -2453 6831 -2447
rect 6627 -2530 6642 -2496
rect 6962 -2549 6977 -2226
rect 6996 -2549 7030 -2226
rect 7076 -2232 7266 -2226
rect 7110 -2239 7144 -2235
rect 7198 -2239 7232 -2235
rect 7104 -2260 7150 -2239
rect 7192 -2260 7238 -2239
rect 7329 -2251 7400 -2226
rect 7461 -2251 7619 -2226
rect 7680 -2251 7715 -2217
rect 7110 -2264 7144 -2260
rect 7198 -2264 7232 -2260
rect 3414 -2587 3432 -2575
rect 3460 -2587 3462 -2576
rect 6996 -2583 7011 -2549
rect 3383 -2590 3432 -2587
rect -824 -2655 -789 -2621
rect -491 -2638 -438 -2602
rect 3383 -2650 3420 -2590
rect 3429 -2650 3432 -2590
rect 3383 -2653 3432 -2650
rect 3471 -2653 3508 -2587
rect 7329 -2602 7399 -2251
rect 7681 -2270 7715 -2251
rect 7511 -2319 7569 -2313
rect 7511 -2353 7523 -2319
rect 7511 -2359 7569 -2353
rect 7511 -2519 7569 -2513
rect 7511 -2553 7523 -2519
rect 7511 -2559 7569 -2553
rect 7329 -2638 7382 -2602
rect 3414 -2665 3432 -2653
rect 7700 -2655 7715 -2270
rect 7734 -2304 7769 -2270
rect 7734 -2655 7768 -2304
rect 7880 -2372 7938 -2366
rect 7880 -2406 7892 -2372
rect 7880 -2412 7938 -2406
rect 7880 -2572 7938 -2566
rect 7880 -2606 7892 -2572
rect 7880 -2612 7938 -2606
rect 187 -2800 200 -2680
rect 2999 -2708 3068 -2687
rect 3098 -2708 3175 -2687
rect 3829 -2708 3892 -2687
rect 7734 -2689 7749 -2655
rect 215 -2828 228 -2708
rect 2971 -2736 3068 -2715
rect 3098 -2736 3175 -2715
rect 3829 -2736 3920 -2715
rect 2619 -2826 4272 -2791
rect 187 -3200 200 -3080
rect 215 -3228 228 -3108
rect 187 -3600 200 -3480
rect 215 -3628 228 -3508
rect 187 -4000 200 -3880
rect 215 -4028 228 -3908
<< nwell >>
rect 3414 1135 3477 1539
rect 2907 989 2908 991
rect 3983 989 3984 991
rect 3414 441 3485 845
<< poly >>
rect 1604 1863 1813 1893
rect 1782 1821 1813 1863
rect 5079 1863 5321 1893
rect 5079 1821 5109 1863
rect 1782 827 1812 1153
rect 5079 827 5109 1153
<< metal1 >>
rect 1876 1947 4986 1980
rect 2907 1935 3984 1947
rect 1546 1834 1556 1886
rect 1608 1834 1618 1886
rect 3414 1876 3478 1935
rect 6891 1921 6948 1980
rect 5253 1834 5263 1886
rect 5315 1834 5325 1886
rect 3326 1529 3414 1663
rect 3497 1533 3507 1585
rect 3559 1533 3569 1585
rect 2849 1417 2859 1469
rect 2911 1417 2921 1469
rect 4003 1433 4013 1485
rect 4065 1433 4075 1485
rect 3414 1135 3483 1255
rect -56 909 0 1071
rect 3414 725 3477 845
rect 1812 385 1878 443
rect 2894 426 2922 534
rect 3970 487 3980 539
rect 4032 487 4042 539
rect 3467 419 3477 471
rect 3529 419 3539 471
rect 3364 303 3416 336
rect 3344 251 3354 303
rect 3406 251 3416 303
rect 0 0 200 200
rect 3414 47 3477 104
rect 6920 59 6948 1921
rect 1906 0 5172 47
rect 6891 0 6948 59
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
<< via1 >>
rect 1556 1834 1608 1886
rect 5263 1834 5315 1886
rect 3507 1533 3559 1585
rect 2859 1417 2911 1469
rect 4013 1433 4065 1485
rect 3980 487 4032 539
rect 3477 419 3529 471
rect 3354 251 3406 303
<< metal2 >>
rect 1556 1886 1608 1896
rect 5263 1886 5315 1896
rect 1608 1834 5263 1852
rect 1556 1824 5315 1834
rect 659 1556 721 1628
rect 3507 1585 3559 1595
rect 6170 1556 6232 1628
rect 3507 1523 3559 1533
rect 3529 1479 3557 1523
rect 2859 1469 3557 1479
rect 2911 1451 3557 1469
rect 4013 1485 4066 1495
rect 4065 1433 4066 1485
rect 4013 1423 4066 1433
rect 2859 1407 2911 1417
rect 316 577 344 1405
rect 4038 605 4066 1423
rect 3501 577 4066 605
rect 291 523 363 577
rect 316 122 344 523
rect 3501 481 3529 577
rect 6547 575 6575 1405
rect 3980 539 4032 549
rect 3477 471 3529 481
rect 659 349 721 424
rect 3477 409 3529 419
rect 3853 487 3980 508
rect 3853 480 4032 487
rect 3853 313 3881 480
rect 3980 477 4032 480
rect 6170 352 6232 424
rect 3354 303 3881 313
rect 3406 285 3881 303
rect 3354 241 3406 251
rect 6547 122 6575 572
rect 316 94 6575 122
use contacto  contacto_0
timestamp 1616018980
transform 1 0 1558 0 1 1830
box 0 4 66 62
use contacto  contacto_1
timestamp 1616018980
transform 1 0 5263 0 1 1830
box 0 4 66 62
use contador1bit  contador1bit_1
timestamp 1624053917
transform 1 0 3337 0 1 -32
box -1604 -4676 5429 1783
use contador1bit  contador1bit_0
timestamp 1624053917
transform -1 0 3554 0 1 -32
box -1604 -4676 5429 1783
use contador1bit  contador1bit_2
timestamp 1624053917
transform 1 0 3337 0 -1 2012
box -1604 -4676 5429 1783
use contador1bit  contador1bit_3
timestamp 1624053917
transform -1 0 3554 0 -1 2012
box -1604 -4676 5429 1783
use contador1bit  x1
timestamp 1624053917
transform 1 0 -140 0 1 568
box -1604 -4676 5429 1783
use contador1bit  x2
timestamp 1624053917
transform 1 0 3274 0 1 568
box -1604 -4676 5429 1783
use contador1bit  x3
timestamp 1624053917
transform 1 0 6688 0 1 568
box -1604 -4676 5429 1783
use contador1bit  x4
timestamp 1624053917
transform 1 0 10102 0 1 568
box -1604 -4676 5429 1783
<< labels >>
rlabel metal1 1812 386 1878 442 1 CLK
rlabel metal2 291 523 363 577 1 CLR
rlabel metal2 659 1556 721 1628 1 Q3
rlabel metal2 6170 1556 6232 1628 1 Q2
rlabel metal2 6170 352 6232 424 1 Q1
rlabel metal2 659 349 721 424 1 Q0
rlabel metal1 2894 426 2922 534 1 CE
rlabel metal1 3326 1529 3414 1663 1 Sout
rlabel metal1 6920 0 6948 1980 1 vss
rlabel metal1 -56 909 0 1071 1 vdd
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q0
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Q2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Q3
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Q1
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 CE
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 CLR
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 Sout
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 vss
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 CLK
port 10 nsew
<< end >>
