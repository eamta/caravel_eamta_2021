magic
tech sky130A
magscale 1 2
timestamp 1615925795
<< pwell >>
rect -637 2040 12265 2068
rect -637 -1147 12467 2040
rect -435 -1175 12467 -1147
<< psubdiff >>
rect -307 1619 -211 1653
rect 12041 1619 12137 1653
rect -307 1557 -273 1619
rect -307 -726 -273 -664
rect 12103 1557 12137 1619
rect 12103 -726 12137 -664
rect -307 -760 -211 -726
rect 12041 -760 12137 -726
<< psubdiffcont >>
rect -211 1619 12041 1653
rect -307 -664 -273 1557
rect 12103 -664 12137 1557
rect -211 -760 12041 -726
<< locali >>
rect -307 1619 -211 1653
rect 12041 1619 12137 1653
rect -307 1557 -273 1619
rect -307 -726 -273 -664
rect 12103 1557 12137 1619
rect 12103 -726 12137 -664
rect -307 -760 -211 -726
rect 12041 -760 12137 -726
<< metal1 >>
rect -7 810 3 1386
rect 55 810 65 1386
rect 111 810 121 1386
rect 173 810 183 1386
rect 229 810 239 1386
rect 291 810 301 1386
rect 347 810 357 1386
rect 409 810 419 1386
rect 465 810 475 1386
rect 527 810 537 1386
rect 583 810 593 1386
rect 645 810 655 1386
rect 701 810 711 1386
rect 763 810 773 1386
rect 819 810 829 1386
rect 881 810 891 1386
rect 937 810 947 1386
rect 999 810 1009 1386
rect 1055 810 1065 1386
rect 1117 810 1127 1386
rect 1173 810 1183 1386
rect 1235 810 1245 1386
rect 1291 810 1301 1386
rect 1353 810 1363 1386
rect 1409 810 1419 1386
rect 1471 810 1481 1386
rect 1527 810 1537 1386
rect 1589 810 1599 1386
rect 1645 810 1655 1386
rect 1707 810 1717 1386
rect 1763 810 1773 1386
rect 1825 810 1835 1386
rect 1881 810 1891 1386
rect 1943 810 1953 1386
rect 1999 810 2009 1386
rect 2061 810 2071 1386
rect 2117 810 2127 1386
rect 2179 810 2189 1386
rect 2235 810 2245 1386
rect 2297 810 2307 1386
rect 2353 810 2363 1386
rect 2415 810 2425 1386
rect 2471 810 2481 1386
rect 2533 810 2543 1386
rect 2589 810 2599 1386
rect 2651 810 2661 1386
rect 2707 810 2717 1386
rect 2769 810 2779 1386
rect 2825 810 2835 1386
rect 2887 810 2897 1386
rect 2943 810 2953 1386
rect 3005 810 3015 1386
rect 3061 810 3071 1386
rect 3123 810 3133 1386
rect 3179 810 3189 1386
rect 3241 810 3251 1386
rect 3297 810 3307 1386
rect 3359 810 3369 1386
rect 3415 810 3425 1386
rect 3477 810 3487 1386
rect 3533 810 3543 1386
rect 3595 810 3605 1386
rect 3651 810 3661 1386
rect 3713 810 3723 1386
rect 3769 810 3779 1386
rect 3831 810 3841 1386
rect 3887 810 3897 1386
rect 3949 810 3959 1386
rect 4005 810 4015 1386
rect 4067 810 4077 1386
rect 4123 810 4133 1386
rect 4185 810 4195 1386
rect 4241 810 4251 1386
rect 4303 810 4313 1386
rect 4359 810 4369 1386
rect 4421 810 4431 1386
rect 4477 810 4487 1386
rect 4539 810 4549 1386
rect 4595 810 4605 1386
rect 4657 810 4667 1386
rect 4713 810 4723 1386
rect 4775 810 4785 1386
rect 4831 810 4841 1386
rect 4893 810 4903 1386
rect 4949 810 4959 1386
rect 5011 810 5021 1386
rect 5067 810 5077 1386
rect 5129 810 5139 1386
rect 5185 810 5195 1386
rect 5247 810 5257 1386
rect 5303 810 5313 1386
rect 5365 810 5375 1386
rect 5421 810 5431 1386
rect 5483 810 5493 1386
rect 5539 810 5549 1386
rect 5601 810 5611 1386
rect 5657 810 5667 1386
rect 5719 810 5729 1386
rect 5775 810 5785 1386
rect 5837 810 5847 1386
rect 5893 810 5903 1386
rect 5955 810 5965 1386
rect 6011 810 6021 1386
rect 6073 810 6083 1386
rect 6129 810 6139 1386
rect 6191 810 6201 1386
rect 6247 810 6257 1386
rect 6309 810 6319 1386
rect 6365 810 6375 1386
rect 6427 810 6437 1386
rect 6483 810 6493 1386
rect 6545 810 6555 1386
rect 6601 810 6611 1386
rect 6663 810 6673 1386
rect 6719 810 6729 1386
rect 6781 810 6791 1386
rect 6837 810 6847 1386
rect 6899 810 6909 1386
rect 6955 810 6965 1386
rect 7017 810 7027 1386
rect 7073 810 7083 1386
rect 7135 810 7145 1386
rect 7191 810 7201 1386
rect 7253 810 7263 1386
rect 7309 810 7319 1386
rect 7371 810 7381 1386
rect 7427 810 7437 1386
rect 7489 810 7499 1386
rect 7545 810 7555 1386
rect 7607 810 7617 1386
rect 7663 810 7673 1386
rect 7725 810 7735 1386
rect 7781 810 7791 1386
rect 7843 810 7853 1386
rect 7899 810 7909 1386
rect 7961 810 7971 1386
rect 8017 810 8027 1386
rect 8079 810 8089 1386
rect 8135 810 8145 1386
rect 8197 810 8207 1386
rect 8253 810 8263 1386
rect 8315 810 8325 1386
rect 8371 810 8381 1386
rect 8433 810 8443 1386
rect 8489 810 8499 1386
rect 8551 810 8561 1386
rect 8607 810 8617 1386
rect 8669 810 8679 1386
rect 8725 810 8735 1386
rect 8787 810 8797 1386
rect 8843 810 8853 1386
rect 8905 810 8915 1386
rect 8961 810 8971 1386
rect 9023 810 9033 1386
rect 9079 810 9089 1386
rect 9141 810 9151 1386
rect 9197 810 9207 1386
rect 9259 810 9269 1386
rect 9315 810 9325 1386
rect 9377 810 9387 1386
rect 9433 810 9443 1386
rect 9495 810 9505 1386
rect 9551 810 9561 1386
rect 9613 810 9623 1386
rect 9669 810 9679 1386
rect 9731 810 9741 1386
rect 9787 810 9797 1386
rect 9849 810 9859 1386
rect 9905 810 9915 1386
rect 9967 810 9977 1386
rect 10023 810 10033 1386
rect 10085 810 10095 1386
rect 10141 810 10151 1386
rect 10203 810 10213 1386
rect 10259 810 10269 1386
rect 10321 810 10331 1386
rect 10377 810 10387 1386
rect 10439 810 10449 1386
rect 10495 810 10505 1386
rect 10557 810 10567 1386
rect 10613 810 10623 1386
rect 10675 810 10685 1386
rect 10731 810 10741 1386
rect 10793 810 10803 1386
rect 10849 810 10859 1386
rect 10911 810 10921 1386
rect 10967 810 10977 1386
rect 11029 810 11039 1386
rect 11085 810 11095 1386
rect 11147 810 11157 1386
rect 11203 810 11213 1386
rect 11265 810 11275 1386
rect 11321 810 11331 1386
rect 11383 810 11393 1386
rect 11439 810 11449 1386
rect 11501 810 11511 1386
rect 11557 810 11567 1386
rect 11619 810 11629 1386
rect 11675 810 11685 1386
rect 11737 810 11747 1386
rect 11793 810 11803 1386
rect 11855 810 11865 1386
rect -115 720 11973 766
rect -115 526 -35 720
rect -115 466 -105 526
rect -45 466 -35 526
rect -115 418 -35 466
rect -115 358 -105 418
rect -45 358 -35 418
rect -115 310 -35 358
rect -115 250 -105 310
rect -45 250 -35 310
rect -115 56 -35 250
rect -7 100 3 676
rect 55 100 65 676
rect 111 100 121 676
rect 173 100 183 676
rect 229 100 239 676
rect 291 100 301 676
rect 347 100 357 676
rect 409 100 419 676
rect 465 100 475 676
rect 527 100 537 676
rect 583 100 593 676
rect 645 100 655 676
rect 701 100 711 676
rect 763 100 773 676
rect 819 100 829 676
rect 881 100 891 676
rect 937 100 947 676
rect 999 100 1009 676
rect 1055 100 1065 676
rect 1117 100 1127 676
rect 1173 100 1183 676
rect 1235 100 1245 676
rect 1291 100 1301 676
rect 1353 100 1363 676
rect 1409 100 1419 676
rect 1471 100 1481 676
rect 1527 100 1537 676
rect 1589 100 1599 676
rect 1645 100 1655 676
rect 1707 100 1717 676
rect 1763 100 1773 676
rect 1825 100 1835 676
rect 1881 100 1891 676
rect 1943 100 1953 676
rect 1999 100 2009 676
rect 2061 100 2071 676
rect 2117 100 2127 676
rect 2179 100 2189 676
rect 2235 100 2245 676
rect 2297 100 2307 676
rect 2353 100 2363 676
rect 2415 100 2425 676
rect 2471 100 2481 676
rect 2533 100 2543 676
rect 2589 100 2599 676
rect 2651 100 2661 676
rect 2707 100 2717 676
rect 2769 100 2779 676
rect 2825 100 2835 676
rect 2887 100 2897 676
rect 2943 100 2953 676
rect 3005 100 3015 676
rect 3061 100 3071 676
rect 3123 100 3133 676
rect 3179 100 3189 676
rect 3241 100 3251 676
rect 3297 100 3307 676
rect 3359 100 3369 676
rect 3415 100 3425 676
rect 3477 100 3487 676
rect 3533 100 3543 676
rect 3595 100 3605 676
rect 3651 100 3661 676
rect 3713 100 3723 676
rect 3769 100 3779 676
rect 3831 100 3841 676
rect 3887 100 3897 676
rect 3949 100 3959 676
rect 4005 100 4015 676
rect 4067 100 4077 676
rect 4123 100 4133 676
rect 4185 100 4195 676
rect 4241 100 4251 676
rect 4303 100 4313 676
rect 4359 100 4369 676
rect 4421 100 4431 676
rect 4477 100 4487 676
rect 4539 100 4549 676
rect 4595 100 4605 676
rect 4657 100 4667 676
rect 4713 100 4723 676
rect 4775 100 4785 676
rect 4831 100 4841 676
rect 4893 100 4903 676
rect 4949 100 4959 676
rect 5011 100 5021 676
rect 5067 100 5077 676
rect 5129 100 5139 676
rect 5185 100 5195 676
rect 5247 100 5257 676
rect 5303 100 5313 676
rect 5365 100 5375 676
rect 5421 100 5431 676
rect 5483 100 5493 676
rect 5539 100 5549 676
rect 5601 100 5611 676
rect 5657 100 5667 676
rect 5719 100 5729 676
rect 5775 100 5785 676
rect 5837 100 5847 676
rect 5893 100 5903 676
rect 5955 100 5965 676
rect 6011 100 6021 676
rect 6073 100 6083 676
rect 6129 100 6139 676
rect 6191 100 6201 676
rect 6247 100 6257 676
rect 6309 100 6319 676
rect 6365 100 6375 676
rect 6427 100 6437 676
rect 6483 100 6493 676
rect 6545 100 6555 676
rect 6601 100 6611 676
rect 6663 100 6673 676
rect 6719 100 6729 676
rect 6781 100 6791 676
rect 6837 100 6847 676
rect 6899 100 6909 676
rect 6955 100 6965 676
rect 7017 100 7027 676
rect 7073 100 7083 676
rect 7135 100 7145 676
rect 7191 100 7201 676
rect 7253 100 7263 676
rect 7309 100 7319 676
rect 7371 100 7381 676
rect 7427 100 7437 676
rect 7489 100 7499 676
rect 7545 100 7555 676
rect 7607 100 7617 676
rect 7663 100 7673 676
rect 7725 100 7735 676
rect 7781 100 7791 676
rect 7843 100 7853 676
rect 7899 100 7909 676
rect 7961 100 7971 676
rect 8017 100 8027 676
rect 8079 100 8089 676
rect 8135 100 8145 676
rect 8197 100 8207 676
rect 8253 100 8263 676
rect 8315 100 8325 676
rect 8371 100 8381 676
rect 8433 100 8443 676
rect 8489 100 8499 676
rect 8551 100 8561 676
rect 8607 100 8617 676
rect 8669 100 8679 676
rect 8725 100 8735 676
rect 8787 100 8797 676
rect 8843 100 8853 676
rect 8905 100 8915 676
rect 8961 100 8971 676
rect 9023 100 9033 676
rect 9079 100 9089 676
rect 9141 100 9151 676
rect 9197 100 9207 676
rect 9259 100 9269 676
rect 9315 100 9325 676
rect 9377 100 9387 676
rect 9433 100 9443 676
rect 9495 100 9505 676
rect 9551 100 9561 676
rect 9613 100 9623 676
rect 9669 100 9679 676
rect 9731 100 9741 676
rect 9787 100 9797 676
rect 9849 100 9859 676
rect 9905 100 9915 676
rect 9967 100 9977 676
rect 10023 100 10033 676
rect 10085 100 10095 676
rect 10141 100 10151 676
rect 10203 100 10213 676
rect 10259 100 10269 676
rect 10321 100 10331 676
rect 10377 100 10387 676
rect 10439 100 10449 676
rect 10495 100 10505 676
rect 10557 100 10567 676
rect 10613 100 10623 676
rect 10675 100 10685 676
rect 10731 100 10741 676
rect 10793 100 10803 676
rect 10849 100 10859 676
rect 10911 100 10921 676
rect 10967 100 10977 676
rect 11029 100 11039 676
rect 11085 100 11095 676
rect 11147 100 11157 676
rect 11203 100 11213 676
rect 11265 100 11275 676
rect 11321 100 11331 676
rect 11383 100 11393 676
rect 11439 100 11449 676
rect 11501 100 11511 676
rect 11557 100 11567 676
rect 11619 100 11629 676
rect 11675 100 11685 676
rect 11737 100 11747 676
rect 11793 100 11803 676
rect 11855 100 11865 676
rect 11893 56 11973 720
rect -115 10 11973 56
rect -7 -610 3 -34
rect 55 -610 65 -34
rect 111 -610 121 -34
rect 173 -610 183 -34
rect 229 -610 239 -34
rect 291 -610 301 -34
rect 347 -610 357 -34
rect 409 -610 419 -34
rect 465 -610 475 -34
rect 527 -610 537 -34
rect 583 -610 593 -34
rect 645 -610 655 -34
rect 701 -610 711 -34
rect 763 -610 773 -34
rect 819 -610 829 -34
rect 881 -610 891 -34
rect 937 -610 947 -34
rect 999 -610 1009 -34
rect 1055 -610 1065 -34
rect 1117 -610 1127 -34
rect 1173 -610 1183 -34
rect 1235 -610 1245 -34
rect 1291 -610 1301 -34
rect 1353 -610 1363 -34
rect 1409 -610 1419 -34
rect 1471 -610 1481 -34
rect 1527 -610 1537 -34
rect 1589 -610 1599 -34
rect 1645 -610 1655 -34
rect 1707 -610 1717 -34
rect 1763 -610 1773 -34
rect 1825 -610 1835 -34
rect 1881 -610 1891 -34
rect 1943 -610 1953 -34
rect 1999 -610 2009 -34
rect 2061 -610 2071 -34
rect 2117 -610 2127 -34
rect 2179 -610 2189 -34
rect 2235 -610 2245 -34
rect 2297 -610 2307 -34
rect 2353 -610 2363 -34
rect 2415 -610 2425 -34
rect 2471 -610 2481 -34
rect 2533 -610 2543 -34
rect 2589 -610 2599 -34
rect 2651 -610 2661 -34
rect 2707 -610 2717 -34
rect 2769 -610 2779 -34
rect 2825 -610 2835 -34
rect 2887 -610 2897 -34
rect 2943 -610 2953 -34
rect 3005 -610 3015 -34
rect 3061 -610 3071 -34
rect 3123 -610 3133 -34
rect 3179 -610 3189 -34
rect 3241 -610 3251 -34
rect 3297 -610 3307 -34
rect 3359 -610 3369 -34
rect 3415 -610 3425 -34
rect 3477 -610 3487 -34
rect 3533 -610 3543 -34
rect 3595 -610 3605 -34
rect 3651 -610 3661 -34
rect 3713 -610 3723 -34
rect 3769 -610 3779 -34
rect 3831 -610 3841 -34
rect 3887 -610 3897 -34
rect 3949 -610 3959 -34
rect 4005 -610 4015 -34
rect 4067 -610 4077 -34
rect 4123 -610 4133 -34
rect 4185 -610 4195 -34
rect 4241 -610 4251 -34
rect 4303 -610 4313 -34
rect 4359 -610 4369 -34
rect 4421 -610 4431 -34
rect 4477 -610 4487 -34
rect 4539 -610 4549 -34
rect 4595 -610 4605 -34
rect 4657 -610 4667 -34
rect 4713 -610 4723 -34
rect 4775 -610 4785 -34
rect 4831 -610 4841 -34
rect 4893 -610 4903 -34
rect 4949 -610 4959 -34
rect 5011 -610 5021 -34
rect 5067 -610 5077 -34
rect 5129 -610 5139 -34
rect 5185 -610 5195 -34
rect 5247 -610 5257 -34
rect 5303 -610 5313 -34
rect 5365 -610 5375 -34
rect 5421 -610 5431 -34
rect 5483 -610 5493 -34
rect 5539 -610 5549 -34
rect 5601 -610 5611 -34
rect 5657 -610 5667 -34
rect 5719 -610 5729 -34
rect 5775 -610 5785 -34
rect 5837 -610 5847 -34
rect 5893 -610 5903 -34
rect 5955 -610 5965 -34
rect 6011 -610 6021 -34
rect 6073 -610 6083 -34
rect 6129 -610 6139 -34
rect 6191 -610 6201 -34
rect 6247 -610 6257 -34
rect 6309 -610 6319 -34
rect 6365 -610 6375 -34
rect 6427 -610 6437 -34
rect 6483 -610 6493 -34
rect 6545 -610 6555 -34
rect 6601 -610 6611 -34
rect 6663 -610 6673 -34
rect 6719 -610 6729 -34
rect 6781 -610 6791 -34
rect 6837 -610 6847 -34
rect 6899 -610 6909 -34
rect 6955 -610 6965 -34
rect 7017 -610 7027 -34
rect 7073 -610 7083 -34
rect 7135 -610 7145 -34
rect 7191 -610 7201 -34
rect 7253 -610 7263 -34
rect 7309 -610 7319 -34
rect 7371 -610 7381 -34
rect 7427 -610 7437 -34
rect 7489 -610 7499 -34
rect 7545 -610 7555 -34
rect 7607 -610 7617 -34
rect 7663 -610 7673 -34
rect 7725 -610 7735 -34
rect 7781 -610 7791 -34
rect 7843 -610 7853 -34
rect 7899 -610 7909 -34
rect 7961 -610 7971 -34
rect 8017 -610 8027 -34
rect 8079 -610 8089 -34
rect 8135 -610 8145 -34
rect 8197 -610 8207 -34
rect 8253 -610 8263 -34
rect 8315 -610 8325 -34
rect 8371 -610 8381 -34
rect 8433 -610 8443 -34
rect 8489 -610 8499 -34
rect 8551 -610 8561 -34
rect 8607 -610 8617 -34
rect 8669 -610 8679 -34
rect 8725 -610 8735 -34
rect 8787 -610 8797 -34
rect 8843 -610 8853 -34
rect 8905 -610 8915 -34
rect 8961 -610 8971 -34
rect 9023 -610 9033 -34
rect 9079 -610 9089 -34
rect 9141 -610 9151 -34
rect 9197 -610 9207 -34
rect 9259 -610 9269 -34
rect 9315 -610 9325 -34
rect 9377 -610 9387 -34
rect 9433 -610 9443 -34
rect 9495 -610 9505 -34
rect 9551 -610 9561 -34
rect 9613 -610 9623 -34
rect 9669 -610 9679 -34
rect 9731 -610 9741 -34
rect 9787 -610 9797 -34
rect 9849 -610 9859 -34
rect 9905 -610 9915 -34
rect 9967 -610 9977 -34
rect 10023 -610 10033 -34
rect 10085 -610 10095 -34
rect 10141 -610 10151 -34
rect 10203 -610 10213 -34
rect 10259 -610 10269 -34
rect 10321 -610 10331 -34
rect 10377 -610 10387 -34
rect 10439 -610 10449 -34
rect 10495 -610 10505 -34
rect 10557 -610 10567 -34
rect 10613 -610 10623 -34
rect 10675 -610 10685 -34
rect 10731 -610 10741 -34
rect 10793 -610 10803 -34
rect 10849 -610 10859 -34
rect 10911 -610 10921 -34
rect 10967 -610 10977 -34
rect 11029 -610 11039 -34
rect 11085 -610 11095 -34
rect 11147 -610 11157 -34
rect 11203 -610 11213 -34
rect 11265 -610 11275 -34
rect 11321 -610 11331 -34
rect 11383 -610 11393 -34
rect 11439 -610 11449 -34
rect 11501 -610 11511 -34
rect 11557 -610 11567 -34
rect 11619 -610 11629 -34
rect 11675 -610 11685 -34
rect 11737 -610 11747 -34
rect 11793 -610 11803 -34
rect 11855 -610 11865 -34
<< via1 >>
rect 3 810 55 1386
rect 121 810 173 1386
rect 239 810 291 1386
rect 357 810 409 1386
rect 475 810 527 1386
rect 593 810 645 1386
rect 711 810 763 1386
rect 829 810 881 1386
rect 947 810 999 1386
rect 1065 810 1117 1386
rect 1183 810 1235 1386
rect 1301 810 1353 1386
rect 1419 810 1471 1386
rect 1537 810 1589 1386
rect 1655 810 1707 1386
rect 1773 810 1825 1386
rect 1891 810 1943 1386
rect 2009 810 2061 1386
rect 2127 810 2179 1386
rect 2245 810 2297 1386
rect 2363 810 2415 1386
rect 2481 810 2533 1386
rect 2599 810 2651 1386
rect 2717 810 2769 1386
rect 2835 810 2887 1386
rect 2953 810 3005 1386
rect 3071 810 3123 1386
rect 3189 810 3241 1386
rect 3307 810 3359 1386
rect 3425 810 3477 1386
rect 3543 810 3595 1386
rect 3661 810 3713 1386
rect 3779 810 3831 1386
rect 3897 810 3949 1386
rect 4015 810 4067 1386
rect 4133 810 4185 1386
rect 4251 810 4303 1386
rect 4369 810 4421 1386
rect 4487 810 4539 1386
rect 4605 810 4657 1386
rect 4723 810 4775 1386
rect 4841 810 4893 1386
rect 4959 810 5011 1386
rect 5077 810 5129 1386
rect 5195 810 5247 1386
rect 5313 810 5365 1386
rect 5431 810 5483 1386
rect 5549 810 5601 1386
rect 5667 810 5719 1386
rect 5785 810 5837 1386
rect 5903 810 5955 1386
rect 6021 810 6073 1386
rect 6139 810 6191 1386
rect 6257 810 6309 1386
rect 6375 810 6427 1386
rect 6493 810 6545 1386
rect 6611 810 6663 1386
rect 6729 810 6781 1386
rect 6847 810 6899 1386
rect 6965 810 7017 1386
rect 7083 810 7135 1386
rect 7201 810 7253 1386
rect 7319 810 7371 1386
rect 7437 810 7489 1386
rect 7555 810 7607 1386
rect 7673 810 7725 1386
rect 7791 810 7843 1386
rect 7909 810 7961 1386
rect 8027 810 8079 1386
rect 8145 810 8197 1386
rect 8263 810 8315 1386
rect 8381 810 8433 1386
rect 8499 810 8551 1386
rect 8617 810 8669 1386
rect 8735 810 8787 1386
rect 8853 810 8905 1386
rect 8971 810 9023 1386
rect 9089 810 9141 1386
rect 9207 810 9259 1386
rect 9325 810 9377 1386
rect 9443 810 9495 1386
rect 9561 810 9613 1386
rect 9679 810 9731 1386
rect 9797 810 9849 1386
rect 9915 810 9967 1386
rect 10033 810 10085 1386
rect 10151 810 10203 1386
rect 10269 810 10321 1386
rect 10387 810 10439 1386
rect 10505 810 10557 1386
rect 10623 810 10675 1386
rect 10741 810 10793 1386
rect 10859 810 10911 1386
rect 10977 810 11029 1386
rect 11095 810 11147 1386
rect 11213 810 11265 1386
rect 11331 810 11383 1386
rect 11449 810 11501 1386
rect 11567 810 11619 1386
rect 11685 810 11737 1386
rect 11803 810 11855 1386
rect -105 466 -45 526
rect -105 358 -45 418
rect -105 250 -45 310
rect 3 100 55 676
rect 121 100 173 676
rect 239 100 291 676
rect 357 100 409 676
rect 475 100 527 676
rect 593 100 645 676
rect 711 100 763 676
rect 829 100 881 676
rect 947 100 999 676
rect 1065 100 1117 676
rect 1183 100 1235 676
rect 1301 100 1353 676
rect 1419 100 1471 676
rect 1537 100 1589 676
rect 1655 100 1707 676
rect 1773 100 1825 676
rect 1891 100 1943 676
rect 2009 100 2061 676
rect 2127 100 2179 676
rect 2245 100 2297 676
rect 2363 100 2415 676
rect 2481 100 2533 676
rect 2599 100 2651 676
rect 2717 100 2769 676
rect 2835 100 2887 676
rect 2953 100 3005 676
rect 3071 100 3123 676
rect 3189 100 3241 676
rect 3307 100 3359 676
rect 3425 100 3477 676
rect 3543 100 3595 676
rect 3661 100 3713 676
rect 3779 100 3831 676
rect 3897 100 3949 676
rect 4015 100 4067 676
rect 4133 100 4185 676
rect 4251 100 4303 676
rect 4369 100 4421 676
rect 4487 100 4539 676
rect 4605 100 4657 676
rect 4723 100 4775 676
rect 4841 100 4893 676
rect 4959 100 5011 676
rect 5077 100 5129 676
rect 5195 100 5247 676
rect 5313 100 5365 676
rect 5431 100 5483 676
rect 5549 100 5601 676
rect 5667 100 5719 676
rect 5785 100 5837 676
rect 5903 100 5955 676
rect 6021 100 6073 676
rect 6139 100 6191 676
rect 6257 100 6309 676
rect 6375 100 6427 676
rect 6493 100 6545 676
rect 6611 100 6663 676
rect 6729 100 6781 676
rect 6847 100 6899 676
rect 6965 100 7017 676
rect 7083 100 7135 676
rect 7201 100 7253 676
rect 7319 100 7371 676
rect 7437 100 7489 676
rect 7555 100 7607 676
rect 7673 100 7725 676
rect 7791 100 7843 676
rect 7909 100 7961 676
rect 8027 100 8079 676
rect 8145 100 8197 676
rect 8263 100 8315 676
rect 8381 100 8433 676
rect 8499 100 8551 676
rect 8617 100 8669 676
rect 8735 100 8787 676
rect 8853 100 8905 676
rect 8971 100 9023 676
rect 9089 100 9141 676
rect 9207 100 9259 676
rect 9325 100 9377 676
rect 9443 100 9495 676
rect 9561 100 9613 676
rect 9679 100 9731 676
rect 9797 100 9849 676
rect 9915 100 9967 676
rect 10033 100 10085 676
rect 10151 100 10203 676
rect 10269 100 10321 676
rect 10387 100 10439 676
rect 10505 100 10557 676
rect 10623 100 10675 676
rect 10741 100 10793 676
rect 10859 100 10911 676
rect 10977 100 11029 676
rect 11095 100 11147 676
rect 11213 100 11265 676
rect 11331 100 11383 676
rect 11449 100 11501 676
rect 11567 100 11619 676
rect 11685 100 11737 676
rect 11803 100 11855 676
rect 3 -610 55 -34
rect 121 -610 173 -34
rect 239 -610 291 -34
rect 357 -610 409 -34
rect 475 -610 527 -34
rect 593 -610 645 -34
rect 711 -610 763 -34
rect 829 -610 881 -34
rect 947 -610 999 -34
rect 1065 -610 1117 -34
rect 1183 -610 1235 -34
rect 1301 -610 1353 -34
rect 1419 -610 1471 -34
rect 1537 -610 1589 -34
rect 1655 -610 1707 -34
rect 1773 -610 1825 -34
rect 1891 -610 1943 -34
rect 2009 -610 2061 -34
rect 2127 -610 2179 -34
rect 2245 -610 2297 -34
rect 2363 -610 2415 -34
rect 2481 -610 2533 -34
rect 2599 -610 2651 -34
rect 2717 -610 2769 -34
rect 2835 -610 2887 -34
rect 2953 -610 3005 -34
rect 3071 -610 3123 -34
rect 3189 -610 3241 -34
rect 3307 -610 3359 -34
rect 3425 -610 3477 -34
rect 3543 -610 3595 -34
rect 3661 -610 3713 -34
rect 3779 -610 3831 -34
rect 3897 -610 3949 -34
rect 4015 -610 4067 -34
rect 4133 -610 4185 -34
rect 4251 -610 4303 -34
rect 4369 -610 4421 -34
rect 4487 -610 4539 -34
rect 4605 -610 4657 -34
rect 4723 -610 4775 -34
rect 4841 -610 4893 -34
rect 4959 -610 5011 -34
rect 5077 -610 5129 -34
rect 5195 -610 5247 -34
rect 5313 -610 5365 -34
rect 5431 -610 5483 -34
rect 5549 -610 5601 -34
rect 5667 -610 5719 -34
rect 5785 -610 5837 -34
rect 5903 -610 5955 -34
rect 6021 -610 6073 -34
rect 6139 -610 6191 -34
rect 6257 -610 6309 -34
rect 6375 -610 6427 -34
rect 6493 -610 6545 -34
rect 6611 -610 6663 -34
rect 6729 -610 6781 -34
rect 6847 -610 6899 -34
rect 6965 -610 7017 -34
rect 7083 -610 7135 -34
rect 7201 -610 7253 -34
rect 7319 -610 7371 -34
rect 7437 -610 7489 -34
rect 7555 -610 7607 -34
rect 7673 -610 7725 -34
rect 7791 -610 7843 -34
rect 7909 -610 7961 -34
rect 8027 -610 8079 -34
rect 8145 -610 8197 -34
rect 8263 -610 8315 -34
rect 8381 -610 8433 -34
rect 8499 -610 8551 -34
rect 8617 -610 8669 -34
rect 8735 -610 8787 -34
rect 8853 -610 8905 -34
rect 8971 -610 9023 -34
rect 9089 -610 9141 -34
rect 9207 -610 9259 -34
rect 9325 -610 9377 -34
rect 9443 -610 9495 -34
rect 9561 -610 9613 -34
rect 9679 -610 9731 -34
rect 9797 -610 9849 -34
rect 9915 -610 9967 -34
rect 10033 -610 10085 -34
rect 10151 -610 10203 -34
rect 10269 -610 10321 -34
rect 10387 -610 10439 -34
rect 10505 -610 10557 -34
rect 10623 -610 10675 -34
rect 10741 -610 10793 -34
rect 10859 -610 10911 -34
rect 10977 -610 11029 -34
rect 11095 -610 11147 -34
rect 11213 -610 11265 -34
rect 11331 -610 11383 -34
rect 11449 -610 11501 -34
rect 11567 -610 11619 -34
rect 11685 -610 11737 -34
rect 11803 -610 11855 -34
<< metal2 >>
rect 109 1534 185 1544
rect 109 1478 119 1534
rect 175 1478 185 1534
rect 109 1468 185 1478
rect 345 1534 421 1544
rect 345 1478 355 1534
rect 411 1478 421 1534
rect 345 1468 421 1478
rect 581 1534 657 1544
rect 581 1478 591 1534
rect 647 1478 657 1534
rect 581 1468 657 1478
rect 817 1534 893 1544
rect 817 1478 827 1534
rect 883 1478 893 1534
rect 817 1468 893 1478
rect 1053 1534 1129 1544
rect 1053 1478 1063 1534
rect 1119 1478 1129 1534
rect 1053 1468 1129 1478
rect 1289 1534 1365 1544
rect 1289 1478 1299 1534
rect 1355 1478 1365 1534
rect 1289 1468 1365 1478
rect 1525 1534 1601 1544
rect 1525 1478 1535 1534
rect 1591 1478 1601 1534
rect 1525 1468 1601 1478
rect 1761 1534 1837 1544
rect 1761 1478 1771 1534
rect 1827 1478 1837 1534
rect 1761 1468 1837 1478
rect 1997 1534 2073 1544
rect 1997 1478 2007 1534
rect 2063 1478 2073 1534
rect 1997 1468 2073 1478
rect 2233 1534 2309 1544
rect 2233 1478 2243 1534
rect 2299 1478 2309 1534
rect 2233 1468 2309 1478
rect 2469 1534 2545 1544
rect 2469 1478 2479 1534
rect 2535 1478 2545 1534
rect 2469 1468 2545 1478
rect 2705 1534 2781 1544
rect 2705 1478 2715 1534
rect 2771 1478 2781 1534
rect 2705 1468 2781 1478
rect 2941 1534 3017 1544
rect 2941 1478 2951 1534
rect 3007 1478 3017 1534
rect 2941 1468 3017 1478
rect 3177 1534 3253 1544
rect 3177 1478 3187 1534
rect 3243 1478 3253 1534
rect 3177 1468 3253 1478
rect 3413 1534 3489 1544
rect 3413 1478 3423 1534
rect 3479 1478 3489 1534
rect 3413 1468 3489 1478
rect 3649 1534 3725 1544
rect 3649 1478 3659 1534
rect 3715 1478 3725 1534
rect 3649 1468 3725 1478
rect 3885 1534 3961 1544
rect 3885 1478 3895 1534
rect 3951 1478 3961 1534
rect 3885 1468 3961 1478
rect 4121 1534 4197 1544
rect 4121 1478 4131 1534
rect 4187 1478 4197 1534
rect 4121 1468 4197 1478
rect 4357 1534 4433 1544
rect 4357 1478 4367 1534
rect 4423 1478 4433 1534
rect 4357 1468 4433 1478
rect 4593 1534 4669 1544
rect 4593 1478 4603 1534
rect 4659 1478 4669 1534
rect 4593 1468 4669 1478
rect 4829 1534 4905 1544
rect 4829 1478 4839 1534
rect 4895 1478 4905 1534
rect 4829 1468 4905 1478
rect 5065 1534 5141 1544
rect 5065 1478 5075 1534
rect 5131 1478 5141 1534
rect 5065 1468 5141 1478
rect 5301 1534 5377 1544
rect 5301 1478 5311 1534
rect 5367 1478 5377 1534
rect 5301 1468 5377 1478
rect 5537 1534 5613 1544
rect 5537 1478 5547 1534
rect 5603 1478 5613 1534
rect 5537 1468 5613 1478
rect 5773 1534 5849 1544
rect 5773 1478 5783 1534
rect 5839 1478 5849 1534
rect 5773 1468 5849 1478
rect 6009 1534 6085 1544
rect 6009 1478 6019 1534
rect 6075 1478 6085 1534
rect 6009 1468 6085 1478
rect 6245 1534 6321 1544
rect 6245 1478 6255 1534
rect 6311 1478 6321 1534
rect 6245 1468 6321 1478
rect 6481 1534 6557 1544
rect 6481 1478 6491 1534
rect 6547 1478 6557 1534
rect 6481 1468 6557 1478
rect 6717 1534 6793 1544
rect 6717 1478 6727 1534
rect 6783 1478 6793 1534
rect 6717 1468 6793 1478
rect 6953 1534 7029 1544
rect 6953 1478 6963 1534
rect 7019 1478 7029 1534
rect 6953 1468 7029 1478
rect 7189 1534 7265 1544
rect 7189 1478 7199 1534
rect 7255 1478 7265 1534
rect 7189 1468 7265 1478
rect 7425 1534 7501 1544
rect 7425 1478 7435 1534
rect 7491 1478 7501 1534
rect 7425 1468 7501 1478
rect 7661 1534 7737 1544
rect 7661 1478 7671 1534
rect 7727 1478 7737 1534
rect 7661 1468 7737 1478
rect 7897 1534 7973 1544
rect 7897 1478 7907 1534
rect 7963 1478 7973 1534
rect 7897 1468 7973 1478
rect 8133 1534 8209 1544
rect 8133 1478 8143 1534
rect 8199 1478 8209 1534
rect 8133 1468 8209 1478
rect 8369 1534 8445 1544
rect 8369 1478 8379 1534
rect 8435 1478 8445 1534
rect 8369 1468 8445 1478
rect 8605 1534 8681 1544
rect 8605 1478 8615 1534
rect 8671 1478 8681 1534
rect 8605 1468 8681 1478
rect 8841 1534 8917 1544
rect 8841 1478 8851 1534
rect 8907 1478 8917 1534
rect 8841 1468 8917 1478
rect 9077 1534 9153 1544
rect 9077 1478 9087 1534
rect 9143 1478 9153 1534
rect 9077 1468 9153 1478
rect 9313 1534 9389 1544
rect 9313 1478 9323 1534
rect 9379 1478 9389 1534
rect 9313 1468 9389 1478
rect 9549 1534 9625 1544
rect 9549 1478 9559 1534
rect 9615 1478 9625 1534
rect 9549 1468 9625 1478
rect 9785 1534 9861 1544
rect 9785 1478 9795 1534
rect 9851 1478 9861 1534
rect 9785 1468 9861 1478
rect 10021 1534 10097 1544
rect 10021 1478 10031 1534
rect 10087 1478 10097 1534
rect 10021 1468 10097 1478
rect 10257 1534 10333 1544
rect 10257 1478 10267 1534
rect 10323 1478 10333 1534
rect 10257 1468 10333 1478
rect 10493 1534 10569 1544
rect 10493 1478 10503 1534
rect 10559 1478 10569 1534
rect 10493 1468 10569 1478
rect 10729 1534 10805 1544
rect 10729 1478 10739 1534
rect 10795 1478 10805 1534
rect 10729 1468 10805 1478
rect 10965 1534 11041 1544
rect 10965 1478 10975 1534
rect 11031 1478 11041 1534
rect 10965 1468 11041 1478
rect 11201 1534 11277 1544
rect 11201 1478 11211 1534
rect 11267 1478 11277 1534
rect 11201 1468 11277 1478
rect 11437 1534 11513 1544
rect 11437 1478 11447 1534
rect 11503 1478 11513 1534
rect 11437 1468 11513 1478
rect 11673 1534 11749 1544
rect 11673 1478 11683 1534
rect 11739 1478 11749 1534
rect 11673 1468 11749 1478
rect 3 1386 55 1396
rect 3 676 55 810
rect -105 526 -45 536
rect -105 456 -45 466
rect -105 418 -45 428
rect -105 348 -45 358
rect -105 310 -45 320
rect -105 240 -45 250
rect 3 -34 55 100
rect 3 -739 55 -610
rect 121 1386 173 1468
rect 121 676 173 810
rect 121 -34 173 100
rect 121 -620 173 -610
rect 239 1386 291 1396
rect 239 676 291 810
rect 239 -34 291 100
rect 239 -739 291 -610
rect 357 1386 409 1468
rect 357 676 409 810
rect 357 -34 409 100
rect 357 -620 409 -610
rect 475 1386 527 1396
rect 475 676 527 810
rect 475 -34 527 100
rect 475 -739 527 -610
rect 593 1386 645 1468
rect 593 676 645 810
rect 593 -34 645 100
rect 593 -620 645 -610
rect 711 1386 763 1396
rect 711 676 763 810
rect 711 -34 763 100
rect 711 -739 763 -610
rect 829 1386 881 1468
rect 829 676 881 810
rect 829 -34 881 100
rect 829 -620 881 -610
rect 947 1386 999 1396
rect 947 676 999 810
rect 947 -34 999 100
rect 947 -739 999 -610
rect 1065 1386 1117 1468
rect 1065 676 1117 810
rect 1065 -34 1117 100
rect 1065 -620 1117 -610
rect 1183 1386 1235 1396
rect 1183 676 1235 810
rect 1183 -34 1235 100
rect 1183 -739 1235 -610
rect 1301 1386 1353 1468
rect 1301 676 1353 810
rect 1301 -34 1353 100
rect 1301 -620 1353 -610
rect 1419 1386 1471 1396
rect 1419 676 1471 810
rect 1419 -34 1471 100
rect 1419 -739 1471 -610
rect 1537 1386 1589 1468
rect 1537 676 1589 810
rect 1537 -34 1589 100
rect 1537 -620 1589 -610
rect 1655 1386 1707 1396
rect 1655 676 1707 810
rect 1655 -34 1707 100
rect 1655 -739 1707 -610
rect 1773 1386 1825 1468
rect 1773 676 1825 810
rect 1773 -34 1825 100
rect 1773 -620 1825 -610
rect 1891 1386 1943 1396
rect 1891 676 1943 810
rect 1891 -34 1943 100
rect 1891 -739 1943 -610
rect 2009 1386 2061 1468
rect 2009 676 2061 810
rect 2009 -34 2061 100
rect 2009 -620 2061 -610
rect 2127 1386 2179 1396
rect 2127 676 2179 810
rect 2127 -34 2179 100
rect 2127 -739 2179 -610
rect 2245 1386 2297 1468
rect 2245 676 2297 810
rect 2245 -34 2297 100
rect 2245 -620 2297 -610
rect 2363 1386 2415 1396
rect 2363 676 2415 810
rect 2363 -34 2415 100
rect 2363 -739 2415 -610
rect 2481 1386 2533 1468
rect 2481 676 2533 810
rect 2481 -34 2533 100
rect 2481 -620 2533 -610
rect 2599 1386 2651 1396
rect 2599 676 2651 810
rect 2599 -34 2651 100
rect 2599 -739 2651 -610
rect 2717 1386 2769 1468
rect 2717 676 2769 810
rect 2717 -34 2769 100
rect 2717 -620 2769 -610
rect 2835 1386 2887 1396
rect 2835 676 2887 810
rect 2835 -34 2887 100
rect 2835 -739 2887 -610
rect 2953 1386 3005 1468
rect 2953 676 3005 810
rect 2953 -34 3005 100
rect 2953 -620 3005 -610
rect 3071 1386 3123 1396
rect 3071 676 3123 810
rect 3071 -34 3123 100
rect 3071 -739 3123 -610
rect 3189 1386 3241 1468
rect 3189 676 3241 810
rect 3189 -34 3241 100
rect 3189 -620 3241 -610
rect 3307 1386 3359 1396
rect 3307 676 3359 810
rect 3307 -34 3359 100
rect 3307 -739 3359 -610
rect 3425 1386 3477 1468
rect 3425 676 3477 810
rect 3425 -34 3477 100
rect 3425 -620 3477 -610
rect 3543 1386 3595 1396
rect 3543 676 3595 810
rect 3543 -34 3595 100
rect 3543 -739 3595 -610
rect 3661 1386 3713 1468
rect 3661 676 3713 810
rect 3661 -34 3713 100
rect 3661 -620 3713 -610
rect 3779 1386 3831 1396
rect 3779 676 3831 810
rect 3779 -34 3831 100
rect 3779 -739 3831 -610
rect 3897 1386 3949 1468
rect 3897 676 3949 810
rect 3897 -34 3949 100
rect 3897 -620 3949 -610
rect 4015 1386 4067 1396
rect 4015 676 4067 810
rect 4015 -34 4067 100
rect 4015 -739 4067 -610
rect 4133 1386 4185 1468
rect 4133 676 4185 810
rect 4133 -34 4185 100
rect 4133 -620 4185 -610
rect 4251 1386 4303 1396
rect 4251 676 4303 810
rect 4251 -34 4303 100
rect 4251 -739 4303 -610
rect 4369 1386 4421 1468
rect 4369 676 4421 810
rect 4369 -34 4421 100
rect 4369 -620 4421 -610
rect 4487 1386 4539 1396
rect 4487 676 4539 810
rect 4487 -34 4539 100
rect 4487 -739 4539 -610
rect 4605 1386 4657 1468
rect 4605 676 4657 810
rect 4605 -34 4657 100
rect 4605 -620 4657 -610
rect 4723 1386 4775 1396
rect 4723 676 4775 810
rect 4723 -34 4775 100
rect 4723 -739 4775 -610
rect 4841 1386 4893 1468
rect 4841 676 4893 810
rect 4841 -34 4893 100
rect 4841 -620 4893 -610
rect 4959 1386 5011 1396
rect 4959 676 5011 810
rect 4959 -34 5011 100
rect 4959 -739 5011 -610
rect 5077 1386 5129 1468
rect 5077 676 5129 810
rect 5077 -34 5129 100
rect 5077 -620 5129 -610
rect 5195 1386 5247 1396
rect 5195 676 5247 810
rect 5195 -34 5247 100
rect 5195 -739 5247 -610
rect 5313 1386 5365 1468
rect 5313 676 5365 810
rect 5313 -34 5365 100
rect 5313 -620 5365 -610
rect 5431 1386 5483 1396
rect 5431 676 5483 810
rect 5431 -34 5483 100
rect 5431 -739 5483 -610
rect 5549 1386 5601 1468
rect 5549 676 5601 810
rect 5549 -34 5601 100
rect 5549 -620 5601 -610
rect 5667 1386 5719 1396
rect 5667 676 5719 810
rect 5667 -34 5719 100
rect 5667 -739 5719 -610
rect 5785 1386 5837 1468
rect 5785 676 5837 810
rect 5785 -34 5837 100
rect 5785 -620 5837 -610
rect 5903 1386 5955 1396
rect 5903 676 5955 810
rect 5903 -34 5955 100
rect 5903 -739 5955 -610
rect 6021 1386 6073 1468
rect 6021 676 6073 810
rect 6021 -34 6073 100
rect 6021 -620 6073 -610
rect 6139 1386 6191 1396
rect 6139 676 6191 810
rect 6139 -34 6191 100
rect 6139 -739 6191 -610
rect 6257 1386 6309 1468
rect 6257 676 6309 810
rect 6257 -34 6309 100
rect 6257 -620 6309 -610
rect 6375 1386 6427 1396
rect 6375 676 6427 810
rect 6375 -34 6427 100
rect 6375 -739 6427 -610
rect 6493 1386 6545 1468
rect 6493 676 6545 810
rect 6493 -34 6545 100
rect 6493 -620 6545 -610
rect 6611 1386 6663 1396
rect 6611 676 6663 810
rect 6611 -34 6663 100
rect 6611 -739 6663 -610
rect 6729 1386 6781 1468
rect 6729 676 6781 810
rect 6729 -34 6781 100
rect 6729 -620 6781 -610
rect 6847 1386 6899 1396
rect 6847 676 6899 810
rect 6847 -34 6899 100
rect 6847 -739 6899 -610
rect 6965 1386 7017 1468
rect 6965 676 7017 810
rect 6965 -34 7017 100
rect 6965 -620 7017 -610
rect 7083 1386 7135 1396
rect 7083 676 7135 810
rect 7083 -34 7135 100
rect 7083 -739 7135 -610
rect 7201 1386 7253 1468
rect 7201 676 7253 810
rect 7201 -34 7253 100
rect 7201 -620 7253 -610
rect 7319 1386 7371 1396
rect 7319 676 7371 810
rect 7319 -34 7371 100
rect 7319 -739 7371 -610
rect 7437 1386 7489 1468
rect 7437 676 7489 810
rect 7437 -34 7489 100
rect 7437 -620 7489 -610
rect 7555 1386 7607 1396
rect 7555 676 7607 810
rect 7555 -34 7607 100
rect 7555 -739 7607 -610
rect 7673 1386 7725 1468
rect 7673 676 7725 810
rect 7673 -34 7725 100
rect 7673 -620 7725 -610
rect 7791 1386 7843 1396
rect 7791 676 7843 810
rect 7791 -34 7843 100
rect 7791 -739 7843 -610
rect 7909 1386 7961 1468
rect 7909 676 7961 810
rect 7909 -34 7961 100
rect 7909 -620 7961 -610
rect 8027 1386 8079 1396
rect 8027 676 8079 810
rect 8027 -34 8079 100
rect 8027 -739 8079 -610
rect 8145 1386 8197 1468
rect 8145 676 8197 810
rect 8145 -34 8197 100
rect 8145 -620 8197 -610
rect 8263 1386 8315 1396
rect 8263 676 8315 810
rect 8263 -34 8315 100
rect 8263 -739 8315 -610
rect 8381 1386 8433 1468
rect 8381 676 8433 810
rect 8381 -34 8433 100
rect 8381 -620 8433 -610
rect 8499 1386 8551 1396
rect 8499 676 8551 810
rect 8499 -34 8551 100
rect 8499 -739 8551 -610
rect 8617 1386 8669 1468
rect 8617 676 8669 810
rect 8617 -34 8669 100
rect 8617 -620 8669 -610
rect 8735 1386 8787 1396
rect 8735 676 8787 810
rect 8735 -34 8787 100
rect 8735 -739 8787 -610
rect 8853 1386 8905 1468
rect 8853 676 8905 810
rect 8853 -34 8905 100
rect 8853 -620 8905 -610
rect 8971 1386 9023 1396
rect 8971 676 9023 810
rect 8971 -34 9023 100
rect 8971 -739 9023 -610
rect 9089 1386 9141 1468
rect 9089 676 9141 810
rect 9089 -34 9141 100
rect 9089 -620 9141 -610
rect 9207 1386 9259 1396
rect 9207 676 9259 810
rect 9207 -34 9259 100
rect 9207 -739 9259 -610
rect 9325 1386 9377 1468
rect 9325 676 9377 810
rect 9325 -34 9377 100
rect 9325 -620 9377 -610
rect 9443 1386 9495 1396
rect 9443 676 9495 810
rect 9443 -34 9495 100
rect 9443 -739 9495 -610
rect 9561 1386 9613 1468
rect 9561 676 9613 810
rect 9561 -34 9613 100
rect 9561 -620 9613 -610
rect 9679 1386 9731 1396
rect 9679 676 9731 810
rect 9679 -34 9731 100
rect 9679 -739 9731 -610
rect 9797 1386 9849 1468
rect 9797 676 9849 810
rect 9797 -34 9849 100
rect 9797 -620 9849 -610
rect 9915 1386 9967 1396
rect 9915 676 9967 810
rect 9915 -34 9967 100
rect 9915 -739 9967 -610
rect 10033 1386 10085 1468
rect 10033 676 10085 810
rect 10033 -34 10085 100
rect 10033 -620 10085 -610
rect 10151 1386 10203 1396
rect 10151 676 10203 810
rect 10151 -34 10203 100
rect 10151 -739 10203 -610
rect 10269 1386 10321 1468
rect 10269 676 10321 810
rect 10269 -34 10321 100
rect 10269 -620 10321 -610
rect 10387 1386 10439 1396
rect 10387 676 10439 810
rect 10387 -34 10439 100
rect 10387 -739 10439 -610
rect 10505 1386 10557 1468
rect 10505 676 10557 810
rect 10505 -34 10557 100
rect 10505 -620 10557 -610
rect 10623 1386 10675 1396
rect 10623 676 10675 810
rect 10623 -34 10675 100
rect 10623 -739 10675 -610
rect 10741 1386 10793 1468
rect 10741 676 10793 810
rect 10741 -34 10793 100
rect 10741 -620 10793 -610
rect 10859 1386 10911 1396
rect 10859 676 10911 810
rect 10859 -34 10911 100
rect 10859 -739 10911 -610
rect 10977 1386 11029 1468
rect 10977 676 11029 810
rect 10977 -34 11029 100
rect 10977 -620 11029 -610
rect 11095 1386 11147 1396
rect 11095 676 11147 810
rect 11095 -34 11147 100
rect 11095 -739 11147 -610
rect 11213 1386 11265 1468
rect 11213 676 11265 810
rect 11213 -34 11265 100
rect 11213 -620 11265 -610
rect 11331 1386 11383 1396
rect 11331 676 11383 810
rect 11331 -34 11383 100
rect 11331 -739 11383 -610
rect 11449 1386 11501 1468
rect 11449 676 11501 810
rect 11449 -34 11501 100
rect 11449 -620 11501 -610
rect 11567 1386 11619 1396
rect 11567 676 11619 810
rect 11567 -34 11619 100
rect 11567 -739 11619 -610
rect 11685 1386 11737 1468
rect 11685 676 11737 810
rect 11685 -34 11737 100
rect 11685 -620 11737 -610
rect 11803 1386 11855 1396
rect 11803 676 11855 810
rect 11803 -34 11855 100
rect 11803 -739 11855 -610
<< via2 >>
rect 119 1478 175 1534
rect 355 1478 411 1534
rect 591 1478 647 1534
rect 827 1478 883 1534
rect 1063 1478 1119 1534
rect 1299 1478 1355 1534
rect 1535 1478 1591 1534
rect 1771 1478 1827 1534
rect 2007 1478 2063 1534
rect 2243 1478 2299 1534
rect 2479 1478 2535 1534
rect 2715 1478 2771 1534
rect 2951 1478 3007 1534
rect 3187 1478 3243 1534
rect 3423 1478 3479 1534
rect 3659 1478 3715 1534
rect 3895 1478 3951 1534
rect 4131 1478 4187 1534
rect 4367 1478 4423 1534
rect 4603 1478 4659 1534
rect 4839 1478 4895 1534
rect 5075 1478 5131 1534
rect 5311 1478 5367 1534
rect 5547 1478 5603 1534
rect 5783 1478 5839 1534
rect 6019 1478 6075 1534
rect 6255 1478 6311 1534
rect 6491 1478 6547 1534
rect 6727 1478 6783 1534
rect 6963 1478 7019 1534
rect 7199 1478 7255 1534
rect 7435 1478 7491 1534
rect 7671 1478 7727 1534
rect 7907 1478 7963 1534
rect 8143 1478 8199 1534
rect 8379 1478 8435 1534
rect 8615 1478 8671 1534
rect 8851 1478 8907 1534
rect 9087 1478 9143 1534
rect 9323 1478 9379 1534
rect 9559 1478 9615 1534
rect 9795 1478 9851 1534
rect 10031 1478 10087 1534
rect 10267 1478 10323 1534
rect 10503 1478 10559 1534
rect 10739 1478 10795 1534
rect 10975 1478 11031 1534
rect 11211 1478 11267 1534
rect 11447 1478 11503 1534
rect 11683 1478 11739 1534
rect -105 466 -45 526
rect -105 358 -45 418
rect -105 250 -45 310
<< metal3 >>
rect 109 1534 11749 1544
rect 109 1478 119 1534
rect 175 1478 355 1534
rect 411 1478 591 1534
rect 647 1478 827 1534
rect 883 1478 1063 1534
rect 1119 1478 1299 1534
rect 1355 1478 1535 1534
rect 1591 1478 1771 1534
rect 1827 1478 2007 1534
rect 2063 1478 2243 1534
rect 2299 1478 2479 1534
rect 2535 1478 2715 1534
rect 2771 1478 2951 1534
rect 3007 1478 3187 1534
rect 3243 1478 3423 1534
rect 3479 1478 3659 1534
rect 3715 1478 3895 1534
rect 3951 1478 4131 1534
rect 4187 1478 4367 1534
rect 4423 1478 4603 1534
rect 4659 1478 4839 1534
rect 4895 1478 5075 1534
rect 5131 1478 5311 1534
rect 5367 1478 5547 1534
rect 5603 1478 5783 1534
rect 5839 1478 6019 1534
rect 6075 1478 6255 1534
rect 6311 1478 6491 1534
rect 6547 1478 6727 1534
rect 6783 1478 6963 1534
rect 7019 1478 7199 1534
rect 7255 1478 7435 1534
rect 7491 1478 7671 1534
rect 7727 1478 7907 1534
rect 7963 1478 8143 1534
rect 8199 1478 8379 1534
rect 8435 1478 8615 1534
rect 8671 1478 8851 1534
rect 8907 1478 9087 1534
rect 9143 1478 9323 1534
rect 9379 1478 9559 1534
rect 9615 1478 9795 1534
rect 9851 1478 10031 1534
rect 10087 1478 10267 1534
rect 10323 1478 10503 1534
rect 10559 1478 10739 1534
rect 10795 1478 10975 1534
rect 11031 1478 11211 1534
rect 11267 1478 11447 1534
rect 11503 1478 11683 1534
rect 11739 1478 11749 1534
rect 109 1468 11749 1478
rect -148 526 -35 536
rect -148 466 -105 526
rect -45 466 -35 526
rect -148 418 -35 466
rect -148 358 -105 418
rect -45 358 -35 418
rect -148 310 -35 358
rect -148 250 -105 310
rect -45 250 -35 310
rect -148 240 -35 250
use sky130_fd_pr__nfet_01v8_F2M6PM  sky130_fd_pr__nfet_01v8_F2M6PM_0
timestamp 1615923543
transform 1 0 5929 0 1 388
box -5929 -388 5929 388
use sky130_fd_pr__nfet_01v8_93MENK  sky130_fd_pr__nfet_01v8_93MENK_0
timestamp 1615923543
transform 1 0 5929 0 1 1067
box -5929 -357 5929 357
use sky130_fd_pr__nfet_01v8_93MENK  sky130_fd_pr__nfet_01v8_93MENK_1
timestamp 1615923543
transform 1 0 5929 0 -1 -291
box -5929 -357 5929 357
<< end >>
