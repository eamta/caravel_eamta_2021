magic
tech sky130A
magscale 1 2
timestamp 1619113446
<< pwell >>
rect -2257 -2691 2257 2691
<< nmos >>
rect -2061 2181 -1701 2481
rect -1643 2181 -1283 2481
rect -1225 2181 -865 2481
rect -807 2181 -447 2481
rect -389 2181 -29 2481
rect 29 2181 389 2481
rect 447 2181 807 2481
rect 865 2181 1225 2481
rect 1283 2181 1643 2481
rect 1701 2181 2061 2481
rect -2061 1663 -1701 1963
rect -1643 1663 -1283 1963
rect -1225 1663 -865 1963
rect -807 1663 -447 1963
rect -389 1663 -29 1963
rect 29 1663 389 1963
rect 447 1663 807 1963
rect 865 1663 1225 1963
rect 1283 1663 1643 1963
rect 1701 1663 2061 1963
rect -2061 1145 -1701 1445
rect -1643 1145 -1283 1445
rect -1225 1145 -865 1445
rect -807 1145 -447 1445
rect -389 1145 -29 1445
rect 29 1145 389 1445
rect 447 1145 807 1445
rect 865 1145 1225 1445
rect 1283 1145 1643 1445
rect 1701 1145 2061 1445
rect -2061 627 -1701 927
rect -1643 627 -1283 927
rect -1225 627 -865 927
rect -807 627 -447 927
rect -389 627 -29 927
rect 29 627 389 927
rect 447 627 807 927
rect 865 627 1225 927
rect 1283 627 1643 927
rect 1701 627 2061 927
rect -2061 109 -1701 409
rect -1643 109 -1283 409
rect -1225 109 -865 409
rect -807 109 -447 409
rect -389 109 -29 409
rect 29 109 389 409
rect 447 109 807 409
rect 865 109 1225 409
rect 1283 109 1643 409
rect 1701 109 2061 409
rect -2061 -409 -1701 -109
rect -1643 -409 -1283 -109
rect -1225 -409 -865 -109
rect -807 -409 -447 -109
rect -389 -409 -29 -109
rect 29 -409 389 -109
rect 447 -409 807 -109
rect 865 -409 1225 -109
rect 1283 -409 1643 -109
rect 1701 -409 2061 -109
rect -2061 -927 -1701 -627
rect -1643 -927 -1283 -627
rect -1225 -927 -865 -627
rect -807 -927 -447 -627
rect -389 -927 -29 -627
rect 29 -927 389 -627
rect 447 -927 807 -627
rect 865 -927 1225 -627
rect 1283 -927 1643 -627
rect 1701 -927 2061 -627
rect -2061 -1445 -1701 -1145
rect -1643 -1445 -1283 -1145
rect -1225 -1445 -865 -1145
rect -807 -1445 -447 -1145
rect -389 -1445 -29 -1145
rect 29 -1445 389 -1145
rect 447 -1445 807 -1145
rect 865 -1445 1225 -1145
rect 1283 -1445 1643 -1145
rect 1701 -1445 2061 -1145
rect -2061 -1963 -1701 -1663
rect -1643 -1963 -1283 -1663
rect -1225 -1963 -865 -1663
rect -807 -1963 -447 -1663
rect -389 -1963 -29 -1663
rect 29 -1963 389 -1663
rect 447 -1963 807 -1663
rect 865 -1963 1225 -1663
rect 1283 -1963 1643 -1663
rect 1701 -1963 2061 -1663
rect -2061 -2481 -1701 -2181
rect -1643 -2481 -1283 -2181
rect -1225 -2481 -865 -2181
rect -807 -2481 -447 -2181
rect -389 -2481 -29 -2181
rect 29 -2481 389 -2181
rect 447 -2481 807 -2181
rect 865 -2481 1225 -2181
rect 1283 -2481 1643 -2181
rect 1701 -2481 2061 -2181
<< ndiff >>
rect -2119 2469 -2061 2481
rect -2119 2193 -2107 2469
rect -2073 2193 -2061 2469
rect -2119 2181 -2061 2193
rect -1701 2469 -1643 2481
rect -1701 2193 -1689 2469
rect -1655 2193 -1643 2469
rect -1701 2181 -1643 2193
rect -1283 2469 -1225 2481
rect -1283 2193 -1271 2469
rect -1237 2193 -1225 2469
rect -1283 2181 -1225 2193
rect -865 2469 -807 2481
rect -865 2193 -853 2469
rect -819 2193 -807 2469
rect -865 2181 -807 2193
rect -447 2469 -389 2481
rect -447 2193 -435 2469
rect -401 2193 -389 2469
rect -447 2181 -389 2193
rect -29 2469 29 2481
rect -29 2193 -17 2469
rect 17 2193 29 2469
rect -29 2181 29 2193
rect 389 2469 447 2481
rect 389 2193 401 2469
rect 435 2193 447 2469
rect 389 2181 447 2193
rect 807 2469 865 2481
rect 807 2193 819 2469
rect 853 2193 865 2469
rect 807 2181 865 2193
rect 1225 2469 1283 2481
rect 1225 2193 1237 2469
rect 1271 2193 1283 2469
rect 1225 2181 1283 2193
rect 1643 2469 1701 2481
rect 1643 2193 1655 2469
rect 1689 2193 1701 2469
rect 1643 2181 1701 2193
rect 2061 2469 2119 2481
rect 2061 2193 2073 2469
rect 2107 2193 2119 2469
rect 2061 2181 2119 2193
rect -2119 1951 -2061 1963
rect -2119 1675 -2107 1951
rect -2073 1675 -2061 1951
rect -2119 1663 -2061 1675
rect -1701 1951 -1643 1963
rect -1701 1675 -1689 1951
rect -1655 1675 -1643 1951
rect -1701 1663 -1643 1675
rect -1283 1951 -1225 1963
rect -1283 1675 -1271 1951
rect -1237 1675 -1225 1951
rect -1283 1663 -1225 1675
rect -865 1951 -807 1963
rect -865 1675 -853 1951
rect -819 1675 -807 1951
rect -865 1663 -807 1675
rect -447 1951 -389 1963
rect -447 1675 -435 1951
rect -401 1675 -389 1951
rect -447 1663 -389 1675
rect -29 1951 29 1963
rect -29 1675 -17 1951
rect 17 1675 29 1951
rect -29 1663 29 1675
rect 389 1951 447 1963
rect 389 1675 401 1951
rect 435 1675 447 1951
rect 389 1663 447 1675
rect 807 1951 865 1963
rect 807 1675 819 1951
rect 853 1675 865 1951
rect 807 1663 865 1675
rect 1225 1951 1283 1963
rect 1225 1675 1237 1951
rect 1271 1675 1283 1951
rect 1225 1663 1283 1675
rect 1643 1951 1701 1963
rect 1643 1675 1655 1951
rect 1689 1675 1701 1951
rect 1643 1663 1701 1675
rect 2061 1951 2119 1963
rect 2061 1675 2073 1951
rect 2107 1675 2119 1951
rect 2061 1663 2119 1675
rect -2119 1433 -2061 1445
rect -2119 1157 -2107 1433
rect -2073 1157 -2061 1433
rect -2119 1145 -2061 1157
rect -1701 1433 -1643 1445
rect -1701 1157 -1689 1433
rect -1655 1157 -1643 1433
rect -1701 1145 -1643 1157
rect -1283 1433 -1225 1445
rect -1283 1157 -1271 1433
rect -1237 1157 -1225 1433
rect -1283 1145 -1225 1157
rect -865 1433 -807 1445
rect -865 1157 -853 1433
rect -819 1157 -807 1433
rect -865 1145 -807 1157
rect -447 1433 -389 1445
rect -447 1157 -435 1433
rect -401 1157 -389 1433
rect -447 1145 -389 1157
rect -29 1433 29 1445
rect -29 1157 -17 1433
rect 17 1157 29 1433
rect -29 1145 29 1157
rect 389 1433 447 1445
rect 389 1157 401 1433
rect 435 1157 447 1433
rect 389 1145 447 1157
rect 807 1433 865 1445
rect 807 1157 819 1433
rect 853 1157 865 1433
rect 807 1145 865 1157
rect 1225 1433 1283 1445
rect 1225 1157 1237 1433
rect 1271 1157 1283 1433
rect 1225 1145 1283 1157
rect 1643 1433 1701 1445
rect 1643 1157 1655 1433
rect 1689 1157 1701 1433
rect 1643 1145 1701 1157
rect 2061 1433 2119 1445
rect 2061 1157 2073 1433
rect 2107 1157 2119 1433
rect 2061 1145 2119 1157
rect -2119 915 -2061 927
rect -2119 639 -2107 915
rect -2073 639 -2061 915
rect -2119 627 -2061 639
rect -1701 915 -1643 927
rect -1701 639 -1689 915
rect -1655 639 -1643 915
rect -1701 627 -1643 639
rect -1283 915 -1225 927
rect -1283 639 -1271 915
rect -1237 639 -1225 915
rect -1283 627 -1225 639
rect -865 915 -807 927
rect -865 639 -853 915
rect -819 639 -807 915
rect -865 627 -807 639
rect -447 915 -389 927
rect -447 639 -435 915
rect -401 639 -389 915
rect -447 627 -389 639
rect -29 915 29 927
rect -29 639 -17 915
rect 17 639 29 915
rect -29 627 29 639
rect 389 915 447 927
rect 389 639 401 915
rect 435 639 447 915
rect 389 627 447 639
rect 807 915 865 927
rect 807 639 819 915
rect 853 639 865 915
rect 807 627 865 639
rect 1225 915 1283 927
rect 1225 639 1237 915
rect 1271 639 1283 915
rect 1225 627 1283 639
rect 1643 915 1701 927
rect 1643 639 1655 915
rect 1689 639 1701 915
rect 1643 627 1701 639
rect 2061 915 2119 927
rect 2061 639 2073 915
rect 2107 639 2119 915
rect 2061 627 2119 639
rect -2119 397 -2061 409
rect -2119 121 -2107 397
rect -2073 121 -2061 397
rect -2119 109 -2061 121
rect -1701 397 -1643 409
rect -1701 121 -1689 397
rect -1655 121 -1643 397
rect -1701 109 -1643 121
rect -1283 397 -1225 409
rect -1283 121 -1271 397
rect -1237 121 -1225 397
rect -1283 109 -1225 121
rect -865 397 -807 409
rect -865 121 -853 397
rect -819 121 -807 397
rect -865 109 -807 121
rect -447 397 -389 409
rect -447 121 -435 397
rect -401 121 -389 397
rect -447 109 -389 121
rect -29 397 29 409
rect -29 121 -17 397
rect 17 121 29 397
rect -29 109 29 121
rect 389 397 447 409
rect 389 121 401 397
rect 435 121 447 397
rect 389 109 447 121
rect 807 397 865 409
rect 807 121 819 397
rect 853 121 865 397
rect 807 109 865 121
rect 1225 397 1283 409
rect 1225 121 1237 397
rect 1271 121 1283 397
rect 1225 109 1283 121
rect 1643 397 1701 409
rect 1643 121 1655 397
rect 1689 121 1701 397
rect 1643 109 1701 121
rect 2061 397 2119 409
rect 2061 121 2073 397
rect 2107 121 2119 397
rect 2061 109 2119 121
rect -2119 -121 -2061 -109
rect -2119 -397 -2107 -121
rect -2073 -397 -2061 -121
rect -2119 -409 -2061 -397
rect -1701 -121 -1643 -109
rect -1701 -397 -1689 -121
rect -1655 -397 -1643 -121
rect -1701 -409 -1643 -397
rect -1283 -121 -1225 -109
rect -1283 -397 -1271 -121
rect -1237 -397 -1225 -121
rect -1283 -409 -1225 -397
rect -865 -121 -807 -109
rect -865 -397 -853 -121
rect -819 -397 -807 -121
rect -865 -409 -807 -397
rect -447 -121 -389 -109
rect -447 -397 -435 -121
rect -401 -397 -389 -121
rect -447 -409 -389 -397
rect -29 -121 29 -109
rect -29 -397 -17 -121
rect 17 -397 29 -121
rect -29 -409 29 -397
rect 389 -121 447 -109
rect 389 -397 401 -121
rect 435 -397 447 -121
rect 389 -409 447 -397
rect 807 -121 865 -109
rect 807 -397 819 -121
rect 853 -397 865 -121
rect 807 -409 865 -397
rect 1225 -121 1283 -109
rect 1225 -397 1237 -121
rect 1271 -397 1283 -121
rect 1225 -409 1283 -397
rect 1643 -121 1701 -109
rect 1643 -397 1655 -121
rect 1689 -397 1701 -121
rect 1643 -409 1701 -397
rect 2061 -121 2119 -109
rect 2061 -397 2073 -121
rect 2107 -397 2119 -121
rect 2061 -409 2119 -397
rect -2119 -639 -2061 -627
rect -2119 -915 -2107 -639
rect -2073 -915 -2061 -639
rect -2119 -927 -2061 -915
rect -1701 -639 -1643 -627
rect -1701 -915 -1689 -639
rect -1655 -915 -1643 -639
rect -1701 -927 -1643 -915
rect -1283 -639 -1225 -627
rect -1283 -915 -1271 -639
rect -1237 -915 -1225 -639
rect -1283 -927 -1225 -915
rect -865 -639 -807 -627
rect -865 -915 -853 -639
rect -819 -915 -807 -639
rect -865 -927 -807 -915
rect -447 -639 -389 -627
rect -447 -915 -435 -639
rect -401 -915 -389 -639
rect -447 -927 -389 -915
rect -29 -639 29 -627
rect -29 -915 -17 -639
rect 17 -915 29 -639
rect -29 -927 29 -915
rect 389 -639 447 -627
rect 389 -915 401 -639
rect 435 -915 447 -639
rect 389 -927 447 -915
rect 807 -639 865 -627
rect 807 -915 819 -639
rect 853 -915 865 -639
rect 807 -927 865 -915
rect 1225 -639 1283 -627
rect 1225 -915 1237 -639
rect 1271 -915 1283 -639
rect 1225 -927 1283 -915
rect 1643 -639 1701 -627
rect 1643 -915 1655 -639
rect 1689 -915 1701 -639
rect 1643 -927 1701 -915
rect 2061 -639 2119 -627
rect 2061 -915 2073 -639
rect 2107 -915 2119 -639
rect 2061 -927 2119 -915
rect -2119 -1157 -2061 -1145
rect -2119 -1433 -2107 -1157
rect -2073 -1433 -2061 -1157
rect -2119 -1445 -2061 -1433
rect -1701 -1157 -1643 -1145
rect -1701 -1433 -1689 -1157
rect -1655 -1433 -1643 -1157
rect -1701 -1445 -1643 -1433
rect -1283 -1157 -1225 -1145
rect -1283 -1433 -1271 -1157
rect -1237 -1433 -1225 -1157
rect -1283 -1445 -1225 -1433
rect -865 -1157 -807 -1145
rect -865 -1433 -853 -1157
rect -819 -1433 -807 -1157
rect -865 -1445 -807 -1433
rect -447 -1157 -389 -1145
rect -447 -1433 -435 -1157
rect -401 -1433 -389 -1157
rect -447 -1445 -389 -1433
rect -29 -1157 29 -1145
rect -29 -1433 -17 -1157
rect 17 -1433 29 -1157
rect -29 -1445 29 -1433
rect 389 -1157 447 -1145
rect 389 -1433 401 -1157
rect 435 -1433 447 -1157
rect 389 -1445 447 -1433
rect 807 -1157 865 -1145
rect 807 -1433 819 -1157
rect 853 -1433 865 -1157
rect 807 -1445 865 -1433
rect 1225 -1157 1283 -1145
rect 1225 -1433 1237 -1157
rect 1271 -1433 1283 -1157
rect 1225 -1445 1283 -1433
rect 1643 -1157 1701 -1145
rect 1643 -1433 1655 -1157
rect 1689 -1433 1701 -1157
rect 1643 -1445 1701 -1433
rect 2061 -1157 2119 -1145
rect 2061 -1433 2073 -1157
rect 2107 -1433 2119 -1157
rect 2061 -1445 2119 -1433
rect -2119 -1675 -2061 -1663
rect -2119 -1951 -2107 -1675
rect -2073 -1951 -2061 -1675
rect -2119 -1963 -2061 -1951
rect -1701 -1675 -1643 -1663
rect -1701 -1951 -1689 -1675
rect -1655 -1951 -1643 -1675
rect -1701 -1963 -1643 -1951
rect -1283 -1675 -1225 -1663
rect -1283 -1951 -1271 -1675
rect -1237 -1951 -1225 -1675
rect -1283 -1963 -1225 -1951
rect -865 -1675 -807 -1663
rect -865 -1951 -853 -1675
rect -819 -1951 -807 -1675
rect -865 -1963 -807 -1951
rect -447 -1675 -389 -1663
rect -447 -1951 -435 -1675
rect -401 -1951 -389 -1675
rect -447 -1963 -389 -1951
rect -29 -1675 29 -1663
rect -29 -1951 -17 -1675
rect 17 -1951 29 -1675
rect -29 -1963 29 -1951
rect 389 -1675 447 -1663
rect 389 -1951 401 -1675
rect 435 -1951 447 -1675
rect 389 -1963 447 -1951
rect 807 -1675 865 -1663
rect 807 -1951 819 -1675
rect 853 -1951 865 -1675
rect 807 -1963 865 -1951
rect 1225 -1675 1283 -1663
rect 1225 -1951 1237 -1675
rect 1271 -1951 1283 -1675
rect 1225 -1963 1283 -1951
rect 1643 -1675 1701 -1663
rect 1643 -1951 1655 -1675
rect 1689 -1951 1701 -1675
rect 1643 -1963 1701 -1951
rect 2061 -1675 2119 -1663
rect 2061 -1951 2073 -1675
rect 2107 -1951 2119 -1675
rect 2061 -1963 2119 -1951
rect -2119 -2193 -2061 -2181
rect -2119 -2469 -2107 -2193
rect -2073 -2469 -2061 -2193
rect -2119 -2481 -2061 -2469
rect -1701 -2193 -1643 -2181
rect -1701 -2469 -1689 -2193
rect -1655 -2469 -1643 -2193
rect -1701 -2481 -1643 -2469
rect -1283 -2193 -1225 -2181
rect -1283 -2469 -1271 -2193
rect -1237 -2469 -1225 -2193
rect -1283 -2481 -1225 -2469
rect -865 -2193 -807 -2181
rect -865 -2469 -853 -2193
rect -819 -2469 -807 -2193
rect -865 -2481 -807 -2469
rect -447 -2193 -389 -2181
rect -447 -2469 -435 -2193
rect -401 -2469 -389 -2193
rect -447 -2481 -389 -2469
rect -29 -2193 29 -2181
rect -29 -2469 -17 -2193
rect 17 -2469 29 -2193
rect -29 -2481 29 -2469
rect 389 -2193 447 -2181
rect 389 -2469 401 -2193
rect 435 -2469 447 -2193
rect 389 -2481 447 -2469
rect 807 -2193 865 -2181
rect 807 -2469 819 -2193
rect 853 -2469 865 -2193
rect 807 -2481 865 -2469
rect 1225 -2193 1283 -2181
rect 1225 -2469 1237 -2193
rect 1271 -2469 1283 -2193
rect 1225 -2481 1283 -2469
rect 1643 -2193 1701 -2181
rect 1643 -2469 1655 -2193
rect 1689 -2469 1701 -2193
rect 1643 -2481 1701 -2469
rect 2061 -2193 2119 -2181
rect 2061 -2469 2073 -2193
rect 2107 -2469 2119 -2193
rect 2061 -2481 2119 -2469
<< ndiffc >>
rect -2107 2193 -2073 2469
rect -1689 2193 -1655 2469
rect -1271 2193 -1237 2469
rect -853 2193 -819 2469
rect -435 2193 -401 2469
rect -17 2193 17 2469
rect 401 2193 435 2469
rect 819 2193 853 2469
rect 1237 2193 1271 2469
rect 1655 2193 1689 2469
rect 2073 2193 2107 2469
rect -2107 1675 -2073 1951
rect -1689 1675 -1655 1951
rect -1271 1675 -1237 1951
rect -853 1675 -819 1951
rect -435 1675 -401 1951
rect -17 1675 17 1951
rect 401 1675 435 1951
rect 819 1675 853 1951
rect 1237 1675 1271 1951
rect 1655 1675 1689 1951
rect 2073 1675 2107 1951
rect -2107 1157 -2073 1433
rect -1689 1157 -1655 1433
rect -1271 1157 -1237 1433
rect -853 1157 -819 1433
rect -435 1157 -401 1433
rect -17 1157 17 1433
rect 401 1157 435 1433
rect 819 1157 853 1433
rect 1237 1157 1271 1433
rect 1655 1157 1689 1433
rect 2073 1157 2107 1433
rect -2107 639 -2073 915
rect -1689 639 -1655 915
rect -1271 639 -1237 915
rect -853 639 -819 915
rect -435 639 -401 915
rect -17 639 17 915
rect 401 639 435 915
rect 819 639 853 915
rect 1237 639 1271 915
rect 1655 639 1689 915
rect 2073 639 2107 915
rect -2107 121 -2073 397
rect -1689 121 -1655 397
rect -1271 121 -1237 397
rect -853 121 -819 397
rect -435 121 -401 397
rect -17 121 17 397
rect 401 121 435 397
rect 819 121 853 397
rect 1237 121 1271 397
rect 1655 121 1689 397
rect 2073 121 2107 397
rect -2107 -397 -2073 -121
rect -1689 -397 -1655 -121
rect -1271 -397 -1237 -121
rect -853 -397 -819 -121
rect -435 -397 -401 -121
rect -17 -397 17 -121
rect 401 -397 435 -121
rect 819 -397 853 -121
rect 1237 -397 1271 -121
rect 1655 -397 1689 -121
rect 2073 -397 2107 -121
rect -2107 -915 -2073 -639
rect -1689 -915 -1655 -639
rect -1271 -915 -1237 -639
rect -853 -915 -819 -639
rect -435 -915 -401 -639
rect -17 -915 17 -639
rect 401 -915 435 -639
rect 819 -915 853 -639
rect 1237 -915 1271 -639
rect 1655 -915 1689 -639
rect 2073 -915 2107 -639
rect -2107 -1433 -2073 -1157
rect -1689 -1433 -1655 -1157
rect -1271 -1433 -1237 -1157
rect -853 -1433 -819 -1157
rect -435 -1433 -401 -1157
rect -17 -1433 17 -1157
rect 401 -1433 435 -1157
rect 819 -1433 853 -1157
rect 1237 -1433 1271 -1157
rect 1655 -1433 1689 -1157
rect 2073 -1433 2107 -1157
rect -2107 -1951 -2073 -1675
rect -1689 -1951 -1655 -1675
rect -1271 -1951 -1237 -1675
rect -853 -1951 -819 -1675
rect -435 -1951 -401 -1675
rect -17 -1951 17 -1675
rect 401 -1951 435 -1675
rect 819 -1951 853 -1675
rect 1237 -1951 1271 -1675
rect 1655 -1951 1689 -1675
rect 2073 -1951 2107 -1675
rect -2107 -2469 -2073 -2193
rect -1689 -2469 -1655 -2193
rect -1271 -2469 -1237 -2193
rect -853 -2469 -819 -2193
rect -435 -2469 -401 -2193
rect -17 -2469 17 -2193
rect 401 -2469 435 -2193
rect 819 -2469 853 -2193
rect 1237 -2469 1271 -2193
rect 1655 -2469 1689 -2193
rect 2073 -2469 2107 -2193
<< psubdiff >>
rect -2221 2621 -2125 2655
rect 2125 2621 2221 2655
rect -2221 2559 -2187 2621
rect 2187 2559 2221 2621
rect -2221 -2621 -2187 -2559
rect 2187 -2621 2221 -2559
rect -2221 -2655 -2125 -2621
rect 2125 -2655 2221 -2621
<< psubdiffcont >>
rect -2125 2621 2125 2655
rect -2221 -2559 -2187 2559
rect 2187 -2559 2221 2559
rect -2125 -2655 2125 -2621
<< poly >>
rect -2061 2553 -1701 2569
rect -2061 2519 -2045 2553
rect -1717 2519 -1701 2553
rect -2061 2481 -1701 2519
rect -1643 2553 -1283 2569
rect -1643 2519 -1627 2553
rect -1299 2519 -1283 2553
rect -1643 2481 -1283 2519
rect -1225 2553 -865 2569
rect -1225 2519 -1209 2553
rect -881 2519 -865 2553
rect -1225 2481 -865 2519
rect -807 2553 -447 2569
rect -807 2519 -791 2553
rect -463 2519 -447 2553
rect -807 2481 -447 2519
rect -389 2553 -29 2569
rect -389 2519 -373 2553
rect -45 2519 -29 2553
rect -389 2481 -29 2519
rect 29 2553 389 2569
rect 29 2519 45 2553
rect 373 2519 389 2553
rect 29 2481 389 2519
rect 447 2553 807 2569
rect 447 2519 463 2553
rect 791 2519 807 2553
rect 447 2481 807 2519
rect 865 2553 1225 2569
rect 865 2519 881 2553
rect 1209 2519 1225 2553
rect 865 2481 1225 2519
rect 1283 2553 1643 2569
rect 1283 2519 1299 2553
rect 1627 2519 1643 2553
rect 1283 2481 1643 2519
rect 1701 2553 2061 2569
rect 1701 2519 1717 2553
rect 2045 2519 2061 2553
rect 1701 2481 2061 2519
rect -2061 2143 -1701 2181
rect -2061 2109 -2045 2143
rect -1717 2109 -1701 2143
rect -2061 2093 -1701 2109
rect -1643 2143 -1283 2181
rect -1643 2109 -1627 2143
rect -1299 2109 -1283 2143
rect -1643 2093 -1283 2109
rect -1225 2143 -865 2181
rect -1225 2109 -1209 2143
rect -881 2109 -865 2143
rect -1225 2093 -865 2109
rect -807 2143 -447 2181
rect -807 2109 -791 2143
rect -463 2109 -447 2143
rect -807 2093 -447 2109
rect -389 2143 -29 2181
rect -389 2109 -373 2143
rect -45 2109 -29 2143
rect -389 2093 -29 2109
rect 29 2143 389 2181
rect 29 2109 45 2143
rect 373 2109 389 2143
rect 29 2093 389 2109
rect 447 2143 807 2181
rect 447 2109 463 2143
rect 791 2109 807 2143
rect 447 2093 807 2109
rect 865 2143 1225 2181
rect 865 2109 881 2143
rect 1209 2109 1225 2143
rect 865 2093 1225 2109
rect 1283 2143 1643 2181
rect 1283 2109 1299 2143
rect 1627 2109 1643 2143
rect 1283 2093 1643 2109
rect 1701 2143 2061 2181
rect 1701 2109 1717 2143
rect 2045 2109 2061 2143
rect 1701 2093 2061 2109
rect -2061 2035 -1701 2051
rect -2061 2001 -2045 2035
rect -1717 2001 -1701 2035
rect -2061 1963 -1701 2001
rect -1643 2035 -1283 2051
rect -1643 2001 -1627 2035
rect -1299 2001 -1283 2035
rect -1643 1963 -1283 2001
rect -1225 2035 -865 2051
rect -1225 2001 -1209 2035
rect -881 2001 -865 2035
rect -1225 1963 -865 2001
rect -807 2035 -447 2051
rect -807 2001 -791 2035
rect -463 2001 -447 2035
rect -807 1963 -447 2001
rect -389 2035 -29 2051
rect -389 2001 -373 2035
rect -45 2001 -29 2035
rect -389 1963 -29 2001
rect 29 2035 389 2051
rect 29 2001 45 2035
rect 373 2001 389 2035
rect 29 1963 389 2001
rect 447 2035 807 2051
rect 447 2001 463 2035
rect 791 2001 807 2035
rect 447 1963 807 2001
rect 865 2035 1225 2051
rect 865 2001 881 2035
rect 1209 2001 1225 2035
rect 865 1963 1225 2001
rect 1283 2035 1643 2051
rect 1283 2001 1299 2035
rect 1627 2001 1643 2035
rect 1283 1963 1643 2001
rect 1701 2035 2061 2051
rect 1701 2001 1717 2035
rect 2045 2001 2061 2035
rect 1701 1963 2061 2001
rect -2061 1625 -1701 1663
rect -2061 1591 -2045 1625
rect -1717 1591 -1701 1625
rect -2061 1575 -1701 1591
rect -1643 1625 -1283 1663
rect -1643 1591 -1627 1625
rect -1299 1591 -1283 1625
rect -1643 1575 -1283 1591
rect -1225 1625 -865 1663
rect -1225 1591 -1209 1625
rect -881 1591 -865 1625
rect -1225 1575 -865 1591
rect -807 1625 -447 1663
rect -807 1591 -791 1625
rect -463 1591 -447 1625
rect -807 1575 -447 1591
rect -389 1625 -29 1663
rect -389 1591 -373 1625
rect -45 1591 -29 1625
rect -389 1575 -29 1591
rect 29 1625 389 1663
rect 29 1591 45 1625
rect 373 1591 389 1625
rect 29 1575 389 1591
rect 447 1625 807 1663
rect 447 1591 463 1625
rect 791 1591 807 1625
rect 447 1575 807 1591
rect 865 1625 1225 1663
rect 865 1591 881 1625
rect 1209 1591 1225 1625
rect 865 1575 1225 1591
rect 1283 1625 1643 1663
rect 1283 1591 1299 1625
rect 1627 1591 1643 1625
rect 1283 1575 1643 1591
rect 1701 1625 2061 1663
rect 1701 1591 1717 1625
rect 2045 1591 2061 1625
rect 1701 1575 2061 1591
rect -2061 1517 -1701 1533
rect -2061 1483 -2045 1517
rect -1717 1483 -1701 1517
rect -2061 1445 -1701 1483
rect -1643 1517 -1283 1533
rect -1643 1483 -1627 1517
rect -1299 1483 -1283 1517
rect -1643 1445 -1283 1483
rect -1225 1517 -865 1533
rect -1225 1483 -1209 1517
rect -881 1483 -865 1517
rect -1225 1445 -865 1483
rect -807 1517 -447 1533
rect -807 1483 -791 1517
rect -463 1483 -447 1517
rect -807 1445 -447 1483
rect -389 1517 -29 1533
rect -389 1483 -373 1517
rect -45 1483 -29 1517
rect -389 1445 -29 1483
rect 29 1517 389 1533
rect 29 1483 45 1517
rect 373 1483 389 1517
rect 29 1445 389 1483
rect 447 1517 807 1533
rect 447 1483 463 1517
rect 791 1483 807 1517
rect 447 1445 807 1483
rect 865 1517 1225 1533
rect 865 1483 881 1517
rect 1209 1483 1225 1517
rect 865 1445 1225 1483
rect 1283 1517 1643 1533
rect 1283 1483 1299 1517
rect 1627 1483 1643 1517
rect 1283 1445 1643 1483
rect 1701 1517 2061 1533
rect 1701 1483 1717 1517
rect 2045 1483 2061 1517
rect 1701 1445 2061 1483
rect -2061 1107 -1701 1145
rect -2061 1073 -2045 1107
rect -1717 1073 -1701 1107
rect -2061 1057 -1701 1073
rect -1643 1107 -1283 1145
rect -1643 1073 -1627 1107
rect -1299 1073 -1283 1107
rect -1643 1057 -1283 1073
rect -1225 1107 -865 1145
rect -1225 1073 -1209 1107
rect -881 1073 -865 1107
rect -1225 1057 -865 1073
rect -807 1107 -447 1145
rect -807 1073 -791 1107
rect -463 1073 -447 1107
rect -807 1057 -447 1073
rect -389 1107 -29 1145
rect -389 1073 -373 1107
rect -45 1073 -29 1107
rect -389 1057 -29 1073
rect 29 1107 389 1145
rect 29 1073 45 1107
rect 373 1073 389 1107
rect 29 1057 389 1073
rect 447 1107 807 1145
rect 447 1073 463 1107
rect 791 1073 807 1107
rect 447 1057 807 1073
rect 865 1107 1225 1145
rect 865 1073 881 1107
rect 1209 1073 1225 1107
rect 865 1057 1225 1073
rect 1283 1107 1643 1145
rect 1283 1073 1299 1107
rect 1627 1073 1643 1107
rect 1283 1057 1643 1073
rect 1701 1107 2061 1145
rect 1701 1073 1717 1107
rect 2045 1073 2061 1107
rect 1701 1057 2061 1073
rect -2061 999 -1701 1015
rect -2061 965 -2045 999
rect -1717 965 -1701 999
rect -2061 927 -1701 965
rect -1643 999 -1283 1015
rect -1643 965 -1627 999
rect -1299 965 -1283 999
rect -1643 927 -1283 965
rect -1225 999 -865 1015
rect -1225 965 -1209 999
rect -881 965 -865 999
rect -1225 927 -865 965
rect -807 999 -447 1015
rect -807 965 -791 999
rect -463 965 -447 999
rect -807 927 -447 965
rect -389 999 -29 1015
rect -389 965 -373 999
rect -45 965 -29 999
rect -389 927 -29 965
rect 29 999 389 1015
rect 29 965 45 999
rect 373 965 389 999
rect 29 927 389 965
rect 447 999 807 1015
rect 447 965 463 999
rect 791 965 807 999
rect 447 927 807 965
rect 865 999 1225 1015
rect 865 965 881 999
rect 1209 965 1225 999
rect 865 927 1225 965
rect 1283 999 1643 1015
rect 1283 965 1299 999
rect 1627 965 1643 999
rect 1283 927 1643 965
rect 1701 999 2061 1015
rect 1701 965 1717 999
rect 2045 965 2061 999
rect 1701 927 2061 965
rect -2061 589 -1701 627
rect -2061 555 -2045 589
rect -1717 555 -1701 589
rect -2061 539 -1701 555
rect -1643 589 -1283 627
rect -1643 555 -1627 589
rect -1299 555 -1283 589
rect -1643 539 -1283 555
rect -1225 589 -865 627
rect -1225 555 -1209 589
rect -881 555 -865 589
rect -1225 539 -865 555
rect -807 589 -447 627
rect -807 555 -791 589
rect -463 555 -447 589
rect -807 539 -447 555
rect -389 589 -29 627
rect -389 555 -373 589
rect -45 555 -29 589
rect -389 539 -29 555
rect 29 589 389 627
rect 29 555 45 589
rect 373 555 389 589
rect 29 539 389 555
rect 447 589 807 627
rect 447 555 463 589
rect 791 555 807 589
rect 447 539 807 555
rect 865 589 1225 627
rect 865 555 881 589
rect 1209 555 1225 589
rect 865 539 1225 555
rect 1283 589 1643 627
rect 1283 555 1299 589
rect 1627 555 1643 589
rect 1283 539 1643 555
rect 1701 589 2061 627
rect 1701 555 1717 589
rect 2045 555 2061 589
rect 1701 539 2061 555
rect -2061 481 -1701 497
rect -2061 447 -2045 481
rect -1717 447 -1701 481
rect -2061 409 -1701 447
rect -1643 481 -1283 497
rect -1643 447 -1627 481
rect -1299 447 -1283 481
rect -1643 409 -1283 447
rect -1225 481 -865 497
rect -1225 447 -1209 481
rect -881 447 -865 481
rect -1225 409 -865 447
rect -807 481 -447 497
rect -807 447 -791 481
rect -463 447 -447 481
rect -807 409 -447 447
rect -389 481 -29 497
rect -389 447 -373 481
rect -45 447 -29 481
rect -389 409 -29 447
rect 29 481 389 497
rect 29 447 45 481
rect 373 447 389 481
rect 29 409 389 447
rect 447 481 807 497
rect 447 447 463 481
rect 791 447 807 481
rect 447 409 807 447
rect 865 481 1225 497
rect 865 447 881 481
rect 1209 447 1225 481
rect 865 409 1225 447
rect 1283 481 1643 497
rect 1283 447 1299 481
rect 1627 447 1643 481
rect 1283 409 1643 447
rect 1701 481 2061 497
rect 1701 447 1717 481
rect 2045 447 2061 481
rect 1701 409 2061 447
rect -2061 71 -1701 109
rect -2061 37 -2045 71
rect -1717 37 -1701 71
rect -2061 21 -1701 37
rect -1643 71 -1283 109
rect -1643 37 -1627 71
rect -1299 37 -1283 71
rect -1643 21 -1283 37
rect -1225 71 -865 109
rect -1225 37 -1209 71
rect -881 37 -865 71
rect -1225 21 -865 37
rect -807 71 -447 109
rect -807 37 -791 71
rect -463 37 -447 71
rect -807 21 -447 37
rect -389 71 -29 109
rect -389 37 -373 71
rect -45 37 -29 71
rect -389 21 -29 37
rect 29 71 389 109
rect 29 37 45 71
rect 373 37 389 71
rect 29 21 389 37
rect 447 71 807 109
rect 447 37 463 71
rect 791 37 807 71
rect 447 21 807 37
rect 865 71 1225 109
rect 865 37 881 71
rect 1209 37 1225 71
rect 865 21 1225 37
rect 1283 71 1643 109
rect 1283 37 1299 71
rect 1627 37 1643 71
rect 1283 21 1643 37
rect 1701 71 2061 109
rect 1701 37 1717 71
rect 2045 37 2061 71
rect 1701 21 2061 37
rect -2061 -37 -1701 -21
rect -2061 -71 -2045 -37
rect -1717 -71 -1701 -37
rect -2061 -109 -1701 -71
rect -1643 -37 -1283 -21
rect -1643 -71 -1627 -37
rect -1299 -71 -1283 -37
rect -1643 -109 -1283 -71
rect -1225 -37 -865 -21
rect -1225 -71 -1209 -37
rect -881 -71 -865 -37
rect -1225 -109 -865 -71
rect -807 -37 -447 -21
rect -807 -71 -791 -37
rect -463 -71 -447 -37
rect -807 -109 -447 -71
rect -389 -37 -29 -21
rect -389 -71 -373 -37
rect -45 -71 -29 -37
rect -389 -109 -29 -71
rect 29 -37 389 -21
rect 29 -71 45 -37
rect 373 -71 389 -37
rect 29 -109 389 -71
rect 447 -37 807 -21
rect 447 -71 463 -37
rect 791 -71 807 -37
rect 447 -109 807 -71
rect 865 -37 1225 -21
rect 865 -71 881 -37
rect 1209 -71 1225 -37
rect 865 -109 1225 -71
rect 1283 -37 1643 -21
rect 1283 -71 1299 -37
rect 1627 -71 1643 -37
rect 1283 -109 1643 -71
rect 1701 -37 2061 -21
rect 1701 -71 1717 -37
rect 2045 -71 2061 -37
rect 1701 -109 2061 -71
rect -2061 -447 -1701 -409
rect -2061 -481 -2045 -447
rect -1717 -481 -1701 -447
rect -2061 -497 -1701 -481
rect -1643 -447 -1283 -409
rect -1643 -481 -1627 -447
rect -1299 -481 -1283 -447
rect -1643 -497 -1283 -481
rect -1225 -447 -865 -409
rect -1225 -481 -1209 -447
rect -881 -481 -865 -447
rect -1225 -497 -865 -481
rect -807 -447 -447 -409
rect -807 -481 -791 -447
rect -463 -481 -447 -447
rect -807 -497 -447 -481
rect -389 -447 -29 -409
rect -389 -481 -373 -447
rect -45 -481 -29 -447
rect -389 -497 -29 -481
rect 29 -447 389 -409
rect 29 -481 45 -447
rect 373 -481 389 -447
rect 29 -497 389 -481
rect 447 -447 807 -409
rect 447 -481 463 -447
rect 791 -481 807 -447
rect 447 -497 807 -481
rect 865 -447 1225 -409
rect 865 -481 881 -447
rect 1209 -481 1225 -447
rect 865 -497 1225 -481
rect 1283 -447 1643 -409
rect 1283 -481 1299 -447
rect 1627 -481 1643 -447
rect 1283 -497 1643 -481
rect 1701 -447 2061 -409
rect 1701 -481 1717 -447
rect 2045 -481 2061 -447
rect 1701 -497 2061 -481
rect -2061 -555 -1701 -539
rect -2061 -589 -2045 -555
rect -1717 -589 -1701 -555
rect -2061 -627 -1701 -589
rect -1643 -555 -1283 -539
rect -1643 -589 -1627 -555
rect -1299 -589 -1283 -555
rect -1643 -627 -1283 -589
rect -1225 -555 -865 -539
rect -1225 -589 -1209 -555
rect -881 -589 -865 -555
rect -1225 -627 -865 -589
rect -807 -555 -447 -539
rect -807 -589 -791 -555
rect -463 -589 -447 -555
rect -807 -627 -447 -589
rect -389 -555 -29 -539
rect -389 -589 -373 -555
rect -45 -589 -29 -555
rect -389 -627 -29 -589
rect 29 -555 389 -539
rect 29 -589 45 -555
rect 373 -589 389 -555
rect 29 -627 389 -589
rect 447 -555 807 -539
rect 447 -589 463 -555
rect 791 -589 807 -555
rect 447 -627 807 -589
rect 865 -555 1225 -539
rect 865 -589 881 -555
rect 1209 -589 1225 -555
rect 865 -627 1225 -589
rect 1283 -555 1643 -539
rect 1283 -589 1299 -555
rect 1627 -589 1643 -555
rect 1283 -627 1643 -589
rect 1701 -555 2061 -539
rect 1701 -589 1717 -555
rect 2045 -589 2061 -555
rect 1701 -627 2061 -589
rect -2061 -965 -1701 -927
rect -2061 -999 -2045 -965
rect -1717 -999 -1701 -965
rect -2061 -1015 -1701 -999
rect -1643 -965 -1283 -927
rect -1643 -999 -1627 -965
rect -1299 -999 -1283 -965
rect -1643 -1015 -1283 -999
rect -1225 -965 -865 -927
rect -1225 -999 -1209 -965
rect -881 -999 -865 -965
rect -1225 -1015 -865 -999
rect -807 -965 -447 -927
rect -807 -999 -791 -965
rect -463 -999 -447 -965
rect -807 -1015 -447 -999
rect -389 -965 -29 -927
rect -389 -999 -373 -965
rect -45 -999 -29 -965
rect -389 -1015 -29 -999
rect 29 -965 389 -927
rect 29 -999 45 -965
rect 373 -999 389 -965
rect 29 -1015 389 -999
rect 447 -965 807 -927
rect 447 -999 463 -965
rect 791 -999 807 -965
rect 447 -1015 807 -999
rect 865 -965 1225 -927
rect 865 -999 881 -965
rect 1209 -999 1225 -965
rect 865 -1015 1225 -999
rect 1283 -965 1643 -927
rect 1283 -999 1299 -965
rect 1627 -999 1643 -965
rect 1283 -1015 1643 -999
rect 1701 -965 2061 -927
rect 1701 -999 1717 -965
rect 2045 -999 2061 -965
rect 1701 -1015 2061 -999
rect -2061 -1073 -1701 -1057
rect -2061 -1107 -2045 -1073
rect -1717 -1107 -1701 -1073
rect -2061 -1145 -1701 -1107
rect -1643 -1073 -1283 -1057
rect -1643 -1107 -1627 -1073
rect -1299 -1107 -1283 -1073
rect -1643 -1145 -1283 -1107
rect -1225 -1073 -865 -1057
rect -1225 -1107 -1209 -1073
rect -881 -1107 -865 -1073
rect -1225 -1145 -865 -1107
rect -807 -1073 -447 -1057
rect -807 -1107 -791 -1073
rect -463 -1107 -447 -1073
rect -807 -1145 -447 -1107
rect -389 -1073 -29 -1057
rect -389 -1107 -373 -1073
rect -45 -1107 -29 -1073
rect -389 -1145 -29 -1107
rect 29 -1073 389 -1057
rect 29 -1107 45 -1073
rect 373 -1107 389 -1073
rect 29 -1145 389 -1107
rect 447 -1073 807 -1057
rect 447 -1107 463 -1073
rect 791 -1107 807 -1073
rect 447 -1145 807 -1107
rect 865 -1073 1225 -1057
rect 865 -1107 881 -1073
rect 1209 -1107 1225 -1073
rect 865 -1145 1225 -1107
rect 1283 -1073 1643 -1057
rect 1283 -1107 1299 -1073
rect 1627 -1107 1643 -1073
rect 1283 -1145 1643 -1107
rect 1701 -1073 2061 -1057
rect 1701 -1107 1717 -1073
rect 2045 -1107 2061 -1073
rect 1701 -1145 2061 -1107
rect -2061 -1483 -1701 -1445
rect -2061 -1517 -2045 -1483
rect -1717 -1517 -1701 -1483
rect -2061 -1533 -1701 -1517
rect -1643 -1483 -1283 -1445
rect -1643 -1517 -1627 -1483
rect -1299 -1517 -1283 -1483
rect -1643 -1533 -1283 -1517
rect -1225 -1483 -865 -1445
rect -1225 -1517 -1209 -1483
rect -881 -1517 -865 -1483
rect -1225 -1533 -865 -1517
rect -807 -1483 -447 -1445
rect -807 -1517 -791 -1483
rect -463 -1517 -447 -1483
rect -807 -1533 -447 -1517
rect -389 -1483 -29 -1445
rect -389 -1517 -373 -1483
rect -45 -1517 -29 -1483
rect -389 -1533 -29 -1517
rect 29 -1483 389 -1445
rect 29 -1517 45 -1483
rect 373 -1517 389 -1483
rect 29 -1533 389 -1517
rect 447 -1483 807 -1445
rect 447 -1517 463 -1483
rect 791 -1517 807 -1483
rect 447 -1533 807 -1517
rect 865 -1483 1225 -1445
rect 865 -1517 881 -1483
rect 1209 -1517 1225 -1483
rect 865 -1533 1225 -1517
rect 1283 -1483 1643 -1445
rect 1283 -1517 1299 -1483
rect 1627 -1517 1643 -1483
rect 1283 -1533 1643 -1517
rect 1701 -1483 2061 -1445
rect 1701 -1517 1717 -1483
rect 2045 -1517 2061 -1483
rect 1701 -1533 2061 -1517
rect -2061 -1591 -1701 -1575
rect -2061 -1625 -2045 -1591
rect -1717 -1625 -1701 -1591
rect -2061 -1663 -1701 -1625
rect -1643 -1591 -1283 -1575
rect -1643 -1625 -1627 -1591
rect -1299 -1625 -1283 -1591
rect -1643 -1663 -1283 -1625
rect -1225 -1591 -865 -1575
rect -1225 -1625 -1209 -1591
rect -881 -1625 -865 -1591
rect -1225 -1663 -865 -1625
rect -807 -1591 -447 -1575
rect -807 -1625 -791 -1591
rect -463 -1625 -447 -1591
rect -807 -1663 -447 -1625
rect -389 -1591 -29 -1575
rect -389 -1625 -373 -1591
rect -45 -1625 -29 -1591
rect -389 -1663 -29 -1625
rect 29 -1591 389 -1575
rect 29 -1625 45 -1591
rect 373 -1625 389 -1591
rect 29 -1663 389 -1625
rect 447 -1591 807 -1575
rect 447 -1625 463 -1591
rect 791 -1625 807 -1591
rect 447 -1663 807 -1625
rect 865 -1591 1225 -1575
rect 865 -1625 881 -1591
rect 1209 -1625 1225 -1591
rect 865 -1663 1225 -1625
rect 1283 -1591 1643 -1575
rect 1283 -1625 1299 -1591
rect 1627 -1625 1643 -1591
rect 1283 -1663 1643 -1625
rect 1701 -1591 2061 -1575
rect 1701 -1625 1717 -1591
rect 2045 -1625 2061 -1591
rect 1701 -1663 2061 -1625
rect -2061 -2001 -1701 -1963
rect -2061 -2035 -2045 -2001
rect -1717 -2035 -1701 -2001
rect -2061 -2051 -1701 -2035
rect -1643 -2001 -1283 -1963
rect -1643 -2035 -1627 -2001
rect -1299 -2035 -1283 -2001
rect -1643 -2051 -1283 -2035
rect -1225 -2001 -865 -1963
rect -1225 -2035 -1209 -2001
rect -881 -2035 -865 -2001
rect -1225 -2051 -865 -2035
rect -807 -2001 -447 -1963
rect -807 -2035 -791 -2001
rect -463 -2035 -447 -2001
rect -807 -2051 -447 -2035
rect -389 -2001 -29 -1963
rect -389 -2035 -373 -2001
rect -45 -2035 -29 -2001
rect -389 -2051 -29 -2035
rect 29 -2001 389 -1963
rect 29 -2035 45 -2001
rect 373 -2035 389 -2001
rect 29 -2051 389 -2035
rect 447 -2001 807 -1963
rect 447 -2035 463 -2001
rect 791 -2035 807 -2001
rect 447 -2051 807 -2035
rect 865 -2001 1225 -1963
rect 865 -2035 881 -2001
rect 1209 -2035 1225 -2001
rect 865 -2051 1225 -2035
rect 1283 -2001 1643 -1963
rect 1283 -2035 1299 -2001
rect 1627 -2035 1643 -2001
rect 1283 -2051 1643 -2035
rect 1701 -2001 2061 -1963
rect 1701 -2035 1717 -2001
rect 2045 -2035 2061 -2001
rect 1701 -2051 2061 -2035
rect -2061 -2109 -1701 -2093
rect -2061 -2143 -2045 -2109
rect -1717 -2143 -1701 -2109
rect -2061 -2181 -1701 -2143
rect -1643 -2109 -1283 -2093
rect -1643 -2143 -1627 -2109
rect -1299 -2143 -1283 -2109
rect -1643 -2181 -1283 -2143
rect -1225 -2109 -865 -2093
rect -1225 -2143 -1209 -2109
rect -881 -2143 -865 -2109
rect -1225 -2181 -865 -2143
rect -807 -2109 -447 -2093
rect -807 -2143 -791 -2109
rect -463 -2143 -447 -2109
rect -807 -2181 -447 -2143
rect -389 -2109 -29 -2093
rect -389 -2143 -373 -2109
rect -45 -2143 -29 -2109
rect -389 -2181 -29 -2143
rect 29 -2109 389 -2093
rect 29 -2143 45 -2109
rect 373 -2143 389 -2109
rect 29 -2181 389 -2143
rect 447 -2109 807 -2093
rect 447 -2143 463 -2109
rect 791 -2143 807 -2109
rect 447 -2181 807 -2143
rect 865 -2109 1225 -2093
rect 865 -2143 881 -2109
rect 1209 -2143 1225 -2109
rect 865 -2181 1225 -2143
rect 1283 -2109 1643 -2093
rect 1283 -2143 1299 -2109
rect 1627 -2143 1643 -2109
rect 1283 -2181 1643 -2143
rect 1701 -2109 2061 -2093
rect 1701 -2143 1717 -2109
rect 2045 -2143 2061 -2109
rect 1701 -2181 2061 -2143
rect -2061 -2519 -1701 -2481
rect -2061 -2553 -2045 -2519
rect -1717 -2553 -1701 -2519
rect -2061 -2569 -1701 -2553
rect -1643 -2519 -1283 -2481
rect -1643 -2553 -1627 -2519
rect -1299 -2553 -1283 -2519
rect -1643 -2569 -1283 -2553
rect -1225 -2519 -865 -2481
rect -1225 -2553 -1209 -2519
rect -881 -2553 -865 -2519
rect -1225 -2569 -865 -2553
rect -807 -2519 -447 -2481
rect -807 -2553 -791 -2519
rect -463 -2553 -447 -2519
rect -807 -2569 -447 -2553
rect -389 -2519 -29 -2481
rect -389 -2553 -373 -2519
rect -45 -2553 -29 -2519
rect -389 -2569 -29 -2553
rect 29 -2519 389 -2481
rect 29 -2553 45 -2519
rect 373 -2553 389 -2519
rect 29 -2569 389 -2553
rect 447 -2519 807 -2481
rect 447 -2553 463 -2519
rect 791 -2553 807 -2519
rect 447 -2569 807 -2553
rect 865 -2519 1225 -2481
rect 865 -2553 881 -2519
rect 1209 -2553 1225 -2519
rect 865 -2569 1225 -2553
rect 1283 -2519 1643 -2481
rect 1283 -2553 1299 -2519
rect 1627 -2553 1643 -2519
rect 1283 -2569 1643 -2553
rect 1701 -2519 2061 -2481
rect 1701 -2553 1717 -2519
rect 2045 -2553 2061 -2519
rect 1701 -2569 2061 -2553
<< polycont >>
rect -2045 2519 -1717 2553
rect -1627 2519 -1299 2553
rect -1209 2519 -881 2553
rect -791 2519 -463 2553
rect -373 2519 -45 2553
rect 45 2519 373 2553
rect 463 2519 791 2553
rect 881 2519 1209 2553
rect 1299 2519 1627 2553
rect 1717 2519 2045 2553
rect -2045 2109 -1717 2143
rect -1627 2109 -1299 2143
rect -1209 2109 -881 2143
rect -791 2109 -463 2143
rect -373 2109 -45 2143
rect 45 2109 373 2143
rect 463 2109 791 2143
rect 881 2109 1209 2143
rect 1299 2109 1627 2143
rect 1717 2109 2045 2143
rect -2045 2001 -1717 2035
rect -1627 2001 -1299 2035
rect -1209 2001 -881 2035
rect -791 2001 -463 2035
rect -373 2001 -45 2035
rect 45 2001 373 2035
rect 463 2001 791 2035
rect 881 2001 1209 2035
rect 1299 2001 1627 2035
rect 1717 2001 2045 2035
rect -2045 1591 -1717 1625
rect -1627 1591 -1299 1625
rect -1209 1591 -881 1625
rect -791 1591 -463 1625
rect -373 1591 -45 1625
rect 45 1591 373 1625
rect 463 1591 791 1625
rect 881 1591 1209 1625
rect 1299 1591 1627 1625
rect 1717 1591 2045 1625
rect -2045 1483 -1717 1517
rect -1627 1483 -1299 1517
rect -1209 1483 -881 1517
rect -791 1483 -463 1517
rect -373 1483 -45 1517
rect 45 1483 373 1517
rect 463 1483 791 1517
rect 881 1483 1209 1517
rect 1299 1483 1627 1517
rect 1717 1483 2045 1517
rect -2045 1073 -1717 1107
rect -1627 1073 -1299 1107
rect -1209 1073 -881 1107
rect -791 1073 -463 1107
rect -373 1073 -45 1107
rect 45 1073 373 1107
rect 463 1073 791 1107
rect 881 1073 1209 1107
rect 1299 1073 1627 1107
rect 1717 1073 2045 1107
rect -2045 965 -1717 999
rect -1627 965 -1299 999
rect -1209 965 -881 999
rect -791 965 -463 999
rect -373 965 -45 999
rect 45 965 373 999
rect 463 965 791 999
rect 881 965 1209 999
rect 1299 965 1627 999
rect 1717 965 2045 999
rect -2045 555 -1717 589
rect -1627 555 -1299 589
rect -1209 555 -881 589
rect -791 555 -463 589
rect -373 555 -45 589
rect 45 555 373 589
rect 463 555 791 589
rect 881 555 1209 589
rect 1299 555 1627 589
rect 1717 555 2045 589
rect -2045 447 -1717 481
rect -1627 447 -1299 481
rect -1209 447 -881 481
rect -791 447 -463 481
rect -373 447 -45 481
rect 45 447 373 481
rect 463 447 791 481
rect 881 447 1209 481
rect 1299 447 1627 481
rect 1717 447 2045 481
rect -2045 37 -1717 71
rect -1627 37 -1299 71
rect -1209 37 -881 71
rect -791 37 -463 71
rect -373 37 -45 71
rect 45 37 373 71
rect 463 37 791 71
rect 881 37 1209 71
rect 1299 37 1627 71
rect 1717 37 2045 71
rect -2045 -71 -1717 -37
rect -1627 -71 -1299 -37
rect -1209 -71 -881 -37
rect -791 -71 -463 -37
rect -373 -71 -45 -37
rect 45 -71 373 -37
rect 463 -71 791 -37
rect 881 -71 1209 -37
rect 1299 -71 1627 -37
rect 1717 -71 2045 -37
rect -2045 -481 -1717 -447
rect -1627 -481 -1299 -447
rect -1209 -481 -881 -447
rect -791 -481 -463 -447
rect -373 -481 -45 -447
rect 45 -481 373 -447
rect 463 -481 791 -447
rect 881 -481 1209 -447
rect 1299 -481 1627 -447
rect 1717 -481 2045 -447
rect -2045 -589 -1717 -555
rect -1627 -589 -1299 -555
rect -1209 -589 -881 -555
rect -791 -589 -463 -555
rect -373 -589 -45 -555
rect 45 -589 373 -555
rect 463 -589 791 -555
rect 881 -589 1209 -555
rect 1299 -589 1627 -555
rect 1717 -589 2045 -555
rect -2045 -999 -1717 -965
rect -1627 -999 -1299 -965
rect -1209 -999 -881 -965
rect -791 -999 -463 -965
rect -373 -999 -45 -965
rect 45 -999 373 -965
rect 463 -999 791 -965
rect 881 -999 1209 -965
rect 1299 -999 1627 -965
rect 1717 -999 2045 -965
rect -2045 -1107 -1717 -1073
rect -1627 -1107 -1299 -1073
rect -1209 -1107 -881 -1073
rect -791 -1107 -463 -1073
rect -373 -1107 -45 -1073
rect 45 -1107 373 -1073
rect 463 -1107 791 -1073
rect 881 -1107 1209 -1073
rect 1299 -1107 1627 -1073
rect 1717 -1107 2045 -1073
rect -2045 -1517 -1717 -1483
rect -1627 -1517 -1299 -1483
rect -1209 -1517 -881 -1483
rect -791 -1517 -463 -1483
rect -373 -1517 -45 -1483
rect 45 -1517 373 -1483
rect 463 -1517 791 -1483
rect 881 -1517 1209 -1483
rect 1299 -1517 1627 -1483
rect 1717 -1517 2045 -1483
rect -2045 -1625 -1717 -1591
rect -1627 -1625 -1299 -1591
rect -1209 -1625 -881 -1591
rect -791 -1625 -463 -1591
rect -373 -1625 -45 -1591
rect 45 -1625 373 -1591
rect 463 -1625 791 -1591
rect 881 -1625 1209 -1591
rect 1299 -1625 1627 -1591
rect 1717 -1625 2045 -1591
rect -2045 -2035 -1717 -2001
rect -1627 -2035 -1299 -2001
rect -1209 -2035 -881 -2001
rect -791 -2035 -463 -2001
rect -373 -2035 -45 -2001
rect 45 -2035 373 -2001
rect 463 -2035 791 -2001
rect 881 -2035 1209 -2001
rect 1299 -2035 1627 -2001
rect 1717 -2035 2045 -2001
rect -2045 -2143 -1717 -2109
rect -1627 -2143 -1299 -2109
rect -1209 -2143 -881 -2109
rect -791 -2143 -463 -2109
rect -373 -2143 -45 -2109
rect 45 -2143 373 -2109
rect 463 -2143 791 -2109
rect 881 -2143 1209 -2109
rect 1299 -2143 1627 -2109
rect 1717 -2143 2045 -2109
rect -2045 -2553 -1717 -2519
rect -1627 -2553 -1299 -2519
rect -1209 -2553 -881 -2519
rect -791 -2553 -463 -2519
rect -373 -2553 -45 -2519
rect 45 -2553 373 -2519
rect 463 -2553 791 -2519
rect 881 -2553 1209 -2519
rect 1299 -2553 1627 -2519
rect 1717 -2553 2045 -2519
<< locali >>
rect -2221 2621 -2125 2655
rect 2125 2621 2221 2655
rect -2221 2559 -2187 2621
rect 2187 2559 2221 2621
rect -2061 2519 -2045 2553
rect -1717 2519 -1701 2553
rect -1643 2519 -1627 2553
rect -1299 2519 -1283 2553
rect -1225 2519 -1209 2553
rect -881 2519 -865 2553
rect -807 2519 -791 2553
rect -463 2519 -447 2553
rect -389 2519 -373 2553
rect -45 2519 -29 2553
rect 29 2519 45 2553
rect 373 2519 389 2553
rect 447 2519 463 2553
rect 791 2519 807 2553
rect 865 2519 881 2553
rect 1209 2519 1225 2553
rect 1283 2519 1299 2553
rect 1627 2519 1643 2553
rect 1701 2519 1717 2553
rect 2045 2519 2061 2553
rect -2107 2469 -2073 2485
rect -2107 2177 -2073 2193
rect -1689 2469 -1655 2485
rect -1689 2177 -1655 2193
rect -1271 2469 -1237 2485
rect -1271 2177 -1237 2193
rect -853 2469 -819 2485
rect -853 2177 -819 2193
rect -435 2469 -401 2485
rect -435 2177 -401 2193
rect -17 2469 17 2485
rect -17 2177 17 2193
rect 401 2469 435 2485
rect 401 2177 435 2193
rect 819 2469 853 2485
rect 819 2177 853 2193
rect 1237 2469 1271 2485
rect 1237 2177 1271 2193
rect 1655 2469 1689 2485
rect 1655 2177 1689 2193
rect 2073 2469 2107 2485
rect 2073 2177 2107 2193
rect -2061 2109 -2045 2143
rect -1717 2109 -1701 2143
rect -1643 2109 -1627 2143
rect -1299 2109 -1283 2143
rect -1225 2109 -1209 2143
rect -881 2109 -865 2143
rect -807 2109 -791 2143
rect -463 2109 -447 2143
rect -389 2109 -373 2143
rect -45 2109 -29 2143
rect 29 2109 45 2143
rect 373 2109 389 2143
rect 447 2109 463 2143
rect 791 2109 807 2143
rect 865 2109 881 2143
rect 1209 2109 1225 2143
rect 1283 2109 1299 2143
rect 1627 2109 1643 2143
rect 1701 2109 1717 2143
rect 2045 2109 2061 2143
rect -2061 2001 -2045 2035
rect -1717 2001 -1701 2035
rect -1643 2001 -1627 2035
rect -1299 2001 -1283 2035
rect -1225 2001 -1209 2035
rect -881 2001 -865 2035
rect -807 2001 -791 2035
rect -463 2001 -447 2035
rect -389 2001 -373 2035
rect -45 2001 -29 2035
rect 29 2001 45 2035
rect 373 2001 389 2035
rect 447 2001 463 2035
rect 791 2001 807 2035
rect 865 2001 881 2035
rect 1209 2001 1225 2035
rect 1283 2001 1299 2035
rect 1627 2001 1643 2035
rect 1701 2001 1717 2035
rect 2045 2001 2061 2035
rect -2107 1951 -2073 1967
rect -2107 1659 -2073 1675
rect -1689 1951 -1655 1967
rect -1689 1659 -1655 1675
rect -1271 1951 -1237 1967
rect -1271 1659 -1237 1675
rect -853 1951 -819 1967
rect -853 1659 -819 1675
rect -435 1951 -401 1967
rect -435 1659 -401 1675
rect -17 1951 17 1967
rect -17 1659 17 1675
rect 401 1951 435 1967
rect 401 1659 435 1675
rect 819 1951 853 1967
rect 819 1659 853 1675
rect 1237 1951 1271 1967
rect 1237 1659 1271 1675
rect 1655 1951 1689 1967
rect 1655 1659 1689 1675
rect 2073 1951 2107 1967
rect 2073 1659 2107 1675
rect -2061 1591 -2045 1625
rect -1717 1591 -1701 1625
rect -1643 1591 -1627 1625
rect -1299 1591 -1283 1625
rect -1225 1591 -1209 1625
rect -881 1591 -865 1625
rect -807 1591 -791 1625
rect -463 1591 -447 1625
rect -389 1591 -373 1625
rect -45 1591 -29 1625
rect 29 1591 45 1625
rect 373 1591 389 1625
rect 447 1591 463 1625
rect 791 1591 807 1625
rect 865 1591 881 1625
rect 1209 1591 1225 1625
rect 1283 1591 1299 1625
rect 1627 1591 1643 1625
rect 1701 1591 1717 1625
rect 2045 1591 2061 1625
rect -2061 1483 -2045 1517
rect -1717 1483 -1701 1517
rect -1643 1483 -1627 1517
rect -1299 1483 -1283 1517
rect -1225 1483 -1209 1517
rect -881 1483 -865 1517
rect -807 1483 -791 1517
rect -463 1483 -447 1517
rect -389 1483 -373 1517
rect -45 1483 -29 1517
rect 29 1483 45 1517
rect 373 1483 389 1517
rect 447 1483 463 1517
rect 791 1483 807 1517
rect 865 1483 881 1517
rect 1209 1483 1225 1517
rect 1283 1483 1299 1517
rect 1627 1483 1643 1517
rect 1701 1483 1717 1517
rect 2045 1483 2061 1517
rect -2107 1433 -2073 1449
rect -2107 1141 -2073 1157
rect -1689 1433 -1655 1449
rect -1689 1141 -1655 1157
rect -1271 1433 -1237 1449
rect -1271 1141 -1237 1157
rect -853 1433 -819 1449
rect -853 1141 -819 1157
rect -435 1433 -401 1449
rect -435 1141 -401 1157
rect -17 1433 17 1449
rect -17 1141 17 1157
rect 401 1433 435 1449
rect 401 1141 435 1157
rect 819 1433 853 1449
rect 819 1141 853 1157
rect 1237 1433 1271 1449
rect 1237 1141 1271 1157
rect 1655 1433 1689 1449
rect 1655 1141 1689 1157
rect 2073 1433 2107 1449
rect 2073 1141 2107 1157
rect -2061 1073 -2045 1107
rect -1717 1073 -1701 1107
rect -1643 1073 -1627 1107
rect -1299 1073 -1283 1107
rect -1225 1073 -1209 1107
rect -881 1073 -865 1107
rect -807 1073 -791 1107
rect -463 1073 -447 1107
rect -389 1073 -373 1107
rect -45 1073 -29 1107
rect 29 1073 45 1107
rect 373 1073 389 1107
rect 447 1073 463 1107
rect 791 1073 807 1107
rect 865 1073 881 1107
rect 1209 1073 1225 1107
rect 1283 1073 1299 1107
rect 1627 1073 1643 1107
rect 1701 1073 1717 1107
rect 2045 1073 2061 1107
rect -2061 965 -2045 999
rect -1717 965 -1701 999
rect -1643 965 -1627 999
rect -1299 965 -1283 999
rect -1225 965 -1209 999
rect -881 965 -865 999
rect -807 965 -791 999
rect -463 965 -447 999
rect -389 965 -373 999
rect -45 965 -29 999
rect 29 965 45 999
rect 373 965 389 999
rect 447 965 463 999
rect 791 965 807 999
rect 865 965 881 999
rect 1209 965 1225 999
rect 1283 965 1299 999
rect 1627 965 1643 999
rect 1701 965 1717 999
rect 2045 965 2061 999
rect -2107 915 -2073 931
rect -2107 623 -2073 639
rect -1689 915 -1655 931
rect -1689 623 -1655 639
rect -1271 915 -1237 931
rect -1271 623 -1237 639
rect -853 915 -819 931
rect -853 623 -819 639
rect -435 915 -401 931
rect -435 623 -401 639
rect -17 915 17 931
rect -17 623 17 639
rect 401 915 435 931
rect 401 623 435 639
rect 819 915 853 931
rect 819 623 853 639
rect 1237 915 1271 931
rect 1237 623 1271 639
rect 1655 915 1689 931
rect 1655 623 1689 639
rect 2073 915 2107 931
rect 2073 623 2107 639
rect -2061 555 -2045 589
rect -1717 555 -1701 589
rect -1643 555 -1627 589
rect -1299 555 -1283 589
rect -1225 555 -1209 589
rect -881 555 -865 589
rect -807 555 -791 589
rect -463 555 -447 589
rect -389 555 -373 589
rect -45 555 -29 589
rect 29 555 45 589
rect 373 555 389 589
rect 447 555 463 589
rect 791 555 807 589
rect 865 555 881 589
rect 1209 555 1225 589
rect 1283 555 1299 589
rect 1627 555 1643 589
rect 1701 555 1717 589
rect 2045 555 2061 589
rect -2061 447 -2045 481
rect -1717 447 -1701 481
rect -1643 447 -1627 481
rect -1299 447 -1283 481
rect -1225 447 -1209 481
rect -881 447 -865 481
rect -807 447 -791 481
rect -463 447 -447 481
rect -389 447 -373 481
rect -45 447 -29 481
rect 29 447 45 481
rect 373 447 389 481
rect 447 447 463 481
rect 791 447 807 481
rect 865 447 881 481
rect 1209 447 1225 481
rect 1283 447 1299 481
rect 1627 447 1643 481
rect 1701 447 1717 481
rect 2045 447 2061 481
rect -2107 397 -2073 413
rect -2107 105 -2073 121
rect -1689 397 -1655 413
rect -1689 105 -1655 121
rect -1271 397 -1237 413
rect -1271 105 -1237 121
rect -853 397 -819 413
rect -853 105 -819 121
rect -435 397 -401 413
rect -435 105 -401 121
rect -17 397 17 413
rect -17 105 17 121
rect 401 397 435 413
rect 401 105 435 121
rect 819 397 853 413
rect 819 105 853 121
rect 1237 397 1271 413
rect 1237 105 1271 121
rect 1655 397 1689 413
rect 1655 105 1689 121
rect 2073 397 2107 413
rect 2073 105 2107 121
rect -2061 37 -2045 71
rect -1717 37 -1701 71
rect -1643 37 -1627 71
rect -1299 37 -1283 71
rect -1225 37 -1209 71
rect -881 37 -865 71
rect -807 37 -791 71
rect -463 37 -447 71
rect -389 37 -373 71
rect -45 37 -29 71
rect 29 37 45 71
rect 373 37 389 71
rect 447 37 463 71
rect 791 37 807 71
rect 865 37 881 71
rect 1209 37 1225 71
rect 1283 37 1299 71
rect 1627 37 1643 71
rect 1701 37 1717 71
rect 2045 37 2061 71
rect -2061 -71 -2045 -37
rect -1717 -71 -1701 -37
rect -1643 -71 -1627 -37
rect -1299 -71 -1283 -37
rect -1225 -71 -1209 -37
rect -881 -71 -865 -37
rect -807 -71 -791 -37
rect -463 -71 -447 -37
rect -389 -71 -373 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 373 -71 389 -37
rect 447 -71 463 -37
rect 791 -71 807 -37
rect 865 -71 881 -37
rect 1209 -71 1225 -37
rect 1283 -71 1299 -37
rect 1627 -71 1643 -37
rect 1701 -71 1717 -37
rect 2045 -71 2061 -37
rect -2107 -121 -2073 -105
rect -2107 -413 -2073 -397
rect -1689 -121 -1655 -105
rect -1689 -413 -1655 -397
rect -1271 -121 -1237 -105
rect -1271 -413 -1237 -397
rect -853 -121 -819 -105
rect -853 -413 -819 -397
rect -435 -121 -401 -105
rect -435 -413 -401 -397
rect -17 -121 17 -105
rect -17 -413 17 -397
rect 401 -121 435 -105
rect 401 -413 435 -397
rect 819 -121 853 -105
rect 819 -413 853 -397
rect 1237 -121 1271 -105
rect 1237 -413 1271 -397
rect 1655 -121 1689 -105
rect 1655 -413 1689 -397
rect 2073 -121 2107 -105
rect 2073 -413 2107 -397
rect -2061 -481 -2045 -447
rect -1717 -481 -1701 -447
rect -1643 -481 -1627 -447
rect -1299 -481 -1283 -447
rect -1225 -481 -1209 -447
rect -881 -481 -865 -447
rect -807 -481 -791 -447
rect -463 -481 -447 -447
rect -389 -481 -373 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 373 -481 389 -447
rect 447 -481 463 -447
rect 791 -481 807 -447
rect 865 -481 881 -447
rect 1209 -481 1225 -447
rect 1283 -481 1299 -447
rect 1627 -481 1643 -447
rect 1701 -481 1717 -447
rect 2045 -481 2061 -447
rect -2061 -589 -2045 -555
rect -1717 -589 -1701 -555
rect -1643 -589 -1627 -555
rect -1299 -589 -1283 -555
rect -1225 -589 -1209 -555
rect -881 -589 -865 -555
rect -807 -589 -791 -555
rect -463 -589 -447 -555
rect -389 -589 -373 -555
rect -45 -589 -29 -555
rect 29 -589 45 -555
rect 373 -589 389 -555
rect 447 -589 463 -555
rect 791 -589 807 -555
rect 865 -589 881 -555
rect 1209 -589 1225 -555
rect 1283 -589 1299 -555
rect 1627 -589 1643 -555
rect 1701 -589 1717 -555
rect 2045 -589 2061 -555
rect -2107 -639 -2073 -623
rect -2107 -931 -2073 -915
rect -1689 -639 -1655 -623
rect -1689 -931 -1655 -915
rect -1271 -639 -1237 -623
rect -1271 -931 -1237 -915
rect -853 -639 -819 -623
rect -853 -931 -819 -915
rect -435 -639 -401 -623
rect -435 -931 -401 -915
rect -17 -639 17 -623
rect -17 -931 17 -915
rect 401 -639 435 -623
rect 401 -931 435 -915
rect 819 -639 853 -623
rect 819 -931 853 -915
rect 1237 -639 1271 -623
rect 1237 -931 1271 -915
rect 1655 -639 1689 -623
rect 1655 -931 1689 -915
rect 2073 -639 2107 -623
rect 2073 -931 2107 -915
rect -2061 -999 -2045 -965
rect -1717 -999 -1701 -965
rect -1643 -999 -1627 -965
rect -1299 -999 -1283 -965
rect -1225 -999 -1209 -965
rect -881 -999 -865 -965
rect -807 -999 -791 -965
rect -463 -999 -447 -965
rect -389 -999 -373 -965
rect -45 -999 -29 -965
rect 29 -999 45 -965
rect 373 -999 389 -965
rect 447 -999 463 -965
rect 791 -999 807 -965
rect 865 -999 881 -965
rect 1209 -999 1225 -965
rect 1283 -999 1299 -965
rect 1627 -999 1643 -965
rect 1701 -999 1717 -965
rect 2045 -999 2061 -965
rect -2061 -1107 -2045 -1073
rect -1717 -1107 -1701 -1073
rect -1643 -1107 -1627 -1073
rect -1299 -1107 -1283 -1073
rect -1225 -1107 -1209 -1073
rect -881 -1107 -865 -1073
rect -807 -1107 -791 -1073
rect -463 -1107 -447 -1073
rect -389 -1107 -373 -1073
rect -45 -1107 -29 -1073
rect 29 -1107 45 -1073
rect 373 -1107 389 -1073
rect 447 -1107 463 -1073
rect 791 -1107 807 -1073
rect 865 -1107 881 -1073
rect 1209 -1107 1225 -1073
rect 1283 -1107 1299 -1073
rect 1627 -1107 1643 -1073
rect 1701 -1107 1717 -1073
rect 2045 -1107 2061 -1073
rect -2107 -1157 -2073 -1141
rect -2107 -1449 -2073 -1433
rect -1689 -1157 -1655 -1141
rect -1689 -1449 -1655 -1433
rect -1271 -1157 -1237 -1141
rect -1271 -1449 -1237 -1433
rect -853 -1157 -819 -1141
rect -853 -1449 -819 -1433
rect -435 -1157 -401 -1141
rect -435 -1449 -401 -1433
rect -17 -1157 17 -1141
rect -17 -1449 17 -1433
rect 401 -1157 435 -1141
rect 401 -1449 435 -1433
rect 819 -1157 853 -1141
rect 819 -1449 853 -1433
rect 1237 -1157 1271 -1141
rect 1237 -1449 1271 -1433
rect 1655 -1157 1689 -1141
rect 1655 -1449 1689 -1433
rect 2073 -1157 2107 -1141
rect 2073 -1449 2107 -1433
rect -2061 -1517 -2045 -1483
rect -1717 -1517 -1701 -1483
rect -1643 -1517 -1627 -1483
rect -1299 -1517 -1283 -1483
rect -1225 -1517 -1209 -1483
rect -881 -1517 -865 -1483
rect -807 -1517 -791 -1483
rect -463 -1517 -447 -1483
rect -389 -1517 -373 -1483
rect -45 -1517 -29 -1483
rect 29 -1517 45 -1483
rect 373 -1517 389 -1483
rect 447 -1517 463 -1483
rect 791 -1517 807 -1483
rect 865 -1517 881 -1483
rect 1209 -1517 1225 -1483
rect 1283 -1517 1299 -1483
rect 1627 -1517 1643 -1483
rect 1701 -1517 1717 -1483
rect 2045 -1517 2061 -1483
rect -2061 -1625 -2045 -1591
rect -1717 -1625 -1701 -1591
rect -1643 -1625 -1627 -1591
rect -1299 -1625 -1283 -1591
rect -1225 -1625 -1209 -1591
rect -881 -1625 -865 -1591
rect -807 -1625 -791 -1591
rect -463 -1625 -447 -1591
rect -389 -1625 -373 -1591
rect -45 -1625 -29 -1591
rect 29 -1625 45 -1591
rect 373 -1625 389 -1591
rect 447 -1625 463 -1591
rect 791 -1625 807 -1591
rect 865 -1625 881 -1591
rect 1209 -1625 1225 -1591
rect 1283 -1625 1299 -1591
rect 1627 -1625 1643 -1591
rect 1701 -1625 1717 -1591
rect 2045 -1625 2061 -1591
rect -2107 -1675 -2073 -1659
rect -2107 -1967 -2073 -1951
rect -1689 -1675 -1655 -1659
rect -1689 -1967 -1655 -1951
rect -1271 -1675 -1237 -1659
rect -1271 -1967 -1237 -1951
rect -853 -1675 -819 -1659
rect -853 -1967 -819 -1951
rect -435 -1675 -401 -1659
rect -435 -1967 -401 -1951
rect -17 -1675 17 -1659
rect -17 -1967 17 -1951
rect 401 -1675 435 -1659
rect 401 -1967 435 -1951
rect 819 -1675 853 -1659
rect 819 -1967 853 -1951
rect 1237 -1675 1271 -1659
rect 1237 -1967 1271 -1951
rect 1655 -1675 1689 -1659
rect 1655 -1967 1689 -1951
rect 2073 -1675 2107 -1659
rect 2073 -1967 2107 -1951
rect -2061 -2035 -2045 -2001
rect -1717 -2035 -1701 -2001
rect -1643 -2035 -1627 -2001
rect -1299 -2035 -1283 -2001
rect -1225 -2035 -1209 -2001
rect -881 -2035 -865 -2001
rect -807 -2035 -791 -2001
rect -463 -2035 -447 -2001
rect -389 -2035 -373 -2001
rect -45 -2035 -29 -2001
rect 29 -2035 45 -2001
rect 373 -2035 389 -2001
rect 447 -2035 463 -2001
rect 791 -2035 807 -2001
rect 865 -2035 881 -2001
rect 1209 -2035 1225 -2001
rect 1283 -2035 1299 -2001
rect 1627 -2035 1643 -2001
rect 1701 -2035 1717 -2001
rect 2045 -2035 2061 -2001
rect -2061 -2143 -2045 -2109
rect -1717 -2143 -1701 -2109
rect -1643 -2143 -1627 -2109
rect -1299 -2143 -1283 -2109
rect -1225 -2143 -1209 -2109
rect -881 -2143 -865 -2109
rect -807 -2143 -791 -2109
rect -463 -2143 -447 -2109
rect -389 -2143 -373 -2109
rect -45 -2143 -29 -2109
rect 29 -2143 45 -2109
rect 373 -2143 389 -2109
rect 447 -2143 463 -2109
rect 791 -2143 807 -2109
rect 865 -2143 881 -2109
rect 1209 -2143 1225 -2109
rect 1283 -2143 1299 -2109
rect 1627 -2143 1643 -2109
rect 1701 -2143 1717 -2109
rect 2045 -2143 2061 -2109
rect -2107 -2193 -2073 -2177
rect -2107 -2485 -2073 -2469
rect -1689 -2193 -1655 -2177
rect -1689 -2485 -1655 -2469
rect -1271 -2193 -1237 -2177
rect -1271 -2485 -1237 -2469
rect -853 -2193 -819 -2177
rect -853 -2485 -819 -2469
rect -435 -2193 -401 -2177
rect -435 -2485 -401 -2469
rect -17 -2193 17 -2177
rect -17 -2485 17 -2469
rect 401 -2193 435 -2177
rect 401 -2485 435 -2469
rect 819 -2193 853 -2177
rect 819 -2485 853 -2469
rect 1237 -2193 1271 -2177
rect 1237 -2485 1271 -2469
rect 1655 -2193 1689 -2177
rect 1655 -2485 1689 -2469
rect 2073 -2193 2107 -2177
rect 2073 -2485 2107 -2469
rect -2061 -2553 -2045 -2519
rect -1717 -2553 -1701 -2519
rect -1643 -2553 -1627 -2519
rect -1299 -2553 -1283 -2519
rect -1225 -2553 -1209 -2519
rect -881 -2553 -865 -2519
rect -807 -2553 -791 -2519
rect -463 -2553 -447 -2519
rect -389 -2553 -373 -2519
rect -45 -2553 -29 -2519
rect 29 -2553 45 -2519
rect 373 -2553 389 -2519
rect 447 -2553 463 -2519
rect 791 -2553 807 -2519
rect 865 -2553 881 -2519
rect 1209 -2553 1225 -2519
rect 1283 -2553 1299 -2519
rect 1627 -2553 1643 -2519
rect 1701 -2553 1717 -2519
rect 2045 -2553 2061 -2519
rect -2221 -2621 -2187 -2559
rect 2187 -2621 2221 -2559
rect -2221 -2655 -2125 -2621
rect 2125 -2655 2221 -2621
<< viali >>
rect -2045 2519 -1717 2553
rect -1627 2519 -1299 2553
rect -1209 2519 -881 2553
rect -791 2519 -463 2553
rect -373 2519 -45 2553
rect 45 2519 373 2553
rect 463 2519 791 2553
rect 881 2519 1209 2553
rect 1299 2519 1627 2553
rect 1717 2519 2045 2553
rect -2107 2193 -2073 2469
rect -1689 2193 -1655 2469
rect -1271 2193 -1237 2469
rect -853 2193 -819 2469
rect -435 2193 -401 2469
rect -17 2193 17 2469
rect 401 2193 435 2469
rect 819 2193 853 2469
rect 1237 2193 1271 2469
rect 1655 2193 1689 2469
rect 2073 2193 2107 2469
rect -2045 2109 -1717 2143
rect -1627 2109 -1299 2143
rect -1209 2109 -881 2143
rect -791 2109 -463 2143
rect -373 2109 -45 2143
rect 45 2109 373 2143
rect 463 2109 791 2143
rect 881 2109 1209 2143
rect 1299 2109 1627 2143
rect 1717 2109 2045 2143
rect -2045 2001 -1717 2035
rect -1627 2001 -1299 2035
rect -1209 2001 -881 2035
rect -791 2001 -463 2035
rect -373 2001 -45 2035
rect 45 2001 373 2035
rect 463 2001 791 2035
rect 881 2001 1209 2035
rect 1299 2001 1627 2035
rect 1717 2001 2045 2035
rect -2107 1675 -2073 1951
rect -1689 1675 -1655 1951
rect -1271 1675 -1237 1951
rect -853 1675 -819 1951
rect -435 1675 -401 1951
rect -17 1675 17 1951
rect 401 1675 435 1951
rect 819 1675 853 1951
rect 1237 1675 1271 1951
rect 1655 1675 1689 1951
rect 2073 1675 2107 1951
rect -2045 1591 -1717 1625
rect -1627 1591 -1299 1625
rect -1209 1591 -881 1625
rect -791 1591 -463 1625
rect -373 1591 -45 1625
rect 45 1591 373 1625
rect 463 1591 791 1625
rect 881 1591 1209 1625
rect 1299 1591 1627 1625
rect 1717 1591 2045 1625
rect -2045 1483 -1717 1517
rect -1627 1483 -1299 1517
rect -1209 1483 -881 1517
rect -791 1483 -463 1517
rect -373 1483 -45 1517
rect 45 1483 373 1517
rect 463 1483 791 1517
rect 881 1483 1209 1517
rect 1299 1483 1627 1517
rect 1717 1483 2045 1517
rect -2107 1157 -2073 1433
rect -1689 1157 -1655 1433
rect -1271 1157 -1237 1433
rect -853 1157 -819 1433
rect -435 1157 -401 1433
rect -17 1157 17 1433
rect 401 1157 435 1433
rect 819 1157 853 1433
rect 1237 1157 1271 1433
rect 1655 1157 1689 1433
rect 2073 1157 2107 1433
rect -2045 1073 -1717 1107
rect -1627 1073 -1299 1107
rect -1209 1073 -881 1107
rect -791 1073 -463 1107
rect -373 1073 -45 1107
rect 45 1073 373 1107
rect 463 1073 791 1107
rect 881 1073 1209 1107
rect 1299 1073 1627 1107
rect 1717 1073 2045 1107
rect -2045 965 -1717 999
rect -1627 965 -1299 999
rect -1209 965 -881 999
rect -791 965 -463 999
rect -373 965 -45 999
rect 45 965 373 999
rect 463 965 791 999
rect 881 965 1209 999
rect 1299 965 1627 999
rect 1717 965 2045 999
rect -2107 639 -2073 915
rect -1689 639 -1655 915
rect -1271 639 -1237 915
rect -853 639 -819 915
rect -435 639 -401 915
rect -17 639 17 915
rect 401 639 435 915
rect 819 639 853 915
rect 1237 639 1271 915
rect 1655 639 1689 915
rect 2073 639 2107 915
rect -2045 555 -1717 589
rect -1627 555 -1299 589
rect -1209 555 -881 589
rect -791 555 -463 589
rect -373 555 -45 589
rect 45 555 373 589
rect 463 555 791 589
rect 881 555 1209 589
rect 1299 555 1627 589
rect 1717 555 2045 589
rect -2045 447 -1717 481
rect -1627 447 -1299 481
rect -1209 447 -881 481
rect -791 447 -463 481
rect -373 447 -45 481
rect 45 447 373 481
rect 463 447 791 481
rect 881 447 1209 481
rect 1299 447 1627 481
rect 1717 447 2045 481
rect -2107 121 -2073 397
rect -1689 121 -1655 397
rect -1271 121 -1237 397
rect -853 121 -819 397
rect -435 121 -401 397
rect -17 121 17 397
rect 401 121 435 397
rect 819 121 853 397
rect 1237 121 1271 397
rect 1655 121 1689 397
rect 2073 121 2107 397
rect -2045 37 -1717 71
rect -1627 37 -1299 71
rect -1209 37 -881 71
rect -791 37 -463 71
rect -373 37 -45 71
rect 45 37 373 71
rect 463 37 791 71
rect 881 37 1209 71
rect 1299 37 1627 71
rect 1717 37 2045 71
rect -2045 -71 -1717 -37
rect -1627 -71 -1299 -37
rect -1209 -71 -881 -37
rect -791 -71 -463 -37
rect -373 -71 -45 -37
rect 45 -71 373 -37
rect 463 -71 791 -37
rect 881 -71 1209 -37
rect 1299 -71 1627 -37
rect 1717 -71 2045 -37
rect -2107 -397 -2073 -121
rect -1689 -397 -1655 -121
rect -1271 -397 -1237 -121
rect -853 -397 -819 -121
rect -435 -397 -401 -121
rect -17 -397 17 -121
rect 401 -397 435 -121
rect 819 -397 853 -121
rect 1237 -397 1271 -121
rect 1655 -397 1689 -121
rect 2073 -397 2107 -121
rect -2045 -481 -1717 -447
rect -1627 -481 -1299 -447
rect -1209 -481 -881 -447
rect -791 -481 -463 -447
rect -373 -481 -45 -447
rect 45 -481 373 -447
rect 463 -481 791 -447
rect 881 -481 1209 -447
rect 1299 -481 1627 -447
rect 1717 -481 2045 -447
rect -2045 -589 -1717 -555
rect -1627 -589 -1299 -555
rect -1209 -589 -881 -555
rect -791 -589 -463 -555
rect -373 -589 -45 -555
rect 45 -589 373 -555
rect 463 -589 791 -555
rect 881 -589 1209 -555
rect 1299 -589 1627 -555
rect 1717 -589 2045 -555
rect -2107 -915 -2073 -639
rect -1689 -915 -1655 -639
rect -1271 -915 -1237 -639
rect -853 -915 -819 -639
rect -435 -915 -401 -639
rect -17 -915 17 -639
rect 401 -915 435 -639
rect 819 -915 853 -639
rect 1237 -915 1271 -639
rect 1655 -915 1689 -639
rect 2073 -915 2107 -639
rect -2045 -999 -1717 -965
rect -1627 -999 -1299 -965
rect -1209 -999 -881 -965
rect -791 -999 -463 -965
rect -373 -999 -45 -965
rect 45 -999 373 -965
rect 463 -999 791 -965
rect 881 -999 1209 -965
rect 1299 -999 1627 -965
rect 1717 -999 2045 -965
rect -2045 -1107 -1717 -1073
rect -1627 -1107 -1299 -1073
rect -1209 -1107 -881 -1073
rect -791 -1107 -463 -1073
rect -373 -1107 -45 -1073
rect 45 -1107 373 -1073
rect 463 -1107 791 -1073
rect 881 -1107 1209 -1073
rect 1299 -1107 1627 -1073
rect 1717 -1107 2045 -1073
rect -2107 -1433 -2073 -1157
rect -1689 -1433 -1655 -1157
rect -1271 -1433 -1237 -1157
rect -853 -1433 -819 -1157
rect -435 -1433 -401 -1157
rect -17 -1433 17 -1157
rect 401 -1433 435 -1157
rect 819 -1433 853 -1157
rect 1237 -1433 1271 -1157
rect 1655 -1433 1689 -1157
rect 2073 -1433 2107 -1157
rect -2045 -1517 -1717 -1483
rect -1627 -1517 -1299 -1483
rect -1209 -1517 -881 -1483
rect -791 -1517 -463 -1483
rect -373 -1517 -45 -1483
rect 45 -1517 373 -1483
rect 463 -1517 791 -1483
rect 881 -1517 1209 -1483
rect 1299 -1517 1627 -1483
rect 1717 -1517 2045 -1483
rect -2045 -1625 -1717 -1591
rect -1627 -1625 -1299 -1591
rect -1209 -1625 -881 -1591
rect -791 -1625 -463 -1591
rect -373 -1625 -45 -1591
rect 45 -1625 373 -1591
rect 463 -1625 791 -1591
rect 881 -1625 1209 -1591
rect 1299 -1625 1627 -1591
rect 1717 -1625 2045 -1591
rect -2107 -1951 -2073 -1675
rect -1689 -1951 -1655 -1675
rect -1271 -1951 -1237 -1675
rect -853 -1951 -819 -1675
rect -435 -1951 -401 -1675
rect -17 -1951 17 -1675
rect 401 -1951 435 -1675
rect 819 -1951 853 -1675
rect 1237 -1951 1271 -1675
rect 1655 -1951 1689 -1675
rect 2073 -1951 2107 -1675
rect -2045 -2035 -1717 -2001
rect -1627 -2035 -1299 -2001
rect -1209 -2035 -881 -2001
rect -791 -2035 -463 -2001
rect -373 -2035 -45 -2001
rect 45 -2035 373 -2001
rect 463 -2035 791 -2001
rect 881 -2035 1209 -2001
rect 1299 -2035 1627 -2001
rect 1717 -2035 2045 -2001
rect -2045 -2143 -1717 -2109
rect -1627 -2143 -1299 -2109
rect -1209 -2143 -881 -2109
rect -791 -2143 -463 -2109
rect -373 -2143 -45 -2109
rect 45 -2143 373 -2109
rect 463 -2143 791 -2109
rect 881 -2143 1209 -2109
rect 1299 -2143 1627 -2109
rect 1717 -2143 2045 -2109
rect -2107 -2469 -2073 -2193
rect -1689 -2469 -1655 -2193
rect -1271 -2469 -1237 -2193
rect -853 -2469 -819 -2193
rect -435 -2469 -401 -2193
rect -17 -2469 17 -2193
rect 401 -2469 435 -2193
rect 819 -2469 853 -2193
rect 1237 -2469 1271 -2193
rect 1655 -2469 1689 -2193
rect 2073 -2469 2107 -2193
rect -2045 -2553 -1717 -2519
rect -1627 -2553 -1299 -2519
rect -1209 -2553 -881 -2519
rect -791 -2553 -463 -2519
rect -373 -2553 -45 -2519
rect 45 -2553 373 -2519
rect 463 -2553 791 -2519
rect 881 -2553 1209 -2519
rect 1299 -2553 1627 -2519
rect 1717 -2553 2045 -2519
<< metal1 >>
rect -2057 2553 -1705 2559
rect -2057 2519 -2045 2553
rect -1717 2519 -1705 2553
rect -2057 2513 -1705 2519
rect -1639 2553 -1287 2559
rect -1639 2519 -1627 2553
rect -1299 2519 -1287 2553
rect -1639 2513 -1287 2519
rect -1221 2553 -869 2559
rect -1221 2519 -1209 2553
rect -881 2519 -869 2553
rect -1221 2513 -869 2519
rect -803 2553 -451 2559
rect -803 2519 -791 2553
rect -463 2519 -451 2553
rect -803 2513 -451 2519
rect -385 2553 -33 2559
rect -385 2519 -373 2553
rect -45 2519 -33 2553
rect -385 2513 -33 2519
rect 33 2553 385 2559
rect 33 2519 45 2553
rect 373 2519 385 2553
rect 33 2513 385 2519
rect 451 2553 803 2559
rect 451 2519 463 2553
rect 791 2519 803 2553
rect 451 2513 803 2519
rect 869 2553 1221 2559
rect 869 2519 881 2553
rect 1209 2519 1221 2553
rect 869 2513 1221 2519
rect 1287 2553 1639 2559
rect 1287 2519 1299 2553
rect 1627 2519 1639 2553
rect 1287 2513 1639 2519
rect 1705 2553 2057 2559
rect 1705 2519 1717 2553
rect 2045 2519 2057 2553
rect 1705 2513 2057 2519
rect -2113 2469 -2067 2481
rect -2113 2193 -2107 2469
rect -2073 2193 -2067 2469
rect -2113 2181 -2067 2193
rect -1695 2469 -1649 2481
rect -1695 2193 -1689 2469
rect -1655 2193 -1649 2469
rect -1695 2181 -1649 2193
rect -1277 2469 -1231 2481
rect -1277 2193 -1271 2469
rect -1237 2193 -1231 2469
rect -1277 2181 -1231 2193
rect -859 2469 -813 2481
rect -859 2193 -853 2469
rect -819 2193 -813 2469
rect -859 2181 -813 2193
rect -441 2469 -395 2481
rect -441 2193 -435 2469
rect -401 2193 -395 2469
rect -441 2181 -395 2193
rect -23 2469 23 2481
rect -23 2193 -17 2469
rect 17 2193 23 2469
rect -23 2181 23 2193
rect 395 2469 441 2481
rect 395 2193 401 2469
rect 435 2193 441 2469
rect 395 2181 441 2193
rect 813 2469 859 2481
rect 813 2193 819 2469
rect 853 2193 859 2469
rect 813 2181 859 2193
rect 1231 2469 1277 2481
rect 1231 2193 1237 2469
rect 1271 2193 1277 2469
rect 1231 2181 1277 2193
rect 1649 2469 1695 2481
rect 1649 2193 1655 2469
rect 1689 2193 1695 2469
rect 1649 2181 1695 2193
rect 2067 2469 2113 2481
rect 2067 2193 2073 2469
rect 2107 2193 2113 2469
rect 2067 2181 2113 2193
rect -2057 2143 -1705 2149
rect -2057 2109 -2045 2143
rect -1717 2109 -1705 2143
rect -2057 2103 -1705 2109
rect -1639 2143 -1287 2149
rect -1639 2109 -1627 2143
rect -1299 2109 -1287 2143
rect -1639 2103 -1287 2109
rect -1221 2143 -869 2149
rect -1221 2109 -1209 2143
rect -881 2109 -869 2143
rect -1221 2103 -869 2109
rect -803 2143 -451 2149
rect -803 2109 -791 2143
rect -463 2109 -451 2143
rect -803 2103 -451 2109
rect -385 2143 -33 2149
rect -385 2109 -373 2143
rect -45 2109 -33 2143
rect -385 2103 -33 2109
rect 33 2143 385 2149
rect 33 2109 45 2143
rect 373 2109 385 2143
rect 33 2103 385 2109
rect 451 2143 803 2149
rect 451 2109 463 2143
rect 791 2109 803 2143
rect 451 2103 803 2109
rect 869 2143 1221 2149
rect 869 2109 881 2143
rect 1209 2109 1221 2143
rect 869 2103 1221 2109
rect 1287 2143 1639 2149
rect 1287 2109 1299 2143
rect 1627 2109 1639 2143
rect 1287 2103 1639 2109
rect 1705 2143 2057 2149
rect 1705 2109 1717 2143
rect 2045 2109 2057 2143
rect 1705 2103 2057 2109
rect -2057 2035 -1705 2041
rect -2057 2001 -2045 2035
rect -1717 2001 -1705 2035
rect -2057 1995 -1705 2001
rect -1639 2035 -1287 2041
rect -1639 2001 -1627 2035
rect -1299 2001 -1287 2035
rect -1639 1995 -1287 2001
rect -1221 2035 -869 2041
rect -1221 2001 -1209 2035
rect -881 2001 -869 2035
rect -1221 1995 -869 2001
rect -803 2035 -451 2041
rect -803 2001 -791 2035
rect -463 2001 -451 2035
rect -803 1995 -451 2001
rect -385 2035 -33 2041
rect -385 2001 -373 2035
rect -45 2001 -33 2035
rect -385 1995 -33 2001
rect 33 2035 385 2041
rect 33 2001 45 2035
rect 373 2001 385 2035
rect 33 1995 385 2001
rect 451 2035 803 2041
rect 451 2001 463 2035
rect 791 2001 803 2035
rect 451 1995 803 2001
rect 869 2035 1221 2041
rect 869 2001 881 2035
rect 1209 2001 1221 2035
rect 869 1995 1221 2001
rect 1287 2035 1639 2041
rect 1287 2001 1299 2035
rect 1627 2001 1639 2035
rect 1287 1995 1639 2001
rect 1705 2035 2057 2041
rect 1705 2001 1717 2035
rect 2045 2001 2057 2035
rect 1705 1995 2057 2001
rect -2113 1951 -2067 1963
rect -2113 1675 -2107 1951
rect -2073 1675 -2067 1951
rect -2113 1663 -2067 1675
rect -1695 1951 -1649 1963
rect -1695 1675 -1689 1951
rect -1655 1675 -1649 1951
rect -1695 1663 -1649 1675
rect -1277 1951 -1231 1963
rect -1277 1675 -1271 1951
rect -1237 1675 -1231 1951
rect -1277 1663 -1231 1675
rect -859 1951 -813 1963
rect -859 1675 -853 1951
rect -819 1675 -813 1951
rect -859 1663 -813 1675
rect -441 1951 -395 1963
rect -441 1675 -435 1951
rect -401 1675 -395 1951
rect -441 1663 -395 1675
rect -23 1951 23 1963
rect -23 1675 -17 1951
rect 17 1675 23 1951
rect -23 1663 23 1675
rect 395 1951 441 1963
rect 395 1675 401 1951
rect 435 1675 441 1951
rect 395 1663 441 1675
rect 813 1951 859 1963
rect 813 1675 819 1951
rect 853 1675 859 1951
rect 813 1663 859 1675
rect 1231 1951 1277 1963
rect 1231 1675 1237 1951
rect 1271 1675 1277 1951
rect 1231 1663 1277 1675
rect 1649 1951 1695 1963
rect 1649 1675 1655 1951
rect 1689 1675 1695 1951
rect 1649 1663 1695 1675
rect 2067 1951 2113 1963
rect 2067 1675 2073 1951
rect 2107 1675 2113 1951
rect 2067 1663 2113 1675
rect -2057 1625 -1705 1631
rect -2057 1591 -2045 1625
rect -1717 1591 -1705 1625
rect -2057 1585 -1705 1591
rect -1639 1625 -1287 1631
rect -1639 1591 -1627 1625
rect -1299 1591 -1287 1625
rect -1639 1585 -1287 1591
rect -1221 1625 -869 1631
rect -1221 1591 -1209 1625
rect -881 1591 -869 1625
rect -1221 1585 -869 1591
rect -803 1625 -451 1631
rect -803 1591 -791 1625
rect -463 1591 -451 1625
rect -803 1585 -451 1591
rect -385 1625 -33 1631
rect -385 1591 -373 1625
rect -45 1591 -33 1625
rect -385 1585 -33 1591
rect 33 1625 385 1631
rect 33 1591 45 1625
rect 373 1591 385 1625
rect 33 1585 385 1591
rect 451 1625 803 1631
rect 451 1591 463 1625
rect 791 1591 803 1625
rect 451 1585 803 1591
rect 869 1625 1221 1631
rect 869 1591 881 1625
rect 1209 1591 1221 1625
rect 869 1585 1221 1591
rect 1287 1625 1639 1631
rect 1287 1591 1299 1625
rect 1627 1591 1639 1625
rect 1287 1585 1639 1591
rect 1705 1625 2057 1631
rect 1705 1591 1717 1625
rect 2045 1591 2057 1625
rect 1705 1585 2057 1591
rect -2057 1517 -1705 1523
rect -2057 1483 -2045 1517
rect -1717 1483 -1705 1517
rect -2057 1477 -1705 1483
rect -1639 1517 -1287 1523
rect -1639 1483 -1627 1517
rect -1299 1483 -1287 1517
rect -1639 1477 -1287 1483
rect -1221 1517 -869 1523
rect -1221 1483 -1209 1517
rect -881 1483 -869 1517
rect -1221 1477 -869 1483
rect -803 1517 -451 1523
rect -803 1483 -791 1517
rect -463 1483 -451 1517
rect -803 1477 -451 1483
rect -385 1517 -33 1523
rect -385 1483 -373 1517
rect -45 1483 -33 1517
rect -385 1477 -33 1483
rect 33 1517 385 1523
rect 33 1483 45 1517
rect 373 1483 385 1517
rect 33 1477 385 1483
rect 451 1517 803 1523
rect 451 1483 463 1517
rect 791 1483 803 1517
rect 451 1477 803 1483
rect 869 1517 1221 1523
rect 869 1483 881 1517
rect 1209 1483 1221 1517
rect 869 1477 1221 1483
rect 1287 1517 1639 1523
rect 1287 1483 1299 1517
rect 1627 1483 1639 1517
rect 1287 1477 1639 1483
rect 1705 1517 2057 1523
rect 1705 1483 1717 1517
rect 2045 1483 2057 1517
rect 1705 1477 2057 1483
rect -2113 1433 -2067 1445
rect -2113 1157 -2107 1433
rect -2073 1157 -2067 1433
rect -2113 1145 -2067 1157
rect -1695 1433 -1649 1445
rect -1695 1157 -1689 1433
rect -1655 1157 -1649 1433
rect -1695 1145 -1649 1157
rect -1277 1433 -1231 1445
rect -1277 1157 -1271 1433
rect -1237 1157 -1231 1433
rect -1277 1145 -1231 1157
rect -859 1433 -813 1445
rect -859 1157 -853 1433
rect -819 1157 -813 1433
rect -859 1145 -813 1157
rect -441 1433 -395 1445
rect -441 1157 -435 1433
rect -401 1157 -395 1433
rect -441 1145 -395 1157
rect -23 1433 23 1445
rect -23 1157 -17 1433
rect 17 1157 23 1433
rect -23 1145 23 1157
rect 395 1433 441 1445
rect 395 1157 401 1433
rect 435 1157 441 1433
rect 395 1145 441 1157
rect 813 1433 859 1445
rect 813 1157 819 1433
rect 853 1157 859 1433
rect 813 1145 859 1157
rect 1231 1433 1277 1445
rect 1231 1157 1237 1433
rect 1271 1157 1277 1433
rect 1231 1145 1277 1157
rect 1649 1433 1695 1445
rect 1649 1157 1655 1433
rect 1689 1157 1695 1433
rect 1649 1145 1695 1157
rect 2067 1433 2113 1445
rect 2067 1157 2073 1433
rect 2107 1157 2113 1433
rect 2067 1145 2113 1157
rect -2057 1107 -1705 1113
rect -2057 1073 -2045 1107
rect -1717 1073 -1705 1107
rect -2057 1067 -1705 1073
rect -1639 1107 -1287 1113
rect -1639 1073 -1627 1107
rect -1299 1073 -1287 1107
rect -1639 1067 -1287 1073
rect -1221 1107 -869 1113
rect -1221 1073 -1209 1107
rect -881 1073 -869 1107
rect -1221 1067 -869 1073
rect -803 1107 -451 1113
rect -803 1073 -791 1107
rect -463 1073 -451 1107
rect -803 1067 -451 1073
rect -385 1107 -33 1113
rect -385 1073 -373 1107
rect -45 1073 -33 1107
rect -385 1067 -33 1073
rect 33 1107 385 1113
rect 33 1073 45 1107
rect 373 1073 385 1107
rect 33 1067 385 1073
rect 451 1107 803 1113
rect 451 1073 463 1107
rect 791 1073 803 1107
rect 451 1067 803 1073
rect 869 1107 1221 1113
rect 869 1073 881 1107
rect 1209 1073 1221 1107
rect 869 1067 1221 1073
rect 1287 1107 1639 1113
rect 1287 1073 1299 1107
rect 1627 1073 1639 1107
rect 1287 1067 1639 1073
rect 1705 1107 2057 1113
rect 1705 1073 1717 1107
rect 2045 1073 2057 1107
rect 1705 1067 2057 1073
rect -2057 999 -1705 1005
rect -2057 965 -2045 999
rect -1717 965 -1705 999
rect -2057 959 -1705 965
rect -1639 999 -1287 1005
rect -1639 965 -1627 999
rect -1299 965 -1287 999
rect -1639 959 -1287 965
rect -1221 999 -869 1005
rect -1221 965 -1209 999
rect -881 965 -869 999
rect -1221 959 -869 965
rect -803 999 -451 1005
rect -803 965 -791 999
rect -463 965 -451 999
rect -803 959 -451 965
rect -385 999 -33 1005
rect -385 965 -373 999
rect -45 965 -33 999
rect -385 959 -33 965
rect 33 999 385 1005
rect 33 965 45 999
rect 373 965 385 999
rect 33 959 385 965
rect 451 999 803 1005
rect 451 965 463 999
rect 791 965 803 999
rect 451 959 803 965
rect 869 999 1221 1005
rect 869 965 881 999
rect 1209 965 1221 999
rect 869 959 1221 965
rect 1287 999 1639 1005
rect 1287 965 1299 999
rect 1627 965 1639 999
rect 1287 959 1639 965
rect 1705 999 2057 1005
rect 1705 965 1717 999
rect 2045 965 2057 999
rect 1705 959 2057 965
rect -2113 915 -2067 927
rect -2113 639 -2107 915
rect -2073 639 -2067 915
rect -2113 627 -2067 639
rect -1695 915 -1649 927
rect -1695 639 -1689 915
rect -1655 639 -1649 915
rect -1695 627 -1649 639
rect -1277 915 -1231 927
rect -1277 639 -1271 915
rect -1237 639 -1231 915
rect -1277 627 -1231 639
rect -859 915 -813 927
rect -859 639 -853 915
rect -819 639 -813 915
rect -859 627 -813 639
rect -441 915 -395 927
rect -441 639 -435 915
rect -401 639 -395 915
rect -441 627 -395 639
rect -23 915 23 927
rect -23 639 -17 915
rect 17 639 23 915
rect -23 627 23 639
rect 395 915 441 927
rect 395 639 401 915
rect 435 639 441 915
rect 395 627 441 639
rect 813 915 859 927
rect 813 639 819 915
rect 853 639 859 915
rect 813 627 859 639
rect 1231 915 1277 927
rect 1231 639 1237 915
rect 1271 639 1277 915
rect 1231 627 1277 639
rect 1649 915 1695 927
rect 1649 639 1655 915
rect 1689 639 1695 915
rect 1649 627 1695 639
rect 2067 915 2113 927
rect 2067 639 2073 915
rect 2107 639 2113 915
rect 2067 627 2113 639
rect -2057 589 -1705 595
rect -2057 555 -2045 589
rect -1717 555 -1705 589
rect -2057 549 -1705 555
rect -1639 589 -1287 595
rect -1639 555 -1627 589
rect -1299 555 -1287 589
rect -1639 549 -1287 555
rect -1221 589 -869 595
rect -1221 555 -1209 589
rect -881 555 -869 589
rect -1221 549 -869 555
rect -803 589 -451 595
rect -803 555 -791 589
rect -463 555 -451 589
rect -803 549 -451 555
rect -385 589 -33 595
rect -385 555 -373 589
rect -45 555 -33 589
rect -385 549 -33 555
rect 33 589 385 595
rect 33 555 45 589
rect 373 555 385 589
rect 33 549 385 555
rect 451 589 803 595
rect 451 555 463 589
rect 791 555 803 589
rect 451 549 803 555
rect 869 589 1221 595
rect 869 555 881 589
rect 1209 555 1221 589
rect 869 549 1221 555
rect 1287 589 1639 595
rect 1287 555 1299 589
rect 1627 555 1639 589
rect 1287 549 1639 555
rect 1705 589 2057 595
rect 1705 555 1717 589
rect 2045 555 2057 589
rect 1705 549 2057 555
rect -2057 481 -1705 487
rect -2057 447 -2045 481
rect -1717 447 -1705 481
rect -2057 441 -1705 447
rect -1639 481 -1287 487
rect -1639 447 -1627 481
rect -1299 447 -1287 481
rect -1639 441 -1287 447
rect -1221 481 -869 487
rect -1221 447 -1209 481
rect -881 447 -869 481
rect -1221 441 -869 447
rect -803 481 -451 487
rect -803 447 -791 481
rect -463 447 -451 481
rect -803 441 -451 447
rect -385 481 -33 487
rect -385 447 -373 481
rect -45 447 -33 481
rect -385 441 -33 447
rect 33 481 385 487
rect 33 447 45 481
rect 373 447 385 481
rect 33 441 385 447
rect 451 481 803 487
rect 451 447 463 481
rect 791 447 803 481
rect 451 441 803 447
rect 869 481 1221 487
rect 869 447 881 481
rect 1209 447 1221 481
rect 869 441 1221 447
rect 1287 481 1639 487
rect 1287 447 1299 481
rect 1627 447 1639 481
rect 1287 441 1639 447
rect 1705 481 2057 487
rect 1705 447 1717 481
rect 2045 447 2057 481
rect 1705 441 2057 447
rect -2113 397 -2067 409
rect -2113 121 -2107 397
rect -2073 121 -2067 397
rect -2113 109 -2067 121
rect -1695 397 -1649 409
rect -1695 121 -1689 397
rect -1655 121 -1649 397
rect -1695 109 -1649 121
rect -1277 397 -1231 409
rect -1277 121 -1271 397
rect -1237 121 -1231 397
rect -1277 109 -1231 121
rect -859 397 -813 409
rect -859 121 -853 397
rect -819 121 -813 397
rect -859 109 -813 121
rect -441 397 -395 409
rect -441 121 -435 397
rect -401 121 -395 397
rect -441 109 -395 121
rect -23 397 23 409
rect -23 121 -17 397
rect 17 121 23 397
rect -23 109 23 121
rect 395 397 441 409
rect 395 121 401 397
rect 435 121 441 397
rect 395 109 441 121
rect 813 397 859 409
rect 813 121 819 397
rect 853 121 859 397
rect 813 109 859 121
rect 1231 397 1277 409
rect 1231 121 1237 397
rect 1271 121 1277 397
rect 1231 109 1277 121
rect 1649 397 1695 409
rect 1649 121 1655 397
rect 1689 121 1695 397
rect 1649 109 1695 121
rect 2067 397 2113 409
rect 2067 121 2073 397
rect 2107 121 2113 397
rect 2067 109 2113 121
rect -2057 71 -1705 77
rect -2057 37 -2045 71
rect -1717 37 -1705 71
rect -2057 31 -1705 37
rect -1639 71 -1287 77
rect -1639 37 -1627 71
rect -1299 37 -1287 71
rect -1639 31 -1287 37
rect -1221 71 -869 77
rect -1221 37 -1209 71
rect -881 37 -869 71
rect -1221 31 -869 37
rect -803 71 -451 77
rect -803 37 -791 71
rect -463 37 -451 71
rect -803 31 -451 37
rect -385 71 -33 77
rect -385 37 -373 71
rect -45 37 -33 71
rect -385 31 -33 37
rect 33 71 385 77
rect 33 37 45 71
rect 373 37 385 71
rect 33 31 385 37
rect 451 71 803 77
rect 451 37 463 71
rect 791 37 803 71
rect 451 31 803 37
rect 869 71 1221 77
rect 869 37 881 71
rect 1209 37 1221 71
rect 869 31 1221 37
rect 1287 71 1639 77
rect 1287 37 1299 71
rect 1627 37 1639 71
rect 1287 31 1639 37
rect 1705 71 2057 77
rect 1705 37 1717 71
rect 2045 37 2057 71
rect 1705 31 2057 37
rect -2057 -37 -1705 -31
rect -2057 -71 -2045 -37
rect -1717 -71 -1705 -37
rect -2057 -77 -1705 -71
rect -1639 -37 -1287 -31
rect -1639 -71 -1627 -37
rect -1299 -71 -1287 -37
rect -1639 -77 -1287 -71
rect -1221 -37 -869 -31
rect -1221 -71 -1209 -37
rect -881 -71 -869 -37
rect -1221 -77 -869 -71
rect -803 -37 -451 -31
rect -803 -71 -791 -37
rect -463 -71 -451 -37
rect -803 -77 -451 -71
rect -385 -37 -33 -31
rect -385 -71 -373 -37
rect -45 -71 -33 -37
rect -385 -77 -33 -71
rect 33 -37 385 -31
rect 33 -71 45 -37
rect 373 -71 385 -37
rect 33 -77 385 -71
rect 451 -37 803 -31
rect 451 -71 463 -37
rect 791 -71 803 -37
rect 451 -77 803 -71
rect 869 -37 1221 -31
rect 869 -71 881 -37
rect 1209 -71 1221 -37
rect 869 -77 1221 -71
rect 1287 -37 1639 -31
rect 1287 -71 1299 -37
rect 1627 -71 1639 -37
rect 1287 -77 1639 -71
rect 1705 -37 2057 -31
rect 1705 -71 1717 -37
rect 2045 -71 2057 -37
rect 1705 -77 2057 -71
rect -2113 -121 -2067 -109
rect -2113 -397 -2107 -121
rect -2073 -397 -2067 -121
rect -2113 -409 -2067 -397
rect -1695 -121 -1649 -109
rect -1695 -397 -1689 -121
rect -1655 -397 -1649 -121
rect -1695 -409 -1649 -397
rect -1277 -121 -1231 -109
rect -1277 -397 -1271 -121
rect -1237 -397 -1231 -121
rect -1277 -409 -1231 -397
rect -859 -121 -813 -109
rect -859 -397 -853 -121
rect -819 -397 -813 -121
rect -859 -409 -813 -397
rect -441 -121 -395 -109
rect -441 -397 -435 -121
rect -401 -397 -395 -121
rect -441 -409 -395 -397
rect -23 -121 23 -109
rect -23 -397 -17 -121
rect 17 -397 23 -121
rect -23 -409 23 -397
rect 395 -121 441 -109
rect 395 -397 401 -121
rect 435 -397 441 -121
rect 395 -409 441 -397
rect 813 -121 859 -109
rect 813 -397 819 -121
rect 853 -397 859 -121
rect 813 -409 859 -397
rect 1231 -121 1277 -109
rect 1231 -397 1237 -121
rect 1271 -397 1277 -121
rect 1231 -409 1277 -397
rect 1649 -121 1695 -109
rect 1649 -397 1655 -121
rect 1689 -397 1695 -121
rect 1649 -409 1695 -397
rect 2067 -121 2113 -109
rect 2067 -397 2073 -121
rect 2107 -397 2113 -121
rect 2067 -409 2113 -397
rect -2057 -447 -1705 -441
rect -2057 -481 -2045 -447
rect -1717 -481 -1705 -447
rect -2057 -487 -1705 -481
rect -1639 -447 -1287 -441
rect -1639 -481 -1627 -447
rect -1299 -481 -1287 -447
rect -1639 -487 -1287 -481
rect -1221 -447 -869 -441
rect -1221 -481 -1209 -447
rect -881 -481 -869 -447
rect -1221 -487 -869 -481
rect -803 -447 -451 -441
rect -803 -481 -791 -447
rect -463 -481 -451 -447
rect -803 -487 -451 -481
rect -385 -447 -33 -441
rect -385 -481 -373 -447
rect -45 -481 -33 -447
rect -385 -487 -33 -481
rect 33 -447 385 -441
rect 33 -481 45 -447
rect 373 -481 385 -447
rect 33 -487 385 -481
rect 451 -447 803 -441
rect 451 -481 463 -447
rect 791 -481 803 -447
rect 451 -487 803 -481
rect 869 -447 1221 -441
rect 869 -481 881 -447
rect 1209 -481 1221 -447
rect 869 -487 1221 -481
rect 1287 -447 1639 -441
rect 1287 -481 1299 -447
rect 1627 -481 1639 -447
rect 1287 -487 1639 -481
rect 1705 -447 2057 -441
rect 1705 -481 1717 -447
rect 2045 -481 2057 -447
rect 1705 -487 2057 -481
rect -2057 -555 -1705 -549
rect -2057 -589 -2045 -555
rect -1717 -589 -1705 -555
rect -2057 -595 -1705 -589
rect -1639 -555 -1287 -549
rect -1639 -589 -1627 -555
rect -1299 -589 -1287 -555
rect -1639 -595 -1287 -589
rect -1221 -555 -869 -549
rect -1221 -589 -1209 -555
rect -881 -589 -869 -555
rect -1221 -595 -869 -589
rect -803 -555 -451 -549
rect -803 -589 -791 -555
rect -463 -589 -451 -555
rect -803 -595 -451 -589
rect -385 -555 -33 -549
rect -385 -589 -373 -555
rect -45 -589 -33 -555
rect -385 -595 -33 -589
rect 33 -555 385 -549
rect 33 -589 45 -555
rect 373 -589 385 -555
rect 33 -595 385 -589
rect 451 -555 803 -549
rect 451 -589 463 -555
rect 791 -589 803 -555
rect 451 -595 803 -589
rect 869 -555 1221 -549
rect 869 -589 881 -555
rect 1209 -589 1221 -555
rect 869 -595 1221 -589
rect 1287 -555 1639 -549
rect 1287 -589 1299 -555
rect 1627 -589 1639 -555
rect 1287 -595 1639 -589
rect 1705 -555 2057 -549
rect 1705 -589 1717 -555
rect 2045 -589 2057 -555
rect 1705 -595 2057 -589
rect -2113 -639 -2067 -627
rect -2113 -915 -2107 -639
rect -2073 -915 -2067 -639
rect -2113 -927 -2067 -915
rect -1695 -639 -1649 -627
rect -1695 -915 -1689 -639
rect -1655 -915 -1649 -639
rect -1695 -927 -1649 -915
rect -1277 -639 -1231 -627
rect -1277 -915 -1271 -639
rect -1237 -915 -1231 -639
rect -1277 -927 -1231 -915
rect -859 -639 -813 -627
rect -859 -915 -853 -639
rect -819 -915 -813 -639
rect -859 -927 -813 -915
rect -441 -639 -395 -627
rect -441 -915 -435 -639
rect -401 -915 -395 -639
rect -441 -927 -395 -915
rect -23 -639 23 -627
rect -23 -915 -17 -639
rect 17 -915 23 -639
rect -23 -927 23 -915
rect 395 -639 441 -627
rect 395 -915 401 -639
rect 435 -915 441 -639
rect 395 -927 441 -915
rect 813 -639 859 -627
rect 813 -915 819 -639
rect 853 -915 859 -639
rect 813 -927 859 -915
rect 1231 -639 1277 -627
rect 1231 -915 1237 -639
rect 1271 -915 1277 -639
rect 1231 -927 1277 -915
rect 1649 -639 1695 -627
rect 1649 -915 1655 -639
rect 1689 -915 1695 -639
rect 1649 -927 1695 -915
rect 2067 -639 2113 -627
rect 2067 -915 2073 -639
rect 2107 -915 2113 -639
rect 2067 -927 2113 -915
rect -2057 -965 -1705 -959
rect -2057 -999 -2045 -965
rect -1717 -999 -1705 -965
rect -2057 -1005 -1705 -999
rect -1639 -965 -1287 -959
rect -1639 -999 -1627 -965
rect -1299 -999 -1287 -965
rect -1639 -1005 -1287 -999
rect -1221 -965 -869 -959
rect -1221 -999 -1209 -965
rect -881 -999 -869 -965
rect -1221 -1005 -869 -999
rect -803 -965 -451 -959
rect -803 -999 -791 -965
rect -463 -999 -451 -965
rect -803 -1005 -451 -999
rect -385 -965 -33 -959
rect -385 -999 -373 -965
rect -45 -999 -33 -965
rect -385 -1005 -33 -999
rect 33 -965 385 -959
rect 33 -999 45 -965
rect 373 -999 385 -965
rect 33 -1005 385 -999
rect 451 -965 803 -959
rect 451 -999 463 -965
rect 791 -999 803 -965
rect 451 -1005 803 -999
rect 869 -965 1221 -959
rect 869 -999 881 -965
rect 1209 -999 1221 -965
rect 869 -1005 1221 -999
rect 1287 -965 1639 -959
rect 1287 -999 1299 -965
rect 1627 -999 1639 -965
rect 1287 -1005 1639 -999
rect 1705 -965 2057 -959
rect 1705 -999 1717 -965
rect 2045 -999 2057 -965
rect 1705 -1005 2057 -999
rect -2057 -1073 -1705 -1067
rect -2057 -1107 -2045 -1073
rect -1717 -1107 -1705 -1073
rect -2057 -1113 -1705 -1107
rect -1639 -1073 -1287 -1067
rect -1639 -1107 -1627 -1073
rect -1299 -1107 -1287 -1073
rect -1639 -1113 -1287 -1107
rect -1221 -1073 -869 -1067
rect -1221 -1107 -1209 -1073
rect -881 -1107 -869 -1073
rect -1221 -1113 -869 -1107
rect -803 -1073 -451 -1067
rect -803 -1107 -791 -1073
rect -463 -1107 -451 -1073
rect -803 -1113 -451 -1107
rect -385 -1073 -33 -1067
rect -385 -1107 -373 -1073
rect -45 -1107 -33 -1073
rect -385 -1113 -33 -1107
rect 33 -1073 385 -1067
rect 33 -1107 45 -1073
rect 373 -1107 385 -1073
rect 33 -1113 385 -1107
rect 451 -1073 803 -1067
rect 451 -1107 463 -1073
rect 791 -1107 803 -1073
rect 451 -1113 803 -1107
rect 869 -1073 1221 -1067
rect 869 -1107 881 -1073
rect 1209 -1107 1221 -1073
rect 869 -1113 1221 -1107
rect 1287 -1073 1639 -1067
rect 1287 -1107 1299 -1073
rect 1627 -1107 1639 -1073
rect 1287 -1113 1639 -1107
rect 1705 -1073 2057 -1067
rect 1705 -1107 1717 -1073
rect 2045 -1107 2057 -1073
rect 1705 -1113 2057 -1107
rect -2113 -1157 -2067 -1145
rect -2113 -1433 -2107 -1157
rect -2073 -1433 -2067 -1157
rect -2113 -1445 -2067 -1433
rect -1695 -1157 -1649 -1145
rect -1695 -1433 -1689 -1157
rect -1655 -1433 -1649 -1157
rect -1695 -1445 -1649 -1433
rect -1277 -1157 -1231 -1145
rect -1277 -1433 -1271 -1157
rect -1237 -1433 -1231 -1157
rect -1277 -1445 -1231 -1433
rect -859 -1157 -813 -1145
rect -859 -1433 -853 -1157
rect -819 -1433 -813 -1157
rect -859 -1445 -813 -1433
rect -441 -1157 -395 -1145
rect -441 -1433 -435 -1157
rect -401 -1433 -395 -1157
rect -441 -1445 -395 -1433
rect -23 -1157 23 -1145
rect -23 -1433 -17 -1157
rect 17 -1433 23 -1157
rect -23 -1445 23 -1433
rect 395 -1157 441 -1145
rect 395 -1433 401 -1157
rect 435 -1433 441 -1157
rect 395 -1445 441 -1433
rect 813 -1157 859 -1145
rect 813 -1433 819 -1157
rect 853 -1433 859 -1157
rect 813 -1445 859 -1433
rect 1231 -1157 1277 -1145
rect 1231 -1433 1237 -1157
rect 1271 -1433 1277 -1157
rect 1231 -1445 1277 -1433
rect 1649 -1157 1695 -1145
rect 1649 -1433 1655 -1157
rect 1689 -1433 1695 -1157
rect 1649 -1445 1695 -1433
rect 2067 -1157 2113 -1145
rect 2067 -1433 2073 -1157
rect 2107 -1433 2113 -1157
rect 2067 -1445 2113 -1433
rect -2057 -1483 -1705 -1477
rect -2057 -1517 -2045 -1483
rect -1717 -1517 -1705 -1483
rect -2057 -1523 -1705 -1517
rect -1639 -1483 -1287 -1477
rect -1639 -1517 -1627 -1483
rect -1299 -1517 -1287 -1483
rect -1639 -1523 -1287 -1517
rect -1221 -1483 -869 -1477
rect -1221 -1517 -1209 -1483
rect -881 -1517 -869 -1483
rect -1221 -1523 -869 -1517
rect -803 -1483 -451 -1477
rect -803 -1517 -791 -1483
rect -463 -1517 -451 -1483
rect -803 -1523 -451 -1517
rect -385 -1483 -33 -1477
rect -385 -1517 -373 -1483
rect -45 -1517 -33 -1483
rect -385 -1523 -33 -1517
rect 33 -1483 385 -1477
rect 33 -1517 45 -1483
rect 373 -1517 385 -1483
rect 33 -1523 385 -1517
rect 451 -1483 803 -1477
rect 451 -1517 463 -1483
rect 791 -1517 803 -1483
rect 451 -1523 803 -1517
rect 869 -1483 1221 -1477
rect 869 -1517 881 -1483
rect 1209 -1517 1221 -1483
rect 869 -1523 1221 -1517
rect 1287 -1483 1639 -1477
rect 1287 -1517 1299 -1483
rect 1627 -1517 1639 -1483
rect 1287 -1523 1639 -1517
rect 1705 -1483 2057 -1477
rect 1705 -1517 1717 -1483
rect 2045 -1517 2057 -1483
rect 1705 -1523 2057 -1517
rect -2057 -1591 -1705 -1585
rect -2057 -1625 -2045 -1591
rect -1717 -1625 -1705 -1591
rect -2057 -1631 -1705 -1625
rect -1639 -1591 -1287 -1585
rect -1639 -1625 -1627 -1591
rect -1299 -1625 -1287 -1591
rect -1639 -1631 -1287 -1625
rect -1221 -1591 -869 -1585
rect -1221 -1625 -1209 -1591
rect -881 -1625 -869 -1591
rect -1221 -1631 -869 -1625
rect -803 -1591 -451 -1585
rect -803 -1625 -791 -1591
rect -463 -1625 -451 -1591
rect -803 -1631 -451 -1625
rect -385 -1591 -33 -1585
rect -385 -1625 -373 -1591
rect -45 -1625 -33 -1591
rect -385 -1631 -33 -1625
rect 33 -1591 385 -1585
rect 33 -1625 45 -1591
rect 373 -1625 385 -1591
rect 33 -1631 385 -1625
rect 451 -1591 803 -1585
rect 451 -1625 463 -1591
rect 791 -1625 803 -1591
rect 451 -1631 803 -1625
rect 869 -1591 1221 -1585
rect 869 -1625 881 -1591
rect 1209 -1625 1221 -1591
rect 869 -1631 1221 -1625
rect 1287 -1591 1639 -1585
rect 1287 -1625 1299 -1591
rect 1627 -1625 1639 -1591
rect 1287 -1631 1639 -1625
rect 1705 -1591 2057 -1585
rect 1705 -1625 1717 -1591
rect 2045 -1625 2057 -1591
rect 1705 -1631 2057 -1625
rect -2113 -1675 -2067 -1663
rect -2113 -1951 -2107 -1675
rect -2073 -1951 -2067 -1675
rect -2113 -1963 -2067 -1951
rect -1695 -1675 -1649 -1663
rect -1695 -1951 -1689 -1675
rect -1655 -1951 -1649 -1675
rect -1695 -1963 -1649 -1951
rect -1277 -1675 -1231 -1663
rect -1277 -1951 -1271 -1675
rect -1237 -1951 -1231 -1675
rect -1277 -1963 -1231 -1951
rect -859 -1675 -813 -1663
rect -859 -1951 -853 -1675
rect -819 -1951 -813 -1675
rect -859 -1963 -813 -1951
rect -441 -1675 -395 -1663
rect -441 -1951 -435 -1675
rect -401 -1951 -395 -1675
rect -441 -1963 -395 -1951
rect -23 -1675 23 -1663
rect -23 -1951 -17 -1675
rect 17 -1951 23 -1675
rect -23 -1963 23 -1951
rect 395 -1675 441 -1663
rect 395 -1951 401 -1675
rect 435 -1951 441 -1675
rect 395 -1963 441 -1951
rect 813 -1675 859 -1663
rect 813 -1951 819 -1675
rect 853 -1951 859 -1675
rect 813 -1963 859 -1951
rect 1231 -1675 1277 -1663
rect 1231 -1951 1237 -1675
rect 1271 -1951 1277 -1675
rect 1231 -1963 1277 -1951
rect 1649 -1675 1695 -1663
rect 1649 -1951 1655 -1675
rect 1689 -1951 1695 -1675
rect 1649 -1963 1695 -1951
rect 2067 -1675 2113 -1663
rect 2067 -1951 2073 -1675
rect 2107 -1951 2113 -1675
rect 2067 -1963 2113 -1951
rect -2057 -2001 -1705 -1995
rect -2057 -2035 -2045 -2001
rect -1717 -2035 -1705 -2001
rect -2057 -2041 -1705 -2035
rect -1639 -2001 -1287 -1995
rect -1639 -2035 -1627 -2001
rect -1299 -2035 -1287 -2001
rect -1639 -2041 -1287 -2035
rect -1221 -2001 -869 -1995
rect -1221 -2035 -1209 -2001
rect -881 -2035 -869 -2001
rect -1221 -2041 -869 -2035
rect -803 -2001 -451 -1995
rect -803 -2035 -791 -2001
rect -463 -2035 -451 -2001
rect -803 -2041 -451 -2035
rect -385 -2001 -33 -1995
rect -385 -2035 -373 -2001
rect -45 -2035 -33 -2001
rect -385 -2041 -33 -2035
rect 33 -2001 385 -1995
rect 33 -2035 45 -2001
rect 373 -2035 385 -2001
rect 33 -2041 385 -2035
rect 451 -2001 803 -1995
rect 451 -2035 463 -2001
rect 791 -2035 803 -2001
rect 451 -2041 803 -2035
rect 869 -2001 1221 -1995
rect 869 -2035 881 -2001
rect 1209 -2035 1221 -2001
rect 869 -2041 1221 -2035
rect 1287 -2001 1639 -1995
rect 1287 -2035 1299 -2001
rect 1627 -2035 1639 -2001
rect 1287 -2041 1639 -2035
rect 1705 -2001 2057 -1995
rect 1705 -2035 1717 -2001
rect 2045 -2035 2057 -2001
rect 1705 -2041 2057 -2035
rect -2057 -2109 -1705 -2103
rect -2057 -2143 -2045 -2109
rect -1717 -2143 -1705 -2109
rect -2057 -2149 -1705 -2143
rect -1639 -2109 -1287 -2103
rect -1639 -2143 -1627 -2109
rect -1299 -2143 -1287 -2109
rect -1639 -2149 -1287 -2143
rect -1221 -2109 -869 -2103
rect -1221 -2143 -1209 -2109
rect -881 -2143 -869 -2109
rect -1221 -2149 -869 -2143
rect -803 -2109 -451 -2103
rect -803 -2143 -791 -2109
rect -463 -2143 -451 -2109
rect -803 -2149 -451 -2143
rect -385 -2109 -33 -2103
rect -385 -2143 -373 -2109
rect -45 -2143 -33 -2109
rect -385 -2149 -33 -2143
rect 33 -2109 385 -2103
rect 33 -2143 45 -2109
rect 373 -2143 385 -2109
rect 33 -2149 385 -2143
rect 451 -2109 803 -2103
rect 451 -2143 463 -2109
rect 791 -2143 803 -2109
rect 451 -2149 803 -2143
rect 869 -2109 1221 -2103
rect 869 -2143 881 -2109
rect 1209 -2143 1221 -2109
rect 869 -2149 1221 -2143
rect 1287 -2109 1639 -2103
rect 1287 -2143 1299 -2109
rect 1627 -2143 1639 -2109
rect 1287 -2149 1639 -2143
rect 1705 -2109 2057 -2103
rect 1705 -2143 1717 -2109
rect 2045 -2143 2057 -2109
rect 1705 -2149 2057 -2143
rect -2113 -2193 -2067 -2181
rect -2113 -2469 -2107 -2193
rect -2073 -2469 -2067 -2193
rect -2113 -2481 -2067 -2469
rect -1695 -2193 -1649 -2181
rect -1695 -2469 -1689 -2193
rect -1655 -2469 -1649 -2193
rect -1695 -2481 -1649 -2469
rect -1277 -2193 -1231 -2181
rect -1277 -2469 -1271 -2193
rect -1237 -2469 -1231 -2193
rect -1277 -2481 -1231 -2469
rect -859 -2193 -813 -2181
rect -859 -2469 -853 -2193
rect -819 -2469 -813 -2193
rect -859 -2481 -813 -2469
rect -441 -2193 -395 -2181
rect -441 -2469 -435 -2193
rect -401 -2469 -395 -2193
rect -441 -2481 -395 -2469
rect -23 -2193 23 -2181
rect -23 -2469 -17 -2193
rect 17 -2469 23 -2193
rect -23 -2481 23 -2469
rect 395 -2193 441 -2181
rect 395 -2469 401 -2193
rect 435 -2469 441 -2193
rect 395 -2481 441 -2469
rect 813 -2193 859 -2181
rect 813 -2469 819 -2193
rect 853 -2469 859 -2193
rect 813 -2481 859 -2469
rect 1231 -2193 1277 -2181
rect 1231 -2469 1237 -2193
rect 1271 -2469 1277 -2193
rect 1231 -2481 1277 -2469
rect 1649 -2193 1695 -2181
rect 1649 -2469 1655 -2193
rect 1689 -2469 1695 -2193
rect 1649 -2481 1695 -2469
rect 2067 -2193 2113 -2181
rect 2067 -2469 2073 -2193
rect 2107 -2469 2113 -2193
rect 2067 -2481 2113 -2469
rect -2057 -2519 -1705 -2513
rect -2057 -2553 -2045 -2519
rect -1717 -2553 -1705 -2519
rect -2057 -2559 -1705 -2553
rect -1639 -2519 -1287 -2513
rect -1639 -2553 -1627 -2519
rect -1299 -2553 -1287 -2519
rect -1639 -2559 -1287 -2553
rect -1221 -2519 -869 -2513
rect -1221 -2553 -1209 -2519
rect -881 -2553 -869 -2519
rect -1221 -2559 -869 -2553
rect -803 -2519 -451 -2513
rect -803 -2553 -791 -2519
rect -463 -2553 -451 -2519
rect -803 -2559 -451 -2553
rect -385 -2519 -33 -2513
rect -385 -2553 -373 -2519
rect -45 -2553 -33 -2519
rect -385 -2559 -33 -2553
rect 33 -2519 385 -2513
rect 33 -2553 45 -2519
rect 373 -2553 385 -2519
rect 33 -2559 385 -2553
rect 451 -2519 803 -2513
rect 451 -2553 463 -2519
rect 791 -2553 803 -2519
rect 451 -2559 803 -2553
rect 869 -2519 1221 -2513
rect 869 -2553 881 -2519
rect 1209 -2553 1221 -2519
rect 869 -2559 1221 -2553
rect 1287 -2519 1639 -2513
rect 1287 -2553 1299 -2519
rect 1627 -2553 1639 -2519
rect 1287 -2559 1639 -2553
rect 1705 -2519 2057 -2513
rect 1705 -2553 1717 -2519
rect 2045 -2553 2057 -2519
rect 1705 -2559 2057 -2553
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2204 -2638 2204 2638
string parameters w 1.5 l 1.8 m 10 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
