magic
tech sky130A
magscale 1 2
timestamp 1619113446
<< error_p >>
rect -1421 2395 -1363 2401
rect -1229 2395 -1171 2401
rect -1037 2395 -979 2401
rect -845 2395 -787 2401
rect -653 2395 -595 2401
rect -461 2395 -403 2401
rect -269 2395 -211 2401
rect -77 2395 -19 2401
rect 115 2395 173 2401
rect 307 2395 365 2401
rect 499 2395 557 2401
rect 691 2395 749 2401
rect 883 2395 941 2401
rect 1075 2395 1133 2401
rect 1267 2395 1325 2401
rect -1421 2361 -1409 2395
rect -1229 2361 -1217 2395
rect -1037 2361 -1025 2395
rect -845 2361 -833 2395
rect -653 2361 -641 2395
rect -461 2361 -449 2395
rect -269 2361 -257 2395
rect -77 2361 -65 2395
rect 115 2361 127 2395
rect 307 2361 319 2395
rect 499 2361 511 2395
rect 691 2361 703 2395
rect 883 2361 895 2395
rect 1075 2361 1087 2395
rect 1267 2361 1279 2395
rect -1421 2355 -1363 2361
rect -1229 2355 -1171 2361
rect -1037 2355 -979 2361
rect -845 2355 -787 2361
rect -653 2355 -595 2361
rect -461 2355 -403 2361
rect -269 2355 -211 2361
rect -77 2355 -19 2361
rect 115 2355 173 2361
rect 307 2355 365 2361
rect 499 2355 557 2361
rect 691 2355 749 2361
rect 883 2355 941 2361
rect 1075 2355 1133 2361
rect 1267 2355 1325 2361
rect -1325 1895 -1267 1901
rect -1133 1895 -1075 1901
rect -941 1895 -883 1901
rect -749 1895 -691 1901
rect -557 1895 -499 1901
rect -365 1895 -307 1901
rect -173 1895 -115 1901
rect 19 1895 77 1901
rect 211 1895 269 1901
rect 403 1895 461 1901
rect 595 1895 653 1901
rect 787 1895 845 1901
rect 979 1895 1037 1901
rect 1171 1895 1229 1901
rect 1363 1895 1421 1901
rect -1325 1861 -1313 1895
rect -1133 1861 -1121 1895
rect -941 1861 -929 1895
rect -749 1861 -737 1895
rect -557 1861 -545 1895
rect -365 1861 -353 1895
rect -173 1861 -161 1895
rect 19 1861 31 1895
rect 211 1861 223 1895
rect 403 1861 415 1895
rect 595 1861 607 1895
rect 787 1861 799 1895
rect 979 1861 991 1895
rect 1171 1861 1183 1895
rect 1363 1861 1375 1895
rect -1325 1855 -1267 1861
rect -1133 1855 -1075 1861
rect -941 1855 -883 1861
rect -749 1855 -691 1861
rect -557 1855 -499 1861
rect -365 1855 -307 1861
rect -173 1855 -115 1861
rect 19 1855 77 1861
rect 211 1855 269 1861
rect 403 1855 461 1861
rect 595 1855 653 1861
rect 787 1855 845 1861
rect 979 1855 1037 1861
rect 1171 1855 1229 1861
rect 1363 1855 1421 1861
rect -1325 1787 -1267 1793
rect -1133 1787 -1075 1793
rect -941 1787 -883 1793
rect -749 1787 -691 1793
rect -557 1787 -499 1793
rect -365 1787 -307 1793
rect -173 1787 -115 1793
rect 19 1787 77 1793
rect 211 1787 269 1793
rect 403 1787 461 1793
rect 595 1787 653 1793
rect 787 1787 845 1793
rect 979 1787 1037 1793
rect 1171 1787 1229 1793
rect 1363 1787 1421 1793
rect -1325 1753 -1313 1787
rect -1133 1753 -1121 1787
rect -941 1753 -929 1787
rect -749 1753 -737 1787
rect -557 1753 -545 1787
rect -365 1753 -353 1787
rect -173 1753 -161 1787
rect 19 1753 31 1787
rect 211 1753 223 1787
rect 403 1753 415 1787
rect 595 1753 607 1787
rect 787 1753 799 1787
rect 979 1753 991 1787
rect 1171 1753 1183 1787
rect 1363 1753 1375 1787
rect -1325 1747 -1267 1753
rect -1133 1747 -1075 1753
rect -941 1747 -883 1753
rect -749 1747 -691 1753
rect -557 1747 -499 1753
rect -365 1747 -307 1753
rect -173 1747 -115 1753
rect 19 1747 77 1753
rect 211 1747 269 1753
rect 403 1747 461 1753
rect 595 1747 653 1753
rect 787 1747 845 1753
rect 979 1747 1037 1753
rect 1171 1747 1229 1753
rect 1363 1747 1421 1753
rect -1421 1287 -1363 1293
rect -1229 1287 -1171 1293
rect -1037 1287 -979 1293
rect -845 1287 -787 1293
rect -653 1287 -595 1293
rect -461 1287 -403 1293
rect -269 1287 -211 1293
rect -77 1287 -19 1293
rect 115 1287 173 1293
rect 307 1287 365 1293
rect 499 1287 557 1293
rect 691 1287 749 1293
rect 883 1287 941 1293
rect 1075 1287 1133 1293
rect 1267 1287 1325 1293
rect -1421 1253 -1409 1287
rect -1229 1253 -1217 1287
rect -1037 1253 -1025 1287
rect -845 1253 -833 1287
rect -653 1253 -641 1287
rect -461 1253 -449 1287
rect -269 1253 -257 1287
rect -77 1253 -65 1287
rect 115 1253 127 1287
rect 307 1253 319 1287
rect 499 1253 511 1287
rect 691 1253 703 1287
rect 883 1253 895 1287
rect 1075 1253 1087 1287
rect 1267 1253 1279 1287
rect -1421 1247 -1363 1253
rect -1229 1247 -1171 1253
rect -1037 1247 -979 1253
rect -845 1247 -787 1253
rect -653 1247 -595 1253
rect -461 1247 -403 1253
rect -269 1247 -211 1253
rect -77 1247 -19 1253
rect 115 1247 173 1253
rect 307 1247 365 1253
rect 499 1247 557 1253
rect 691 1247 749 1253
rect 883 1247 941 1253
rect 1075 1247 1133 1253
rect 1267 1247 1325 1253
rect -1421 1179 -1363 1185
rect -1229 1179 -1171 1185
rect -1037 1179 -979 1185
rect -845 1179 -787 1185
rect -653 1179 -595 1185
rect -461 1179 -403 1185
rect -269 1179 -211 1185
rect -77 1179 -19 1185
rect 115 1179 173 1185
rect 307 1179 365 1185
rect 499 1179 557 1185
rect 691 1179 749 1185
rect 883 1179 941 1185
rect 1075 1179 1133 1185
rect 1267 1179 1325 1185
rect -1421 1145 -1409 1179
rect -1229 1145 -1217 1179
rect -1037 1145 -1025 1179
rect -845 1145 -833 1179
rect -653 1145 -641 1179
rect -461 1145 -449 1179
rect -269 1145 -257 1179
rect -77 1145 -65 1179
rect 115 1145 127 1179
rect 307 1145 319 1179
rect 499 1145 511 1179
rect 691 1145 703 1179
rect 883 1145 895 1179
rect 1075 1145 1087 1179
rect 1267 1145 1279 1179
rect -1421 1139 -1363 1145
rect -1229 1139 -1171 1145
rect -1037 1139 -979 1145
rect -845 1139 -787 1145
rect -653 1139 -595 1145
rect -461 1139 -403 1145
rect -269 1139 -211 1145
rect -77 1139 -19 1145
rect 115 1139 173 1145
rect 307 1139 365 1145
rect 499 1139 557 1145
rect 691 1139 749 1145
rect 883 1139 941 1145
rect 1075 1139 1133 1145
rect 1267 1139 1325 1145
rect -1325 679 -1267 685
rect -1133 679 -1075 685
rect -941 679 -883 685
rect -749 679 -691 685
rect -557 679 -499 685
rect -365 679 -307 685
rect -173 679 -115 685
rect 19 679 77 685
rect 211 679 269 685
rect 403 679 461 685
rect 595 679 653 685
rect 787 679 845 685
rect 979 679 1037 685
rect 1171 679 1229 685
rect 1363 679 1421 685
rect -1325 645 -1313 679
rect -1133 645 -1121 679
rect -941 645 -929 679
rect -749 645 -737 679
rect -557 645 -545 679
rect -365 645 -353 679
rect -173 645 -161 679
rect 19 645 31 679
rect 211 645 223 679
rect 403 645 415 679
rect 595 645 607 679
rect 787 645 799 679
rect 979 645 991 679
rect 1171 645 1183 679
rect 1363 645 1375 679
rect -1325 639 -1267 645
rect -1133 639 -1075 645
rect -941 639 -883 645
rect -749 639 -691 645
rect -557 639 -499 645
rect -365 639 -307 645
rect -173 639 -115 645
rect 19 639 77 645
rect 211 639 269 645
rect 403 639 461 645
rect 595 639 653 645
rect 787 639 845 645
rect 979 639 1037 645
rect 1171 639 1229 645
rect 1363 639 1421 645
rect -1325 571 -1267 577
rect -1133 571 -1075 577
rect -941 571 -883 577
rect -749 571 -691 577
rect -557 571 -499 577
rect -365 571 -307 577
rect -173 571 -115 577
rect 19 571 77 577
rect 211 571 269 577
rect 403 571 461 577
rect 595 571 653 577
rect 787 571 845 577
rect 979 571 1037 577
rect 1171 571 1229 577
rect 1363 571 1421 577
rect -1325 537 -1313 571
rect -1133 537 -1121 571
rect -941 537 -929 571
rect -749 537 -737 571
rect -557 537 -545 571
rect -365 537 -353 571
rect -173 537 -161 571
rect 19 537 31 571
rect 211 537 223 571
rect 403 537 415 571
rect 595 537 607 571
rect 787 537 799 571
rect 979 537 991 571
rect 1171 537 1183 571
rect 1363 537 1375 571
rect -1325 531 -1267 537
rect -1133 531 -1075 537
rect -941 531 -883 537
rect -749 531 -691 537
rect -557 531 -499 537
rect -365 531 -307 537
rect -173 531 -115 537
rect 19 531 77 537
rect 211 531 269 537
rect 403 531 461 537
rect 595 531 653 537
rect 787 531 845 537
rect 979 531 1037 537
rect 1171 531 1229 537
rect 1363 531 1421 537
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect -1325 -537 -1267 -531
rect -1133 -537 -1075 -531
rect -941 -537 -883 -531
rect -749 -537 -691 -531
rect -557 -537 -499 -531
rect -365 -537 -307 -531
rect -173 -537 -115 -531
rect 19 -537 77 -531
rect 211 -537 269 -531
rect 403 -537 461 -531
rect 595 -537 653 -531
rect 787 -537 845 -531
rect 979 -537 1037 -531
rect 1171 -537 1229 -531
rect 1363 -537 1421 -531
rect -1325 -571 -1313 -537
rect -1133 -571 -1121 -537
rect -941 -571 -929 -537
rect -749 -571 -737 -537
rect -557 -571 -545 -537
rect -365 -571 -353 -537
rect -173 -571 -161 -537
rect 19 -571 31 -537
rect 211 -571 223 -537
rect 403 -571 415 -537
rect 595 -571 607 -537
rect 787 -571 799 -537
rect 979 -571 991 -537
rect 1171 -571 1183 -537
rect 1363 -571 1375 -537
rect -1325 -577 -1267 -571
rect -1133 -577 -1075 -571
rect -941 -577 -883 -571
rect -749 -577 -691 -571
rect -557 -577 -499 -571
rect -365 -577 -307 -571
rect -173 -577 -115 -571
rect 19 -577 77 -571
rect 211 -577 269 -571
rect 403 -577 461 -571
rect 595 -577 653 -571
rect 787 -577 845 -571
rect 979 -577 1037 -571
rect 1171 -577 1229 -571
rect 1363 -577 1421 -571
rect -1325 -645 -1267 -639
rect -1133 -645 -1075 -639
rect -941 -645 -883 -639
rect -749 -645 -691 -639
rect -557 -645 -499 -639
rect -365 -645 -307 -639
rect -173 -645 -115 -639
rect 19 -645 77 -639
rect 211 -645 269 -639
rect 403 -645 461 -639
rect 595 -645 653 -639
rect 787 -645 845 -639
rect 979 -645 1037 -639
rect 1171 -645 1229 -639
rect 1363 -645 1421 -639
rect -1325 -679 -1313 -645
rect -1133 -679 -1121 -645
rect -941 -679 -929 -645
rect -749 -679 -737 -645
rect -557 -679 -545 -645
rect -365 -679 -353 -645
rect -173 -679 -161 -645
rect 19 -679 31 -645
rect 211 -679 223 -645
rect 403 -679 415 -645
rect 595 -679 607 -645
rect 787 -679 799 -645
rect 979 -679 991 -645
rect 1171 -679 1183 -645
rect 1363 -679 1375 -645
rect -1325 -685 -1267 -679
rect -1133 -685 -1075 -679
rect -941 -685 -883 -679
rect -749 -685 -691 -679
rect -557 -685 -499 -679
rect -365 -685 -307 -679
rect -173 -685 -115 -679
rect 19 -685 77 -679
rect 211 -685 269 -679
rect 403 -685 461 -679
rect 595 -685 653 -679
rect 787 -685 845 -679
rect 979 -685 1037 -679
rect 1171 -685 1229 -679
rect 1363 -685 1421 -679
rect -1421 -1145 -1363 -1139
rect -1229 -1145 -1171 -1139
rect -1037 -1145 -979 -1139
rect -845 -1145 -787 -1139
rect -653 -1145 -595 -1139
rect -461 -1145 -403 -1139
rect -269 -1145 -211 -1139
rect -77 -1145 -19 -1139
rect 115 -1145 173 -1139
rect 307 -1145 365 -1139
rect 499 -1145 557 -1139
rect 691 -1145 749 -1139
rect 883 -1145 941 -1139
rect 1075 -1145 1133 -1139
rect 1267 -1145 1325 -1139
rect -1421 -1179 -1409 -1145
rect -1229 -1179 -1217 -1145
rect -1037 -1179 -1025 -1145
rect -845 -1179 -833 -1145
rect -653 -1179 -641 -1145
rect -461 -1179 -449 -1145
rect -269 -1179 -257 -1145
rect -77 -1179 -65 -1145
rect 115 -1179 127 -1145
rect 307 -1179 319 -1145
rect 499 -1179 511 -1145
rect 691 -1179 703 -1145
rect 883 -1179 895 -1145
rect 1075 -1179 1087 -1145
rect 1267 -1179 1279 -1145
rect -1421 -1185 -1363 -1179
rect -1229 -1185 -1171 -1179
rect -1037 -1185 -979 -1179
rect -845 -1185 -787 -1179
rect -653 -1185 -595 -1179
rect -461 -1185 -403 -1179
rect -269 -1185 -211 -1179
rect -77 -1185 -19 -1179
rect 115 -1185 173 -1179
rect 307 -1185 365 -1179
rect 499 -1185 557 -1179
rect 691 -1185 749 -1179
rect 883 -1185 941 -1179
rect 1075 -1185 1133 -1179
rect 1267 -1185 1325 -1179
rect -1421 -1253 -1363 -1247
rect -1229 -1253 -1171 -1247
rect -1037 -1253 -979 -1247
rect -845 -1253 -787 -1247
rect -653 -1253 -595 -1247
rect -461 -1253 -403 -1247
rect -269 -1253 -211 -1247
rect -77 -1253 -19 -1247
rect 115 -1253 173 -1247
rect 307 -1253 365 -1247
rect 499 -1253 557 -1247
rect 691 -1253 749 -1247
rect 883 -1253 941 -1247
rect 1075 -1253 1133 -1247
rect 1267 -1253 1325 -1247
rect -1421 -1287 -1409 -1253
rect -1229 -1287 -1217 -1253
rect -1037 -1287 -1025 -1253
rect -845 -1287 -833 -1253
rect -653 -1287 -641 -1253
rect -461 -1287 -449 -1253
rect -269 -1287 -257 -1253
rect -77 -1287 -65 -1253
rect 115 -1287 127 -1253
rect 307 -1287 319 -1253
rect 499 -1287 511 -1253
rect 691 -1287 703 -1253
rect 883 -1287 895 -1253
rect 1075 -1287 1087 -1253
rect 1267 -1287 1279 -1253
rect -1421 -1293 -1363 -1287
rect -1229 -1293 -1171 -1287
rect -1037 -1293 -979 -1287
rect -845 -1293 -787 -1287
rect -653 -1293 -595 -1287
rect -461 -1293 -403 -1287
rect -269 -1293 -211 -1287
rect -77 -1293 -19 -1287
rect 115 -1293 173 -1287
rect 307 -1293 365 -1287
rect 499 -1293 557 -1287
rect 691 -1293 749 -1287
rect 883 -1293 941 -1287
rect 1075 -1293 1133 -1287
rect 1267 -1293 1325 -1287
rect -1325 -1753 -1267 -1747
rect -1133 -1753 -1075 -1747
rect -941 -1753 -883 -1747
rect -749 -1753 -691 -1747
rect -557 -1753 -499 -1747
rect -365 -1753 -307 -1747
rect -173 -1753 -115 -1747
rect 19 -1753 77 -1747
rect 211 -1753 269 -1747
rect 403 -1753 461 -1747
rect 595 -1753 653 -1747
rect 787 -1753 845 -1747
rect 979 -1753 1037 -1747
rect 1171 -1753 1229 -1747
rect 1363 -1753 1421 -1747
rect -1325 -1787 -1313 -1753
rect -1133 -1787 -1121 -1753
rect -941 -1787 -929 -1753
rect -749 -1787 -737 -1753
rect -557 -1787 -545 -1753
rect -365 -1787 -353 -1753
rect -173 -1787 -161 -1753
rect 19 -1787 31 -1753
rect 211 -1787 223 -1753
rect 403 -1787 415 -1753
rect 595 -1787 607 -1753
rect 787 -1787 799 -1753
rect 979 -1787 991 -1753
rect 1171 -1787 1183 -1753
rect 1363 -1787 1375 -1753
rect -1325 -1793 -1267 -1787
rect -1133 -1793 -1075 -1787
rect -941 -1793 -883 -1787
rect -749 -1793 -691 -1787
rect -557 -1793 -499 -1787
rect -365 -1793 -307 -1787
rect -173 -1793 -115 -1787
rect 19 -1793 77 -1787
rect 211 -1793 269 -1787
rect 403 -1793 461 -1787
rect 595 -1793 653 -1787
rect 787 -1793 845 -1787
rect 979 -1793 1037 -1787
rect 1171 -1793 1229 -1787
rect 1363 -1793 1421 -1787
rect -1325 -1861 -1267 -1855
rect -1133 -1861 -1075 -1855
rect -941 -1861 -883 -1855
rect -749 -1861 -691 -1855
rect -557 -1861 -499 -1855
rect -365 -1861 -307 -1855
rect -173 -1861 -115 -1855
rect 19 -1861 77 -1855
rect 211 -1861 269 -1855
rect 403 -1861 461 -1855
rect 595 -1861 653 -1855
rect 787 -1861 845 -1855
rect 979 -1861 1037 -1855
rect 1171 -1861 1229 -1855
rect 1363 -1861 1421 -1855
rect -1325 -1895 -1313 -1861
rect -1133 -1895 -1121 -1861
rect -941 -1895 -929 -1861
rect -749 -1895 -737 -1861
rect -557 -1895 -545 -1861
rect -365 -1895 -353 -1861
rect -173 -1895 -161 -1861
rect 19 -1895 31 -1861
rect 211 -1895 223 -1861
rect 403 -1895 415 -1861
rect 595 -1895 607 -1861
rect 787 -1895 799 -1861
rect 979 -1895 991 -1861
rect 1171 -1895 1183 -1861
rect 1363 -1895 1375 -1861
rect -1325 -1901 -1267 -1895
rect -1133 -1901 -1075 -1895
rect -941 -1901 -883 -1895
rect -749 -1901 -691 -1895
rect -557 -1901 -499 -1895
rect -365 -1901 -307 -1895
rect -173 -1901 -115 -1895
rect 19 -1901 77 -1895
rect 211 -1901 269 -1895
rect 403 -1901 461 -1895
rect 595 -1901 653 -1895
rect 787 -1901 845 -1895
rect 979 -1901 1037 -1895
rect 1171 -1901 1229 -1895
rect 1363 -1901 1421 -1895
rect -1421 -2361 -1363 -2355
rect -1229 -2361 -1171 -2355
rect -1037 -2361 -979 -2355
rect -845 -2361 -787 -2355
rect -653 -2361 -595 -2355
rect -461 -2361 -403 -2355
rect -269 -2361 -211 -2355
rect -77 -2361 -19 -2355
rect 115 -2361 173 -2355
rect 307 -2361 365 -2355
rect 499 -2361 557 -2355
rect 691 -2361 749 -2355
rect 883 -2361 941 -2355
rect 1075 -2361 1133 -2355
rect 1267 -2361 1325 -2355
rect -1421 -2395 -1409 -2361
rect -1229 -2395 -1217 -2361
rect -1037 -2395 -1025 -2361
rect -845 -2395 -833 -2361
rect -653 -2395 -641 -2361
rect -461 -2395 -449 -2361
rect -269 -2395 -257 -2361
rect -77 -2395 -65 -2361
rect 115 -2395 127 -2361
rect 307 -2395 319 -2361
rect 499 -2395 511 -2361
rect 691 -2395 703 -2361
rect 883 -2395 895 -2361
rect 1075 -2395 1087 -2361
rect 1267 -2395 1279 -2361
rect -1421 -2401 -1363 -2395
rect -1229 -2401 -1171 -2395
rect -1037 -2401 -979 -2395
rect -845 -2401 -787 -2395
rect -653 -2401 -595 -2395
rect -461 -2401 -403 -2395
rect -269 -2401 -211 -2395
rect -77 -2401 -19 -2395
rect 115 -2401 173 -2395
rect 307 -2401 365 -2395
rect 499 -2401 557 -2395
rect 691 -2401 749 -2395
rect 883 -2401 941 -2395
rect 1075 -2401 1133 -2395
rect 1267 -2401 1325 -2395
<< pwell >>
rect -1607 -2533 1607 2533
<< nmos >>
rect -1407 1933 -1377 2323
rect -1311 1933 -1281 2323
rect -1215 1933 -1185 2323
rect -1119 1933 -1089 2323
rect -1023 1933 -993 2323
rect -927 1933 -897 2323
rect -831 1933 -801 2323
rect -735 1933 -705 2323
rect -639 1933 -609 2323
rect -543 1933 -513 2323
rect -447 1933 -417 2323
rect -351 1933 -321 2323
rect -255 1933 -225 2323
rect -159 1933 -129 2323
rect -63 1933 -33 2323
rect 33 1933 63 2323
rect 129 1933 159 2323
rect 225 1933 255 2323
rect 321 1933 351 2323
rect 417 1933 447 2323
rect 513 1933 543 2323
rect 609 1933 639 2323
rect 705 1933 735 2323
rect 801 1933 831 2323
rect 897 1933 927 2323
rect 993 1933 1023 2323
rect 1089 1933 1119 2323
rect 1185 1933 1215 2323
rect 1281 1933 1311 2323
rect 1377 1933 1407 2323
rect -1407 1325 -1377 1715
rect -1311 1325 -1281 1715
rect -1215 1325 -1185 1715
rect -1119 1325 -1089 1715
rect -1023 1325 -993 1715
rect -927 1325 -897 1715
rect -831 1325 -801 1715
rect -735 1325 -705 1715
rect -639 1325 -609 1715
rect -543 1325 -513 1715
rect -447 1325 -417 1715
rect -351 1325 -321 1715
rect -255 1325 -225 1715
rect -159 1325 -129 1715
rect -63 1325 -33 1715
rect 33 1325 63 1715
rect 129 1325 159 1715
rect 225 1325 255 1715
rect 321 1325 351 1715
rect 417 1325 447 1715
rect 513 1325 543 1715
rect 609 1325 639 1715
rect 705 1325 735 1715
rect 801 1325 831 1715
rect 897 1325 927 1715
rect 993 1325 1023 1715
rect 1089 1325 1119 1715
rect 1185 1325 1215 1715
rect 1281 1325 1311 1715
rect 1377 1325 1407 1715
rect -1407 717 -1377 1107
rect -1311 717 -1281 1107
rect -1215 717 -1185 1107
rect -1119 717 -1089 1107
rect -1023 717 -993 1107
rect -927 717 -897 1107
rect -831 717 -801 1107
rect -735 717 -705 1107
rect -639 717 -609 1107
rect -543 717 -513 1107
rect -447 717 -417 1107
rect -351 717 -321 1107
rect -255 717 -225 1107
rect -159 717 -129 1107
rect -63 717 -33 1107
rect 33 717 63 1107
rect 129 717 159 1107
rect 225 717 255 1107
rect 321 717 351 1107
rect 417 717 447 1107
rect 513 717 543 1107
rect 609 717 639 1107
rect 705 717 735 1107
rect 801 717 831 1107
rect 897 717 927 1107
rect 993 717 1023 1107
rect 1089 717 1119 1107
rect 1185 717 1215 1107
rect 1281 717 1311 1107
rect 1377 717 1407 1107
rect -1407 109 -1377 499
rect -1311 109 -1281 499
rect -1215 109 -1185 499
rect -1119 109 -1089 499
rect -1023 109 -993 499
rect -927 109 -897 499
rect -831 109 -801 499
rect -735 109 -705 499
rect -639 109 -609 499
rect -543 109 -513 499
rect -447 109 -417 499
rect -351 109 -321 499
rect -255 109 -225 499
rect -159 109 -129 499
rect -63 109 -33 499
rect 33 109 63 499
rect 129 109 159 499
rect 225 109 255 499
rect 321 109 351 499
rect 417 109 447 499
rect 513 109 543 499
rect 609 109 639 499
rect 705 109 735 499
rect 801 109 831 499
rect 897 109 927 499
rect 993 109 1023 499
rect 1089 109 1119 499
rect 1185 109 1215 499
rect 1281 109 1311 499
rect 1377 109 1407 499
rect -1407 -499 -1377 -109
rect -1311 -499 -1281 -109
rect -1215 -499 -1185 -109
rect -1119 -499 -1089 -109
rect -1023 -499 -993 -109
rect -927 -499 -897 -109
rect -831 -499 -801 -109
rect -735 -499 -705 -109
rect -639 -499 -609 -109
rect -543 -499 -513 -109
rect -447 -499 -417 -109
rect -351 -499 -321 -109
rect -255 -499 -225 -109
rect -159 -499 -129 -109
rect -63 -499 -33 -109
rect 33 -499 63 -109
rect 129 -499 159 -109
rect 225 -499 255 -109
rect 321 -499 351 -109
rect 417 -499 447 -109
rect 513 -499 543 -109
rect 609 -499 639 -109
rect 705 -499 735 -109
rect 801 -499 831 -109
rect 897 -499 927 -109
rect 993 -499 1023 -109
rect 1089 -499 1119 -109
rect 1185 -499 1215 -109
rect 1281 -499 1311 -109
rect 1377 -499 1407 -109
rect -1407 -1107 -1377 -717
rect -1311 -1107 -1281 -717
rect -1215 -1107 -1185 -717
rect -1119 -1107 -1089 -717
rect -1023 -1107 -993 -717
rect -927 -1107 -897 -717
rect -831 -1107 -801 -717
rect -735 -1107 -705 -717
rect -639 -1107 -609 -717
rect -543 -1107 -513 -717
rect -447 -1107 -417 -717
rect -351 -1107 -321 -717
rect -255 -1107 -225 -717
rect -159 -1107 -129 -717
rect -63 -1107 -33 -717
rect 33 -1107 63 -717
rect 129 -1107 159 -717
rect 225 -1107 255 -717
rect 321 -1107 351 -717
rect 417 -1107 447 -717
rect 513 -1107 543 -717
rect 609 -1107 639 -717
rect 705 -1107 735 -717
rect 801 -1107 831 -717
rect 897 -1107 927 -717
rect 993 -1107 1023 -717
rect 1089 -1107 1119 -717
rect 1185 -1107 1215 -717
rect 1281 -1107 1311 -717
rect 1377 -1107 1407 -717
rect -1407 -1715 -1377 -1325
rect -1311 -1715 -1281 -1325
rect -1215 -1715 -1185 -1325
rect -1119 -1715 -1089 -1325
rect -1023 -1715 -993 -1325
rect -927 -1715 -897 -1325
rect -831 -1715 -801 -1325
rect -735 -1715 -705 -1325
rect -639 -1715 -609 -1325
rect -543 -1715 -513 -1325
rect -447 -1715 -417 -1325
rect -351 -1715 -321 -1325
rect -255 -1715 -225 -1325
rect -159 -1715 -129 -1325
rect -63 -1715 -33 -1325
rect 33 -1715 63 -1325
rect 129 -1715 159 -1325
rect 225 -1715 255 -1325
rect 321 -1715 351 -1325
rect 417 -1715 447 -1325
rect 513 -1715 543 -1325
rect 609 -1715 639 -1325
rect 705 -1715 735 -1325
rect 801 -1715 831 -1325
rect 897 -1715 927 -1325
rect 993 -1715 1023 -1325
rect 1089 -1715 1119 -1325
rect 1185 -1715 1215 -1325
rect 1281 -1715 1311 -1325
rect 1377 -1715 1407 -1325
rect -1407 -2323 -1377 -1933
rect -1311 -2323 -1281 -1933
rect -1215 -2323 -1185 -1933
rect -1119 -2323 -1089 -1933
rect -1023 -2323 -993 -1933
rect -927 -2323 -897 -1933
rect -831 -2323 -801 -1933
rect -735 -2323 -705 -1933
rect -639 -2323 -609 -1933
rect -543 -2323 -513 -1933
rect -447 -2323 -417 -1933
rect -351 -2323 -321 -1933
rect -255 -2323 -225 -1933
rect -159 -2323 -129 -1933
rect -63 -2323 -33 -1933
rect 33 -2323 63 -1933
rect 129 -2323 159 -1933
rect 225 -2323 255 -1933
rect 321 -2323 351 -1933
rect 417 -2323 447 -1933
rect 513 -2323 543 -1933
rect 609 -2323 639 -1933
rect 705 -2323 735 -1933
rect 801 -2323 831 -1933
rect 897 -2323 927 -1933
rect 993 -2323 1023 -1933
rect 1089 -2323 1119 -1933
rect 1185 -2323 1215 -1933
rect 1281 -2323 1311 -1933
rect 1377 -2323 1407 -1933
<< ndiff >>
rect -1469 2311 -1407 2323
rect -1469 1945 -1457 2311
rect -1423 1945 -1407 2311
rect -1469 1933 -1407 1945
rect -1377 2311 -1311 2323
rect -1377 1945 -1361 2311
rect -1327 1945 -1311 2311
rect -1377 1933 -1311 1945
rect -1281 2311 -1215 2323
rect -1281 1945 -1265 2311
rect -1231 1945 -1215 2311
rect -1281 1933 -1215 1945
rect -1185 2311 -1119 2323
rect -1185 1945 -1169 2311
rect -1135 1945 -1119 2311
rect -1185 1933 -1119 1945
rect -1089 2311 -1023 2323
rect -1089 1945 -1073 2311
rect -1039 1945 -1023 2311
rect -1089 1933 -1023 1945
rect -993 2311 -927 2323
rect -993 1945 -977 2311
rect -943 1945 -927 2311
rect -993 1933 -927 1945
rect -897 2311 -831 2323
rect -897 1945 -881 2311
rect -847 1945 -831 2311
rect -897 1933 -831 1945
rect -801 2311 -735 2323
rect -801 1945 -785 2311
rect -751 1945 -735 2311
rect -801 1933 -735 1945
rect -705 2311 -639 2323
rect -705 1945 -689 2311
rect -655 1945 -639 2311
rect -705 1933 -639 1945
rect -609 2311 -543 2323
rect -609 1945 -593 2311
rect -559 1945 -543 2311
rect -609 1933 -543 1945
rect -513 2311 -447 2323
rect -513 1945 -497 2311
rect -463 1945 -447 2311
rect -513 1933 -447 1945
rect -417 2311 -351 2323
rect -417 1945 -401 2311
rect -367 1945 -351 2311
rect -417 1933 -351 1945
rect -321 2311 -255 2323
rect -321 1945 -305 2311
rect -271 1945 -255 2311
rect -321 1933 -255 1945
rect -225 2311 -159 2323
rect -225 1945 -209 2311
rect -175 1945 -159 2311
rect -225 1933 -159 1945
rect -129 2311 -63 2323
rect -129 1945 -113 2311
rect -79 1945 -63 2311
rect -129 1933 -63 1945
rect -33 2311 33 2323
rect -33 1945 -17 2311
rect 17 1945 33 2311
rect -33 1933 33 1945
rect 63 2311 129 2323
rect 63 1945 79 2311
rect 113 1945 129 2311
rect 63 1933 129 1945
rect 159 2311 225 2323
rect 159 1945 175 2311
rect 209 1945 225 2311
rect 159 1933 225 1945
rect 255 2311 321 2323
rect 255 1945 271 2311
rect 305 1945 321 2311
rect 255 1933 321 1945
rect 351 2311 417 2323
rect 351 1945 367 2311
rect 401 1945 417 2311
rect 351 1933 417 1945
rect 447 2311 513 2323
rect 447 1945 463 2311
rect 497 1945 513 2311
rect 447 1933 513 1945
rect 543 2311 609 2323
rect 543 1945 559 2311
rect 593 1945 609 2311
rect 543 1933 609 1945
rect 639 2311 705 2323
rect 639 1945 655 2311
rect 689 1945 705 2311
rect 639 1933 705 1945
rect 735 2311 801 2323
rect 735 1945 751 2311
rect 785 1945 801 2311
rect 735 1933 801 1945
rect 831 2311 897 2323
rect 831 1945 847 2311
rect 881 1945 897 2311
rect 831 1933 897 1945
rect 927 2311 993 2323
rect 927 1945 943 2311
rect 977 1945 993 2311
rect 927 1933 993 1945
rect 1023 2311 1089 2323
rect 1023 1945 1039 2311
rect 1073 1945 1089 2311
rect 1023 1933 1089 1945
rect 1119 2311 1185 2323
rect 1119 1945 1135 2311
rect 1169 1945 1185 2311
rect 1119 1933 1185 1945
rect 1215 2311 1281 2323
rect 1215 1945 1231 2311
rect 1265 1945 1281 2311
rect 1215 1933 1281 1945
rect 1311 2311 1377 2323
rect 1311 1945 1327 2311
rect 1361 1945 1377 2311
rect 1311 1933 1377 1945
rect 1407 2311 1469 2323
rect 1407 1945 1423 2311
rect 1457 1945 1469 2311
rect 1407 1933 1469 1945
rect -1469 1703 -1407 1715
rect -1469 1337 -1457 1703
rect -1423 1337 -1407 1703
rect -1469 1325 -1407 1337
rect -1377 1703 -1311 1715
rect -1377 1337 -1361 1703
rect -1327 1337 -1311 1703
rect -1377 1325 -1311 1337
rect -1281 1703 -1215 1715
rect -1281 1337 -1265 1703
rect -1231 1337 -1215 1703
rect -1281 1325 -1215 1337
rect -1185 1703 -1119 1715
rect -1185 1337 -1169 1703
rect -1135 1337 -1119 1703
rect -1185 1325 -1119 1337
rect -1089 1703 -1023 1715
rect -1089 1337 -1073 1703
rect -1039 1337 -1023 1703
rect -1089 1325 -1023 1337
rect -993 1703 -927 1715
rect -993 1337 -977 1703
rect -943 1337 -927 1703
rect -993 1325 -927 1337
rect -897 1703 -831 1715
rect -897 1337 -881 1703
rect -847 1337 -831 1703
rect -897 1325 -831 1337
rect -801 1703 -735 1715
rect -801 1337 -785 1703
rect -751 1337 -735 1703
rect -801 1325 -735 1337
rect -705 1703 -639 1715
rect -705 1337 -689 1703
rect -655 1337 -639 1703
rect -705 1325 -639 1337
rect -609 1703 -543 1715
rect -609 1337 -593 1703
rect -559 1337 -543 1703
rect -609 1325 -543 1337
rect -513 1703 -447 1715
rect -513 1337 -497 1703
rect -463 1337 -447 1703
rect -513 1325 -447 1337
rect -417 1703 -351 1715
rect -417 1337 -401 1703
rect -367 1337 -351 1703
rect -417 1325 -351 1337
rect -321 1703 -255 1715
rect -321 1337 -305 1703
rect -271 1337 -255 1703
rect -321 1325 -255 1337
rect -225 1703 -159 1715
rect -225 1337 -209 1703
rect -175 1337 -159 1703
rect -225 1325 -159 1337
rect -129 1703 -63 1715
rect -129 1337 -113 1703
rect -79 1337 -63 1703
rect -129 1325 -63 1337
rect -33 1703 33 1715
rect -33 1337 -17 1703
rect 17 1337 33 1703
rect -33 1325 33 1337
rect 63 1703 129 1715
rect 63 1337 79 1703
rect 113 1337 129 1703
rect 63 1325 129 1337
rect 159 1703 225 1715
rect 159 1337 175 1703
rect 209 1337 225 1703
rect 159 1325 225 1337
rect 255 1703 321 1715
rect 255 1337 271 1703
rect 305 1337 321 1703
rect 255 1325 321 1337
rect 351 1703 417 1715
rect 351 1337 367 1703
rect 401 1337 417 1703
rect 351 1325 417 1337
rect 447 1703 513 1715
rect 447 1337 463 1703
rect 497 1337 513 1703
rect 447 1325 513 1337
rect 543 1703 609 1715
rect 543 1337 559 1703
rect 593 1337 609 1703
rect 543 1325 609 1337
rect 639 1703 705 1715
rect 639 1337 655 1703
rect 689 1337 705 1703
rect 639 1325 705 1337
rect 735 1703 801 1715
rect 735 1337 751 1703
rect 785 1337 801 1703
rect 735 1325 801 1337
rect 831 1703 897 1715
rect 831 1337 847 1703
rect 881 1337 897 1703
rect 831 1325 897 1337
rect 927 1703 993 1715
rect 927 1337 943 1703
rect 977 1337 993 1703
rect 927 1325 993 1337
rect 1023 1703 1089 1715
rect 1023 1337 1039 1703
rect 1073 1337 1089 1703
rect 1023 1325 1089 1337
rect 1119 1703 1185 1715
rect 1119 1337 1135 1703
rect 1169 1337 1185 1703
rect 1119 1325 1185 1337
rect 1215 1703 1281 1715
rect 1215 1337 1231 1703
rect 1265 1337 1281 1703
rect 1215 1325 1281 1337
rect 1311 1703 1377 1715
rect 1311 1337 1327 1703
rect 1361 1337 1377 1703
rect 1311 1325 1377 1337
rect 1407 1703 1469 1715
rect 1407 1337 1423 1703
rect 1457 1337 1469 1703
rect 1407 1325 1469 1337
rect -1469 1095 -1407 1107
rect -1469 729 -1457 1095
rect -1423 729 -1407 1095
rect -1469 717 -1407 729
rect -1377 1095 -1311 1107
rect -1377 729 -1361 1095
rect -1327 729 -1311 1095
rect -1377 717 -1311 729
rect -1281 1095 -1215 1107
rect -1281 729 -1265 1095
rect -1231 729 -1215 1095
rect -1281 717 -1215 729
rect -1185 1095 -1119 1107
rect -1185 729 -1169 1095
rect -1135 729 -1119 1095
rect -1185 717 -1119 729
rect -1089 1095 -1023 1107
rect -1089 729 -1073 1095
rect -1039 729 -1023 1095
rect -1089 717 -1023 729
rect -993 1095 -927 1107
rect -993 729 -977 1095
rect -943 729 -927 1095
rect -993 717 -927 729
rect -897 1095 -831 1107
rect -897 729 -881 1095
rect -847 729 -831 1095
rect -897 717 -831 729
rect -801 1095 -735 1107
rect -801 729 -785 1095
rect -751 729 -735 1095
rect -801 717 -735 729
rect -705 1095 -639 1107
rect -705 729 -689 1095
rect -655 729 -639 1095
rect -705 717 -639 729
rect -609 1095 -543 1107
rect -609 729 -593 1095
rect -559 729 -543 1095
rect -609 717 -543 729
rect -513 1095 -447 1107
rect -513 729 -497 1095
rect -463 729 -447 1095
rect -513 717 -447 729
rect -417 1095 -351 1107
rect -417 729 -401 1095
rect -367 729 -351 1095
rect -417 717 -351 729
rect -321 1095 -255 1107
rect -321 729 -305 1095
rect -271 729 -255 1095
rect -321 717 -255 729
rect -225 1095 -159 1107
rect -225 729 -209 1095
rect -175 729 -159 1095
rect -225 717 -159 729
rect -129 1095 -63 1107
rect -129 729 -113 1095
rect -79 729 -63 1095
rect -129 717 -63 729
rect -33 1095 33 1107
rect -33 729 -17 1095
rect 17 729 33 1095
rect -33 717 33 729
rect 63 1095 129 1107
rect 63 729 79 1095
rect 113 729 129 1095
rect 63 717 129 729
rect 159 1095 225 1107
rect 159 729 175 1095
rect 209 729 225 1095
rect 159 717 225 729
rect 255 1095 321 1107
rect 255 729 271 1095
rect 305 729 321 1095
rect 255 717 321 729
rect 351 1095 417 1107
rect 351 729 367 1095
rect 401 729 417 1095
rect 351 717 417 729
rect 447 1095 513 1107
rect 447 729 463 1095
rect 497 729 513 1095
rect 447 717 513 729
rect 543 1095 609 1107
rect 543 729 559 1095
rect 593 729 609 1095
rect 543 717 609 729
rect 639 1095 705 1107
rect 639 729 655 1095
rect 689 729 705 1095
rect 639 717 705 729
rect 735 1095 801 1107
rect 735 729 751 1095
rect 785 729 801 1095
rect 735 717 801 729
rect 831 1095 897 1107
rect 831 729 847 1095
rect 881 729 897 1095
rect 831 717 897 729
rect 927 1095 993 1107
rect 927 729 943 1095
rect 977 729 993 1095
rect 927 717 993 729
rect 1023 1095 1089 1107
rect 1023 729 1039 1095
rect 1073 729 1089 1095
rect 1023 717 1089 729
rect 1119 1095 1185 1107
rect 1119 729 1135 1095
rect 1169 729 1185 1095
rect 1119 717 1185 729
rect 1215 1095 1281 1107
rect 1215 729 1231 1095
rect 1265 729 1281 1095
rect 1215 717 1281 729
rect 1311 1095 1377 1107
rect 1311 729 1327 1095
rect 1361 729 1377 1095
rect 1311 717 1377 729
rect 1407 1095 1469 1107
rect 1407 729 1423 1095
rect 1457 729 1469 1095
rect 1407 717 1469 729
rect -1469 487 -1407 499
rect -1469 121 -1457 487
rect -1423 121 -1407 487
rect -1469 109 -1407 121
rect -1377 487 -1311 499
rect -1377 121 -1361 487
rect -1327 121 -1311 487
rect -1377 109 -1311 121
rect -1281 487 -1215 499
rect -1281 121 -1265 487
rect -1231 121 -1215 487
rect -1281 109 -1215 121
rect -1185 487 -1119 499
rect -1185 121 -1169 487
rect -1135 121 -1119 487
rect -1185 109 -1119 121
rect -1089 487 -1023 499
rect -1089 121 -1073 487
rect -1039 121 -1023 487
rect -1089 109 -1023 121
rect -993 487 -927 499
rect -993 121 -977 487
rect -943 121 -927 487
rect -993 109 -927 121
rect -897 487 -831 499
rect -897 121 -881 487
rect -847 121 -831 487
rect -897 109 -831 121
rect -801 487 -735 499
rect -801 121 -785 487
rect -751 121 -735 487
rect -801 109 -735 121
rect -705 487 -639 499
rect -705 121 -689 487
rect -655 121 -639 487
rect -705 109 -639 121
rect -609 487 -543 499
rect -609 121 -593 487
rect -559 121 -543 487
rect -609 109 -543 121
rect -513 487 -447 499
rect -513 121 -497 487
rect -463 121 -447 487
rect -513 109 -447 121
rect -417 487 -351 499
rect -417 121 -401 487
rect -367 121 -351 487
rect -417 109 -351 121
rect -321 487 -255 499
rect -321 121 -305 487
rect -271 121 -255 487
rect -321 109 -255 121
rect -225 487 -159 499
rect -225 121 -209 487
rect -175 121 -159 487
rect -225 109 -159 121
rect -129 487 -63 499
rect -129 121 -113 487
rect -79 121 -63 487
rect -129 109 -63 121
rect -33 487 33 499
rect -33 121 -17 487
rect 17 121 33 487
rect -33 109 33 121
rect 63 487 129 499
rect 63 121 79 487
rect 113 121 129 487
rect 63 109 129 121
rect 159 487 225 499
rect 159 121 175 487
rect 209 121 225 487
rect 159 109 225 121
rect 255 487 321 499
rect 255 121 271 487
rect 305 121 321 487
rect 255 109 321 121
rect 351 487 417 499
rect 351 121 367 487
rect 401 121 417 487
rect 351 109 417 121
rect 447 487 513 499
rect 447 121 463 487
rect 497 121 513 487
rect 447 109 513 121
rect 543 487 609 499
rect 543 121 559 487
rect 593 121 609 487
rect 543 109 609 121
rect 639 487 705 499
rect 639 121 655 487
rect 689 121 705 487
rect 639 109 705 121
rect 735 487 801 499
rect 735 121 751 487
rect 785 121 801 487
rect 735 109 801 121
rect 831 487 897 499
rect 831 121 847 487
rect 881 121 897 487
rect 831 109 897 121
rect 927 487 993 499
rect 927 121 943 487
rect 977 121 993 487
rect 927 109 993 121
rect 1023 487 1089 499
rect 1023 121 1039 487
rect 1073 121 1089 487
rect 1023 109 1089 121
rect 1119 487 1185 499
rect 1119 121 1135 487
rect 1169 121 1185 487
rect 1119 109 1185 121
rect 1215 487 1281 499
rect 1215 121 1231 487
rect 1265 121 1281 487
rect 1215 109 1281 121
rect 1311 487 1377 499
rect 1311 121 1327 487
rect 1361 121 1377 487
rect 1311 109 1377 121
rect 1407 487 1469 499
rect 1407 121 1423 487
rect 1457 121 1469 487
rect 1407 109 1469 121
rect -1469 -121 -1407 -109
rect -1469 -487 -1457 -121
rect -1423 -487 -1407 -121
rect -1469 -499 -1407 -487
rect -1377 -121 -1311 -109
rect -1377 -487 -1361 -121
rect -1327 -487 -1311 -121
rect -1377 -499 -1311 -487
rect -1281 -121 -1215 -109
rect -1281 -487 -1265 -121
rect -1231 -487 -1215 -121
rect -1281 -499 -1215 -487
rect -1185 -121 -1119 -109
rect -1185 -487 -1169 -121
rect -1135 -487 -1119 -121
rect -1185 -499 -1119 -487
rect -1089 -121 -1023 -109
rect -1089 -487 -1073 -121
rect -1039 -487 -1023 -121
rect -1089 -499 -1023 -487
rect -993 -121 -927 -109
rect -993 -487 -977 -121
rect -943 -487 -927 -121
rect -993 -499 -927 -487
rect -897 -121 -831 -109
rect -897 -487 -881 -121
rect -847 -487 -831 -121
rect -897 -499 -831 -487
rect -801 -121 -735 -109
rect -801 -487 -785 -121
rect -751 -487 -735 -121
rect -801 -499 -735 -487
rect -705 -121 -639 -109
rect -705 -487 -689 -121
rect -655 -487 -639 -121
rect -705 -499 -639 -487
rect -609 -121 -543 -109
rect -609 -487 -593 -121
rect -559 -487 -543 -121
rect -609 -499 -543 -487
rect -513 -121 -447 -109
rect -513 -487 -497 -121
rect -463 -487 -447 -121
rect -513 -499 -447 -487
rect -417 -121 -351 -109
rect -417 -487 -401 -121
rect -367 -487 -351 -121
rect -417 -499 -351 -487
rect -321 -121 -255 -109
rect -321 -487 -305 -121
rect -271 -487 -255 -121
rect -321 -499 -255 -487
rect -225 -121 -159 -109
rect -225 -487 -209 -121
rect -175 -487 -159 -121
rect -225 -499 -159 -487
rect -129 -121 -63 -109
rect -129 -487 -113 -121
rect -79 -487 -63 -121
rect -129 -499 -63 -487
rect -33 -121 33 -109
rect -33 -487 -17 -121
rect 17 -487 33 -121
rect -33 -499 33 -487
rect 63 -121 129 -109
rect 63 -487 79 -121
rect 113 -487 129 -121
rect 63 -499 129 -487
rect 159 -121 225 -109
rect 159 -487 175 -121
rect 209 -487 225 -121
rect 159 -499 225 -487
rect 255 -121 321 -109
rect 255 -487 271 -121
rect 305 -487 321 -121
rect 255 -499 321 -487
rect 351 -121 417 -109
rect 351 -487 367 -121
rect 401 -487 417 -121
rect 351 -499 417 -487
rect 447 -121 513 -109
rect 447 -487 463 -121
rect 497 -487 513 -121
rect 447 -499 513 -487
rect 543 -121 609 -109
rect 543 -487 559 -121
rect 593 -487 609 -121
rect 543 -499 609 -487
rect 639 -121 705 -109
rect 639 -487 655 -121
rect 689 -487 705 -121
rect 639 -499 705 -487
rect 735 -121 801 -109
rect 735 -487 751 -121
rect 785 -487 801 -121
rect 735 -499 801 -487
rect 831 -121 897 -109
rect 831 -487 847 -121
rect 881 -487 897 -121
rect 831 -499 897 -487
rect 927 -121 993 -109
rect 927 -487 943 -121
rect 977 -487 993 -121
rect 927 -499 993 -487
rect 1023 -121 1089 -109
rect 1023 -487 1039 -121
rect 1073 -487 1089 -121
rect 1023 -499 1089 -487
rect 1119 -121 1185 -109
rect 1119 -487 1135 -121
rect 1169 -487 1185 -121
rect 1119 -499 1185 -487
rect 1215 -121 1281 -109
rect 1215 -487 1231 -121
rect 1265 -487 1281 -121
rect 1215 -499 1281 -487
rect 1311 -121 1377 -109
rect 1311 -487 1327 -121
rect 1361 -487 1377 -121
rect 1311 -499 1377 -487
rect 1407 -121 1469 -109
rect 1407 -487 1423 -121
rect 1457 -487 1469 -121
rect 1407 -499 1469 -487
rect -1469 -729 -1407 -717
rect -1469 -1095 -1457 -729
rect -1423 -1095 -1407 -729
rect -1469 -1107 -1407 -1095
rect -1377 -729 -1311 -717
rect -1377 -1095 -1361 -729
rect -1327 -1095 -1311 -729
rect -1377 -1107 -1311 -1095
rect -1281 -729 -1215 -717
rect -1281 -1095 -1265 -729
rect -1231 -1095 -1215 -729
rect -1281 -1107 -1215 -1095
rect -1185 -729 -1119 -717
rect -1185 -1095 -1169 -729
rect -1135 -1095 -1119 -729
rect -1185 -1107 -1119 -1095
rect -1089 -729 -1023 -717
rect -1089 -1095 -1073 -729
rect -1039 -1095 -1023 -729
rect -1089 -1107 -1023 -1095
rect -993 -729 -927 -717
rect -993 -1095 -977 -729
rect -943 -1095 -927 -729
rect -993 -1107 -927 -1095
rect -897 -729 -831 -717
rect -897 -1095 -881 -729
rect -847 -1095 -831 -729
rect -897 -1107 -831 -1095
rect -801 -729 -735 -717
rect -801 -1095 -785 -729
rect -751 -1095 -735 -729
rect -801 -1107 -735 -1095
rect -705 -729 -639 -717
rect -705 -1095 -689 -729
rect -655 -1095 -639 -729
rect -705 -1107 -639 -1095
rect -609 -729 -543 -717
rect -609 -1095 -593 -729
rect -559 -1095 -543 -729
rect -609 -1107 -543 -1095
rect -513 -729 -447 -717
rect -513 -1095 -497 -729
rect -463 -1095 -447 -729
rect -513 -1107 -447 -1095
rect -417 -729 -351 -717
rect -417 -1095 -401 -729
rect -367 -1095 -351 -729
rect -417 -1107 -351 -1095
rect -321 -729 -255 -717
rect -321 -1095 -305 -729
rect -271 -1095 -255 -729
rect -321 -1107 -255 -1095
rect -225 -729 -159 -717
rect -225 -1095 -209 -729
rect -175 -1095 -159 -729
rect -225 -1107 -159 -1095
rect -129 -729 -63 -717
rect -129 -1095 -113 -729
rect -79 -1095 -63 -729
rect -129 -1107 -63 -1095
rect -33 -729 33 -717
rect -33 -1095 -17 -729
rect 17 -1095 33 -729
rect -33 -1107 33 -1095
rect 63 -729 129 -717
rect 63 -1095 79 -729
rect 113 -1095 129 -729
rect 63 -1107 129 -1095
rect 159 -729 225 -717
rect 159 -1095 175 -729
rect 209 -1095 225 -729
rect 159 -1107 225 -1095
rect 255 -729 321 -717
rect 255 -1095 271 -729
rect 305 -1095 321 -729
rect 255 -1107 321 -1095
rect 351 -729 417 -717
rect 351 -1095 367 -729
rect 401 -1095 417 -729
rect 351 -1107 417 -1095
rect 447 -729 513 -717
rect 447 -1095 463 -729
rect 497 -1095 513 -729
rect 447 -1107 513 -1095
rect 543 -729 609 -717
rect 543 -1095 559 -729
rect 593 -1095 609 -729
rect 543 -1107 609 -1095
rect 639 -729 705 -717
rect 639 -1095 655 -729
rect 689 -1095 705 -729
rect 639 -1107 705 -1095
rect 735 -729 801 -717
rect 735 -1095 751 -729
rect 785 -1095 801 -729
rect 735 -1107 801 -1095
rect 831 -729 897 -717
rect 831 -1095 847 -729
rect 881 -1095 897 -729
rect 831 -1107 897 -1095
rect 927 -729 993 -717
rect 927 -1095 943 -729
rect 977 -1095 993 -729
rect 927 -1107 993 -1095
rect 1023 -729 1089 -717
rect 1023 -1095 1039 -729
rect 1073 -1095 1089 -729
rect 1023 -1107 1089 -1095
rect 1119 -729 1185 -717
rect 1119 -1095 1135 -729
rect 1169 -1095 1185 -729
rect 1119 -1107 1185 -1095
rect 1215 -729 1281 -717
rect 1215 -1095 1231 -729
rect 1265 -1095 1281 -729
rect 1215 -1107 1281 -1095
rect 1311 -729 1377 -717
rect 1311 -1095 1327 -729
rect 1361 -1095 1377 -729
rect 1311 -1107 1377 -1095
rect 1407 -729 1469 -717
rect 1407 -1095 1423 -729
rect 1457 -1095 1469 -729
rect 1407 -1107 1469 -1095
rect -1469 -1337 -1407 -1325
rect -1469 -1703 -1457 -1337
rect -1423 -1703 -1407 -1337
rect -1469 -1715 -1407 -1703
rect -1377 -1337 -1311 -1325
rect -1377 -1703 -1361 -1337
rect -1327 -1703 -1311 -1337
rect -1377 -1715 -1311 -1703
rect -1281 -1337 -1215 -1325
rect -1281 -1703 -1265 -1337
rect -1231 -1703 -1215 -1337
rect -1281 -1715 -1215 -1703
rect -1185 -1337 -1119 -1325
rect -1185 -1703 -1169 -1337
rect -1135 -1703 -1119 -1337
rect -1185 -1715 -1119 -1703
rect -1089 -1337 -1023 -1325
rect -1089 -1703 -1073 -1337
rect -1039 -1703 -1023 -1337
rect -1089 -1715 -1023 -1703
rect -993 -1337 -927 -1325
rect -993 -1703 -977 -1337
rect -943 -1703 -927 -1337
rect -993 -1715 -927 -1703
rect -897 -1337 -831 -1325
rect -897 -1703 -881 -1337
rect -847 -1703 -831 -1337
rect -897 -1715 -831 -1703
rect -801 -1337 -735 -1325
rect -801 -1703 -785 -1337
rect -751 -1703 -735 -1337
rect -801 -1715 -735 -1703
rect -705 -1337 -639 -1325
rect -705 -1703 -689 -1337
rect -655 -1703 -639 -1337
rect -705 -1715 -639 -1703
rect -609 -1337 -543 -1325
rect -609 -1703 -593 -1337
rect -559 -1703 -543 -1337
rect -609 -1715 -543 -1703
rect -513 -1337 -447 -1325
rect -513 -1703 -497 -1337
rect -463 -1703 -447 -1337
rect -513 -1715 -447 -1703
rect -417 -1337 -351 -1325
rect -417 -1703 -401 -1337
rect -367 -1703 -351 -1337
rect -417 -1715 -351 -1703
rect -321 -1337 -255 -1325
rect -321 -1703 -305 -1337
rect -271 -1703 -255 -1337
rect -321 -1715 -255 -1703
rect -225 -1337 -159 -1325
rect -225 -1703 -209 -1337
rect -175 -1703 -159 -1337
rect -225 -1715 -159 -1703
rect -129 -1337 -63 -1325
rect -129 -1703 -113 -1337
rect -79 -1703 -63 -1337
rect -129 -1715 -63 -1703
rect -33 -1337 33 -1325
rect -33 -1703 -17 -1337
rect 17 -1703 33 -1337
rect -33 -1715 33 -1703
rect 63 -1337 129 -1325
rect 63 -1703 79 -1337
rect 113 -1703 129 -1337
rect 63 -1715 129 -1703
rect 159 -1337 225 -1325
rect 159 -1703 175 -1337
rect 209 -1703 225 -1337
rect 159 -1715 225 -1703
rect 255 -1337 321 -1325
rect 255 -1703 271 -1337
rect 305 -1703 321 -1337
rect 255 -1715 321 -1703
rect 351 -1337 417 -1325
rect 351 -1703 367 -1337
rect 401 -1703 417 -1337
rect 351 -1715 417 -1703
rect 447 -1337 513 -1325
rect 447 -1703 463 -1337
rect 497 -1703 513 -1337
rect 447 -1715 513 -1703
rect 543 -1337 609 -1325
rect 543 -1703 559 -1337
rect 593 -1703 609 -1337
rect 543 -1715 609 -1703
rect 639 -1337 705 -1325
rect 639 -1703 655 -1337
rect 689 -1703 705 -1337
rect 639 -1715 705 -1703
rect 735 -1337 801 -1325
rect 735 -1703 751 -1337
rect 785 -1703 801 -1337
rect 735 -1715 801 -1703
rect 831 -1337 897 -1325
rect 831 -1703 847 -1337
rect 881 -1703 897 -1337
rect 831 -1715 897 -1703
rect 927 -1337 993 -1325
rect 927 -1703 943 -1337
rect 977 -1703 993 -1337
rect 927 -1715 993 -1703
rect 1023 -1337 1089 -1325
rect 1023 -1703 1039 -1337
rect 1073 -1703 1089 -1337
rect 1023 -1715 1089 -1703
rect 1119 -1337 1185 -1325
rect 1119 -1703 1135 -1337
rect 1169 -1703 1185 -1337
rect 1119 -1715 1185 -1703
rect 1215 -1337 1281 -1325
rect 1215 -1703 1231 -1337
rect 1265 -1703 1281 -1337
rect 1215 -1715 1281 -1703
rect 1311 -1337 1377 -1325
rect 1311 -1703 1327 -1337
rect 1361 -1703 1377 -1337
rect 1311 -1715 1377 -1703
rect 1407 -1337 1469 -1325
rect 1407 -1703 1423 -1337
rect 1457 -1703 1469 -1337
rect 1407 -1715 1469 -1703
rect -1469 -1945 -1407 -1933
rect -1469 -2311 -1457 -1945
rect -1423 -2311 -1407 -1945
rect -1469 -2323 -1407 -2311
rect -1377 -1945 -1311 -1933
rect -1377 -2311 -1361 -1945
rect -1327 -2311 -1311 -1945
rect -1377 -2323 -1311 -2311
rect -1281 -1945 -1215 -1933
rect -1281 -2311 -1265 -1945
rect -1231 -2311 -1215 -1945
rect -1281 -2323 -1215 -2311
rect -1185 -1945 -1119 -1933
rect -1185 -2311 -1169 -1945
rect -1135 -2311 -1119 -1945
rect -1185 -2323 -1119 -2311
rect -1089 -1945 -1023 -1933
rect -1089 -2311 -1073 -1945
rect -1039 -2311 -1023 -1945
rect -1089 -2323 -1023 -2311
rect -993 -1945 -927 -1933
rect -993 -2311 -977 -1945
rect -943 -2311 -927 -1945
rect -993 -2323 -927 -2311
rect -897 -1945 -831 -1933
rect -897 -2311 -881 -1945
rect -847 -2311 -831 -1945
rect -897 -2323 -831 -2311
rect -801 -1945 -735 -1933
rect -801 -2311 -785 -1945
rect -751 -2311 -735 -1945
rect -801 -2323 -735 -2311
rect -705 -1945 -639 -1933
rect -705 -2311 -689 -1945
rect -655 -2311 -639 -1945
rect -705 -2323 -639 -2311
rect -609 -1945 -543 -1933
rect -609 -2311 -593 -1945
rect -559 -2311 -543 -1945
rect -609 -2323 -543 -2311
rect -513 -1945 -447 -1933
rect -513 -2311 -497 -1945
rect -463 -2311 -447 -1945
rect -513 -2323 -447 -2311
rect -417 -1945 -351 -1933
rect -417 -2311 -401 -1945
rect -367 -2311 -351 -1945
rect -417 -2323 -351 -2311
rect -321 -1945 -255 -1933
rect -321 -2311 -305 -1945
rect -271 -2311 -255 -1945
rect -321 -2323 -255 -2311
rect -225 -1945 -159 -1933
rect -225 -2311 -209 -1945
rect -175 -2311 -159 -1945
rect -225 -2323 -159 -2311
rect -129 -1945 -63 -1933
rect -129 -2311 -113 -1945
rect -79 -2311 -63 -1945
rect -129 -2323 -63 -2311
rect -33 -1945 33 -1933
rect -33 -2311 -17 -1945
rect 17 -2311 33 -1945
rect -33 -2323 33 -2311
rect 63 -1945 129 -1933
rect 63 -2311 79 -1945
rect 113 -2311 129 -1945
rect 63 -2323 129 -2311
rect 159 -1945 225 -1933
rect 159 -2311 175 -1945
rect 209 -2311 225 -1945
rect 159 -2323 225 -2311
rect 255 -1945 321 -1933
rect 255 -2311 271 -1945
rect 305 -2311 321 -1945
rect 255 -2323 321 -2311
rect 351 -1945 417 -1933
rect 351 -2311 367 -1945
rect 401 -2311 417 -1945
rect 351 -2323 417 -2311
rect 447 -1945 513 -1933
rect 447 -2311 463 -1945
rect 497 -2311 513 -1945
rect 447 -2323 513 -2311
rect 543 -1945 609 -1933
rect 543 -2311 559 -1945
rect 593 -2311 609 -1945
rect 543 -2323 609 -2311
rect 639 -1945 705 -1933
rect 639 -2311 655 -1945
rect 689 -2311 705 -1945
rect 639 -2323 705 -2311
rect 735 -1945 801 -1933
rect 735 -2311 751 -1945
rect 785 -2311 801 -1945
rect 735 -2323 801 -2311
rect 831 -1945 897 -1933
rect 831 -2311 847 -1945
rect 881 -2311 897 -1945
rect 831 -2323 897 -2311
rect 927 -1945 993 -1933
rect 927 -2311 943 -1945
rect 977 -2311 993 -1945
rect 927 -2323 993 -2311
rect 1023 -1945 1089 -1933
rect 1023 -2311 1039 -1945
rect 1073 -2311 1089 -1945
rect 1023 -2323 1089 -2311
rect 1119 -1945 1185 -1933
rect 1119 -2311 1135 -1945
rect 1169 -2311 1185 -1945
rect 1119 -2323 1185 -2311
rect 1215 -1945 1281 -1933
rect 1215 -2311 1231 -1945
rect 1265 -2311 1281 -1945
rect 1215 -2323 1281 -2311
rect 1311 -1945 1377 -1933
rect 1311 -2311 1327 -1945
rect 1361 -2311 1377 -1945
rect 1311 -2323 1377 -2311
rect 1407 -1945 1469 -1933
rect 1407 -2311 1423 -1945
rect 1457 -2311 1469 -1945
rect 1407 -2323 1469 -2311
<< ndiffc >>
rect -1457 1945 -1423 2311
rect -1361 1945 -1327 2311
rect -1265 1945 -1231 2311
rect -1169 1945 -1135 2311
rect -1073 1945 -1039 2311
rect -977 1945 -943 2311
rect -881 1945 -847 2311
rect -785 1945 -751 2311
rect -689 1945 -655 2311
rect -593 1945 -559 2311
rect -497 1945 -463 2311
rect -401 1945 -367 2311
rect -305 1945 -271 2311
rect -209 1945 -175 2311
rect -113 1945 -79 2311
rect -17 1945 17 2311
rect 79 1945 113 2311
rect 175 1945 209 2311
rect 271 1945 305 2311
rect 367 1945 401 2311
rect 463 1945 497 2311
rect 559 1945 593 2311
rect 655 1945 689 2311
rect 751 1945 785 2311
rect 847 1945 881 2311
rect 943 1945 977 2311
rect 1039 1945 1073 2311
rect 1135 1945 1169 2311
rect 1231 1945 1265 2311
rect 1327 1945 1361 2311
rect 1423 1945 1457 2311
rect -1457 1337 -1423 1703
rect -1361 1337 -1327 1703
rect -1265 1337 -1231 1703
rect -1169 1337 -1135 1703
rect -1073 1337 -1039 1703
rect -977 1337 -943 1703
rect -881 1337 -847 1703
rect -785 1337 -751 1703
rect -689 1337 -655 1703
rect -593 1337 -559 1703
rect -497 1337 -463 1703
rect -401 1337 -367 1703
rect -305 1337 -271 1703
rect -209 1337 -175 1703
rect -113 1337 -79 1703
rect -17 1337 17 1703
rect 79 1337 113 1703
rect 175 1337 209 1703
rect 271 1337 305 1703
rect 367 1337 401 1703
rect 463 1337 497 1703
rect 559 1337 593 1703
rect 655 1337 689 1703
rect 751 1337 785 1703
rect 847 1337 881 1703
rect 943 1337 977 1703
rect 1039 1337 1073 1703
rect 1135 1337 1169 1703
rect 1231 1337 1265 1703
rect 1327 1337 1361 1703
rect 1423 1337 1457 1703
rect -1457 729 -1423 1095
rect -1361 729 -1327 1095
rect -1265 729 -1231 1095
rect -1169 729 -1135 1095
rect -1073 729 -1039 1095
rect -977 729 -943 1095
rect -881 729 -847 1095
rect -785 729 -751 1095
rect -689 729 -655 1095
rect -593 729 -559 1095
rect -497 729 -463 1095
rect -401 729 -367 1095
rect -305 729 -271 1095
rect -209 729 -175 1095
rect -113 729 -79 1095
rect -17 729 17 1095
rect 79 729 113 1095
rect 175 729 209 1095
rect 271 729 305 1095
rect 367 729 401 1095
rect 463 729 497 1095
rect 559 729 593 1095
rect 655 729 689 1095
rect 751 729 785 1095
rect 847 729 881 1095
rect 943 729 977 1095
rect 1039 729 1073 1095
rect 1135 729 1169 1095
rect 1231 729 1265 1095
rect 1327 729 1361 1095
rect 1423 729 1457 1095
rect -1457 121 -1423 487
rect -1361 121 -1327 487
rect -1265 121 -1231 487
rect -1169 121 -1135 487
rect -1073 121 -1039 487
rect -977 121 -943 487
rect -881 121 -847 487
rect -785 121 -751 487
rect -689 121 -655 487
rect -593 121 -559 487
rect -497 121 -463 487
rect -401 121 -367 487
rect -305 121 -271 487
rect -209 121 -175 487
rect -113 121 -79 487
rect -17 121 17 487
rect 79 121 113 487
rect 175 121 209 487
rect 271 121 305 487
rect 367 121 401 487
rect 463 121 497 487
rect 559 121 593 487
rect 655 121 689 487
rect 751 121 785 487
rect 847 121 881 487
rect 943 121 977 487
rect 1039 121 1073 487
rect 1135 121 1169 487
rect 1231 121 1265 487
rect 1327 121 1361 487
rect 1423 121 1457 487
rect -1457 -487 -1423 -121
rect -1361 -487 -1327 -121
rect -1265 -487 -1231 -121
rect -1169 -487 -1135 -121
rect -1073 -487 -1039 -121
rect -977 -487 -943 -121
rect -881 -487 -847 -121
rect -785 -487 -751 -121
rect -689 -487 -655 -121
rect -593 -487 -559 -121
rect -497 -487 -463 -121
rect -401 -487 -367 -121
rect -305 -487 -271 -121
rect -209 -487 -175 -121
rect -113 -487 -79 -121
rect -17 -487 17 -121
rect 79 -487 113 -121
rect 175 -487 209 -121
rect 271 -487 305 -121
rect 367 -487 401 -121
rect 463 -487 497 -121
rect 559 -487 593 -121
rect 655 -487 689 -121
rect 751 -487 785 -121
rect 847 -487 881 -121
rect 943 -487 977 -121
rect 1039 -487 1073 -121
rect 1135 -487 1169 -121
rect 1231 -487 1265 -121
rect 1327 -487 1361 -121
rect 1423 -487 1457 -121
rect -1457 -1095 -1423 -729
rect -1361 -1095 -1327 -729
rect -1265 -1095 -1231 -729
rect -1169 -1095 -1135 -729
rect -1073 -1095 -1039 -729
rect -977 -1095 -943 -729
rect -881 -1095 -847 -729
rect -785 -1095 -751 -729
rect -689 -1095 -655 -729
rect -593 -1095 -559 -729
rect -497 -1095 -463 -729
rect -401 -1095 -367 -729
rect -305 -1095 -271 -729
rect -209 -1095 -175 -729
rect -113 -1095 -79 -729
rect -17 -1095 17 -729
rect 79 -1095 113 -729
rect 175 -1095 209 -729
rect 271 -1095 305 -729
rect 367 -1095 401 -729
rect 463 -1095 497 -729
rect 559 -1095 593 -729
rect 655 -1095 689 -729
rect 751 -1095 785 -729
rect 847 -1095 881 -729
rect 943 -1095 977 -729
rect 1039 -1095 1073 -729
rect 1135 -1095 1169 -729
rect 1231 -1095 1265 -729
rect 1327 -1095 1361 -729
rect 1423 -1095 1457 -729
rect -1457 -1703 -1423 -1337
rect -1361 -1703 -1327 -1337
rect -1265 -1703 -1231 -1337
rect -1169 -1703 -1135 -1337
rect -1073 -1703 -1039 -1337
rect -977 -1703 -943 -1337
rect -881 -1703 -847 -1337
rect -785 -1703 -751 -1337
rect -689 -1703 -655 -1337
rect -593 -1703 -559 -1337
rect -497 -1703 -463 -1337
rect -401 -1703 -367 -1337
rect -305 -1703 -271 -1337
rect -209 -1703 -175 -1337
rect -113 -1703 -79 -1337
rect -17 -1703 17 -1337
rect 79 -1703 113 -1337
rect 175 -1703 209 -1337
rect 271 -1703 305 -1337
rect 367 -1703 401 -1337
rect 463 -1703 497 -1337
rect 559 -1703 593 -1337
rect 655 -1703 689 -1337
rect 751 -1703 785 -1337
rect 847 -1703 881 -1337
rect 943 -1703 977 -1337
rect 1039 -1703 1073 -1337
rect 1135 -1703 1169 -1337
rect 1231 -1703 1265 -1337
rect 1327 -1703 1361 -1337
rect 1423 -1703 1457 -1337
rect -1457 -2311 -1423 -1945
rect -1361 -2311 -1327 -1945
rect -1265 -2311 -1231 -1945
rect -1169 -2311 -1135 -1945
rect -1073 -2311 -1039 -1945
rect -977 -2311 -943 -1945
rect -881 -2311 -847 -1945
rect -785 -2311 -751 -1945
rect -689 -2311 -655 -1945
rect -593 -2311 -559 -1945
rect -497 -2311 -463 -1945
rect -401 -2311 -367 -1945
rect -305 -2311 -271 -1945
rect -209 -2311 -175 -1945
rect -113 -2311 -79 -1945
rect -17 -2311 17 -1945
rect 79 -2311 113 -1945
rect 175 -2311 209 -1945
rect 271 -2311 305 -1945
rect 367 -2311 401 -1945
rect 463 -2311 497 -1945
rect 559 -2311 593 -1945
rect 655 -2311 689 -1945
rect 751 -2311 785 -1945
rect 847 -2311 881 -1945
rect 943 -2311 977 -1945
rect 1039 -2311 1073 -1945
rect 1135 -2311 1169 -1945
rect 1231 -2311 1265 -1945
rect 1327 -2311 1361 -1945
rect 1423 -2311 1457 -1945
<< psubdiff >>
rect -1571 2463 -1475 2497
rect 1475 2463 1571 2497
rect -1571 2401 -1537 2463
rect 1537 2401 1571 2463
rect -1571 -2463 -1537 -2401
rect 1537 -2463 1571 -2401
rect -1571 -2497 -1475 -2463
rect 1475 -2497 1571 -2463
<< psubdiffcont >>
rect -1475 2463 1475 2497
rect -1571 -2401 -1537 2401
rect 1537 -2401 1571 2401
rect -1475 -2497 1475 -2463
<< poly >>
rect -1425 2395 -1359 2411
rect -1425 2361 -1409 2395
rect -1375 2361 -1359 2395
rect -1425 2345 -1359 2361
rect -1233 2395 -1167 2411
rect -1233 2361 -1217 2395
rect -1183 2361 -1167 2395
rect -1407 2323 -1377 2345
rect -1311 2323 -1281 2349
rect -1233 2345 -1167 2361
rect -1041 2395 -975 2411
rect -1041 2361 -1025 2395
rect -991 2361 -975 2395
rect -1215 2323 -1185 2345
rect -1119 2323 -1089 2349
rect -1041 2345 -975 2361
rect -849 2395 -783 2411
rect -849 2361 -833 2395
rect -799 2361 -783 2395
rect -1023 2323 -993 2345
rect -927 2323 -897 2349
rect -849 2345 -783 2361
rect -657 2395 -591 2411
rect -657 2361 -641 2395
rect -607 2361 -591 2395
rect -831 2323 -801 2345
rect -735 2323 -705 2349
rect -657 2345 -591 2361
rect -465 2395 -399 2411
rect -465 2361 -449 2395
rect -415 2361 -399 2395
rect -639 2323 -609 2345
rect -543 2323 -513 2349
rect -465 2345 -399 2361
rect -273 2395 -207 2411
rect -273 2361 -257 2395
rect -223 2361 -207 2395
rect -447 2323 -417 2345
rect -351 2323 -321 2349
rect -273 2345 -207 2361
rect -81 2395 -15 2411
rect -81 2361 -65 2395
rect -31 2361 -15 2395
rect -255 2323 -225 2345
rect -159 2323 -129 2349
rect -81 2345 -15 2361
rect 111 2395 177 2411
rect 111 2361 127 2395
rect 161 2361 177 2395
rect -63 2323 -33 2345
rect 33 2323 63 2349
rect 111 2345 177 2361
rect 303 2395 369 2411
rect 303 2361 319 2395
rect 353 2361 369 2395
rect 129 2323 159 2345
rect 225 2323 255 2349
rect 303 2345 369 2361
rect 495 2395 561 2411
rect 495 2361 511 2395
rect 545 2361 561 2395
rect 321 2323 351 2345
rect 417 2323 447 2349
rect 495 2345 561 2361
rect 687 2395 753 2411
rect 687 2361 703 2395
rect 737 2361 753 2395
rect 513 2323 543 2345
rect 609 2323 639 2349
rect 687 2345 753 2361
rect 879 2395 945 2411
rect 879 2361 895 2395
rect 929 2361 945 2395
rect 705 2323 735 2345
rect 801 2323 831 2349
rect 879 2345 945 2361
rect 1071 2395 1137 2411
rect 1071 2361 1087 2395
rect 1121 2361 1137 2395
rect 897 2323 927 2345
rect 993 2323 1023 2349
rect 1071 2345 1137 2361
rect 1263 2395 1329 2411
rect 1263 2361 1279 2395
rect 1313 2361 1329 2395
rect 1089 2323 1119 2345
rect 1185 2323 1215 2349
rect 1263 2345 1329 2361
rect 1281 2323 1311 2345
rect 1377 2323 1407 2349
rect -1407 1907 -1377 1933
rect -1311 1911 -1281 1933
rect -1329 1895 -1263 1911
rect -1215 1907 -1185 1933
rect -1119 1911 -1089 1933
rect -1329 1861 -1313 1895
rect -1279 1861 -1263 1895
rect -1329 1845 -1263 1861
rect -1137 1895 -1071 1911
rect -1023 1907 -993 1933
rect -927 1911 -897 1933
rect -1137 1861 -1121 1895
rect -1087 1861 -1071 1895
rect -1137 1845 -1071 1861
rect -945 1895 -879 1911
rect -831 1907 -801 1933
rect -735 1911 -705 1933
rect -945 1861 -929 1895
rect -895 1861 -879 1895
rect -945 1845 -879 1861
rect -753 1895 -687 1911
rect -639 1907 -609 1933
rect -543 1911 -513 1933
rect -753 1861 -737 1895
rect -703 1861 -687 1895
rect -753 1845 -687 1861
rect -561 1895 -495 1911
rect -447 1907 -417 1933
rect -351 1911 -321 1933
rect -561 1861 -545 1895
rect -511 1861 -495 1895
rect -561 1845 -495 1861
rect -369 1895 -303 1911
rect -255 1907 -225 1933
rect -159 1911 -129 1933
rect -369 1861 -353 1895
rect -319 1861 -303 1895
rect -369 1845 -303 1861
rect -177 1895 -111 1911
rect -63 1907 -33 1933
rect 33 1911 63 1933
rect -177 1861 -161 1895
rect -127 1861 -111 1895
rect -177 1845 -111 1861
rect 15 1895 81 1911
rect 129 1907 159 1933
rect 225 1911 255 1933
rect 15 1861 31 1895
rect 65 1861 81 1895
rect 15 1845 81 1861
rect 207 1895 273 1911
rect 321 1907 351 1933
rect 417 1911 447 1933
rect 207 1861 223 1895
rect 257 1861 273 1895
rect 207 1845 273 1861
rect 399 1895 465 1911
rect 513 1907 543 1933
rect 609 1911 639 1933
rect 399 1861 415 1895
rect 449 1861 465 1895
rect 399 1845 465 1861
rect 591 1895 657 1911
rect 705 1907 735 1933
rect 801 1911 831 1933
rect 591 1861 607 1895
rect 641 1861 657 1895
rect 591 1845 657 1861
rect 783 1895 849 1911
rect 897 1907 927 1933
rect 993 1911 1023 1933
rect 783 1861 799 1895
rect 833 1861 849 1895
rect 783 1845 849 1861
rect 975 1895 1041 1911
rect 1089 1907 1119 1933
rect 1185 1911 1215 1933
rect 975 1861 991 1895
rect 1025 1861 1041 1895
rect 975 1845 1041 1861
rect 1167 1895 1233 1911
rect 1281 1907 1311 1933
rect 1377 1911 1407 1933
rect 1167 1861 1183 1895
rect 1217 1861 1233 1895
rect 1167 1845 1233 1861
rect 1359 1895 1425 1911
rect 1359 1861 1375 1895
rect 1409 1861 1425 1895
rect 1359 1845 1425 1861
rect -1329 1787 -1263 1803
rect -1329 1753 -1313 1787
rect -1279 1753 -1263 1787
rect -1407 1715 -1377 1741
rect -1329 1737 -1263 1753
rect -1137 1787 -1071 1803
rect -1137 1753 -1121 1787
rect -1087 1753 -1071 1787
rect -1311 1715 -1281 1737
rect -1215 1715 -1185 1741
rect -1137 1737 -1071 1753
rect -945 1787 -879 1803
rect -945 1753 -929 1787
rect -895 1753 -879 1787
rect -1119 1715 -1089 1737
rect -1023 1715 -993 1741
rect -945 1737 -879 1753
rect -753 1787 -687 1803
rect -753 1753 -737 1787
rect -703 1753 -687 1787
rect -927 1715 -897 1737
rect -831 1715 -801 1741
rect -753 1737 -687 1753
rect -561 1787 -495 1803
rect -561 1753 -545 1787
rect -511 1753 -495 1787
rect -735 1715 -705 1737
rect -639 1715 -609 1741
rect -561 1737 -495 1753
rect -369 1787 -303 1803
rect -369 1753 -353 1787
rect -319 1753 -303 1787
rect -543 1715 -513 1737
rect -447 1715 -417 1741
rect -369 1737 -303 1753
rect -177 1787 -111 1803
rect -177 1753 -161 1787
rect -127 1753 -111 1787
rect -351 1715 -321 1737
rect -255 1715 -225 1741
rect -177 1737 -111 1753
rect 15 1787 81 1803
rect 15 1753 31 1787
rect 65 1753 81 1787
rect -159 1715 -129 1737
rect -63 1715 -33 1741
rect 15 1737 81 1753
rect 207 1787 273 1803
rect 207 1753 223 1787
rect 257 1753 273 1787
rect 33 1715 63 1737
rect 129 1715 159 1741
rect 207 1737 273 1753
rect 399 1787 465 1803
rect 399 1753 415 1787
rect 449 1753 465 1787
rect 225 1715 255 1737
rect 321 1715 351 1741
rect 399 1737 465 1753
rect 591 1787 657 1803
rect 591 1753 607 1787
rect 641 1753 657 1787
rect 417 1715 447 1737
rect 513 1715 543 1741
rect 591 1737 657 1753
rect 783 1787 849 1803
rect 783 1753 799 1787
rect 833 1753 849 1787
rect 609 1715 639 1737
rect 705 1715 735 1741
rect 783 1737 849 1753
rect 975 1787 1041 1803
rect 975 1753 991 1787
rect 1025 1753 1041 1787
rect 801 1715 831 1737
rect 897 1715 927 1741
rect 975 1737 1041 1753
rect 1167 1787 1233 1803
rect 1167 1753 1183 1787
rect 1217 1753 1233 1787
rect 993 1715 1023 1737
rect 1089 1715 1119 1741
rect 1167 1737 1233 1753
rect 1359 1787 1425 1803
rect 1359 1753 1375 1787
rect 1409 1753 1425 1787
rect 1185 1715 1215 1737
rect 1281 1715 1311 1741
rect 1359 1737 1425 1753
rect 1377 1715 1407 1737
rect -1407 1303 -1377 1325
rect -1425 1287 -1359 1303
rect -1311 1299 -1281 1325
rect -1215 1303 -1185 1325
rect -1425 1253 -1409 1287
rect -1375 1253 -1359 1287
rect -1425 1237 -1359 1253
rect -1233 1287 -1167 1303
rect -1119 1299 -1089 1325
rect -1023 1303 -993 1325
rect -1233 1253 -1217 1287
rect -1183 1253 -1167 1287
rect -1233 1237 -1167 1253
rect -1041 1287 -975 1303
rect -927 1299 -897 1325
rect -831 1303 -801 1325
rect -1041 1253 -1025 1287
rect -991 1253 -975 1287
rect -1041 1237 -975 1253
rect -849 1287 -783 1303
rect -735 1299 -705 1325
rect -639 1303 -609 1325
rect -849 1253 -833 1287
rect -799 1253 -783 1287
rect -849 1237 -783 1253
rect -657 1287 -591 1303
rect -543 1299 -513 1325
rect -447 1303 -417 1325
rect -657 1253 -641 1287
rect -607 1253 -591 1287
rect -657 1237 -591 1253
rect -465 1287 -399 1303
rect -351 1299 -321 1325
rect -255 1303 -225 1325
rect -465 1253 -449 1287
rect -415 1253 -399 1287
rect -465 1237 -399 1253
rect -273 1287 -207 1303
rect -159 1299 -129 1325
rect -63 1303 -33 1325
rect -273 1253 -257 1287
rect -223 1253 -207 1287
rect -273 1237 -207 1253
rect -81 1287 -15 1303
rect 33 1299 63 1325
rect 129 1303 159 1325
rect -81 1253 -65 1287
rect -31 1253 -15 1287
rect -81 1237 -15 1253
rect 111 1287 177 1303
rect 225 1299 255 1325
rect 321 1303 351 1325
rect 111 1253 127 1287
rect 161 1253 177 1287
rect 111 1237 177 1253
rect 303 1287 369 1303
rect 417 1299 447 1325
rect 513 1303 543 1325
rect 303 1253 319 1287
rect 353 1253 369 1287
rect 303 1237 369 1253
rect 495 1287 561 1303
rect 609 1299 639 1325
rect 705 1303 735 1325
rect 495 1253 511 1287
rect 545 1253 561 1287
rect 495 1237 561 1253
rect 687 1287 753 1303
rect 801 1299 831 1325
rect 897 1303 927 1325
rect 687 1253 703 1287
rect 737 1253 753 1287
rect 687 1237 753 1253
rect 879 1287 945 1303
rect 993 1299 1023 1325
rect 1089 1303 1119 1325
rect 879 1253 895 1287
rect 929 1253 945 1287
rect 879 1237 945 1253
rect 1071 1287 1137 1303
rect 1185 1299 1215 1325
rect 1281 1303 1311 1325
rect 1071 1253 1087 1287
rect 1121 1253 1137 1287
rect 1071 1237 1137 1253
rect 1263 1287 1329 1303
rect 1377 1299 1407 1325
rect 1263 1253 1279 1287
rect 1313 1253 1329 1287
rect 1263 1237 1329 1253
rect -1425 1179 -1359 1195
rect -1425 1145 -1409 1179
rect -1375 1145 -1359 1179
rect -1425 1129 -1359 1145
rect -1233 1179 -1167 1195
rect -1233 1145 -1217 1179
rect -1183 1145 -1167 1179
rect -1407 1107 -1377 1129
rect -1311 1107 -1281 1133
rect -1233 1129 -1167 1145
rect -1041 1179 -975 1195
rect -1041 1145 -1025 1179
rect -991 1145 -975 1179
rect -1215 1107 -1185 1129
rect -1119 1107 -1089 1133
rect -1041 1129 -975 1145
rect -849 1179 -783 1195
rect -849 1145 -833 1179
rect -799 1145 -783 1179
rect -1023 1107 -993 1129
rect -927 1107 -897 1133
rect -849 1129 -783 1145
rect -657 1179 -591 1195
rect -657 1145 -641 1179
rect -607 1145 -591 1179
rect -831 1107 -801 1129
rect -735 1107 -705 1133
rect -657 1129 -591 1145
rect -465 1179 -399 1195
rect -465 1145 -449 1179
rect -415 1145 -399 1179
rect -639 1107 -609 1129
rect -543 1107 -513 1133
rect -465 1129 -399 1145
rect -273 1179 -207 1195
rect -273 1145 -257 1179
rect -223 1145 -207 1179
rect -447 1107 -417 1129
rect -351 1107 -321 1133
rect -273 1129 -207 1145
rect -81 1179 -15 1195
rect -81 1145 -65 1179
rect -31 1145 -15 1179
rect -255 1107 -225 1129
rect -159 1107 -129 1133
rect -81 1129 -15 1145
rect 111 1179 177 1195
rect 111 1145 127 1179
rect 161 1145 177 1179
rect -63 1107 -33 1129
rect 33 1107 63 1133
rect 111 1129 177 1145
rect 303 1179 369 1195
rect 303 1145 319 1179
rect 353 1145 369 1179
rect 129 1107 159 1129
rect 225 1107 255 1133
rect 303 1129 369 1145
rect 495 1179 561 1195
rect 495 1145 511 1179
rect 545 1145 561 1179
rect 321 1107 351 1129
rect 417 1107 447 1133
rect 495 1129 561 1145
rect 687 1179 753 1195
rect 687 1145 703 1179
rect 737 1145 753 1179
rect 513 1107 543 1129
rect 609 1107 639 1133
rect 687 1129 753 1145
rect 879 1179 945 1195
rect 879 1145 895 1179
rect 929 1145 945 1179
rect 705 1107 735 1129
rect 801 1107 831 1133
rect 879 1129 945 1145
rect 1071 1179 1137 1195
rect 1071 1145 1087 1179
rect 1121 1145 1137 1179
rect 897 1107 927 1129
rect 993 1107 1023 1133
rect 1071 1129 1137 1145
rect 1263 1179 1329 1195
rect 1263 1145 1279 1179
rect 1313 1145 1329 1179
rect 1089 1107 1119 1129
rect 1185 1107 1215 1133
rect 1263 1129 1329 1145
rect 1281 1107 1311 1129
rect 1377 1107 1407 1133
rect -1407 691 -1377 717
rect -1311 695 -1281 717
rect -1329 679 -1263 695
rect -1215 691 -1185 717
rect -1119 695 -1089 717
rect -1329 645 -1313 679
rect -1279 645 -1263 679
rect -1329 629 -1263 645
rect -1137 679 -1071 695
rect -1023 691 -993 717
rect -927 695 -897 717
rect -1137 645 -1121 679
rect -1087 645 -1071 679
rect -1137 629 -1071 645
rect -945 679 -879 695
rect -831 691 -801 717
rect -735 695 -705 717
rect -945 645 -929 679
rect -895 645 -879 679
rect -945 629 -879 645
rect -753 679 -687 695
rect -639 691 -609 717
rect -543 695 -513 717
rect -753 645 -737 679
rect -703 645 -687 679
rect -753 629 -687 645
rect -561 679 -495 695
rect -447 691 -417 717
rect -351 695 -321 717
rect -561 645 -545 679
rect -511 645 -495 679
rect -561 629 -495 645
rect -369 679 -303 695
rect -255 691 -225 717
rect -159 695 -129 717
rect -369 645 -353 679
rect -319 645 -303 679
rect -369 629 -303 645
rect -177 679 -111 695
rect -63 691 -33 717
rect 33 695 63 717
rect -177 645 -161 679
rect -127 645 -111 679
rect -177 629 -111 645
rect 15 679 81 695
rect 129 691 159 717
rect 225 695 255 717
rect 15 645 31 679
rect 65 645 81 679
rect 15 629 81 645
rect 207 679 273 695
rect 321 691 351 717
rect 417 695 447 717
rect 207 645 223 679
rect 257 645 273 679
rect 207 629 273 645
rect 399 679 465 695
rect 513 691 543 717
rect 609 695 639 717
rect 399 645 415 679
rect 449 645 465 679
rect 399 629 465 645
rect 591 679 657 695
rect 705 691 735 717
rect 801 695 831 717
rect 591 645 607 679
rect 641 645 657 679
rect 591 629 657 645
rect 783 679 849 695
rect 897 691 927 717
rect 993 695 1023 717
rect 783 645 799 679
rect 833 645 849 679
rect 783 629 849 645
rect 975 679 1041 695
rect 1089 691 1119 717
rect 1185 695 1215 717
rect 975 645 991 679
rect 1025 645 1041 679
rect 975 629 1041 645
rect 1167 679 1233 695
rect 1281 691 1311 717
rect 1377 695 1407 717
rect 1167 645 1183 679
rect 1217 645 1233 679
rect 1167 629 1233 645
rect 1359 679 1425 695
rect 1359 645 1375 679
rect 1409 645 1425 679
rect 1359 629 1425 645
rect -1329 571 -1263 587
rect -1329 537 -1313 571
rect -1279 537 -1263 571
rect -1407 499 -1377 525
rect -1329 521 -1263 537
rect -1137 571 -1071 587
rect -1137 537 -1121 571
rect -1087 537 -1071 571
rect -1311 499 -1281 521
rect -1215 499 -1185 525
rect -1137 521 -1071 537
rect -945 571 -879 587
rect -945 537 -929 571
rect -895 537 -879 571
rect -1119 499 -1089 521
rect -1023 499 -993 525
rect -945 521 -879 537
rect -753 571 -687 587
rect -753 537 -737 571
rect -703 537 -687 571
rect -927 499 -897 521
rect -831 499 -801 525
rect -753 521 -687 537
rect -561 571 -495 587
rect -561 537 -545 571
rect -511 537 -495 571
rect -735 499 -705 521
rect -639 499 -609 525
rect -561 521 -495 537
rect -369 571 -303 587
rect -369 537 -353 571
rect -319 537 -303 571
rect -543 499 -513 521
rect -447 499 -417 525
rect -369 521 -303 537
rect -177 571 -111 587
rect -177 537 -161 571
rect -127 537 -111 571
rect -351 499 -321 521
rect -255 499 -225 525
rect -177 521 -111 537
rect 15 571 81 587
rect 15 537 31 571
rect 65 537 81 571
rect -159 499 -129 521
rect -63 499 -33 525
rect 15 521 81 537
rect 207 571 273 587
rect 207 537 223 571
rect 257 537 273 571
rect 33 499 63 521
rect 129 499 159 525
rect 207 521 273 537
rect 399 571 465 587
rect 399 537 415 571
rect 449 537 465 571
rect 225 499 255 521
rect 321 499 351 525
rect 399 521 465 537
rect 591 571 657 587
rect 591 537 607 571
rect 641 537 657 571
rect 417 499 447 521
rect 513 499 543 525
rect 591 521 657 537
rect 783 571 849 587
rect 783 537 799 571
rect 833 537 849 571
rect 609 499 639 521
rect 705 499 735 525
rect 783 521 849 537
rect 975 571 1041 587
rect 975 537 991 571
rect 1025 537 1041 571
rect 801 499 831 521
rect 897 499 927 525
rect 975 521 1041 537
rect 1167 571 1233 587
rect 1167 537 1183 571
rect 1217 537 1233 571
rect 993 499 1023 521
rect 1089 499 1119 525
rect 1167 521 1233 537
rect 1359 571 1425 587
rect 1359 537 1375 571
rect 1409 537 1425 571
rect 1185 499 1215 521
rect 1281 499 1311 525
rect 1359 521 1425 537
rect 1377 499 1407 521
rect -1407 87 -1377 109
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect -1407 -525 -1377 -499
rect -1311 -521 -1281 -499
rect -1329 -537 -1263 -521
rect -1215 -525 -1185 -499
rect -1119 -521 -1089 -499
rect -1329 -571 -1313 -537
rect -1279 -571 -1263 -537
rect -1329 -587 -1263 -571
rect -1137 -537 -1071 -521
rect -1023 -525 -993 -499
rect -927 -521 -897 -499
rect -1137 -571 -1121 -537
rect -1087 -571 -1071 -537
rect -1137 -587 -1071 -571
rect -945 -537 -879 -521
rect -831 -525 -801 -499
rect -735 -521 -705 -499
rect -945 -571 -929 -537
rect -895 -571 -879 -537
rect -945 -587 -879 -571
rect -753 -537 -687 -521
rect -639 -525 -609 -499
rect -543 -521 -513 -499
rect -753 -571 -737 -537
rect -703 -571 -687 -537
rect -753 -587 -687 -571
rect -561 -537 -495 -521
rect -447 -525 -417 -499
rect -351 -521 -321 -499
rect -561 -571 -545 -537
rect -511 -571 -495 -537
rect -561 -587 -495 -571
rect -369 -537 -303 -521
rect -255 -525 -225 -499
rect -159 -521 -129 -499
rect -369 -571 -353 -537
rect -319 -571 -303 -537
rect -369 -587 -303 -571
rect -177 -537 -111 -521
rect -63 -525 -33 -499
rect 33 -521 63 -499
rect -177 -571 -161 -537
rect -127 -571 -111 -537
rect -177 -587 -111 -571
rect 15 -537 81 -521
rect 129 -525 159 -499
rect 225 -521 255 -499
rect 15 -571 31 -537
rect 65 -571 81 -537
rect 15 -587 81 -571
rect 207 -537 273 -521
rect 321 -525 351 -499
rect 417 -521 447 -499
rect 207 -571 223 -537
rect 257 -571 273 -537
rect 207 -587 273 -571
rect 399 -537 465 -521
rect 513 -525 543 -499
rect 609 -521 639 -499
rect 399 -571 415 -537
rect 449 -571 465 -537
rect 399 -587 465 -571
rect 591 -537 657 -521
rect 705 -525 735 -499
rect 801 -521 831 -499
rect 591 -571 607 -537
rect 641 -571 657 -537
rect 591 -587 657 -571
rect 783 -537 849 -521
rect 897 -525 927 -499
rect 993 -521 1023 -499
rect 783 -571 799 -537
rect 833 -571 849 -537
rect 783 -587 849 -571
rect 975 -537 1041 -521
rect 1089 -525 1119 -499
rect 1185 -521 1215 -499
rect 975 -571 991 -537
rect 1025 -571 1041 -537
rect 975 -587 1041 -571
rect 1167 -537 1233 -521
rect 1281 -525 1311 -499
rect 1377 -521 1407 -499
rect 1167 -571 1183 -537
rect 1217 -571 1233 -537
rect 1167 -587 1233 -571
rect 1359 -537 1425 -521
rect 1359 -571 1375 -537
rect 1409 -571 1425 -537
rect 1359 -587 1425 -571
rect -1329 -645 -1263 -629
rect -1329 -679 -1313 -645
rect -1279 -679 -1263 -645
rect -1407 -717 -1377 -691
rect -1329 -695 -1263 -679
rect -1137 -645 -1071 -629
rect -1137 -679 -1121 -645
rect -1087 -679 -1071 -645
rect -1311 -717 -1281 -695
rect -1215 -717 -1185 -691
rect -1137 -695 -1071 -679
rect -945 -645 -879 -629
rect -945 -679 -929 -645
rect -895 -679 -879 -645
rect -1119 -717 -1089 -695
rect -1023 -717 -993 -691
rect -945 -695 -879 -679
rect -753 -645 -687 -629
rect -753 -679 -737 -645
rect -703 -679 -687 -645
rect -927 -717 -897 -695
rect -831 -717 -801 -691
rect -753 -695 -687 -679
rect -561 -645 -495 -629
rect -561 -679 -545 -645
rect -511 -679 -495 -645
rect -735 -717 -705 -695
rect -639 -717 -609 -691
rect -561 -695 -495 -679
rect -369 -645 -303 -629
rect -369 -679 -353 -645
rect -319 -679 -303 -645
rect -543 -717 -513 -695
rect -447 -717 -417 -691
rect -369 -695 -303 -679
rect -177 -645 -111 -629
rect -177 -679 -161 -645
rect -127 -679 -111 -645
rect -351 -717 -321 -695
rect -255 -717 -225 -691
rect -177 -695 -111 -679
rect 15 -645 81 -629
rect 15 -679 31 -645
rect 65 -679 81 -645
rect -159 -717 -129 -695
rect -63 -717 -33 -691
rect 15 -695 81 -679
rect 207 -645 273 -629
rect 207 -679 223 -645
rect 257 -679 273 -645
rect 33 -717 63 -695
rect 129 -717 159 -691
rect 207 -695 273 -679
rect 399 -645 465 -629
rect 399 -679 415 -645
rect 449 -679 465 -645
rect 225 -717 255 -695
rect 321 -717 351 -691
rect 399 -695 465 -679
rect 591 -645 657 -629
rect 591 -679 607 -645
rect 641 -679 657 -645
rect 417 -717 447 -695
rect 513 -717 543 -691
rect 591 -695 657 -679
rect 783 -645 849 -629
rect 783 -679 799 -645
rect 833 -679 849 -645
rect 609 -717 639 -695
rect 705 -717 735 -691
rect 783 -695 849 -679
rect 975 -645 1041 -629
rect 975 -679 991 -645
rect 1025 -679 1041 -645
rect 801 -717 831 -695
rect 897 -717 927 -691
rect 975 -695 1041 -679
rect 1167 -645 1233 -629
rect 1167 -679 1183 -645
rect 1217 -679 1233 -645
rect 993 -717 1023 -695
rect 1089 -717 1119 -691
rect 1167 -695 1233 -679
rect 1359 -645 1425 -629
rect 1359 -679 1375 -645
rect 1409 -679 1425 -645
rect 1185 -717 1215 -695
rect 1281 -717 1311 -691
rect 1359 -695 1425 -679
rect 1377 -717 1407 -695
rect -1407 -1129 -1377 -1107
rect -1425 -1145 -1359 -1129
rect -1311 -1133 -1281 -1107
rect -1215 -1129 -1185 -1107
rect -1425 -1179 -1409 -1145
rect -1375 -1179 -1359 -1145
rect -1425 -1195 -1359 -1179
rect -1233 -1145 -1167 -1129
rect -1119 -1133 -1089 -1107
rect -1023 -1129 -993 -1107
rect -1233 -1179 -1217 -1145
rect -1183 -1179 -1167 -1145
rect -1233 -1195 -1167 -1179
rect -1041 -1145 -975 -1129
rect -927 -1133 -897 -1107
rect -831 -1129 -801 -1107
rect -1041 -1179 -1025 -1145
rect -991 -1179 -975 -1145
rect -1041 -1195 -975 -1179
rect -849 -1145 -783 -1129
rect -735 -1133 -705 -1107
rect -639 -1129 -609 -1107
rect -849 -1179 -833 -1145
rect -799 -1179 -783 -1145
rect -849 -1195 -783 -1179
rect -657 -1145 -591 -1129
rect -543 -1133 -513 -1107
rect -447 -1129 -417 -1107
rect -657 -1179 -641 -1145
rect -607 -1179 -591 -1145
rect -657 -1195 -591 -1179
rect -465 -1145 -399 -1129
rect -351 -1133 -321 -1107
rect -255 -1129 -225 -1107
rect -465 -1179 -449 -1145
rect -415 -1179 -399 -1145
rect -465 -1195 -399 -1179
rect -273 -1145 -207 -1129
rect -159 -1133 -129 -1107
rect -63 -1129 -33 -1107
rect -273 -1179 -257 -1145
rect -223 -1179 -207 -1145
rect -273 -1195 -207 -1179
rect -81 -1145 -15 -1129
rect 33 -1133 63 -1107
rect 129 -1129 159 -1107
rect -81 -1179 -65 -1145
rect -31 -1179 -15 -1145
rect -81 -1195 -15 -1179
rect 111 -1145 177 -1129
rect 225 -1133 255 -1107
rect 321 -1129 351 -1107
rect 111 -1179 127 -1145
rect 161 -1179 177 -1145
rect 111 -1195 177 -1179
rect 303 -1145 369 -1129
rect 417 -1133 447 -1107
rect 513 -1129 543 -1107
rect 303 -1179 319 -1145
rect 353 -1179 369 -1145
rect 303 -1195 369 -1179
rect 495 -1145 561 -1129
rect 609 -1133 639 -1107
rect 705 -1129 735 -1107
rect 495 -1179 511 -1145
rect 545 -1179 561 -1145
rect 495 -1195 561 -1179
rect 687 -1145 753 -1129
rect 801 -1133 831 -1107
rect 897 -1129 927 -1107
rect 687 -1179 703 -1145
rect 737 -1179 753 -1145
rect 687 -1195 753 -1179
rect 879 -1145 945 -1129
rect 993 -1133 1023 -1107
rect 1089 -1129 1119 -1107
rect 879 -1179 895 -1145
rect 929 -1179 945 -1145
rect 879 -1195 945 -1179
rect 1071 -1145 1137 -1129
rect 1185 -1133 1215 -1107
rect 1281 -1129 1311 -1107
rect 1071 -1179 1087 -1145
rect 1121 -1179 1137 -1145
rect 1071 -1195 1137 -1179
rect 1263 -1145 1329 -1129
rect 1377 -1133 1407 -1107
rect 1263 -1179 1279 -1145
rect 1313 -1179 1329 -1145
rect 1263 -1195 1329 -1179
rect -1425 -1253 -1359 -1237
rect -1425 -1287 -1409 -1253
rect -1375 -1287 -1359 -1253
rect -1425 -1303 -1359 -1287
rect -1233 -1253 -1167 -1237
rect -1233 -1287 -1217 -1253
rect -1183 -1287 -1167 -1253
rect -1407 -1325 -1377 -1303
rect -1311 -1325 -1281 -1299
rect -1233 -1303 -1167 -1287
rect -1041 -1253 -975 -1237
rect -1041 -1287 -1025 -1253
rect -991 -1287 -975 -1253
rect -1215 -1325 -1185 -1303
rect -1119 -1325 -1089 -1299
rect -1041 -1303 -975 -1287
rect -849 -1253 -783 -1237
rect -849 -1287 -833 -1253
rect -799 -1287 -783 -1253
rect -1023 -1325 -993 -1303
rect -927 -1325 -897 -1299
rect -849 -1303 -783 -1287
rect -657 -1253 -591 -1237
rect -657 -1287 -641 -1253
rect -607 -1287 -591 -1253
rect -831 -1325 -801 -1303
rect -735 -1325 -705 -1299
rect -657 -1303 -591 -1287
rect -465 -1253 -399 -1237
rect -465 -1287 -449 -1253
rect -415 -1287 -399 -1253
rect -639 -1325 -609 -1303
rect -543 -1325 -513 -1299
rect -465 -1303 -399 -1287
rect -273 -1253 -207 -1237
rect -273 -1287 -257 -1253
rect -223 -1287 -207 -1253
rect -447 -1325 -417 -1303
rect -351 -1325 -321 -1299
rect -273 -1303 -207 -1287
rect -81 -1253 -15 -1237
rect -81 -1287 -65 -1253
rect -31 -1287 -15 -1253
rect -255 -1325 -225 -1303
rect -159 -1325 -129 -1299
rect -81 -1303 -15 -1287
rect 111 -1253 177 -1237
rect 111 -1287 127 -1253
rect 161 -1287 177 -1253
rect -63 -1325 -33 -1303
rect 33 -1325 63 -1299
rect 111 -1303 177 -1287
rect 303 -1253 369 -1237
rect 303 -1287 319 -1253
rect 353 -1287 369 -1253
rect 129 -1325 159 -1303
rect 225 -1325 255 -1299
rect 303 -1303 369 -1287
rect 495 -1253 561 -1237
rect 495 -1287 511 -1253
rect 545 -1287 561 -1253
rect 321 -1325 351 -1303
rect 417 -1325 447 -1299
rect 495 -1303 561 -1287
rect 687 -1253 753 -1237
rect 687 -1287 703 -1253
rect 737 -1287 753 -1253
rect 513 -1325 543 -1303
rect 609 -1325 639 -1299
rect 687 -1303 753 -1287
rect 879 -1253 945 -1237
rect 879 -1287 895 -1253
rect 929 -1287 945 -1253
rect 705 -1325 735 -1303
rect 801 -1325 831 -1299
rect 879 -1303 945 -1287
rect 1071 -1253 1137 -1237
rect 1071 -1287 1087 -1253
rect 1121 -1287 1137 -1253
rect 897 -1325 927 -1303
rect 993 -1325 1023 -1299
rect 1071 -1303 1137 -1287
rect 1263 -1253 1329 -1237
rect 1263 -1287 1279 -1253
rect 1313 -1287 1329 -1253
rect 1089 -1325 1119 -1303
rect 1185 -1325 1215 -1299
rect 1263 -1303 1329 -1287
rect 1281 -1325 1311 -1303
rect 1377 -1325 1407 -1299
rect -1407 -1741 -1377 -1715
rect -1311 -1737 -1281 -1715
rect -1329 -1753 -1263 -1737
rect -1215 -1741 -1185 -1715
rect -1119 -1737 -1089 -1715
rect -1329 -1787 -1313 -1753
rect -1279 -1787 -1263 -1753
rect -1329 -1803 -1263 -1787
rect -1137 -1753 -1071 -1737
rect -1023 -1741 -993 -1715
rect -927 -1737 -897 -1715
rect -1137 -1787 -1121 -1753
rect -1087 -1787 -1071 -1753
rect -1137 -1803 -1071 -1787
rect -945 -1753 -879 -1737
rect -831 -1741 -801 -1715
rect -735 -1737 -705 -1715
rect -945 -1787 -929 -1753
rect -895 -1787 -879 -1753
rect -945 -1803 -879 -1787
rect -753 -1753 -687 -1737
rect -639 -1741 -609 -1715
rect -543 -1737 -513 -1715
rect -753 -1787 -737 -1753
rect -703 -1787 -687 -1753
rect -753 -1803 -687 -1787
rect -561 -1753 -495 -1737
rect -447 -1741 -417 -1715
rect -351 -1737 -321 -1715
rect -561 -1787 -545 -1753
rect -511 -1787 -495 -1753
rect -561 -1803 -495 -1787
rect -369 -1753 -303 -1737
rect -255 -1741 -225 -1715
rect -159 -1737 -129 -1715
rect -369 -1787 -353 -1753
rect -319 -1787 -303 -1753
rect -369 -1803 -303 -1787
rect -177 -1753 -111 -1737
rect -63 -1741 -33 -1715
rect 33 -1737 63 -1715
rect -177 -1787 -161 -1753
rect -127 -1787 -111 -1753
rect -177 -1803 -111 -1787
rect 15 -1753 81 -1737
rect 129 -1741 159 -1715
rect 225 -1737 255 -1715
rect 15 -1787 31 -1753
rect 65 -1787 81 -1753
rect 15 -1803 81 -1787
rect 207 -1753 273 -1737
rect 321 -1741 351 -1715
rect 417 -1737 447 -1715
rect 207 -1787 223 -1753
rect 257 -1787 273 -1753
rect 207 -1803 273 -1787
rect 399 -1753 465 -1737
rect 513 -1741 543 -1715
rect 609 -1737 639 -1715
rect 399 -1787 415 -1753
rect 449 -1787 465 -1753
rect 399 -1803 465 -1787
rect 591 -1753 657 -1737
rect 705 -1741 735 -1715
rect 801 -1737 831 -1715
rect 591 -1787 607 -1753
rect 641 -1787 657 -1753
rect 591 -1803 657 -1787
rect 783 -1753 849 -1737
rect 897 -1741 927 -1715
rect 993 -1737 1023 -1715
rect 783 -1787 799 -1753
rect 833 -1787 849 -1753
rect 783 -1803 849 -1787
rect 975 -1753 1041 -1737
rect 1089 -1741 1119 -1715
rect 1185 -1737 1215 -1715
rect 975 -1787 991 -1753
rect 1025 -1787 1041 -1753
rect 975 -1803 1041 -1787
rect 1167 -1753 1233 -1737
rect 1281 -1741 1311 -1715
rect 1377 -1737 1407 -1715
rect 1167 -1787 1183 -1753
rect 1217 -1787 1233 -1753
rect 1167 -1803 1233 -1787
rect 1359 -1753 1425 -1737
rect 1359 -1787 1375 -1753
rect 1409 -1787 1425 -1753
rect 1359 -1803 1425 -1787
rect -1329 -1861 -1263 -1845
rect -1329 -1895 -1313 -1861
rect -1279 -1895 -1263 -1861
rect -1407 -1933 -1377 -1907
rect -1329 -1911 -1263 -1895
rect -1137 -1861 -1071 -1845
rect -1137 -1895 -1121 -1861
rect -1087 -1895 -1071 -1861
rect -1311 -1933 -1281 -1911
rect -1215 -1933 -1185 -1907
rect -1137 -1911 -1071 -1895
rect -945 -1861 -879 -1845
rect -945 -1895 -929 -1861
rect -895 -1895 -879 -1861
rect -1119 -1933 -1089 -1911
rect -1023 -1933 -993 -1907
rect -945 -1911 -879 -1895
rect -753 -1861 -687 -1845
rect -753 -1895 -737 -1861
rect -703 -1895 -687 -1861
rect -927 -1933 -897 -1911
rect -831 -1933 -801 -1907
rect -753 -1911 -687 -1895
rect -561 -1861 -495 -1845
rect -561 -1895 -545 -1861
rect -511 -1895 -495 -1861
rect -735 -1933 -705 -1911
rect -639 -1933 -609 -1907
rect -561 -1911 -495 -1895
rect -369 -1861 -303 -1845
rect -369 -1895 -353 -1861
rect -319 -1895 -303 -1861
rect -543 -1933 -513 -1911
rect -447 -1933 -417 -1907
rect -369 -1911 -303 -1895
rect -177 -1861 -111 -1845
rect -177 -1895 -161 -1861
rect -127 -1895 -111 -1861
rect -351 -1933 -321 -1911
rect -255 -1933 -225 -1907
rect -177 -1911 -111 -1895
rect 15 -1861 81 -1845
rect 15 -1895 31 -1861
rect 65 -1895 81 -1861
rect -159 -1933 -129 -1911
rect -63 -1933 -33 -1907
rect 15 -1911 81 -1895
rect 207 -1861 273 -1845
rect 207 -1895 223 -1861
rect 257 -1895 273 -1861
rect 33 -1933 63 -1911
rect 129 -1933 159 -1907
rect 207 -1911 273 -1895
rect 399 -1861 465 -1845
rect 399 -1895 415 -1861
rect 449 -1895 465 -1861
rect 225 -1933 255 -1911
rect 321 -1933 351 -1907
rect 399 -1911 465 -1895
rect 591 -1861 657 -1845
rect 591 -1895 607 -1861
rect 641 -1895 657 -1861
rect 417 -1933 447 -1911
rect 513 -1933 543 -1907
rect 591 -1911 657 -1895
rect 783 -1861 849 -1845
rect 783 -1895 799 -1861
rect 833 -1895 849 -1861
rect 609 -1933 639 -1911
rect 705 -1933 735 -1907
rect 783 -1911 849 -1895
rect 975 -1861 1041 -1845
rect 975 -1895 991 -1861
rect 1025 -1895 1041 -1861
rect 801 -1933 831 -1911
rect 897 -1933 927 -1907
rect 975 -1911 1041 -1895
rect 1167 -1861 1233 -1845
rect 1167 -1895 1183 -1861
rect 1217 -1895 1233 -1861
rect 993 -1933 1023 -1911
rect 1089 -1933 1119 -1907
rect 1167 -1911 1233 -1895
rect 1359 -1861 1425 -1845
rect 1359 -1895 1375 -1861
rect 1409 -1895 1425 -1861
rect 1185 -1933 1215 -1911
rect 1281 -1933 1311 -1907
rect 1359 -1911 1425 -1895
rect 1377 -1933 1407 -1911
rect -1407 -2345 -1377 -2323
rect -1425 -2361 -1359 -2345
rect -1311 -2349 -1281 -2323
rect -1215 -2345 -1185 -2323
rect -1425 -2395 -1409 -2361
rect -1375 -2395 -1359 -2361
rect -1425 -2411 -1359 -2395
rect -1233 -2361 -1167 -2345
rect -1119 -2349 -1089 -2323
rect -1023 -2345 -993 -2323
rect -1233 -2395 -1217 -2361
rect -1183 -2395 -1167 -2361
rect -1233 -2411 -1167 -2395
rect -1041 -2361 -975 -2345
rect -927 -2349 -897 -2323
rect -831 -2345 -801 -2323
rect -1041 -2395 -1025 -2361
rect -991 -2395 -975 -2361
rect -1041 -2411 -975 -2395
rect -849 -2361 -783 -2345
rect -735 -2349 -705 -2323
rect -639 -2345 -609 -2323
rect -849 -2395 -833 -2361
rect -799 -2395 -783 -2361
rect -849 -2411 -783 -2395
rect -657 -2361 -591 -2345
rect -543 -2349 -513 -2323
rect -447 -2345 -417 -2323
rect -657 -2395 -641 -2361
rect -607 -2395 -591 -2361
rect -657 -2411 -591 -2395
rect -465 -2361 -399 -2345
rect -351 -2349 -321 -2323
rect -255 -2345 -225 -2323
rect -465 -2395 -449 -2361
rect -415 -2395 -399 -2361
rect -465 -2411 -399 -2395
rect -273 -2361 -207 -2345
rect -159 -2349 -129 -2323
rect -63 -2345 -33 -2323
rect -273 -2395 -257 -2361
rect -223 -2395 -207 -2361
rect -273 -2411 -207 -2395
rect -81 -2361 -15 -2345
rect 33 -2349 63 -2323
rect 129 -2345 159 -2323
rect -81 -2395 -65 -2361
rect -31 -2395 -15 -2361
rect -81 -2411 -15 -2395
rect 111 -2361 177 -2345
rect 225 -2349 255 -2323
rect 321 -2345 351 -2323
rect 111 -2395 127 -2361
rect 161 -2395 177 -2361
rect 111 -2411 177 -2395
rect 303 -2361 369 -2345
rect 417 -2349 447 -2323
rect 513 -2345 543 -2323
rect 303 -2395 319 -2361
rect 353 -2395 369 -2361
rect 303 -2411 369 -2395
rect 495 -2361 561 -2345
rect 609 -2349 639 -2323
rect 705 -2345 735 -2323
rect 495 -2395 511 -2361
rect 545 -2395 561 -2361
rect 495 -2411 561 -2395
rect 687 -2361 753 -2345
rect 801 -2349 831 -2323
rect 897 -2345 927 -2323
rect 687 -2395 703 -2361
rect 737 -2395 753 -2361
rect 687 -2411 753 -2395
rect 879 -2361 945 -2345
rect 993 -2349 1023 -2323
rect 1089 -2345 1119 -2323
rect 879 -2395 895 -2361
rect 929 -2395 945 -2361
rect 879 -2411 945 -2395
rect 1071 -2361 1137 -2345
rect 1185 -2349 1215 -2323
rect 1281 -2345 1311 -2323
rect 1071 -2395 1087 -2361
rect 1121 -2395 1137 -2361
rect 1071 -2411 1137 -2395
rect 1263 -2361 1329 -2345
rect 1377 -2349 1407 -2323
rect 1263 -2395 1279 -2361
rect 1313 -2395 1329 -2361
rect 1263 -2411 1329 -2395
<< polycont >>
rect -1409 2361 -1375 2395
rect -1217 2361 -1183 2395
rect -1025 2361 -991 2395
rect -833 2361 -799 2395
rect -641 2361 -607 2395
rect -449 2361 -415 2395
rect -257 2361 -223 2395
rect -65 2361 -31 2395
rect 127 2361 161 2395
rect 319 2361 353 2395
rect 511 2361 545 2395
rect 703 2361 737 2395
rect 895 2361 929 2395
rect 1087 2361 1121 2395
rect 1279 2361 1313 2395
rect -1313 1861 -1279 1895
rect -1121 1861 -1087 1895
rect -929 1861 -895 1895
rect -737 1861 -703 1895
rect -545 1861 -511 1895
rect -353 1861 -319 1895
rect -161 1861 -127 1895
rect 31 1861 65 1895
rect 223 1861 257 1895
rect 415 1861 449 1895
rect 607 1861 641 1895
rect 799 1861 833 1895
rect 991 1861 1025 1895
rect 1183 1861 1217 1895
rect 1375 1861 1409 1895
rect -1313 1753 -1279 1787
rect -1121 1753 -1087 1787
rect -929 1753 -895 1787
rect -737 1753 -703 1787
rect -545 1753 -511 1787
rect -353 1753 -319 1787
rect -161 1753 -127 1787
rect 31 1753 65 1787
rect 223 1753 257 1787
rect 415 1753 449 1787
rect 607 1753 641 1787
rect 799 1753 833 1787
rect 991 1753 1025 1787
rect 1183 1753 1217 1787
rect 1375 1753 1409 1787
rect -1409 1253 -1375 1287
rect -1217 1253 -1183 1287
rect -1025 1253 -991 1287
rect -833 1253 -799 1287
rect -641 1253 -607 1287
rect -449 1253 -415 1287
rect -257 1253 -223 1287
rect -65 1253 -31 1287
rect 127 1253 161 1287
rect 319 1253 353 1287
rect 511 1253 545 1287
rect 703 1253 737 1287
rect 895 1253 929 1287
rect 1087 1253 1121 1287
rect 1279 1253 1313 1287
rect -1409 1145 -1375 1179
rect -1217 1145 -1183 1179
rect -1025 1145 -991 1179
rect -833 1145 -799 1179
rect -641 1145 -607 1179
rect -449 1145 -415 1179
rect -257 1145 -223 1179
rect -65 1145 -31 1179
rect 127 1145 161 1179
rect 319 1145 353 1179
rect 511 1145 545 1179
rect 703 1145 737 1179
rect 895 1145 929 1179
rect 1087 1145 1121 1179
rect 1279 1145 1313 1179
rect -1313 645 -1279 679
rect -1121 645 -1087 679
rect -929 645 -895 679
rect -737 645 -703 679
rect -545 645 -511 679
rect -353 645 -319 679
rect -161 645 -127 679
rect 31 645 65 679
rect 223 645 257 679
rect 415 645 449 679
rect 607 645 641 679
rect 799 645 833 679
rect 991 645 1025 679
rect 1183 645 1217 679
rect 1375 645 1409 679
rect -1313 537 -1279 571
rect -1121 537 -1087 571
rect -929 537 -895 571
rect -737 537 -703 571
rect -545 537 -511 571
rect -353 537 -319 571
rect -161 537 -127 571
rect 31 537 65 571
rect 223 537 257 571
rect 415 537 449 571
rect 607 537 641 571
rect 799 537 833 571
rect 991 537 1025 571
rect 1183 537 1217 571
rect 1375 537 1409 571
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect -1313 -571 -1279 -537
rect -1121 -571 -1087 -537
rect -929 -571 -895 -537
rect -737 -571 -703 -537
rect -545 -571 -511 -537
rect -353 -571 -319 -537
rect -161 -571 -127 -537
rect 31 -571 65 -537
rect 223 -571 257 -537
rect 415 -571 449 -537
rect 607 -571 641 -537
rect 799 -571 833 -537
rect 991 -571 1025 -537
rect 1183 -571 1217 -537
rect 1375 -571 1409 -537
rect -1313 -679 -1279 -645
rect -1121 -679 -1087 -645
rect -929 -679 -895 -645
rect -737 -679 -703 -645
rect -545 -679 -511 -645
rect -353 -679 -319 -645
rect -161 -679 -127 -645
rect 31 -679 65 -645
rect 223 -679 257 -645
rect 415 -679 449 -645
rect 607 -679 641 -645
rect 799 -679 833 -645
rect 991 -679 1025 -645
rect 1183 -679 1217 -645
rect 1375 -679 1409 -645
rect -1409 -1179 -1375 -1145
rect -1217 -1179 -1183 -1145
rect -1025 -1179 -991 -1145
rect -833 -1179 -799 -1145
rect -641 -1179 -607 -1145
rect -449 -1179 -415 -1145
rect -257 -1179 -223 -1145
rect -65 -1179 -31 -1145
rect 127 -1179 161 -1145
rect 319 -1179 353 -1145
rect 511 -1179 545 -1145
rect 703 -1179 737 -1145
rect 895 -1179 929 -1145
rect 1087 -1179 1121 -1145
rect 1279 -1179 1313 -1145
rect -1409 -1287 -1375 -1253
rect -1217 -1287 -1183 -1253
rect -1025 -1287 -991 -1253
rect -833 -1287 -799 -1253
rect -641 -1287 -607 -1253
rect -449 -1287 -415 -1253
rect -257 -1287 -223 -1253
rect -65 -1287 -31 -1253
rect 127 -1287 161 -1253
rect 319 -1287 353 -1253
rect 511 -1287 545 -1253
rect 703 -1287 737 -1253
rect 895 -1287 929 -1253
rect 1087 -1287 1121 -1253
rect 1279 -1287 1313 -1253
rect -1313 -1787 -1279 -1753
rect -1121 -1787 -1087 -1753
rect -929 -1787 -895 -1753
rect -737 -1787 -703 -1753
rect -545 -1787 -511 -1753
rect -353 -1787 -319 -1753
rect -161 -1787 -127 -1753
rect 31 -1787 65 -1753
rect 223 -1787 257 -1753
rect 415 -1787 449 -1753
rect 607 -1787 641 -1753
rect 799 -1787 833 -1753
rect 991 -1787 1025 -1753
rect 1183 -1787 1217 -1753
rect 1375 -1787 1409 -1753
rect -1313 -1895 -1279 -1861
rect -1121 -1895 -1087 -1861
rect -929 -1895 -895 -1861
rect -737 -1895 -703 -1861
rect -545 -1895 -511 -1861
rect -353 -1895 -319 -1861
rect -161 -1895 -127 -1861
rect 31 -1895 65 -1861
rect 223 -1895 257 -1861
rect 415 -1895 449 -1861
rect 607 -1895 641 -1861
rect 799 -1895 833 -1861
rect 991 -1895 1025 -1861
rect 1183 -1895 1217 -1861
rect 1375 -1895 1409 -1861
rect -1409 -2395 -1375 -2361
rect -1217 -2395 -1183 -2361
rect -1025 -2395 -991 -2361
rect -833 -2395 -799 -2361
rect -641 -2395 -607 -2361
rect -449 -2395 -415 -2361
rect -257 -2395 -223 -2361
rect -65 -2395 -31 -2361
rect 127 -2395 161 -2361
rect 319 -2395 353 -2361
rect 511 -2395 545 -2361
rect 703 -2395 737 -2361
rect 895 -2395 929 -2361
rect 1087 -2395 1121 -2361
rect 1279 -2395 1313 -2361
<< locali >>
rect -1571 2463 -1475 2497
rect 1475 2463 1571 2497
rect -1571 2401 -1537 2463
rect 1537 2401 1571 2463
rect -1425 2361 -1409 2395
rect -1375 2361 -1359 2395
rect -1233 2361 -1217 2395
rect -1183 2361 -1167 2395
rect -1041 2361 -1025 2395
rect -991 2361 -975 2395
rect -849 2361 -833 2395
rect -799 2361 -783 2395
rect -657 2361 -641 2395
rect -607 2361 -591 2395
rect -465 2361 -449 2395
rect -415 2361 -399 2395
rect -273 2361 -257 2395
rect -223 2361 -207 2395
rect -81 2361 -65 2395
rect -31 2361 -15 2395
rect 111 2361 127 2395
rect 161 2361 177 2395
rect 303 2361 319 2395
rect 353 2361 369 2395
rect 495 2361 511 2395
rect 545 2361 561 2395
rect 687 2361 703 2395
rect 737 2361 753 2395
rect 879 2361 895 2395
rect 929 2361 945 2395
rect 1071 2361 1087 2395
rect 1121 2361 1137 2395
rect 1263 2361 1279 2395
rect 1313 2361 1329 2395
rect -1457 2311 -1423 2327
rect -1457 1929 -1423 1945
rect -1361 2311 -1327 2327
rect -1361 1929 -1327 1945
rect -1265 2311 -1231 2327
rect -1265 1929 -1231 1945
rect -1169 2311 -1135 2327
rect -1169 1929 -1135 1945
rect -1073 2311 -1039 2327
rect -1073 1929 -1039 1945
rect -977 2311 -943 2327
rect -977 1929 -943 1945
rect -881 2311 -847 2327
rect -881 1929 -847 1945
rect -785 2311 -751 2327
rect -785 1929 -751 1945
rect -689 2311 -655 2327
rect -689 1929 -655 1945
rect -593 2311 -559 2327
rect -593 1929 -559 1945
rect -497 2311 -463 2327
rect -497 1929 -463 1945
rect -401 2311 -367 2327
rect -401 1929 -367 1945
rect -305 2311 -271 2327
rect -305 1929 -271 1945
rect -209 2311 -175 2327
rect -209 1929 -175 1945
rect -113 2311 -79 2327
rect -113 1929 -79 1945
rect -17 2311 17 2327
rect -17 1929 17 1945
rect 79 2311 113 2327
rect 79 1929 113 1945
rect 175 2311 209 2327
rect 175 1929 209 1945
rect 271 2311 305 2327
rect 271 1929 305 1945
rect 367 2311 401 2327
rect 367 1929 401 1945
rect 463 2311 497 2327
rect 463 1929 497 1945
rect 559 2311 593 2327
rect 559 1929 593 1945
rect 655 2311 689 2327
rect 655 1929 689 1945
rect 751 2311 785 2327
rect 751 1929 785 1945
rect 847 2311 881 2327
rect 847 1929 881 1945
rect 943 2311 977 2327
rect 943 1929 977 1945
rect 1039 2311 1073 2327
rect 1039 1929 1073 1945
rect 1135 2311 1169 2327
rect 1135 1929 1169 1945
rect 1231 2311 1265 2327
rect 1231 1929 1265 1945
rect 1327 2311 1361 2327
rect 1327 1929 1361 1945
rect 1423 2311 1457 2327
rect 1423 1929 1457 1945
rect -1329 1861 -1313 1895
rect -1279 1861 -1263 1895
rect -1137 1861 -1121 1895
rect -1087 1861 -1071 1895
rect -945 1861 -929 1895
rect -895 1861 -879 1895
rect -753 1861 -737 1895
rect -703 1861 -687 1895
rect -561 1861 -545 1895
rect -511 1861 -495 1895
rect -369 1861 -353 1895
rect -319 1861 -303 1895
rect -177 1861 -161 1895
rect -127 1861 -111 1895
rect 15 1861 31 1895
rect 65 1861 81 1895
rect 207 1861 223 1895
rect 257 1861 273 1895
rect 399 1861 415 1895
rect 449 1861 465 1895
rect 591 1861 607 1895
rect 641 1861 657 1895
rect 783 1861 799 1895
rect 833 1861 849 1895
rect 975 1861 991 1895
rect 1025 1861 1041 1895
rect 1167 1861 1183 1895
rect 1217 1861 1233 1895
rect 1359 1861 1375 1895
rect 1409 1861 1425 1895
rect -1329 1753 -1313 1787
rect -1279 1753 -1263 1787
rect -1137 1753 -1121 1787
rect -1087 1753 -1071 1787
rect -945 1753 -929 1787
rect -895 1753 -879 1787
rect -753 1753 -737 1787
rect -703 1753 -687 1787
rect -561 1753 -545 1787
rect -511 1753 -495 1787
rect -369 1753 -353 1787
rect -319 1753 -303 1787
rect -177 1753 -161 1787
rect -127 1753 -111 1787
rect 15 1753 31 1787
rect 65 1753 81 1787
rect 207 1753 223 1787
rect 257 1753 273 1787
rect 399 1753 415 1787
rect 449 1753 465 1787
rect 591 1753 607 1787
rect 641 1753 657 1787
rect 783 1753 799 1787
rect 833 1753 849 1787
rect 975 1753 991 1787
rect 1025 1753 1041 1787
rect 1167 1753 1183 1787
rect 1217 1753 1233 1787
rect 1359 1753 1375 1787
rect 1409 1753 1425 1787
rect -1457 1703 -1423 1719
rect -1457 1321 -1423 1337
rect -1361 1703 -1327 1719
rect -1361 1321 -1327 1337
rect -1265 1703 -1231 1719
rect -1265 1321 -1231 1337
rect -1169 1703 -1135 1719
rect -1169 1321 -1135 1337
rect -1073 1703 -1039 1719
rect -1073 1321 -1039 1337
rect -977 1703 -943 1719
rect -977 1321 -943 1337
rect -881 1703 -847 1719
rect -881 1321 -847 1337
rect -785 1703 -751 1719
rect -785 1321 -751 1337
rect -689 1703 -655 1719
rect -689 1321 -655 1337
rect -593 1703 -559 1719
rect -593 1321 -559 1337
rect -497 1703 -463 1719
rect -497 1321 -463 1337
rect -401 1703 -367 1719
rect -401 1321 -367 1337
rect -305 1703 -271 1719
rect -305 1321 -271 1337
rect -209 1703 -175 1719
rect -209 1321 -175 1337
rect -113 1703 -79 1719
rect -113 1321 -79 1337
rect -17 1703 17 1719
rect -17 1321 17 1337
rect 79 1703 113 1719
rect 79 1321 113 1337
rect 175 1703 209 1719
rect 175 1321 209 1337
rect 271 1703 305 1719
rect 271 1321 305 1337
rect 367 1703 401 1719
rect 367 1321 401 1337
rect 463 1703 497 1719
rect 463 1321 497 1337
rect 559 1703 593 1719
rect 559 1321 593 1337
rect 655 1703 689 1719
rect 655 1321 689 1337
rect 751 1703 785 1719
rect 751 1321 785 1337
rect 847 1703 881 1719
rect 847 1321 881 1337
rect 943 1703 977 1719
rect 943 1321 977 1337
rect 1039 1703 1073 1719
rect 1039 1321 1073 1337
rect 1135 1703 1169 1719
rect 1135 1321 1169 1337
rect 1231 1703 1265 1719
rect 1231 1321 1265 1337
rect 1327 1703 1361 1719
rect 1327 1321 1361 1337
rect 1423 1703 1457 1719
rect 1423 1321 1457 1337
rect -1425 1253 -1409 1287
rect -1375 1253 -1359 1287
rect -1233 1253 -1217 1287
rect -1183 1253 -1167 1287
rect -1041 1253 -1025 1287
rect -991 1253 -975 1287
rect -849 1253 -833 1287
rect -799 1253 -783 1287
rect -657 1253 -641 1287
rect -607 1253 -591 1287
rect -465 1253 -449 1287
rect -415 1253 -399 1287
rect -273 1253 -257 1287
rect -223 1253 -207 1287
rect -81 1253 -65 1287
rect -31 1253 -15 1287
rect 111 1253 127 1287
rect 161 1253 177 1287
rect 303 1253 319 1287
rect 353 1253 369 1287
rect 495 1253 511 1287
rect 545 1253 561 1287
rect 687 1253 703 1287
rect 737 1253 753 1287
rect 879 1253 895 1287
rect 929 1253 945 1287
rect 1071 1253 1087 1287
rect 1121 1253 1137 1287
rect 1263 1253 1279 1287
rect 1313 1253 1329 1287
rect -1425 1145 -1409 1179
rect -1375 1145 -1359 1179
rect -1233 1145 -1217 1179
rect -1183 1145 -1167 1179
rect -1041 1145 -1025 1179
rect -991 1145 -975 1179
rect -849 1145 -833 1179
rect -799 1145 -783 1179
rect -657 1145 -641 1179
rect -607 1145 -591 1179
rect -465 1145 -449 1179
rect -415 1145 -399 1179
rect -273 1145 -257 1179
rect -223 1145 -207 1179
rect -81 1145 -65 1179
rect -31 1145 -15 1179
rect 111 1145 127 1179
rect 161 1145 177 1179
rect 303 1145 319 1179
rect 353 1145 369 1179
rect 495 1145 511 1179
rect 545 1145 561 1179
rect 687 1145 703 1179
rect 737 1145 753 1179
rect 879 1145 895 1179
rect 929 1145 945 1179
rect 1071 1145 1087 1179
rect 1121 1145 1137 1179
rect 1263 1145 1279 1179
rect 1313 1145 1329 1179
rect -1457 1095 -1423 1111
rect -1457 713 -1423 729
rect -1361 1095 -1327 1111
rect -1361 713 -1327 729
rect -1265 1095 -1231 1111
rect -1265 713 -1231 729
rect -1169 1095 -1135 1111
rect -1169 713 -1135 729
rect -1073 1095 -1039 1111
rect -1073 713 -1039 729
rect -977 1095 -943 1111
rect -977 713 -943 729
rect -881 1095 -847 1111
rect -881 713 -847 729
rect -785 1095 -751 1111
rect -785 713 -751 729
rect -689 1095 -655 1111
rect -689 713 -655 729
rect -593 1095 -559 1111
rect -593 713 -559 729
rect -497 1095 -463 1111
rect -497 713 -463 729
rect -401 1095 -367 1111
rect -401 713 -367 729
rect -305 1095 -271 1111
rect -305 713 -271 729
rect -209 1095 -175 1111
rect -209 713 -175 729
rect -113 1095 -79 1111
rect -113 713 -79 729
rect -17 1095 17 1111
rect -17 713 17 729
rect 79 1095 113 1111
rect 79 713 113 729
rect 175 1095 209 1111
rect 175 713 209 729
rect 271 1095 305 1111
rect 271 713 305 729
rect 367 1095 401 1111
rect 367 713 401 729
rect 463 1095 497 1111
rect 463 713 497 729
rect 559 1095 593 1111
rect 559 713 593 729
rect 655 1095 689 1111
rect 655 713 689 729
rect 751 1095 785 1111
rect 751 713 785 729
rect 847 1095 881 1111
rect 847 713 881 729
rect 943 1095 977 1111
rect 943 713 977 729
rect 1039 1095 1073 1111
rect 1039 713 1073 729
rect 1135 1095 1169 1111
rect 1135 713 1169 729
rect 1231 1095 1265 1111
rect 1231 713 1265 729
rect 1327 1095 1361 1111
rect 1327 713 1361 729
rect 1423 1095 1457 1111
rect 1423 713 1457 729
rect -1329 645 -1313 679
rect -1279 645 -1263 679
rect -1137 645 -1121 679
rect -1087 645 -1071 679
rect -945 645 -929 679
rect -895 645 -879 679
rect -753 645 -737 679
rect -703 645 -687 679
rect -561 645 -545 679
rect -511 645 -495 679
rect -369 645 -353 679
rect -319 645 -303 679
rect -177 645 -161 679
rect -127 645 -111 679
rect 15 645 31 679
rect 65 645 81 679
rect 207 645 223 679
rect 257 645 273 679
rect 399 645 415 679
rect 449 645 465 679
rect 591 645 607 679
rect 641 645 657 679
rect 783 645 799 679
rect 833 645 849 679
rect 975 645 991 679
rect 1025 645 1041 679
rect 1167 645 1183 679
rect 1217 645 1233 679
rect 1359 645 1375 679
rect 1409 645 1425 679
rect -1329 537 -1313 571
rect -1279 537 -1263 571
rect -1137 537 -1121 571
rect -1087 537 -1071 571
rect -945 537 -929 571
rect -895 537 -879 571
rect -753 537 -737 571
rect -703 537 -687 571
rect -561 537 -545 571
rect -511 537 -495 571
rect -369 537 -353 571
rect -319 537 -303 571
rect -177 537 -161 571
rect -127 537 -111 571
rect 15 537 31 571
rect 65 537 81 571
rect 207 537 223 571
rect 257 537 273 571
rect 399 537 415 571
rect 449 537 465 571
rect 591 537 607 571
rect 641 537 657 571
rect 783 537 799 571
rect 833 537 849 571
rect 975 537 991 571
rect 1025 537 1041 571
rect 1167 537 1183 571
rect 1217 537 1233 571
rect 1359 537 1375 571
rect 1409 537 1425 571
rect -1457 487 -1423 503
rect -1457 105 -1423 121
rect -1361 487 -1327 503
rect -1361 105 -1327 121
rect -1265 487 -1231 503
rect -1265 105 -1231 121
rect -1169 487 -1135 503
rect -1169 105 -1135 121
rect -1073 487 -1039 503
rect -1073 105 -1039 121
rect -977 487 -943 503
rect -977 105 -943 121
rect -881 487 -847 503
rect -881 105 -847 121
rect -785 487 -751 503
rect -785 105 -751 121
rect -689 487 -655 503
rect -689 105 -655 121
rect -593 487 -559 503
rect -593 105 -559 121
rect -497 487 -463 503
rect -497 105 -463 121
rect -401 487 -367 503
rect -401 105 -367 121
rect -305 487 -271 503
rect -305 105 -271 121
rect -209 487 -175 503
rect -209 105 -175 121
rect -113 487 -79 503
rect -113 105 -79 121
rect -17 487 17 503
rect -17 105 17 121
rect 79 487 113 503
rect 79 105 113 121
rect 175 487 209 503
rect 175 105 209 121
rect 271 487 305 503
rect 271 105 305 121
rect 367 487 401 503
rect 367 105 401 121
rect 463 487 497 503
rect 463 105 497 121
rect 559 487 593 503
rect 559 105 593 121
rect 655 487 689 503
rect 655 105 689 121
rect 751 487 785 503
rect 751 105 785 121
rect 847 487 881 503
rect 847 105 881 121
rect 943 487 977 503
rect 943 105 977 121
rect 1039 487 1073 503
rect 1039 105 1073 121
rect 1135 487 1169 503
rect 1135 105 1169 121
rect 1231 487 1265 503
rect 1231 105 1265 121
rect 1327 487 1361 503
rect 1327 105 1361 121
rect 1423 487 1457 503
rect 1423 105 1457 121
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect -1457 -121 -1423 -105
rect -1457 -503 -1423 -487
rect -1361 -121 -1327 -105
rect -1361 -503 -1327 -487
rect -1265 -121 -1231 -105
rect -1265 -503 -1231 -487
rect -1169 -121 -1135 -105
rect -1169 -503 -1135 -487
rect -1073 -121 -1039 -105
rect -1073 -503 -1039 -487
rect -977 -121 -943 -105
rect -977 -503 -943 -487
rect -881 -121 -847 -105
rect -881 -503 -847 -487
rect -785 -121 -751 -105
rect -785 -503 -751 -487
rect -689 -121 -655 -105
rect -689 -503 -655 -487
rect -593 -121 -559 -105
rect -593 -503 -559 -487
rect -497 -121 -463 -105
rect -497 -503 -463 -487
rect -401 -121 -367 -105
rect -401 -503 -367 -487
rect -305 -121 -271 -105
rect -305 -503 -271 -487
rect -209 -121 -175 -105
rect -209 -503 -175 -487
rect -113 -121 -79 -105
rect -113 -503 -79 -487
rect -17 -121 17 -105
rect -17 -503 17 -487
rect 79 -121 113 -105
rect 79 -503 113 -487
rect 175 -121 209 -105
rect 175 -503 209 -487
rect 271 -121 305 -105
rect 271 -503 305 -487
rect 367 -121 401 -105
rect 367 -503 401 -487
rect 463 -121 497 -105
rect 463 -503 497 -487
rect 559 -121 593 -105
rect 559 -503 593 -487
rect 655 -121 689 -105
rect 655 -503 689 -487
rect 751 -121 785 -105
rect 751 -503 785 -487
rect 847 -121 881 -105
rect 847 -503 881 -487
rect 943 -121 977 -105
rect 943 -503 977 -487
rect 1039 -121 1073 -105
rect 1039 -503 1073 -487
rect 1135 -121 1169 -105
rect 1135 -503 1169 -487
rect 1231 -121 1265 -105
rect 1231 -503 1265 -487
rect 1327 -121 1361 -105
rect 1327 -503 1361 -487
rect 1423 -121 1457 -105
rect 1423 -503 1457 -487
rect -1329 -571 -1313 -537
rect -1279 -571 -1263 -537
rect -1137 -571 -1121 -537
rect -1087 -571 -1071 -537
rect -945 -571 -929 -537
rect -895 -571 -879 -537
rect -753 -571 -737 -537
rect -703 -571 -687 -537
rect -561 -571 -545 -537
rect -511 -571 -495 -537
rect -369 -571 -353 -537
rect -319 -571 -303 -537
rect -177 -571 -161 -537
rect -127 -571 -111 -537
rect 15 -571 31 -537
rect 65 -571 81 -537
rect 207 -571 223 -537
rect 257 -571 273 -537
rect 399 -571 415 -537
rect 449 -571 465 -537
rect 591 -571 607 -537
rect 641 -571 657 -537
rect 783 -571 799 -537
rect 833 -571 849 -537
rect 975 -571 991 -537
rect 1025 -571 1041 -537
rect 1167 -571 1183 -537
rect 1217 -571 1233 -537
rect 1359 -571 1375 -537
rect 1409 -571 1425 -537
rect -1329 -679 -1313 -645
rect -1279 -679 -1263 -645
rect -1137 -679 -1121 -645
rect -1087 -679 -1071 -645
rect -945 -679 -929 -645
rect -895 -679 -879 -645
rect -753 -679 -737 -645
rect -703 -679 -687 -645
rect -561 -679 -545 -645
rect -511 -679 -495 -645
rect -369 -679 -353 -645
rect -319 -679 -303 -645
rect -177 -679 -161 -645
rect -127 -679 -111 -645
rect 15 -679 31 -645
rect 65 -679 81 -645
rect 207 -679 223 -645
rect 257 -679 273 -645
rect 399 -679 415 -645
rect 449 -679 465 -645
rect 591 -679 607 -645
rect 641 -679 657 -645
rect 783 -679 799 -645
rect 833 -679 849 -645
rect 975 -679 991 -645
rect 1025 -679 1041 -645
rect 1167 -679 1183 -645
rect 1217 -679 1233 -645
rect 1359 -679 1375 -645
rect 1409 -679 1425 -645
rect -1457 -729 -1423 -713
rect -1457 -1111 -1423 -1095
rect -1361 -729 -1327 -713
rect -1361 -1111 -1327 -1095
rect -1265 -729 -1231 -713
rect -1265 -1111 -1231 -1095
rect -1169 -729 -1135 -713
rect -1169 -1111 -1135 -1095
rect -1073 -729 -1039 -713
rect -1073 -1111 -1039 -1095
rect -977 -729 -943 -713
rect -977 -1111 -943 -1095
rect -881 -729 -847 -713
rect -881 -1111 -847 -1095
rect -785 -729 -751 -713
rect -785 -1111 -751 -1095
rect -689 -729 -655 -713
rect -689 -1111 -655 -1095
rect -593 -729 -559 -713
rect -593 -1111 -559 -1095
rect -497 -729 -463 -713
rect -497 -1111 -463 -1095
rect -401 -729 -367 -713
rect -401 -1111 -367 -1095
rect -305 -729 -271 -713
rect -305 -1111 -271 -1095
rect -209 -729 -175 -713
rect -209 -1111 -175 -1095
rect -113 -729 -79 -713
rect -113 -1111 -79 -1095
rect -17 -729 17 -713
rect -17 -1111 17 -1095
rect 79 -729 113 -713
rect 79 -1111 113 -1095
rect 175 -729 209 -713
rect 175 -1111 209 -1095
rect 271 -729 305 -713
rect 271 -1111 305 -1095
rect 367 -729 401 -713
rect 367 -1111 401 -1095
rect 463 -729 497 -713
rect 463 -1111 497 -1095
rect 559 -729 593 -713
rect 559 -1111 593 -1095
rect 655 -729 689 -713
rect 655 -1111 689 -1095
rect 751 -729 785 -713
rect 751 -1111 785 -1095
rect 847 -729 881 -713
rect 847 -1111 881 -1095
rect 943 -729 977 -713
rect 943 -1111 977 -1095
rect 1039 -729 1073 -713
rect 1039 -1111 1073 -1095
rect 1135 -729 1169 -713
rect 1135 -1111 1169 -1095
rect 1231 -729 1265 -713
rect 1231 -1111 1265 -1095
rect 1327 -729 1361 -713
rect 1327 -1111 1361 -1095
rect 1423 -729 1457 -713
rect 1423 -1111 1457 -1095
rect -1425 -1179 -1409 -1145
rect -1375 -1179 -1359 -1145
rect -1233 -1179 -1217 -1145
rect -1183 -1179 -1167 -1145
rect -1041 -1179 -1025 -1145
rect -991 -1179 -975 -1145
rect -849 -1179 -833 -1145
rect -799 -1179 -783 -1145
rect -657 -1179 -641 -1145
rect -607 -1179 -591 -1145
rect -465 -1179 -449 -1145
rect -415 -1179 -399 -1145
rect -273 -1179 -257 -1145
rect -223 -1179 -207 -1145
rect -81 -1179 -65 -1145
rect -31 -1179 -15 -1145
rect 111 -1179 127 -1145
rect 161 -1179 177 -1145
rect 303 -1179 319 -1145
rect 353 -1179 369 -1145
rect 495 -1179 511 -1145
rect 545 -1179 561 -1145
rect 687 -1179 703 -1145
rect 737 -1179 753 -1145
rect 879 -1179 895 -1145
rect 929 -1179 945 -1145
rect 1071 -1179 1087 -1145
rect 1121 -1179 1137 -1145
rect 1263 -1179 1279 -1145
rect 1313 -1179 1329 -1145
rect -1425 -1287 -1409 -1253
rect -1375 -1287 -1359 -1253
rect -1233 -1287 -1217 -1253
rect -1183 -1287 -1167 -1253
rect -1041 -1287 -1025 -1253
rect -991 -1287 -975 -1253
rect -849 -1287 -833 -1253
rect -799 -1287 -783 -1253
rect -657 -1287 -641 -1253
rect -607 -1287 -591 -1253
rect -465 -1287 -449 -1253
rect -415 -1287 -399 -1253
rect -273 -1287 -257 -1253
rect -223 -1287 -207 -1253
rect -81 -1287 -65 -1253
rect -31 -1287 -15 -1253
rect 111 -1287 127 -1253
rect 161 -1287 177 -1253
rect 303 -1287 319 -1253
rect 353 -1287 369 -1253
rect 495 -1287 511 -1253
rect 545 -1287 561 -1253
rect 687 -1287 703 -1253
rect 737 -1287 753 -1253
rect 879 -1287 895 -1253
rect 929 -1287 945 -1253
rect 1071 -1287 1087 -1253
rect 1121 -1287 1137 -1253
rect 1263 -1287 1279 -1253
rect 1313 -1287 1329 -1253
rect -1457 -1337 -1423 -1321
rect -1457 -1719 -1423 -1703
rect -1361 -1337 -1327 -1321
rect -1361 -1719 -1327 -1703
rect -1265 -1337 -1231 -1321
rect -1265 -1719 -1231 -1703
rect -1169 -1337 -1135 -1321
rect -1169 -1719 -1135 -1703
rect -1073 -1337 -1039 -1321
rect -1073 -1719 -1039 -1703
rect -977 -1337 -943 -1321
rect -977 -1719 -943 -1703
rect -881 -1337 -847 -1321
rect -881 -1719 -847 -1703
rect -785 -1337 -751 -1321
rect -785 -1719 -751 -1703
rect -689 -1337 -655 -1321
rect -689 -1719 -655 -1703
rect -593 -1337 -559 -1321
rect -593 -1719 -559 -1703
rect -497 -1337 -463 -1321
rect -497 -1719 -463 -1703
rect -401 -1337 -367 -1321
rect -401 -1719 -367 -1703
rect -305 -1337 -271 -1321
rect -305 -1719 -271 -1703
rect -209 -1337 -175 -1321
rect -209 -1719 -175 -1703
rect -113 -1337 -79 -1321
rect -113 -1719 -79 -1703
rect -17 -1337 17 -1321
rect -17 -1719 17 -1703
rect 79 -1337 113 -1321
rect 79 -1719 113 -1703
rect 175 -1337 209 -1321
rect 175 -1719 209 -1703
rect 271 -1337 305 -1321
rect 271 -1719 305 -1703
rect 367 -1337 401 -1321
rect 367 -1719 401 -1703
rect 463 -1337 497 -1321
rect 463 -1719 497 -1703
rect 559 -1337 593 -1321
rect 559 -1719 593 -1703
rect 655 -1337 689 -1321
rect 655 -1719 689 -1703
rect 751 -1337 785 -1321
rect 751 -1719 785 -1703
rect 847 -1337 881 -1321
rect 847 -1719 881 -1703
rect 943 -1337 977 -1321
rect 943 -1719 977 -1703
rect 1039 -1337 1073 -1321
rect 1039 -1719 1073 -1703
rect 1135 -1337 1169 -1321
rect 1135 -1719 1169 -1703
rect 1231 -1337 1265 -1321
rect 1231 -1719 1265 -1703
rect 1327 -1337 1361 -1321
rect 1327 -1719 1361 -1703
rect 1423 -1337 1457 -1321
rect 1423 -1719 1457 -1703
rect -1329 -1787 -1313 -1753
rect -1279 -1787 -1263 -1753
rect -1137 -1787 -1121 -1753
rect -1087 -1787 -1071 -1753
rect -945 -1787 -929 -1753
rect -895 -1787 -879 -1753
rect -753 -1787 -737 -1753
rect -703 -1787 -687 -1753
rect -561 -1787 -545 -1753
rect -511 -1787 -495 -1753
rect -369 -1787 -353 -1753
rect -319 -1787 -303 -1753
rect -177 -1787 -161 -1753
rect -127 -1787 -111 -1753
rect 15 -1787 31 -1753
rect 65 -1787 81 -1753
rect 207 -1787 223 -1753
rect 257 -1787 273 -1753
rect 399 -1787 415 -1753
rect 449 -1787 465 -1753
rect 591 -1787 607 -1753
rect 641 -1787 657 -1753
rect 783 -1787 799 -1753
rect 833 -1787 849 -1753
rect 975 -1787 991 -1753
rect 1025 -1787 1041 -1753
rect 1167 -1787 1183 -1753
rect 1217 -1787 1233 -1753
rect 1359 -1787 1375 -1753
rect 1409 -1787 1425 -1753
rect -1329 -1895 -1313 -1861
rect -1279 -1895 -1263 -1861
rect -1137 -1895 -1121 -1861
rect -1087 -1895 -1071 -1861
rect -945 -1895 -929 -1861
rect -895 -1895 -879 -1861
rect -753 -1895 -737 -1861
rect -703 -1895 -687 -1861
rect -561 -1895 -545 -1861
rect -511 -1895 -495 -1861
rect -369 -1895 -353 -1861
rect -319 -1895 -303 -1861
rect -177 -1895 -161 -1861
rect -127 -1895 -111 -1861
rect 15 -1895 31 -1861
rect 65 -1895 81 -1861
rect 207 -1895 223 -1861
rect 257 -1895 273 -1861
rect 399 -1895 415 -1861
rect 449 -1895 465 -1861
rect 591 -1895 607 -1861
rect 641 -1895 657 -1861
rect 783 -1895 799 -1861
rect 833 -1895 849 -1861
rect 975 -1895 991 -1861
rect 1025 -1895 1041 -1861
rect 1167 -1895 1183 -1861
rect 1217 -1895 1233 -1861
rect 1359 -1895 1375 -1861
rect 1409 -1895 1425 -1861
rect -1457 -1945 -1423 -1929
rect -1457 -2327 -1423 -2311
rect -1361 -1945 -1327 -1929
rect -1361 -2327 -1327 -2311
rect -1265 -1945 -1231 -1929
rect -1265 -2327 -1231 -2311
rect -1169 -1945 -1135 -1929
rect -1169 -2327 -1135 -2311
rect -1073 -1945 -1039 -1929
rect -1073 -2327 -1039 -2311
rect -977 -1945 -943 -1929
rect -977 -2327 -943 -2311
rect -881 -1945 -847 -1929
rect -881 -2327 -847 -2311
rect -785 -1945 -751 -1929
rect -785 -2327 -751 -2311
rect -689 -1945 -655 -1929
rect -689 -2327 -655 -2311
rect -593 -1945 -559 -1929
rect -593 -2327 -559 -2311
rect -497 -1945 -463 -1929
rect -497 -2327 -463 -2311
rect -401 -1945 -367 -1929
rect -401 -2327 -367 -2311
rect -305 -1945 -271 -1929
rect -305 -2327 -271 -2311
rect -209 -1945 -175 -1929
rect -209 -2327 -175 -2311
rect -113 -1945 -79 -1929
rect -113 -2327 -79 -2311
rect -17 -1945 17 -1929
rect -17 -2327 17 -2311
rect 79 -1945 113 -1929
rect 79 -2327 113 -2311
rect 175 -1945 209 -1929
rect 175 -2327 209 -2311
rect 271 -1945 305 -1929
rect 271 -2327 305 -2311
rect 367 -1945 401 -1929
rect 367 -2327 401 -2311
rect 463 -1945 497 -1929
rect 463 -2327 497 -2311
rect 559 -1945 593 -1929
rect 559 -2327 593 -2311
rect 655 -1945 689 -1929
rect 655 -2327 689 -2311
rect 751 -1945 785 -1929
rect 751 -2327 785 -2311
rect 847 -1945 881 -1929
rect 847 -2327 881 -2311
rect 943 -1945 977 -1929
rect 943 -2327 977 -2311
rect 1039 -1945 1073 -1929
rect 1039 -2327 1073 -2311
rect 1135 -1945 1169 -1929
rect 1135 -2327 1169 -2311
rect 1231 -1945 1265 -1929
rect 1231 -2327 1265 -2311
rect 1327 -1945 1361 -1929
rect 1327 -2327 1361 -2311
rect 1423 -1945 1457 -1929
rect 1423 -2327 1457 -2311
rect -1425 -2395 -1409 -2361
rect -1375 -2395 -1359 -2361
rect -1233 -2395 -1217 -2361
rect -1183 -2395 -1167 -2361
rect -1041 -2395 -1025 -2361
rect -991 -2395 -975 -2361
rect -849 -2395 -833 -2361
rect -799 -2395 -783 -2361
rect -657 -2395 -641 -2361
rect -607 -2395 -591 -2361
rect -465 -2395 -449 -2361
rect -415 -2395 -399 -2361
rect -273 -2395 -257 -2361
rect -223 -2395 -207 -2361
rect -81 -2395 -65 -2361
rect -31 -2395 -15 -2361
rect 111 -2395 127 -2361
rect 161 -2395 177 -2361
rect 303 -2395 319 -2361
rect 353 -2395 369 -2361
rect 495 -2395 511 -2361
rect 545 -2395 561 -2361
rect 687 -2395 703 -2361
rect 737 -2395 753 -2361
rect 879 -2395 895 -2361
rect 929 -2395 945 -2361
rect 1071 -2395 1087 -2361
rect 1121 -2395 1137 -2361
rect 1263 -2395 1279 -2361
rect 1313 -2395 1329 -2361
rect -1571 -2463 -1537 -2401
rect 1537 -2463 1571 -2401
rect -1571 -2497 -1475 -2463
rect 1475 -2497 1571 -2463
<< viali >>
rect -1409 2361 -1375 2395
rect -1217 2361 -1183 2395
rect -1025 2361 -991 2395
rect -833 2361 -799 2395
rect -641 2361 -607 2395
rect -449 2361 -415 2395
rect -257 2361 -223 2395
rect -65 2361 -31 2395
rect 127 2361 161 2395
rect 319 2361 353 2395
rect 511 2361 545 2395
rect 703 2361 737 2395
rect 895 2361 929 2395
rect 1087 2361 1121 2395
rect 1279 2361 1313 2395
rect -1457 1945 -1423 2311
rect -1361 1945 -1327 2311
rect -1265 1945 -1231 2311
rect -1169 1945 -1135 2311
rect -1073 1945 -1039 2311
rect -977 1945 -943 2311
rect -881 1945 -847 2311
rect -785 1945 -751 2311
rect -689 1945 -655 2311
rect -593 1945 -559 2311
rect -497 1945 -463 2311
rect -401 1945 -367 2311
rect -305 1945 -271 2311
rect -209 1945 -175 2311
rect -113 1945 -79 2311
rect -17 1945 17 2311
rect 79 1945 113 2311
rect 175 1945 209 2311
rect 271 1945 305 2311
rect 367 1945 401 2311
rect 463 1945 497 2311
rect 559 1945 593 2311
rect 655 1945 689 2311
rect 751 1945 785 2311
rect 847 1945 881 2311
rect 943 1945 977 2311
rect 1039 1945 1073 2311
rect 1135 1945 1169 2311
rect 1231 1945 1265 2311
rect 1327 1945 1361 2311
rect 1423 1945 1457 2311
rect -1313 1861 -1279 1895
rect -1121 1861 -1087 1895
rect -929 1861 -895 1895
rect -737 1861 -703 1895
rect -545 1861 -511 1895
rect -353 1861 -319 1895
rect -161 1861 -127 1895
rect 31 1861 65 1895
rect 223 1861 257 1895
rect 415 1861 449 1895
rect 607 1861 641 1895
rect 799 1861 833 1895
rect 991 1861 1025 1895
rect 1183 1861 1217 1895
rect 1375 1861 1409 1895
rect -1313 1753 -1279 1787
rect -1121 1753 -1087 1787
rect -929 1753 -895 1787
rect -737 1753 -703 1787
rect -545 1753 -511 1787
rect -353 1753 -319 1787
rect -161 1753 -127 1787
rect 31 1753 65 1787
rect 223 1753 257 1787
rect 415 1753 449 1787
rect 607 1753 641 1787
rect 799 1753 833 1787
rect 991 1753 1025 1787
rect 1183 1753 1217 1787
rect 1375 1753 1409 1787
rect -1457 1337 -1423 1703
rect -1361 1337 -1327 1703
rect -1265 1337 -1231 1703
rect -1169 1337 -1135 1703
rect -1073 1337 -1039 1703
rect -977 1337 -943 1703
rect -881 1337 -847 1703
rect -785 1337 -751 1703
rect -689 1337 -655 1703
rect -593 1337 -559 1703
rect -497 1337 -463 1703
rect -401 1337 -367 1703
rect -305 1337 -271 1703
rect -209 1337 -175 1703
rect -113 1337 -79 1703
rect -17 1337 17 1703
rect 79 1337 113 1703
rect 175 1337 209 1703
rect 271 1337 305 1703
rect 367 1337 401 1703
rect 463 1337 497 1703
rect 559 1337 593 1703
rect 655 1337 689 1703
rect 751 1337 785 1703
rect 847 1337 881 1703
rect 943 1337 977 1703
rect 1039 1337 1073 1703
rect 1135 1337 1169 1703
rect 1231 1337 1265 1703
rect 1327 1337 1361 1703
rect 1423 1337 1457 1703
rect -1409 1253 -1375 1287
rect -1217 1253 -1183 1287
rect -1025 1253 -991 1287
rect -833 1253 -799 1287
rect -641 1253 -607 1287
rect -449 1253 -415 1287
rect -257 1253 -223 1287
rect -65 1253 -31 1287
rect 127 1253 161 1287
rect 319 1253 353 1287
rect 511 1253 545 1287
rect 703 1253 737 1287
rect 895 1253 929 1287
rect 1087 1253 1121 1287
rect 1279 1253 1313 1287
rect -1409 1145 -1375 1179
rect -1217 1145 -1183 1179
rect -1025 1145 -991 1179
rect -833 1145 -799 1179
rect -641 1145 -607 1179
rect -449 1145 -415 1179
rect -257 1145 -223 1179
rect -65 1145 -31 1179
rect 127 1145 161 1179
rect 319 1145 353 1179
rect 511 1145 545 1179
rect 703 1145 737 1179
rect 895 1145 929 1179
rect 1087 1145 1121 1179
rect 1279 1145 1313 1179
rect -1457 729 -1423 1095
rect -1361 729 -1327 1095
rect -1265 729 -1231 1095
rect -1169 729 -1135 1095
rect -1073 729 -1039 1095
rect -977 729 -943 1095
rect -881 729 -847 1095
rect -785 729 -751 1095
rect -689 729 -655 1095
rect -593 729 -559 1095
rect -497 729 -463 1095
rect -401 729 -367 1095
rect -305 729 -271 1095
rect -209 729 -175 1095
rect -113 729 -79 1095
rect -17 729 17 1095
rect 79 729 113 1095
rect 175 729 209 1095
rect 271 729 305 1095
rect 367 729 401 1095
rect 463 729 497 1095
rect 559 729 593 1095
rect 655 729 689 1095
rect 751 729 785 1095
rect 847 729 881 1095
rect 943 729 977 1095
rect 1039 729 1073 1095
rect 1135 729 1169 1095
rect 1231 729 1265 1095
rect 1327 729 1361 1095
rect 1423 729 1457 1095
rect -1313 645 -1279 679
rect -1121 645 -1087 679
rect -929 645 -895 679
rect -737 645 -703 679
rect -545 645 -511 679
rect -353 645 -319 679
rect -161 645 -127 679
rect 31 645 65 679
rect 223 645 257 679
rect 415 645 449 679
rect 607 645 641 679
rect 799 645 833 679
rect 991 645 1025 679
rect 1183 645 1217 679
rect 1375 645 1409 679
rect -1313 537 -1279 571
rect -1121 537 -1087 571
rect -929 537 -895 571
rect -737 537 -703 571
rect -545 537 -511 571
rect -353 537 -319 571
rect -161 537 -127 571
rect 31 537 65 571
rect 223 537 257 571
rect 415 537 449 571
rect 607 537 641 571
rect 799 537 833 571
rect 991 537 1025 571
rect 1183 537 1217 571
rect 1375 537 1409 571
rect -1457 121 -1423 487
rect -1361 121 -1327 487
rect -1265 121 -1231 487
rect -1169 121 -1135 487
rect -1073 121 -1039 487
rect -977 121 -943 487
rect -881 121 -847 487
rect -785 121 -751 487
rect -689 121 -655 487
rect -593 121 -559 487
rect -497 121 -463 487
rect -401 121 -367 487
rect -305 121 -271 487
rect -209 121 -175 487
rect -113 121 -79 487
rect -17 121 17 487
rect 79 121 113 487
rect 175 121 209 487
rect 271 121 305 487
rect 367 121 401 487
rect 463 121 497 487
rect 559 121 593 487
rect 655 121 689 487
rect 751 121 785 487
rect 847 121 881 487
rect 943 121 977 487
rect 1039 121 1073 487
rect 1135 121 1169 487
rect 1231 121 1265 487
rect 1327 121 1361 487
rect 1423 121 1457 487
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect -1457 -487 -1423 -121
rect -1361 -487 -1327 -121
rect -1265 -487 -1231 -121
rect -1169 -487 -1135 -121
rect -1073 -487 -1039 -121
rect -977 -487 -943 -121
rect -881 -487 -847 -121
rect -785 -487 -751 -121
rect -689 -487 -655 -121
rect -593 -487 -559 -121
rect -497 -487 -463 -121
rect -401 -487 -367 -121
rect -305 -487 -271 -121
rect -209 -487 -175 -121
rect -113 -487 -79 -121
rect -17 -487 17 -121
rect 79 -487 113 -121
rect 175 -487 209 -121
rect 271 -487 305 -121
rect 367 -487 401 -121
rect 463 -487 497 -121
rect 559 -487 593 -121
rect 655 -487 689 -121
rect 751 -487 785 -121
rect 847 -487 881 -121
rect 943 -487 977 -121
rect 1039 -487 1073 -121
rect 1135 -487 1169 -121
rect 1231 -487 1265 -121
rect 1327 -487 1361 -121
rect 1423 -487 1457 -121
rect -1313 -571 -1279 -537
rect -1121 -571 -1087 -537
rect -929 -571 -895 -537
rect -737 -571 -703 -537
rect -545 -571 -511 -537
rect -353 -571 -319 -537
rect -161 -571 -127 -537
rect 31 -571 65 -537
rect 223 -571 257 -537
rect 415 -571 449 -537
rect 607 -571 641 -537
rect 799 -571 833 -537
rect 991 -571 1025 -537
rect 1183 -571 1217 -537
rect 1375 -571 1409 -537
rect -1313 -679 -1279 -645
rect -1121 -679 -1087 -645
rect -929 -679 -895 -645
rect -737 -679 -703 -645
rect -545 -679 -511 -645
rect -353 -679 -319 -645
rect -161 -679 -127 -645
rect 31 -679 65 -645
rect 223 -679 257 -645
rect 415 -679 449 -645
rect 607 -679 641 -645
rect 799 -679 833 -645
rect 991 -679 1025 -645
rect 1183 -679 1217 -645
rect 1375 -679 1409 -645
rect -1457 -1095 -1423 -729
rect -1361 -1095 -1327 -729
rect -1265 -1095 -1231 -729
rect -1169 -1095 -1135 -729
rect -1073 -1095 -1039 -729
rect -977 -1095 -943 -729
rect -881 -1095 -847 -729
rect -785 -1095 -751 -729
rect -689 -1095 -655 -729
rect -593 -1095 -559 -729
rect -497 -1095 -463 -729
rect -401 -1095 -367 -729
rect -305 -1095 -271 -729
rect -209 -1095 -175 -729
rect -113 -1095 -79 -729
rect -17 -1095 17 -729
rect 79 -1095 113 -729
rect 175 -1095 209 -729
rect 271 -1095 305 -729
rect 367 -1095 401 -729
rect 463 -1095 497 -729
rect 559 -1095 593 -729
rect 655 -1095 689 -729
rect 751 -1095 785 -729
rect 847 -1095 881 -729
rect 943 -1095 977 -729
rect 1039 -1095 1073 -729
rect 1135 -1095 1169 -729
rect 1231 -1095 1265 -729
rect 1327 -1095 1361 -729
rect 1423 -1095 1457 -729
rect -1409 -1179 -1375 -1145
rect -1217 -1179 -1183 -1145
rect -1025 -1179 -991 -1145
rect -833 -1179 -799 -1145
rect -641 -1179 -607 -1145
rect -449 -1179 -415 -1145
rect -257 -1179 -223 -1145
rect -65 -1179 -31 -1145
rect 127 -1179 161 -1145
rect 319 -1179 353 -1145
rect 511 -1179 545 -1145
rect 703 -1179 737 -1145
rect 895 -1179 929 -1145
rect 1087 -1179 1121 -1145
rect 1279 -1179 1313 -1145
rect -1409 -1287 -1375 -1253
rect -1217 -1287 -1183 -1253
rect -1025 -1287 -991 -1253
rect -833 -1287 -799 -1253
rect -641 -1287 -607 -1253
rect -449 -1287 -415 -1253
rect -257 -1287 -223 -1253
rect -65 -1287 -31 -1253
rect 127 -1287 161 -1253
rect 319 -1287 353 -1253
rect 511 -1287 545 -1253
rect 703 -1287 737 -1253
rect 895 -1287 929 -1253
rect 1087 -1287 1121 -1253
rect 1279 -1287 1313 -1253
rect -1457 -1703 -1423 -1337
rect -1361 -1703 -1327 -1337
rect -1265 -1703 -1231 -1337
rect -1169 -1703 -1135 -1337
rect -1073 -1703 -1039 -1337
rect -977 -1703 -943 -1337
rect -881 -1703 -847 -1337
rect -785 -1703 -751 -1337
rect -689 -1703 -655 -1337
rect -593 -1703 -559 -1337
rect -497 -1703 -463 -1337
rect -401 -1703 -367 -1337
rect -305 -1703 -271 -1337
rect -209 -1703 -175 -1337
rect -113 -1703 -79 -1337
rect -17 -1703 17 -1337
rect 79 -1703 113 -1337
rect 175 -1703 209 -1337
rect 271 -1703 305 -1337
rect 367 -1703 401 -1337
rect 463 -1703 497 -1337
rect 559 -1703 593 -1337
rect 655 -1703 689 -1337
rect 751 -1703 785 -1337
rect 847 -1703 881 -1337
rect 943 -1703 977 -1337
rect 1039 -1703 1073 -1337
rect 1135 -1703 1169 -1337
rect 1231 -1703 1265 -1337
rect 1327 -1703 1361 -1337
rect 1423 -1703 1457 -1337
rect -1313 -1787 -1279 -1753
rect -1121 -1787 -1087 -1753
rect -929 -1787 -895 -1753
rect -737 -1787 -703 -1753
rect -545 -1787 -511 -1753
rect -353 -1787 -319 -1753
rect -161 -1787 -127 -1753
rect 31 -1787 65 -1753
rect 223 -1787 257 -1753
rect 415 -1787 449 -1753
rect 607 -1787 641 -1753
rect 799 -1787 833 -1753
rect 991 -1787 1025 -1753
rect 1183 -1787 1217 -1753
rect 1375 -1787 1409 -1753
rect -1313 -1895 -1279 -1861
rect -1121 -1895 -1087 -1861
rect -929 -1895 -895 -1861
rect -737 -1895 -703 -1861
rect -545 -1895 -511 -1861
rect -353 -1895 -319 -1861
rect -161 -1895 -127 -1861
rect 31 -1895 65 -1861
rect 223 -1895 257 -1861
rect 415 -1895 449 -1861
rect 607 -1895 641 -1861
rect 799 -1895 833 -1861
rect 991 -1895 1025 -1861
rect 1183 -1895 1217 -1861
rect 1375 -1895 1409 -1861
rect -1457 -2311 -1423 -1945
rect -1361 -2311 -1327 -1945
rect -1265 -2311 -1231 -1945
rect -1169 -2311 -1135 -1945
rect -1073 -2311 -1039 -1945
rect -977 -2311 -943 -1945
rect -881 -2311 -847 -1945
rect -785 -2311 -751 -1945
rect -689 -2311 -655 -1945
rect -593 -2311 -559 -1945
rect -497 -2311 -463 -1945
rect -401 -2311 -367 -1945
rect -305 -2311 -271 -1945
rect -209 -2311 -175 -1945
rect -113 -2311 -79 -1945
rect -17 -2311 17 -1945
rect 79 -2311 113 -1945
rect 175 -2311 209 -1945
rect 271 -2311 305 -1945
rect 367 -2311 401 -1945
rect 463 -2311 497 -1945
rect 559 -2311 593 -1945
rect 655 -2311 689 -1945
rect 751 -2311 785 -1945
rect 847 -2311 881 -1945
rect 943 -2311 977 -1945
rect 1039 -2311 1073 -1945
rect 1135 -2311 1169 -1945
rect 1231 -2311 1265 -1945
rect 1327 -2311 1361 -1945
rect 1423 -2311 1457 -1945
rect -1409 -2395 -1375 -2361
rect -1217 -2395 -1183 -2361
rect -1025 -2395 -991 -2361
rect -833 -2395 -799 -2361
rect -641 -2395 -607 -2361
rect -449 -2395 -415 -2361
rect -257 -2395 -223 -2361
rect -65 -2395 -31 -2361
rect 127 -2395 161 -2361
rect 319 -2395 353 -2361
rect 511 -2395 545 -2361
rect 703 -2395 737 -2361
rect 895 -2395 929 -2361
rect 1087 -2395 1121 -2361
rect 1279 -2395 1313 -2361
<< metal1 >>
rect -1421 2395 -1363 2401
rect -1421 2361 -1409 2395
rect -1375 2361 -1363 2395
rect -1421 2355 -1363 2361
rect -1229 2395 -1171 2401
rect -1229 2361 -1217 2395
rect -1183 2361 -1171 2395
rect -1229 2355 -1171 2361
rect -1037 2395 -979 2401
rect -1037 2361 -1025 2395
rect -991 2361 -979 2395
rect -1037 2355 -979 2361
rect -845 2395 -787 2401
rect -845 2361 -833 2395
rect -799 2361 -787 2395
rect -845 2355 -787 2361
rect -653 2395 -595 2401
rect -653 2361 -641 2395
rect -607 2361 -595 2395
rect -653 2355 -595 2361
rect -461 2395 -403 2401
rect -461 2361 -449 2395
rect -415 2361 -403 2395
rect -461 2355 -403 2361
rect -269 2395 -211 2401
rect -269 2361 -257 2395
rect -223 2361 -211 2395
rect -269 2355 -211 2361
rect -77 2395 -19 2401
rect -77 2361 -65 2395
rect -31 2361 -19 2395
rect -77 2355 -19 2361
rect 115 2395 173 2401
rect 115 2361 127 2395
rect 161 2361 173 2395
rect 115 2355 173 2361
rect 307 2395 365 2401
rect 307 2361 319 2395
rect 353 2361 365 2395
rect 307 2355 365 2361
rect 499 2395 557 2401
rect 499 2361 511 2395
rect 545 2361 557 2395
rect 499 2355 557 2361
rect 691 2395 749 2401
rect 691 2361 703 2395
rect 737 2361 749 2395
rect 691 2355 749 2361
rect 883 2395 941 2401
rect 883 2361 895 2395
rect 929 2361 941 2395
rect 883 2355 941 2361
rect 1075 2395 1133 2401
rect 1075 2361 1087 2395
rect 1121 2361 1133 2395
rect 1075 2355 1133 2361
rect 1267 2395 1325 2401
rect 1267 2361 1279 2395
rect 1313 2361 1325 2395
rect 1267 2355 1325 2361
rect -1463 2311 -1417 2323
rect -1463 1945 -1457 2311
rect -1423 1945 -1417 2311
rect -1463 1933 -1417 1945
rect -1367 2311 -1321 2323
rect -1367 1945 -1361 2311
rect -1327 1945 -1321 2311
rect -1367 1933 -1321 1945
rect -1271 2311 -1225 2323
rect -1271 1945 -1265 2311
rect -1231 1945 -1225 2311
rect -1271 1933 -1225 1945
rect -1175 2311 -1129 2323
rect -1175 1945 -1169 2311
rect -1135 1945 -1129 2311
rect -1175 1933 -1129 1945
rect -1079 2311 -1033 2323
rect -1079 1945 -1073 2311
rect -1039 1945 -1033 2311
rect -1079 1933 -1033 1945
rect -983 2311 -937 2323
rect -983 1945 -977 2311
rect -943 1945 -937 2311
rect -983 1933 -937 1945
rect -887 2311 -841 2323
rect -887 1945 -881 2311
rect -847 1945 -841 2311
rect -887 1933 -841 1945
rect -791 2311 -745 2323
rect -791 1945 -785 2311
rect -751 1945 -745 2311
rect -791 1933 -745 1945
rect -695 2311 -649 2323
rect -695 1945 -689 2311
rect -655 1945 -649 2311
rect -695 1933 -649 1945
rect -599 2311 -553 2323
rect -599 1945 -593 2311
rect -559 1945 -553 2311
rect -599 1933 -553 1945
rect -503 2311 -457 2323
rect -503 1945 -497 2311
rect -463 1945 -457 2311
rect -503 1933 -457 1945
rect -407 2311 -361 2323
rect -407 1945 -401 2311
rect -367 1945 -361 2311
rect -407 1933 -361 1945
rect -311 2311 -265 2323
rect -311 1945 -305 2311
rect -271 1945 -265 2311
rect -311 1933 -265 1945
rect -215 2311 -169 2323
rect -215 1945 -209 2311
rect -175 1945 -169 2311
rect -215 1933 -169 1945
rect -119 2311 -73 2323
rect -119 1945 -113 2311
rect -79 1945 -73 2311
rect -119 1933 -73 1945
rect -23 2311 23 2323
rect -23 1945 -17 2311
rect 17 1945 23 2311
rect -23 1933 23 1945
rect 73 2311 119 2323
rect 73 1945 79 2311
rect 113 1945 119 2311
rect 73 1933 119 1945
rect 169 2311 215 2323
rect 169 1945 175 2311
rect 209 1945 215 2311
rect 169 1933 215 1945
rect 265 2311 311 2323
rect 265 1945 271 2311
rect 305 1945 311 2311
rect 265 1933 311 1945
rect 361 2311 407 2323
rect 361 1945 367 2311
rect 401 1945 407 2311
rect 361 1933 407 1945
rect 457 2311 503 2323
rect 457 1945 463 2311
rect 497 1945 503 2311
rect 457 1933 503 1945
rect 553 2311 599 2323
rect 553 1945 559 2311
rect 593 1945 599 2311
rect 553 1933 599 1945
rect 649 2311 695 2323
rect 649 1945 655 2311
rect 689 1945 695 2311
rect 649 1933 695 1945
rect 745 2311 791 2323
rect 745 1945 751 2311
rect 785 1945 791 2311
rect 745 1933 791 1945
rect 841 2311 887 2323
rect 841 1945 847 2311
rect 881 1945 887 2311
rect 841 1933 887 1945
rect 937 2311 983 2323
rect 937 1945 943 2311
rect 977 1945 983 2311
rect 937 1933 983 1945
rect 1033 2311 1079 2323
rect 1033 1945 1039 2311
rect 1073 1945 1079 2311
rect 1033 1933 1079 1945
rect 1129 2311 1175 2323
rect 1129 1945 1135 2311
rect 1169 1945 1175 2311
rect 1129 1933 1175 1945
rect 1225 2311 1271 2323
rect 1225 1945 1231 2311
rect 1265 1945 1271 2311
rect 1225 1933 1271 1945
rect 1321 2311 1367 2323
rect 1321 1945 1327 2311
rect 1361 1945 1367 2311
rect 1321 1933 1367 1945
rect 1417 2311 1463 2323
rect 1417 1945 1423 2311
rect 1457 1945 1463 2311
rect 1417 1933 1463 1945
rect -1325 1895 -1267 1901
rect -1325 1861 -1313 1895
rect -1279 1861 -1267 1895
rect -1325 1855 -1267 1861
rect -1133 1895 -1075 1901
rect -1133 1861 -1121 1895
rect -1087 1861 -1075 1895
rect -1133 1855 -1075 1861
rect -941 1895 -883 1901
rect -941 1861 -929 1895
rect -895 1861 -883 1895
rect -941 1855 -883 1861
rect -749 1895 -691 1901
rect -749 1861 -737 1895
rect -703 1861 -691 1895
rect -749 1855 -691 1861
rect -557 1895 -499 1901
rect -557 1861 -545 1895
rect -511 1861 -499 1895
rect -557 1855 -499 1861
rect -365 1895 -307 1901
rect -365 1861 -353 1895
rect -319 1861 -307 1895
rect -365 1855 -307 1861
rect -173 1895 -115 1901
rect -173 1861 -161 1895
rect -127 1861 -115 1895
rect -173 1855 -115 1861
rect 19 1895 77 1901
rect 19 1861 31 1895
rect 65 1861 77 1895
rect 19 1855 77 1861
rect 211 1895 269 1901
rect 211 1861 223 1895
rect 257 1861 269 1895
rect 211 1855 269 1861
rect 403 1895 461 1901
rect 403 1861 415 1895
rect 449 1861 461 1895
rect 403 1855 461 1861
rect 595 1895 653 1901
rect 595 1861 607 1895
rect 641 1861 653 1895
rect 595 1855 653 1861
rect 787 1895 845 1901
rect 787 1861 799 1895
rect 833 1861 845 1895
rect 787 1855 845 1861
rect 979 1895 1037 1901
rect 979 1861 991 1895
rect 1025 1861 1037 1895
rect 979 1855 1037 1861
rect 1171 1895 1229 1901
rect 1171 1861 1183 1895
rect 1217 1861 1229 1895
rect 1171 1855 1229 1861
rect 1363 1895 1421 1901
rect 1363 1861 1375 1895
rect 1409 1861 1421 1895
rect 1363 1855 1421 1861
rect -1325 1787 -1267 1793
rect -1325 1753 -1313 1787
rect -1279 1753 -1267 1787
rect -1325 1747 -1267 1753
rect -1133 1787 -1075 1793
rect -1133 1753 -1121 1787
rect -1087 1753 -1075 1787
rect -1133 1747 -1075 1753
rect -941 1787 -883 1793
rect -941 1753 -929 1787
rect -895 1753 -883 1787
rect -941 1747 -883 1753
rect -749 1787 -691 1793
rect -749 1753 -737 1787
rect -703 1753 -691 1787
rect -749 1747 -691 1753
rect -557 1787 -499 1793
rect -557 1753 -545 1787
rect -511 1753 -499 1787
rect -557 1747 -499 1753
rect -365 1787 -307 1793
rect -365 1753 -353 1787
rect -319 1753 -307 1787
rect -365 1747 -307 1753
rect -173 1787 -115 1793
rect -173 1753 -161 1787
rect -127 1753 -115 1787
rect -173 1747 -115 1753
rect 19 1787 77 1793
rect 19 1753 31 1787
rect 65 1753 77 1787
rect 19 1747 77 1753
rect 211 1787 269 1793
rect 211 1753 223 1787
rect 257 1753 269 1787
rect 211 1747 269 1753
rect 403 1787 461 1793
rect 403 1753 415 1787
rect 449 1753 461 1787
rect 403 1747 461 1753
rect 595 1787 653 1793
rect 595 1753 607 1787
rect 641 1753 653 1787
rect 595 1747 653 1753
rect 787 1787 845 1793
rect 787 1753 799 1787
rect 833 1753 845 1787
rect 787 1747 845 1753
rect 979 1787 1037 1793
rect 979 1753 991 1787
rect 1025 1753 1037 1787
rect 979 1747 1037 1753
rect 1171 1787 1229 1793
rect 1171 1753 1183 1787
rect 1217 1753 1229 1787
rect 1171 1747 1229 1753
rect 1363 1787 1421 1793
rect 1363 1753 1375 1787
rect 1409 1753 1421 1787
rect 1363 1747 1421 1753
rect -1463 1703 -1417 1715
rect -1463 1337 -1457 1703
rect -1423 1337 -1417 1703
rect -1463 1325 -1417 1337
rect -1367 1703 -1321 1715
rect -1367 1337 -1361 1703
rect -1327 1337 -1321 1703
rect -1367 1325 -1321 1337
rect -1271 1703 -1225 1715
rect -1271 1337 -1265 1703
rect -1231 1337 -1225 1703
rect -1271 1325 -1225 1337
rect -1175 1703 -1129 1715
rect -1175 1337 -1169 1703
rect -1135 1337 -1129 1703
rect -1175 1325 -1129 1337
rect -1079 1703 -1033 1715
rect -1079 1337 -1073 1703
rect -1039 1337 -1033 1703
rect -1079 1325 -1033 1337
rect -983 1703 -937 1715
rect -983 1337 -977 1703
rect -943 1337 -937 1703
rect -983 1325 -937 1337
rect -887 1703 -841 1715
rect -887 1337 -881 1703
rect -847 1337 -841 1703
rect -887 1325 -841 1337
rect -791 1703 -745 1715
rect -791 1337 -785 1703
rect -751 1337 -745 1703
rect -791 1325 -745 1337
rect -695 1703 -649 1715
rect -695 1337 -689 1703
rect -655 1337 -649 1703
rect -695 1325 -649 1337
rect -599 1703 -553 1715
rect -599 1337 -593 1703
rect -559 1337 -553 1703
rect -599 1325 -553 1337
rect -503 1703 -457 1715
rect -503 1337 -497 1703
rect -463 1337 -457 1703
rect -503 1325 -457 1337
rect -407 1703 -361 1715
rect -407 1337 -401 1703
rect -367 1337 -361 1703
rect -407 1325 -361 1337
rect -311 1703 -265 1715
rect -311 1337 -305 1703
rect -271 1337 -265 1703
rect -311 1325 -265 1337
rect -215 1703 -169 1715
rect -215 1337 -209 1703
rect -175 1337 -169 1703
rect -215 1325 -169 1337
rect -119 1703 -73 1715
rect -119 1337 -113 1703
rect -79 1337 -73 1703
rect -119 1325 -73 1337
rect -23 1703 23 1715
rect -23 1337 -17 1703
rect 17 1337 23 1703
rect -23 1325 23 1337
rect 73 1703 119 1715
rect 73 1337 79 1703
rect 113 1337 119 1703
rect 73 1325 119 1337
rect 169 1703 215 1715
rect 169 1337 175 1703
rect 209 1337 215 1703
rect 169 1325 215 1337
rect 265 1703 311 1715
rect 265 1337 271 1703
rect 305 1337 311 1703
rect 265 1325 311 1337
rect 361 1703 407 1715
rect 361 1337 367 1703
rect 401 1337 407 1703
rect 361 1325 407 1337
rect 457 1703 503 1715
rect 457 1337 463 1703
rect 497 1337 503 1703
rect 457 1325 503 1337
rect 553 1703 599 1715
rect 553 1337 559 1703
rect 593 1337 599 1703
rect 553 1325 599 1337
rect 649 1703 695 1715
rect 649 1337 655 1703
rect 689 1337 695 1703
rect 649 1325 695 1337
rect 745 1703 791 1715
rect 745 1337 751 1703
rect 785 1337 791 1703
rect 745 1325 791 1337
rect 841 1703 887 1715
rect 841 1337 847 1703
rect 881 1337 887 1703
rect 841 1325 887 1337
rect 937 1703 983 1715
rect 937 1337 943 1703
rect 977 1337 983 1703
rect 937 1325 983 1337
rect 1033 1703 1079 1715
rect 1033 1337 1039 1703
rect 1073 1337 1079 1703
rect 1033 1325 1079 1337
rect 1129 1703 1175 1715
rect 1129 1337 1135 1703
rect 1169 1337 1175 1703
rect 1129 1325 1175 1337
rect 1225 1703 1271 1715
rect 1225 1337 1231 1703
rect 1265 1337 1271 1703
rect 1225 1325 1271 1337
rect 1321 1703 1367 1715
rect 1321 1337 1327 1703
rect 1361 1337 1367 1703
rect 1321 1325 1367 1337
rect 1417 1703 1463 1715
rect 1417 1337 1423 1703
rect 1457 1337 1463 1703
rect 1417 1325 1463 1337
rect -1421 1287 -1363 1293
rect -1421 1253 -1409 1287
rect -1375 1253 -1363 1287
rect -1421 1247 -1363 1253
rect -1229 1287 -1171 1293
rect -1229 1253 -1217 1287
rect -1183 1253 -1171 1287
rect -1229 1247 -1171 1253
rect -1037 1287 -979 1293
rect -1037 1253 -1025 1287
rect -991 1253 -979 1287
rect -1037 1247 -979 1253
rect -845 1287 -787 1293
rect -845 1253 -833 1287
rect -799 1253 -787 1287
rect -845 1247 -787 1253
rect -653 1287 -595 1293
rect -653 1253 -641 1287
rect -607 1253 -595 1287
rect -653 1247 -595 1253
rect -461 1287 -403 1293
rect -461 1253 -449 1287
rect -415 1253 -403 1287
rect -461 1247 -403 1253
rect -269 1287 -211 1293
rect -269 1253 -257 1287
rect -223 1253 -211 1287
rect -269 1247 -211 1253
rect -77 1287 -19 1293
rect -77 1253 -65 1287
rect -31 1253 -19 1287
rect -77 1247 -19 1253
rect 115 1287 173 1293
rect 115 1253 127 1287
rect 161 1253 173 1287
rect 115 1247 173 1253
rect 307 1287 365 1293
rect 307 1253 319 1287
rect 353 1253 365 1287
rect 307 1247 365 1253
rect 499 1287 557 1293
rect 499 1253 511 1287
rect 545 1253 557 1287
rect 499 1247 557 1253
rect 691 1287 749 1293
rect 691 1253 703 1287
rect 737 1253 749 1287
rect 691 1247 749 1253
rect 883 1287 941 1293
rect 883 1253 895 1287
rect 929 1253 941 1287
rect 883 1247 941 1253
rect 1075 1287 1133 1293
rect 1075 1253 1087 1287
rect 1121 1253 1133 1287
rect 1075 1247 1133 1253
rect 1267 1287 1325 1293
rect 1267 1253 1279 1287
rect 1313 1253 1325 1287
rect 1267 1247 1325 1253
rect -1421 1179 -1363 1185
rect -1421 1145 -1409 1179
rect -1375 1145 -1363 1179
rect -1421 1139 -1363 1145
rect -1229 1179 -1171 1185
rect -1229 1145 -1217 1179
rect -1183 1145 -1171 1179
rect -1229 1139 -1171 1145
rect -1037 1179 -979 1185
rect -1037 1145 -1025 1179
rect -991 1145 -979 1179
rect -1037 1139 -979 1145
rect -845 1179 -787 1185
rect -845 1145 -833 1179
rect -799 1145 -787 1179
rect -845 1139 -787 1145
rect -653 1179 -595 1185
rect -653 1145 -641 1179
rect -607 1145 -595 1179
rect -653 1139 -595 1145
rect -461 1179 -403 1185
rect -461 1145 -449 1179
rect -415 1145 -403 1179
rect -461 1139 -403 1145
rect -269 1179 -211 1185
rect -269 1145 -257 1179
rect -223 1145 -211 1179
rect -269 1139 -211 1145
rect -77 1179 -19 1185
rect -77 1145 -65 1179
rect -31 1145 -19 1179
rect -77 1139 -19 1145
rect 115 1179 173 1185
rect 115 1145 127 1179
rect 161 1145 173 1179
rect 115 1139 173 1145
rect 307 1179 365 1185
rect 307 1145 319 1179
rect 353 1145 365 1179
rect 307 1139 365 1145
rect 499 1179 557 1185
rect 499 1145 511 1179
rect 545 1145 557 1179
rect 499 1139 557 1145
rect 691 1179 749 1185
rect 691 1145 703 1179
rect 737 1145 749 1179
rect 691 1139 749 1145
rect 883 1179 941 1185
rect 883 1145 895 1179
rect 929 1145 941 1179
rect 883 1139 941 1145
rect 1075 1179 1133 1185
rect 1075 1145 1087 1179
rect 1121 1145 1133 1179
rect 1075 1139 1133 1145
rect 1267 1179 1325 1185
rect 1267 1145 1279 1179
rect 1313 1145 1325 1179
rect 1267 1139 1325 1145
rect -1463 1095 -1417 1107
rect -1463 729 -1457 1095
rect -1423 729 -1417 1095
rect -1463 717 -1417 729
rect -1367 1095 -1321 1107
rect -1367 729 -1361 1095
rect -1327 729 -1321 1095
rect -1367 717 -1321 729
rect -1271 1095 -1225 1107
rect -1271 729 -1265 1095
rect -1231 729 -1225 1095
rect -1271 717 -1225 729
rect -1175 1095 -1129 1107
rect -1175 729 -1169 1095
rect -1135 729 -1129 1095
rect -1175 717 -1129 729
rect -1079 1095 -1033 1107
rect -1079 729 -1073 1095
rect -1039 729 -1033 1095
rect -1079 717 -1033 729
rect -983 1095 -937 1107
rect -983 729 -977 1095
rect -943 729 -937 1095
rect -983 717 -937 729
rect -887 1095 -841 1107
rect -887 729 -881 1095
rect -847 729 -841 1095
rect -887 717 -841 729
rect -791 1095 -745 1107
rect -791 729 -785 1095
rect -751 729 -745 1095
rect -791 717 -745 729
rect -695 1095 -649 1107
rect -695 729 -689 1095
rect -655 729 -649 1095
rect -695 717 -649 729
rect -599 1095 -553 1107
rect -599 729 -593 1095
rect -559 729 -553 1095
rect -599 717 -553 729
rect -503 1095 -457 1107
rect -503 729 -497 1095
rect -463 729 -457 1095
rect -503 717 -457 729
rect -407 1095 -361 1107
rect -407 729 -401 1095
rect -367 729 -361 1095
rect -407 717 -361 729
rect -311 1095 -265 1107
rect -311 729 -305 1095
rect -271 729 -265 1095
rect -311 717 -265 729
rect -215 1095 -169 1107
rect -215 729 -209 1095
rect -175 729 -169 1095
rect -215 717 -169 729
rect -119 1095 -73 1107
rect -119 729 -113 1095
rect -79 729 -73 1095
rect -119 717 -73 729
rect -23 1095 23 1107
rect -23 729 -17 1095
rect 17 729 23 1095
rect -23 717 23 729
rect 73 1095 119 1107
rect 73 729 79 1095
rect 113 729 119 1095
rect 73 717 119 729
rect 169 1095 215 1107
rect 169 729 175 1095
rect 209 729 215 1095
rect 169 717 215 729
rect 265 1095 311 1107
rect 265 729 271 1095
rect 305 729 311 1095
rect 265 717 311 729
rect 361 1095 407 1107
rect 361 729 367 1095
rect 401 729 407 1095
rect 361 717 407 729
rect 457 1095 503 1107
rect 457 729 463 1095
rect 497 729 503 1095
rect 457 717 503 729
rect 553 1095 599 1107
rect 553 729 559 1095
rect 593 729 599 1095
rect 553 717 599 729
rect 649 1095 695 1107
rect 649 729 655 1095
rect 689 729 695 1095
rect 649 717 695 729
rect 745 1095 791 1107
rect 745 729 751 1095
rect 785 729 791 1095
rect 745 717 791 729
rect 841 1095 887 1107
rect 841 729 847 1095
rect 881 729 887 1095
rect 841 717 887 729
rect 937 1095 983 1107
rect 937 729 943 1095
rect 977 729 983 1095
rect 937 717 983 729
rect 1033 1095 1079 1107
rect 1033 729 1039 1095
rect 1073 729 1079 1095
rect 1033 717 1079 729
rect 1129 1095 1175 1107
rect 1129 729 1135 1095
rect 1169 729 1175 1095
rect 1129 717 1175 729
rect 1225 1095 1271 1107
rect 1225 729 1231 1095
rect 1265 729 1271 1095
rect 1225 717 1271 729
rect 1321 1095 1367 1107
rect 1321 729 1327 1095
rect 1361 729 1367 1095
rect 1321 717 1367 729
rect 1417 1095 1463 1107
rect 1417 729 1423 1095
rect 1457 729 1463 1095
rect 1417 717 1463 729
rect -1325 679 -1267 685
rect -1325 645 -1313 679
rect -1279 645 -1267 679
rect -1325 639 -1267 645
rect -1133 679 -1075 685
rect -1133 645 -1121 679
rect -1087 645 -1075 679
rect -1133 639 -1075 645
rect -941 679 -883 685
rect -941 645 -929 679
rect -895 645 -883 679
rect -941 639 -883 645
rect -749 679 -691 685
rect -749 645 -737 679
rect -703 645 -691 679
rect -749 639 -691 645
rect -557 679 -499 685
rect -557 645 -545 679
rect -511 645 -499 679
rect -557 639 -499 645
rect -365 679 -307 685
rect -365 645 -353 679
rect -319 645 -307 679
rect -365 639 -307 645
rect -173 679 -115 685
rect -173 645 -161 679
rect -127 645 -115 679
rect -173 639 -115 645
rect 19 679 77 685
rect 19 645 31 679
rect 65 645 77 679
rect 19 639 77 645
rect 211 679 269 685
rect 211 645 223 679
rect 257 645 269 679
rect 211 639 269 645
rect 403 679 461 685
rect 403 645 415 679
rect 449 645 461 679
rect 403 639 461 645
rect 595 679 653 685
rect 595 645 607 679
rect 641 645 653 679
rect 595 639 653 645
rect 787 679 845 685
rect 787 645 799 679
rect 833 645 845 679
rect 787 639 845 645
rect 979 679 1037 685
rect 979 645 991 679
rect 1025 645 1037 679
rect 979 639 1037 645
rect 1171 679 1229 685
rect 1171 645 1183 679
rect 1217 645 1229 679
rect 1171 639 1229 645
rect 1363 679 1421 685
rect 1363 645 1375 679
rect 1409 645 1421 679
rect 1363 639 1421 645
rect -1325 571 -1267 577
rect -1325 537 -1313 571
rect -1279 537 -1267 571
rect -1325 531 -1267 537
rect -1133 571 -1075 577
rect -1133 537 -1121 571
rect -1087 537 -1075 571
rect -1133 531 -1075 537
rect -941 571 -883 577
rect -941 537 -929 571
rect -895 537 -883 571
rect -941 531 -883 537
rect -749 571 -691 577
rect -749 537 -737 571
rect -703 537 -691 571
rect -749 531 -691 537
rect -557 571 -499 577
rect -557 537 -545 571
rect -511 537 -499 571
rect -557 531 -499 537
rect -365 571 -307 577
rect -365 537 -353 571
rect -319 537 -307 571
rect -365 531 -307 537
rect -173 571 -115 577
rect -173 537 -161 571
rect -127 537 -115 571
rect -173 531 -115 537
rect 19 571 77 577
rect 19 537 31 571
rect 65 537 77 571
rect 19 531 77 537
rect 211 571 269 577
rect 211 537 223 571
rect 257 537 269 571
rect 211 531 269 537
rect 403 571 461 577
rect 403 537 415 571
rect 449 537 461 571
rect 403 531 461 537
rect 595 571 653 577
rect 595 537 607 571
rect 641 537 653 571
rect 595 531 653 537
rect 787 571 845 577
rect 787 537 799 571
rect 833 537 845 571
rect 787 531 845 537
rect 979 571 1037 577
rect 979 537 991 571
rect 1025 537 1037 571
rect 979 531 1037 537
rect 1171 571 1229 577
rect 1171 537 1183 571
rect 1217 537 1229 571
rect 1171 531 1229 537
rect 1363 571 1421 577
rect 1363 537 1375 571
rect 1409 537 1421 571
rect 1363 531 1421 537
rect -1463 487 -1417 499
rect -1463 121 -1457 487
rect -1423 121 -1417 487
rect -1463 109 -1417 121
rect -1367 487 -1321 499
rect -1367 121 -1361 487
rect -1327 121 -1321 487
rect -1367 109 -1321 121
rect -1271 487 -1225 499
rect -1271 121 -1265 487
rect -1231 121 -1225 487
rect -1271 109 -1225 121
rect -1175 487 -1129 499
rect -1175 121 -1169 487
rect -1135 121 -1129 487
rect -1175 109 -1129 121
rect -1079 487 -1033 499
rect -1079 121 -1073 487
rect -1039 121 -1033 487
rect -1079 109 -1033 121
rect -983 487 -937 499
rect -983 121 -977 487
rect -943 121 -937 487
rect -983 109 -937 121
rect -887 487 -841 499
rect -887 121 -881 487
rect -847 121 -841 487
rect -887 109 -841 121
rect -791 487 -745 499
rect -791 121 -785 487
rect -751 121 -745 487
rect -791 109 -745 121
rect -695 487 -649 499
rect -695 121 -689 487
rect -655 121 -649 487
rect -695 109 -649 121
rect -599 487 -553 499
rect -599 121 -593 487
rect -559 121 -553 487
rect -599 109 -553 121
rect -503 487 -457 499
rect -503 121 -497 487
rect -463 121 -457 487
rect -503 109 -457 121
rect -407 487 -361 499
rect -407 121 -401 487
rect -367 121 -361 487
rect -407 109 -361 121
rect -311 487 -265 499
rect -311 121 -305 487
rect -271 121 -265 487
rect -311 109 -265 121
rect -215 487 -169 499
rect -215 121 -209 487
rect -175 121 -169 487
rect -215 109 -169 121
rect -119 487 -73 499
rect -119 121 -113 487
rect -79 121 -73 487
rect -119 109 -73 121
rect -23 487 23 499
rect -23 121 -17 487
rect 17 121 23 487
rect -23 109 23 121
rect 73 487 119 499
rect 73 121 79 487
rect 113 121 119 487
rect 73 109 119 121
rect 169 487 215 499
rect 169 121 175 487
rect 209 121 215 487
rect 169 109 215 121
rect 265 487 311 499
rect 265 121 271 487
rect 305 121 311 487
rect 265 109 311 121
rect 361 487 407 499
rect 361 121 367 487
rect 401 121 407 487
rect 361 109 407 121
rect 457 487 503 499
rect 457 121 463 487
rect 497 121 503 487
rect 457 109 503 121
rect 553 487 599 499
rect 553 121 559 487
rect 593 121 599 487
rect 553 109 599 121
rect 649 487 695 499
rect 649 121 655 487
rect 689 121 695 487
rect 649 109 695 121
rect 745 487 791 499
rect 745 121 751 487
rect 785 121 791 487
rect 745 109 791 121
rect 841 487 887 499
rect 841 121 847 487
rect 881 121 887 487
rect 841 109 887 121
rect 937 487 983 499
rect 937 121 943 487
rect 977 121 983 487
rect 937 109 983 121
rect 1033 487 1079 499
rect 1033 121 1039 487
rect 1073 121 1079 487
rect 1033 109 1079 121
rect 1129 487 1175 499
rect 1129 121 1135 487
rect 1169 121 1175 487
rect 1129 109 1175 121
rect 1225 487 1271 499
rect 1225 121 1231 487
rect 1265 121 1271 487
rect 1225 109 1271 121
rect 1321 487 1367 499
rect 1321 121 1327 487
rect 1361 121 1367 487
rect 1321 109 1367 121
rect 1417 487 1463 499
rect 1417 121 1423 487
rect 1457 121 1463 487
rect 1417 109 1463 121
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect -1463 -121 -1417 -109
rect -1463 -487 -1457 -121
rect -1423 -487 -1417 -121
rect -1463 -499 -1417 -487
rect -1367 -121 -1321 -109
rect -1367 -487 -1361 -121
rect -1327 -487 -1321 -121
rect -1367 -499 -1321 -487
rect -1271 -121 -1225 -109
rect -1271 -487 -1265 -121
rect -1231 -487 -1225 -121
rect -1271 -499 -1225 -487
rect -1175 -121 -1129 -109
rect -1175 -487 -1169 -121
rect -1135 -487 -1129 -121
rect -1175 -499 -1129 -487
rect -1079 -121 -1033 -109
rect -1079 -487 -1073 -121
rect -1039 -487 -1033 -121
rect -1079 -499 -1033 -487
rect -983 -121 -937 -109
rect -983 -487 -977 -121
rect -943 -487 -937 -121
rect -983 -499 -937 -487
rect -887 -121 -841 -109
rect -887 -487 -881 -121
rect -847 -487 -841 -121
rect -887 -499 -841 -487
rect -791 -121 -745 -109
rect -791 -487 -785 -121
rect -751 -487 -745 -121
rect -791 -499 -745 -487
rect -695 -121 -649 -109
rect -695 -487 -689 -121
rect -655 -487 -649 -121
rect -695 -499 -649 -487
rect -599 -121 -553 -109
rect -599 -487 -593 -121
rect -559 -487 -553 -121
rect -599 -499 -553 -487
rect -503 -121 -457 -109
rect -503 -487 -497 -121
rect -463 -487 -457 -121
rect -503 -499 -457 -487
rect -407 -121 -361 -109
rect -407 -487 -401 -121
rect -367 -487 -361 -121
rect -407 -499 -361 -487
rect -311 -121 -265 -109
rect -311 -487 -305 -121
rect -271 -487 -265 -121
rect -311 -499 -265 -487
rect -215 -121 -169 -109
rect -215 -487 -209 -121
rect -175 -487 -169 -121
rect -215 -499 -169 -487
rect -119 -121 -73 -109
rect -119 -487 -113 -121
rect -79 -487 -73 -121
rect -119 -499 -73 -487
rect -23 -121 23 -109
rect -23 -487 -17 -121
rect 17 -487 23 -121
rect -23 -499 23 -487
rect 73 -121 119 -109
rect 73 -487 79 -121
rect 113 -487 119 -121
rect 73 -499 119 -487
rect 169 -121 215 -109
rect 169 -487 175 -121
rect 209 -487 215 -121
rect 169 -499 215 -487
rect 265 -121 311 -109
rect 265 -487 271 -121
rect 305 -487 311 -121
rect 265 -499 311 -487
rect 361 -121 407 -109
rect 361 -487 367 -121
rect 401 -487 407 -121
rect 361 -499 407 -487
rect 457 -121 503 -109
rect 457 -487 463 -121
rect 497 -487 503 -121
rect 457 -499 503 -487
rect 553 -121 599 -109
rect 553 -487 559 -121
rect 593 -487 599 -121
rect 553 -499 599 -487
rect 649 -121 695 -109
rect 649 -487 655 -121
rect 689 -487 695 -121
rect 649 -499 695 -487
rect 745 -121 791 -109
rect 745 -487 751 -121
rect 785 -487 791 -121
rect 745 -499 791 -487
rect 841 -121 887 -109
rect 841 -487 847 -121
rect 881 -487 887 -121
rect 841 -499 887 -487
rect 937 -121 983 -109
rect 937 -487 943 -121
rect 977 -487 983 -121
rect 937 -499 983 -487
rect 1033 -121 1079 -109
rect 1033 -487 1039 -121
rect 1073 -487 1079 -121
rect 1033 -499 1079 -487
rect 1129 -121 1175 -109
rect 1129 -487 1135 -121
rect 1169 -487 1175 -121
rect 1129 -499 1175 -487
rect 1225 -121 1271 -109
rect 1225 -487 1231 -121
rect 1265 -487 1271 -121
rect 1225 -499 1271 -487
rect 1321 -121 1367 -109
rect 1321 -487 1327 -121
rect 1361 -487 1367 -121
rect 1321 -499 1367 -487
rect 1417 -121 1463 -109
rect 1417 -487 1423 -121
rect 1457 -487 1463 -121
rect 1417 -499 1463 -487
rect -1325 -537 -1267 -531
rect -1325 -571 -1313 -537
rect -1279 -571 -1267 -537
rect -1325 -577 -1267 -571
rect -1133 -537 -1075 -531
rect -1133 -571 -1121 -537
rect -1087 -571 -1075 -537
rect -1133 -577 -1075 -571
rect -941 -537 -883 -531
rect -941 -571 -929 -537
rect -895 -571 -883 -537
rect -941 -577 -883 -571
rect -749 -537 -691 -531
rect -749 -571 -737 -537
rect -703 -571 -691 -537
rect -749 -577 -691 -571
rect -557 -537 -499 -531
rect -557 -571 -545 -537
rect -511 -571 -499 -537
rect -557 -577 -499 -571
rect -365 -537 -307 -531
rect -365 -571 -353 -537
rect -319 -571 -307 -537
rect -365 -577 -307 -571
rect -173 -537 -115 -531
rect -173 -571 -161 -537
rect -127 -571 -115 -537
rect -173 -577 -115 -571
rect 19 -537 77 -531
rect 19 -571 31 -537
rect 65 -571 77 -537
rect 19 -577 77 -571
rect 211 -537 269 -531
rect 211 -571 223 -537
rect 257 -571 269 -537
rect 211 -577 269 -571
rect 403 -537 461 -531
rect 403 -571 415 -537
rect 449 -571 461 -537
rect 403 -577 461 -571
rect 595 -537 653 -531
rect 595 -571 607 -537
rect 641 -571 653 -537
rect 595 -577 653 -571
rect 787 -537 845 -531
rect 787 -571 799 -537
rect 833 -571 845 -537
rect 787 -577 845 -571
rect 979 -537 1037 -531
rect 979 -571 991 -537
rect 1025 -571 1037 -537
rect 979 -577 1037 -571
rect 1171 -537 1229 -531
rect 1171 -571 1183 -537
rect 1217 -571 1229 -537
rect 1171 -577 1229 -571
rect 1363 -537 1421 -531
rect 1363 -571 1375 -537
rect 1409 -571 1421 -537
rect 1363 -577 1421 -571
rect -1325 -645 -1267 -639
rect -1325 -679 -1313 -645
rect -1279 -679 -1267 -645
rect -1325 -685 -1267 -679
rect -1133 -645 -1075 -639
rect -1133 -679 -1121 -645
rect -1087 -679 -1075 -645
rect -1133 -685 -1075 -679
rect -941 -645 -883 -639
rect -941 -679 -929 -645
rect -895 -679 -883 -645
rect -941 -685 -883 -679
rect -749 -645 -691 -639
rect -749 -679 -737 -645
rect -703 -679 -691 -645
rect -749 -685 -691 -679
rect -557 -645 -499 -639
rect -557 -679 -545 -645
rect -511 -679 -499 -645
rect -557 -685 -499 -679
rect -365 -645 -307 -639
rect -365 -679 -353 -645
rect -319 -679 -307 -645
rect -365 -685 -307 -679
rect -173 -645 -115 -639
rect -173 -679 -161 -645
rect -127 -679 -115 -645
rect -173 -685 -115 -679
rect 19 -645 77 -639
rect 19 -679 31 -645
rect 65 -679 77 -645
rect 19 -685 77 -679
rect 211 -645 269 -639
rect 211 -679 223 -645
rect 257 -679 269 -645
rect 211 -685 269 -679
rect 403 -645 461 -639
rect 403 -679 415 -645
rect 449 -679 461 -645
rect 403 -685 461 -679
rect 595 -645 653 -639
rect 595 -679 607 -645
rect 641 -679 653 -645
rect 595 -685 653 -679
rect 787 -645 845 -639
rect 787 -679 799 -645
rect 833 -679 845 -645
rect 787 -685 845 -679
rect 979 -645 1037 -639
rect 979 -679 991 -645
rect 1025 -679 1037 -645
rect 979 -685 1037 -679
rect 1171 -645 1229 -639
rect 1171 -679 1183 -645
rect 1217 -679 1229 -645
rect 1171 -685 1229 -679
rect 1363 -645 1421 -639
rect 1363 -679 1375 -645
rect 1409 -679 1421 -645
rect 1363 -685 1421 -679
rect -1463 -729 -1417 -717
rect -1463 -1095 -1457 -729
rect -1423 -1095 -1417 -729
rect -1463 -1107 -1417 -1095
rect -1367 -729 -1321 -717
rect -1367 -1095 -1361 -729
rect -1327 -1095 -1321 -729
rect -1367 -1107 -1321 -1095
rect -1271 -729 -1225 -717
rect -1271 -1095 -1265 -729
rect -1231 -1095 -1225 -729
rect -1271 -1107 -1225 -1095
rect -1175 -729 -1129 -717
rect -1175 -1095 -1169 -729
rect -1135 -1095 -1129 -729
rect -1175 -1107 -1129 -1095
rect -1079 -729 -1033 -717
rect -1079 -1095 -1073 -729
rect -1039 -1095 -1033 -729
rect -1079 -1107 -1033 -1095
rect -983 -729 -937 -717
rect -983 -1095 -977 -729
rect -943 -1095 -937 -729
rect -983 -1107 -937 -1095
rect -887 -729 -841 -717
rect -887 -1095 -881 -729
rect -847 -1095 -841 -729
rect -887 -1107 -841 -1095
rect -791 -729 -745 -717
rect -791 -1095 -785 -729
rect -751 -1095 -745 -729
rect -791 -1107 -745 -1095
rect -695 -729 -649 -717
rect -695 -1095 -689 -729
rect -655 -1095 -649 -729
rect -695 -1107 -649 -1095
rect -599 -729 -553 -717
rect -599 -1095 -593 -729
rect -559 -1095 -553 -729
rect -599 -1107 -553 -1095
rect -503 -729 -457 -717
rect -503 -1095 -497 -729
rect -463 -1095 -457 -729
rect -503 -1107 -457 -1095
rect -407 -729 -361 -717
rect -407 -1095 -401 -729
rect -367 -1095 -361 -729
rect -407 -1107 -361 -1095
rect -311 -729 -265 -717
rect -311 -1095 -305 -729
rect -271 -1095 -265 -729
rect -311 -1107 -265 -1095
rect -215 -729 -169 -717
rect -215 -1095 -209 -729
rect -175 -1095 -169 -729
rect -215 -1107 -169 -1095
rect -119 -729 -73 -717
rect -119 -1095 -113 -729
rect -79 -1095 -73 -729
rect -119 -1107 -73 -1095
rect -23 -729 23 -717
rect -23 -1095 -17 -729
rect 17 -1095 23 -729
rect -23 -1107 23 -1095
rect 73 -729 119 -717
rect 73 -1095 79 -729
rect 113 -1095 119 -729
rect 73 -1107 119 -1095
rect 169 -729 215 -717
rect 169 -1095 175 -729
rect 209 -1095 215 -729
rect 169 -1107 215 -1095
rect 265 -729 311 -717
rect 265 -1095 271 -729
rect 305 -1095 311 -729
rect 265 -1107 311 -1095
rect 361 -729 407 -717
rect 361 -1095 367 -729
rect 401 -1095 407 -729
rect 361 -1107 407 -1095
rect 457 -729 503 -717
rect 457 -1095 463 -729
rect 497 -1095 503 -729
rect 457 -1107 503 -1095
rect 553 -729 599 -717
rect 553 -1095 559 -729
rect 593 -1095 599 -729
rect 553 -1107 599 -1095
rect 649 -729 695 -717
rect 649 -1095 655 -729
rect 689 -1095 695 -729
rect 649 -1107 695 -1095
rect 745 -729 791 -717
rect 745 -1095 751 -729
rect 785 -1095 791 -729
rect 745 -1107 791 -1095
rect 841 -729 887 -717
rect 841 -1095 847 -729
rect 881 -1095 887 -729
rect 841 -1107 887 -1095
rect 937 -729 983 -717
rect 937 -1095 943 -729
rect 977 -1095 983 -729
rect 937 -1107 983 -1095
rect 1033 -729 1079 -717
rect 1033 -1095 1039 -729
rect 1073 -1095 1079 -729
rect 1033 -1107 1079 -1095
rect 1129 -729 1175 -717
rect 1129 -1095 1135 -729
rect 1169 -1095 1175 -729
rect 1129 -1107 1175 -1095
rect 1225 -729 1271 -717
rect 1225 -1095 1231 -729
rect 1265 -1095 1271 -729
rect 1225 -1107 1271 -1095
rect 1321 -729 1367 -717
rect 1321 -1095 1327 -729
rect 1361 -1095 1367 -729
rect 1321 -1107 1367 -1095
rect 1417 -729 1463 -717
rect 1417 -1095 1423 -729
rect 1457 -1095 1463 -729
rect 1417 -1107 1463 -1095
rect -1421 -1145 -1363 -1139
rect -1421 -1179 -1409 -1145
rect -1375 -1179 -1363 -1145
rect -1421 -1185 -1363 -1179
rect -1229 -1145 -1171 -1139
rect -1229 -1179 -1217 -1145
rect -1183 -1179 -1171 -1145
rect -1229 -1185 -1171 -1179
rect -1037 -1145 -979 -1139
rect -1037 -1179 -1025 -1145
rect -991 -1179 -979 -1145
rect -1037 -1185 -979 -1179
rect -845 -1145 -787 -1139
rect -845 -1179 -833 -1145
rect -799 -1179 -787 -1145
rect -845 -1185 -787 -1179
rect -653 -1145 -595 -1139
rect -653 -1179 -641 -1145
rect -607 -1179 -595 -1145
rect -653 -1185 -595 -1179
rect -461 -1145 -403 -1139
rect -461 -1179 -449 -1145
rect -415 -1179 -403 -1145
rect -461 -1185 -403 -1179
rect -269 -1145 -211 -1139
rect -269 -1179 -257 -1145
rect -223 -1179 -211 -1145
rect -269 -1185 -211 -1179
rect -77 -1145 -19 -1139
rect -77 -1179 -65 -1145
rect -31 -1179 -19 -1145
rect -77 -1185 -19 -1179
rect 115 -1145 173 -1139
rect 115 -1179 127 -1145
rect 161 -1179 173 -1145
rect 115 -1185 173 -1179
rect 307 -1145 365 -1139
rect 307 -1179 319 -1145
rect 353 -1179 365 -1145
rect 307 -1185 365 -1179
rect 499 -1145 557 -1139
rect 499 -1179 511 -1145
rect 545 -1179 557 -1145
rect 499 -1185 557 -1179
rect 691 -1145 749 -1139
rect 691 -1179 703 -1145
rect 737 -1179 749 -1145
rect 691 -1185 749 -1179
rect 883 -1145 941 -1139
rect 883 -1179 895 -1145
rect 929 -1179 941 -1145
rect 883 -1185 941 -1179
rect 1075 -1145 1133 -1139
rect 1075 -1179 1087 -1145
rect 1121 -1179 1133 -1145
rect 1075 -1185 1133 -1179
rect 1267 -1145 1325 -1139
rect 1267 -1179 1279 -1145
rect 1313 -1179 1325 -1145
rect 1267 -1185 1325 -1179
rect -1421 -1253 -1363 -1247
rect -1421 -1287 -1409 -1253
rect -1375 -1287 -1363 -1253
rect -1421 -1293 -1363 -1287
rect -1229 -1253 -1171 -1247
rect -1229 -1287 -1217 -1253
rect -1183 -1287 -1171 -1253
rect -1229 -1293 -1171 -1287
rect -1037 -1253 -979 -1247
rect -1037 -1287 -1025 -1253
rect -991 -1287 -979 -1253
rect -1037 -1293 -979 -1287
rect -845 -1253 -787 -1247
rect -845 -1287 -833 -1253
rect -799 -1287 -787 -1253
rect -845 -1293 -787 -1287
rect -653 -1253 -595 -1247
rect -653 -1287 -641 -1253
rect -607 -1287 -595 -1253
rect -653 -1293 -595 -1287
rect -461 -1253 -403 -1247
rect -461 -1287 -449 -1253
rect -415 -1287 -403 -1253
rect -461 -1293 -403 -1287
rect -269 -1253 -211 -1247
rect -269 -1287 -257 -1253
rect -223 -1287 -211 -1253
rect -269 -1293 -211 -1287
rect -77 -1253 -19 -1247
rect -77 -1287 -65 -1253
rect -31 -1287 -19 -1253
rect -77 -1293 -19 -1287
rect 115 -1253 173 -1247
rect 115 -1287 127 -1253
rect 161 -1287 173 -1253
rect 115 -1293 173 -1287
rect 307 -1253 365 -1247
rect 307 -1287 319 -1253
rect 353 -1287 365 -1253
rect 307 -1293 365 -1287
rect 499 -1253 557 -1247
rect 499 -1287 511 -1253
rect 545 -1287 557 -1253
rect 499 -1293 557 -1287
rect 691 -1253 749 -1247
rect 691 -1287 703 -1253
rect 737 -1287 749 -1253
rect 691 -1293 749 -1287
rect 883 -1253 941 -1247
rect 883 -1287 895 -1253
rect 929 -1287 941 -1253
rect 883 -1293 941 -1287
rect 1075 -1253 1133 -1247
rect 1075 -1287 1087 -1253
rect 1121 -1287 1133 -1253
rect 1075 -1293 1133 -1287
rect 1267 -1253 1325 -1247
rect 1267 -1287 1279 -1253
rect 1313 -1287 1325 -1253
rect 1267 -1293 1325 -1287
rect -1463 -1337 -1417 -1325
rect -1463 -1703 -1457 -1337
rect -1423 -1703 -1417 -1337
rect -1463 -1715 -1417 -1703
rect -1367 -1337 -1321 -1325
rect -1367 -1703 -1361 -1337
rect -1327 -1703 -1321 -1337
rect -1367 -1715 -1321 -1703
rect -1271 -1337 -1225 -1325
rect -1271 -1703 -1265 -1337
rect -1231 -1703 -1225 -1337
rect -1271 -1715 -1225 -1703
rect -1175 -1337 -1129 -1325
rect -1175 -1703 -1169 -1337
rect -1135 -1703 -1129 -1337
rect -1175 -1715 -1129 -1703
rect -1079 -1337 -1033 -1325
rect -1079 -1703 -1073 -1337
rect -1039 -1703 -1033 -1337
rect -1079 -1715 -1033 -1703
rect -983 -1337 -937 -1325
rect -983 -1703 -977 -1337
rect -943 -1703 -937 -1337
rect -983 -1715 -937 -1703
rect -887 -1337 -841 -1325
rect -887 -1703 -881 -1337
rect -847 -1703 -841 -1337
rect -887 -1715 -841 -1703
rect -791 -1337 -745 -1325
rect -791 -1703 -785 -1337
rect -751 -1703 -745 -1337
rect -791 -1715 -745 -1703
rect -695 -1337 -649 -1325
rect -695 -1703 -689 -1337
rect -655 -1703 -649 -1337
rect -695 -1715 -649 -1703
rect -599 -1337 -553 -1325
rect -599 -1703 -593 -1337
rect -559 -1703 -553 -1337
rect -599 -1715 -553 -1703
rect -503 -1337 -457 -1325
rect -503 -1703 -497 -1337
rect -463 -1703 -457 -1337
rect -503 -1715 -457 -1703
rect -407 -1337 -361 -1325
rect -407 -1703 -401 -1337
rect -367 -1703 -361 -1337
rect -407 -1715 -361 -1703
rect -311 -1337 -265 -1325
rect -311 -1703 -305 -1337
rect -271 -1703 -265 -1337
rect -311 -1715 -265 -1703
rect -215 -1337 -169 -1325
rect -215 -1703 -209 -1337
rect -175 -1703 -169 -1337
rect -215 -1715 -169 -1703
rect -119 -1337 -73 -1325
rect -119 -1703 -113 -1337
rect -79 -1703 -73 -1337
rect -119 -1715 -73 -1703
rect -23 -1337 23 -1325
rect -23 -1703 -17 -1337
rect 17 -1703 23 -1337
rect -23 -1715 23 -1703
rect 73 -1337 119 -1325
rect 73 -1703 79 -1337
rect 113 -1703 119 -1337
rect 73 -1715 119 -1703
rect 169 -1337 215 -1325
rect 169 -1703 175 -1337
rect 209 -1703 215 -1337
rect 169 -1715 215 -1703
rect 265 -1337 311 -1325
rect 265 -1703 271 -1337
rect 305 -1703 311 -1337
rect 265 -1715 311 -1703
rect 361 -1337 407 -1325
rect 361 -1703 367 -1337
rect 401 -1703 407 -1337
rect 361 -1715 407 -1703
rect 457 -1337 503 -1325
rect 457 -1703 463 -1337
rect 497 -1703 503 -1337
rect 457 -1715 503 -1703
rect 553 -1337 599 -1325
rect 553 -1703 559 -1337
rect 593 -1703 599 -1337
rect 553 -1715 599 -1703
rect 649 -1337 695 -1325
rect 649 -1703 655 -1337
rect 689 -1703 695 -1337
rect 649 -1715 695 -1703
rect 745 -1337 791 -1325
rect 745 -1703 751 -1337
rect 785 -1703 791 -1337
rect 745 -1715 791 -1703
rect 841 -1337 887 -1325
rect 841 -1703 847 -1337
rect 881 -1703 887 -1337
rect 841 -1715 887 -1703
rect 937 -1337 983 -1325
rect 937 -1703 943 -1337
rect 977 -1703 983 -1337
rect 937 -1715 983 -1703
rect 1033 -1337 1079 -1325
rect 1033 -1703 1039 -1337
rect 1073 -1703 1079 -1337
rect 1033 -1715 1079 -1703
rect 1129 -1337 1175 -1325
rect 1129 -1703 1135 -1337
rect 1169 -1703 1175 -1337
rect 1129 -1715 1175 -1703
rect 1225 -1337 1271 -1325
rect 1225 -1703 1231 -1337
rect 1265 -1703 1271 -1337
rect 1225 -1715 1271 -1703
rect 1321 -1337 1367 -1325
rect 1321 -1703 1327 -1337
rect 1361 -1703 1367 -1337
rect 1321 -1715 1367 -1703
rect 1417 -1337 1463 -1325
rect 1417 -1703 1423 -1337
rect 1457 -1703 1463 -1337
rect 1417 -1715 1463 -1703
rect -1325 -1753 -1267 -1747
rect -1325 -1787 -1313 -1753
rect -1279 -1787 -1267 -1753
rect -1325 -1793 -1267 -1787
rect -1133 -1753 -1075 -1747
rect -1133 -1787 -1121 -1753
rect -1087 -1787 -1075 -1753
rect -1133 -1793 -1075 -1787
rect -941 -1753 -883 -1747
rect -941 -1787 -929 -1753
rect -895 -1787 -883 -1753
rect -941 -1793 -883 -1787
rect -749 -1753 -691 -1747
rect -749 -1787 -737 -1753
rect -703 -1787 -691 -1753
rect -749 -1793 -691 -1787
rect -557 -1753 -499 -1747
rect -557 -1787 -545 -1753
rect -511 -1787 -499 -1753
rect -557 -1793 -499 -1787
rect -365 -1753 -307 -1747
rect -365 -1787 -353 -1753
rect -319 -1787 -307 -1753
rect -365 -1793 -307 -1787
rect -173 -1753 -115 -1747
rect -173 -1787 -161 -1753
rect -127 -1787 -115 -1753
rect -173 -1793 -115 -1787
rect 19 -1753 77 -1747
rect 19 -1787 31 -1753
rect 65 -1787 77 -1753
rect 19 -1793 77 -1787
rect 211 -1753 269 -1747
rect 211 -1787 223 -1753
rect 257 -1787 269 -1753
rect 211 -1793 269 -1787
rect 403 -1753 461 -1747
rect 403 -1787 415 -1753
rect 449 -1787 461 -1753
rect 403 -1793 461 -1787
rect 595 -1753 653 -1747
rect 595 -1787 607 -1753
rect 641 -1787 653 -1753
rect 595 -1793 653 -1787
rect 787 -1753 845 -1747
rect 787 -1787 799 -1753
rect 833 -1787 845 -1753
rect 787 -1793 845 -1787
rect 979 -1753 1037 -1747
rect 979 -1787 991 -1753
rect 1025 -1787 1037 -1753
rect 979 -1793 1037 -1787
rect 1171 -1753 1229 -1747
rect 1171 -1787 1183 -1753
rect 1217 -1787 1229 -1753
rect 1171 -1793 1229 -1787
rect 1363 -1753 1421 -1747
rect 1363 -1787 1375 -1753
rect 1409 -1787 1421 -1753
rect 1363 -1793 1421 -1787
rect -1325 -1861 -1267 -1855
rect -1325 -1895 -1313 -1861
rect -1279 -1895 -1267 -1861
rect -1325 -1901 -1267 -1895
rect -1133 -1861 -1075 -1855
rect -1133 -1895 -1121 -1861
rect -1087 -1895 -1075 -1861
rect -1133 -1901 -1075 -1895
rect -941 -1861 -883 -1855
rect -941 -1895 -929 -1861
rect -895 -1895 -883 -1861
rect -941 -1901 -883 -1895
rect -749 -1861 -691 -1855
rect -749 -1895 -737 -1861
rect -703 -1895 -691 -1861
rect -749 -1901 -691 -1895
rect -557 -1861 -499 -1855
rect -557 -1895 -545 -1861
rect -511 -1895 -499 -1861
rect -557 -1901 -499 -1895
rect -365 -1861 -307 -1855
rect -365 -1895 -353 -1861
rect -319 -1895 -307 -1861
rect -365 -1901 -307 -1895
rect -173 -1861 -115 -1855
rect -173 -1895 -161 -1861
rect -127 -1895 -115 -1861
rect -173 -1901 -115 -1895
rect 19 -1861 77 -1855
rect 19 -1895 31 -1861
rect 65 -1895 77 -1861
rect 19 -1901 77 -1895
rect 211 -1861 269 -1855
rect 211 -1895 223 -1861
rect 257 -1895 269 -1861
rect 211 -1901 269 -1895
rect 403 -1861 461 -1855
rect 403 -1895 415 -1861
rect 449 -1895 461 -1861
rect 403 -1901 461 -1895
rect 595 -1861 653 -1855
rect 595 -1895 607 -1861
rect 641 -1895 653 -1861
rect 595 -1901 653 -1895
rect 787 -1861 845 -1855
rect 787 -1895 799 -1861
rect 833 -1895 845 -1861
rect 787 -1901 845 -1895
rect 979 -1861 1037 -1855
rect 979 -1895 991 -1861
rect 1025 -1895 1037 -1861
rect 979 -1901 1037 -1895
rect 1171 -1861 1229 -1855
rect 1171 -1895 1183 -1861
rect 1217 -1895 1229 -1861
rect 1171 -1901 1229 -1895
rect 1363 -1861 1421 -1855
rect 1363 -1895 1375 -1861
rect 1409 -1895 1421 -1861
rect 1363 -1901 1421 -1895
rect -1463 -1945 -1417 -1933
rect -1463 -2311 -1457 -1945
rect -1423 -2311 -1417 -1945
rect -1463 -2323 -1417 -2311
rect -1367 -1945 -1321 -1933
rect -1367 -2311 -1361 -1945
rect -1327 -2311 -1321 -1945
rect -1367 -2323 -1321 -2311
rect -1271 -1945 -1225 -1933
rect -1271 -2311 -1265 -1945
rect -1231 -2311 -1225 -1945
rect -1271 -2323 -1225 -2311
rect -1175 -1945 -1129 -1933
rect -1175 -2311 -1169 -1945
rect -1135 -2311 -1129 -1945
rect -1175 -2323 -1129 -2311
rect -1079 -1945 -1033 -1933
rect -1079 -2311 -1073 -1945
rect -1039 -2311 -1033 -1945
rect -1079 -2323 -1033 -2311
rect -983 -1945 -937 -1933
rect -983 -2311 -977 -1945
rect -943 -2311 -937 -1945
rect -983 -2323 -937 -2311
rect -887 -1945 -841 -1933
rect -887 -2311 -881 -1945
rect -847 -2311 -841 -1945
rect -887 -2323 -841 -2311
rect -791 -1945 -745 -1933
rect -791 -2311 -785 -1945
rect -751 -2311 -745 -1945
rect -791 -2323 -745 -2311
rect -695 -1945 -649 -1933
rect -695 -2311 -689 -1945
rect -655 -2311 -649 -1945
rect -695 -2323 -649 -2311
rect -599 -1945 -553 -1933
rect -599 -2311 -593 -1945
rect -559 -2311 -553 -1945
rect -599 -2323 -553 -2311
rect -503 -1945 -457 -1933
rect -503 -2311 -497 -1945
rect -463 -2311 -457 -1945
rect -503 -2323 -457 -2311
rect -407 -1945 -361 -1933
rect -407 -2311 -401 -1945
rect -367 -2311 -361 -1945
rect -407 -2323 -361 -2311
rect -311 -1945 -265 -1933
rect -311 -2311 -305 -1945
rect -271 -2311 -265 -1945
rect -311 -2323 -265 -2311
rect -215 -1945 -169 -1933
rect -215 -2311 -209 -1945
rect -175 -2311 -169 -1945
rect -215 -2323 -169 -2311
rect -119 -1945 -73 -1933
rect -119 -2311 -113 -1945
rect -79 -2311 -73 -1945
rect -119 -2323 -73 -2311
rect -23 -1945 23 -1933
rect -23 -2311 -17 -1945
rect 17 -2311 23 -1945
rect -23 -2323 23 -2311
rect 73 -1945 119 -1933
rect 73 -2311 79 -1945
rect 113 -2311 119 -1945
rect 73 -2323 119 -2311
rect 169 -1945 215 -1933
rect 169 -2311 175 -1945
rect 209 -2311 215 -1945
rect 169 -2323 215 -2311
rect 265 -1945 311 -1933
rect 265 -2311 271 -1945
rect 305 -2311 311 -1945
rect 265 -2323 311 -2311
rect 361 -1945 407 -1933
rect 361 -2311 367 -1945
rect 401 -2311 407 -1945
rect 361 -2323 407 -2311
rect 457 -1945 503 -1933
rect 457 -2311 463 -1945
rect 497 -2311 503 -1945
rect 457 -2323 503 -2311
rect 553 -1945 599 -1933
rect 553 -2311 559 -1945
rect 593 -2311 599 -1945
rect 553 -2323 599 -2311
rect 649 -1945 695 -1933
rect 649 -2311 655 -1945
rect 689 -2311 695 -1945
rect 649 -2323 695 -2311
rect 745 -1945 791 -1933
rect 745 -2311 751 -1945
rect 785 -2311 791 -1945
rect 745 -2323 791 -2311
rect 841 -1945 887 -1933
rect 841 -2311 847 -1945
rect 881 -2311 887 -1945
rect 841 -2323 887 -2311
rect 937 -1945 983 -1933
rect 937 -2311 943 -1945
rect 977 -2311 983 -1945
rect 937 -2323 983 -2311
rect 1033 -1945 1079 -1933
rect 1033 -2311 1039 -1945
rect 1073 -2311 1079 -1945
rect 1033 -2323 1079 -2311
rect 1129 -1945 1175 -1933
rect 1129 -2311 1135 -1945
rect 1169 -2311 1175 -1945
rect 1129 -2323 1175 -2311
rect 1225 -1945 1271 -1933
rect 1225 -2311 1231 -1945
rect 1265 -2311 1271 -1945
rect 1225 -2323 1271 -2311
rect 1321 -1945 1367 -1933
rect 1321 -2311 1327 -1945
rect 1361 -2311 1367 -1945
rect 1321 -2323 1367 -2311
rect 1417 -1945 1463 -1933
rect 1417 -2311 1423 -1945
rect 1457 -2311 1463 -1945
rect 1417 -2323 1463 -2311
rect -1421 -2361 -1363 -2355
rect -1421 -2395 -1409 -2361
rect -1375 -2395 -1363 -2361
rect -1421 -2401 -1363 -2395
rect -1229 -2361 -1171 -2355
rect -1229 -2395 -1217 -2361
rect -1183 -2395 -1171 -2361
rect -1229 -2401 -1171 -2395
rect -1037 -2361 -979 -2355
rect -1037 -2395 -1025 -2361
rect -991 -2395 -979 -2361
rect -1037 -2401 -979 -2395
rect -845 -2361 -787 -2355
rect -845 -2395 -833 -2361
rect -799 -2395 -787 -2361
rect -845 -2401 -787 -2395
rect -653 -2361 -595 -2355
rect -653 -2395 -641 -2361
rect -607 -2395 -595 -2361
rect -653 -2401 -595 -2395
rect -461 -2361 -403 -2355
rect -461 -2395 -449 -2361
rect -415 -2395 -403 -2361
rect -461 -2401 -403 -2395
rect -269 -2361 -211 -2355
rect -269 -2395 -257 -2361
rect -223 -2395 -211 -2361
rect -269 -2401 -211 -2395
rect -77 -2361 -19 -2355
rect -77 -2395 -65 -2361
rect -31 -2395 -19 -2361
rect -77 -2401 -19 -2395
rect 115 -2361 173 -2355
rect 115 -2395 127 -2361
rect 161 -2395 173 -2361
rect 115 -2401 173 -2395
rect 307 -2361 365 -2355
rect 307 -2395 319 -2361
rect 353 -2395 365 -2361
rect 307 -2401 365 -2395
rect 499 -2361 557 -2355
rect 499 -2395 511 -2361
rect 545 -2395 557 -2361
rect 499 -2401 557 -2395
rect 691 -2361 749 -2355
rect 691 -2395 703 -2361
rect 737 -2395 749 -2361
rect 691 -2401 749 -2395
rect 883 -2361 941 -2355
rect 883 -2395 895 -2361
rect 929 -2395 941 -2361
rect 883 -2401 941 -2395
rect 1075 -2361 1133 -2355
rect 1075 -2395 1087 -2361
rect 1121 -2395 1133 -2361
rect 1075 -2401 1133 -2395
rect 1267 -2361 1325 -2355
rect 1267 -2395 1279 -2361
rect 1313 -2395 1325 -2361
rect 1267 -2401 1325 -2395
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1554 -2480 1554 2480
string parameters w 1.95 l 0.150 m 8 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
