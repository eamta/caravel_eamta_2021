magic
tech sky130A
magscale 1 2
timestamp 1622937437
<< error_p >>
rect -927 1131 -865 1137
rect -799 1131 -737 1137
rect -671 1131 -609 1137
rect -543 1131 -481 1137
rect -415 1131 -353 1137
rect -287 1131 -225 1137
rect -159 1131 -97 1137
rect -31 1131 31 1137
rect 97 1131 159 1137
rect 225 1131 287 1137
rect 353 1131 415 1137
rect 481 1131 543 1137
rect 609 1131 671 1137
rect 737 1131 799 1137
rect 865 1131 927 1137
rect -927 1097 -915 1131
rect -799 1097 -787 1131
rect -671 1097 -659 1131
rect -543 1097 -531 1131
rect -415 1097 -403 1131
rect -287 1097 -275 1131
rect -159 1097 -147 1131
rect -31 1097 -19 1131
rect 97 1097 109 1131
rect 225 1097 237 1131
rect 353 1097 365 1131
rect 481 1097 493 1131
rect 609 1097 621 1131
rect 737 1097 749 1131
rect 865 1097 877 1131
rect -927 1091 -865 1097
rect -799 1091 -737 1097
rect -671 1091 -609 1097
rect -543 1091 -481 1097
rect -415 1091 -353 1097
rect -287 1091 -225 1097
rect -159 1091 -97 1097
rect -31 1091 31 1097
rect 97 1091 159 1097
rect 225 1091 287 1097
rect 353 1091 415 1097
rect 481 1091 543 1097
rect 609 1091 671 1097
rect 737 1091 799 1097
rect 865 1091 927 1097
rect -927 -1097 -865 -1091
rect -799 -1097 -737 -1091
rect -671 -1097 -609 -1091
rect -543 -1097 -481 -1091
rect -415 -1097 -353 -1091
rect -287 -1097 -225 -1091
rect -159 -1097 -97 -1091
rect -31 -1097 31 -1091
rect 97 -1097 159 -1091
rect 225 -1097 287 -1091
rect 353 -1097 415 -1091
rect 481 -1097 543 -1091
rect 609 -1097 671 -1091
rect 737 -1097 799 -1091
rect 865 -1097 927 -1091
rect -927 -1131 -915 -1097
rect -799 -1131 -787 -1097
rect -671 -1131 -659 -1097
rect -543 -1131 -531 -1097
rect -415 -1131 -403 -1097
rect -287 -1131 -275 -1097
rect -159 -1131 -147 -1097
rect -31 -1131 -19 -1097
rect 97 -1131 109 -1097
rect 225 -1131 237 -1097
rect 353 -1131 365 -1097
rect 481 -1131 493 -1097
rect 609 -1131 621 -1097
rect 737 -1131 749 -1097
rect 865 -1131 877 -1097
rect -927 -1137 -865 -1131
rect -799 -1137 -737 -1131
rect -671 -1137 -609 -1131
rect -543 -1137 -481 -1131
rect -415 -1137 -353 -1131
rect -287 -1137 -225 -1131
rect -159 -1137 -97 -1131
rect -31 -1137 31 -1131
rect 97 -1137 159 -1131
rect 225 -1137 287 -1131
rect 353 -1137 415 -1131
rect 481 -1137 543 -1131
rect 609 -1137 671 -1131
rect 737 -1137 799 -1131
rect 865 -1137 927 -1131
<< nwell >>
rect -1127 -1269 1127 1269
<< pmos >>
rect -931 -1050 -861 1050
rect -803 -1050 -733 1050
rect -675 -1050 -605 1050
rect -547 -1050 -477 1050
rect -419 -1050 -349 1050
rect -291 -1050 -221 1050
rect -163 -1050 -93 1050
rect -35 -1050 35 1050
rect 93 -1050 163 1050
rect 221 -1050 291 1050
rect 349 -1050 419 1050
rect 477 -1050 547 1050
rect 605 -1050 675 1050
rect 733 -1050 803 1050
rect 861 -1050 931 1050
<< pdiff >>
rect -989 1038 -931 1050
rect -989 -1038 -977 1038
rect -943 -1038 -931 1038
rect -989 -1050 -931 -1038
rect -861 1038 -803 1050
rect -861 -1038 -849 1038
rect -815 -1038 -803 1038
rect -861 -1050 -803 -1038
rect -733 1038 -675 1050
rect -733 -1038 -721 1038
rect -687 -1038 -675 1038
rect -733 -1050 -675 -1038
rect -605 1038 -547 1050
rect -605 -1038 -593 1038
rect -559 -1038 -547 1038
rect -605 -1050 -547 -1038
rect -477 1038 -419 1050
rect -477 -1038 -465 1038
rect -431 -1038 -419 1038
rect -477 -1050 -419 -1038
rect -349 1038 -291 1050
rect -349 -1038 -337 1038
rect -303 -1038 -291 1038
rect -349 -1050 -291 -1038
rect -221 1038 -163 1050
rect -221 -1038 -209 1038
rect -175 -1038 -163 1038
rect -221 -1050 -163 -1038
rect -93 1038 -35 1050
rect -93 -1038 -81 1038
rect -47 -1038 -35 1038
rect -93 -1050 -35 -1038
rect 35 1038 93 1050
rect 35 -1038 47 1038
rect 81 -1038 93 1038
rect 35 -1050 93 -1038
rect 163 1038 221 1050
rect 163 -1038 175 1038
rect 209 -1038 221 1038
rect 163 -1050 221 -1038
rect 291 1038 349 1050
rect 291 -1038 303 1038
rect 337 -1038 349 1038
rect 291 -1050 349 -1038
rect 419 1038 477 1050
rect 419 -1038 431 1038
rect 465 -1038 477 1038
rect 419 -1050 477 -1038
rect 547 1038 605 1050
rect 547 -1038 559 1038
rect 593 -1038 605 1038
rect 547 -1050 605 -1038
rect 675 1038 733 1050
rect 675 -1038 687 1038
rect 721 -1038 733 1038
rect 675 -1050 733 -1038
rect 803 1038 861 1050
rect 803 -1038 815 1038
rect 849 -1038 861 1038
rect 803 -1050 861 -1038
rect 931 1038 989 1050
rect 931 -1038 943 1038
rect 977 -1038 989 1038
rect 931 -1050 989 -1038
<< pdiffc >>
rect -977 -1038 -943 1038
rect -849 -1038 -815 1038
rect -721 -1038 -687 1038
rect -593 -1038 -559 1038
rect -465 -1038 -431 1038
rect -337 -1038 -303 1038
rect -209 -1038 -175 1038
rect -81 -1038 -47 1038
rect 47 -1038 81 1038
rect 175 -1038 209 1038
rect 303 -1038 337 1038
rect 431 -1038 465 1038
rect 559 -1038 593 1038
rect 687 -1038 721 1038
rect 815 -1038 849 1038
rect 943 -1038 977 1038
<< nsubdiff >>
rect -1091 1199 -995 1233
rect 995 1199 1091 1233
rect -1091 1137 -1057 1199
rect 1057 1137 1091 1199
rect -1091 -1199 -1057 -1137
rect 1057 -1199 1091 -1137
rect -1091 -1233 -995 -1199
rect 995 -1233 1091 -1199
<< nsubdiffcont >>
rect -995 1199 995 1233
rect -1091 -1137 -1057 1137
rect 1057 -1137 1091 1137
rect -995 -1233 995 -1199
<< poly >>
rect -931 1131 -861 1147
rect -931 1097 -915 1131
rect -877 1097 -861 1131
rect -931 1050 -861 1097
rect -803 1131 -733 1147
rect -803 1097 -787 1131
rect -749 1097 -733 1131
rect -803 1050 -733 1097
rect -675 1131 -605 1147
rect -675 1097 -659 1131
rect -621 1097 -605 1131
rect -675 1050 -605 1097
rect -547 1131 -477 1147
rect -547 1097 -531 1131
rect -493 1097 -477 1131
rect -547 1050 -477 1097
rect -419 1131 -349 1147
rect -419 1097 -403 1131
rect -365 1097 -349 1131
rect -419 1050 -349 1097
rect -291 1131 -221 1147
rect -291 1097 -275 1131
rect -237 1097 -221 1131
rect -291 1050 -221 1097
rect -163 1131 -93 1147
rect -163 1097 -147 1131
rect -109 1097 -93 1131
rect -163 1050 -93 1097
rect -35 1131 35 1147
rect -35 1097 -19 1131
rect 19 1097 35 1131
rect -35 1050 35 1097
rect 93 1131 163 1147
rect 93 1097 109 1131
rect 147 1097 163 1131
rect 93 1050 163 1097
rect 221 1131 291 1147
rect 221 1097 237 1131
rect 275 1097 291 1131
rect 221 1050 291 1097
rect 349 1131 419 1147
rect 349 1097 365 1131
rect 403 1097 419 1131
rect 349 1050 419 1097
rect 477 1131 547 1147
rect 477 1097 493 1131
rect 531 1097 547 1131
rect 477 1050 547 1097
rect 605 1131 675 1147
rect 605 1097 621 1131
rect 659 1097 675 1131
rect 605 1050 675 1097
rect 733 1131 803 1147
rect 733 1097 749 1131
rect 787 1097 803 1131
rect 733 1050 803 1097
rect 861 1131 931 1147
rect 861 1097 877 1131
rect 915 1097 931 1131
rect 861 1050 931 1097
rect -931 -1097 -861 -1050
rect -931 -1131 -915 -1097
rect -877 -1131 -861 -1097
rect -931 -1147 -861 -1131
rect -803 -1097 -733 -1050
rect -803 -1131 -787 -1097
rect -749 -1131 -733 -1097
rect -803 -1147 -733 -1131
rect -675 -1097 -605 -1050
rect -675 -1131 -659 -1097
rect -621 -1131 -605 -1097
rect -675 -1147 -605 -1131
rect -547 -1097 -477 -1050
rect -547 -1131 -531 -1097
rect -493 -1131 -477 -1097
rect -547 -1147 -477 -1131
rect -419 -1097 -349 -1050
rect -419 -1131 -403 -1097
rect -365 -1131 -349 -1097
rect -419 -1147 -349 -1131
rect -291 -1097 -221 -1050
rect -291 -1131 -275 -1097
rect -237 -1131 -221 -1097
rect -291 -1147 -221 -1131
rect -163 -1097 -93 -1050
rect -163 -1131 -147 -1097
rect -109 -1131 -93 -1097
rect -163 -1147 -93 -1131
rect -35 -1097 35 -1050
rect -35 -1131 -19 -1097
rect 19 -1131 35 -1097
rect -35 -1147 35 -1131
rect 93 -1097 163 -1050
rect 93 -1131 109 -1097
rect 147 -1131 163 -1097
rect 93 -1147 163 -1131
rect 221 -1097 291 -1050
rect 221 -1131 237 -1097
rect 275 -1131 291 -1097
rect 221 -1147 291 -1131
rect 349 -1097 419 -1050
rect 349 -1131 365 -1097
rect 403 -1131 419 -1097
rect 349 -1147 419 -1131
rect 477 -1097 547 -1050
rect 477 -1131 493 -1097
rect 531 -1131 547 -1097
rect 477 -1147 547 -1131
rect 605 -1097 675 -1050
rect 605 -1131 621 -1097
rect 659 -1131 675 -1097
rect 605 -1147 675 -1131
rect 733 -1097 803 -1050
rect 733 -1131 749 -1097
rect 787 -1131 803 -1097
rect 733 -1147 803 -1131
rect 861 -1097 931 -1050
rect 861 -1131 877 -1097
rect 915 -1131 931 -1097
rect 861 -1147 931 -1131
<< polycont >>
rect -915 1097 -877 1131
rect -787 1097 -749 1131
rect -659 1097 -621 1131
rect -531 1097 -493 1131
rect -403 1097 -365 1131
rect -275 1097 -237 1131
rect -147 1097 -109 1131
rect -19 1097 19 1131
rect 109 1097 147 1131
rect 237 1097 275 1131
rect 365 1097 403 1131
rect 493 1097 531 1131
rect 621 1097 659 1131
rect 749 1097 787 1131
rect 877 1097 915 1131
rect -915 -1131 -877 -1097
rect -787 -1131 -749 -1097
rect -659 -1131 -621 -1097
rect -531 -1131 -493 -1097
rect -403 -1131 -365 -1097
rect -275 -1131 -237 -1097
rect -147 -1131 -109 -1097
rect -19 -1131 19 -1097
rect 109 -1131 147 -1097
rect 237 -1131 275 -1097
rect 365 -1131 403 -1097
rect 493 -1131 531 -1097
rect 621 -1131 659 -1097
rect 749 -1131 787 -1097
rect 877 -1131 915 -1097
<< locali >>
rect -1091 1199 -995 1233
rect 995 1199 1091 1233
rect -1091 1137 -1057 1199
rect 1057 1137 1091 1199
rect -931 1097 -915 1131
rect -877 1097 -861 1131
rect -803 1097 -787 1131
rect -749 1097 -733 1131
rect -675 1097 -659 1131
rect -621 1097 -605 1131
rect -547 1097 -531 1131
rect -493 1097 -477 1131
rect -419 1097 -403 1131
rect -365 1097 -349 1131
rect -291 1097 -275 1131
rect -237 1097 -221 1131
rect -163 1097 -147 1131
rect -109 1097 -93 1131
rect -35 1097 -19 1131
rect 19 1097 35 1131
rect 93 1097 109 1131
rect 147 1097 163 1131
rect 221 1097 237 1131
rect 275 1097 291 1131
rect 349 1097 365 1131
rect 403 1097 419 1131
rect 477 1097 493 1131
rect 531 1097 547 1131
rect 605 1097 621 1131
rect 659 1097 675 1131
rect 733 1097 749 1131
rect 787 1097 803 1131
rect 861 1097 877 1131
rect 915 1097 931 1131
rect -977 1038 -943 1054
rect -977 -1054 -943 -1038
rect -849 1038 -815 1054
rect -849 -1054 -815 -1038
rect -721 1038 -687 1054
rect -721 -1054 -687 -1038
rect -593 1038 -559 1054
rect -593 -1054 -559 -1038
rect -465 1038 -431 1054
rect -465 -1054 -431 -1038
rect -337 1038 -303 1054
rect -337 -1054 -303 -1038
rect -209 1038 -175 1054
rect -209 -1054 -175 -1038
rect -81 1038 -47 1054
rect -81 -1054 -47 -1038
rect 47 1038 81 1054
rect 47 -1054 81 -1038
rect 175 1038 209 1054
rect 175 -1054 209 -1038
rect 303 1038 337 1054
rect 303 -1054 337 -1038
rect 431 1038 465 1054
rect 431 -1054 465 -1038
rect 559 1038 593 1054
rect 559 -1054 593 -1038
rect 687 1038 721 1054
rect 687 -1054 721 -1038
rect 815 1038 849 1054
rect 815 -1054 849 -1038
rect 943 1038 977 1054
rect 943 -1054 977 -1038
rect -931 -1131 -915 -1097
rect -877 -1131 -861 -1097
rect -803 -1131 -787 -1097
rect -749 -1131 -733 -1097
rect -675 -1131 -659 -1097
rect -621 -1131 -605 -1097
rect -547 -1131 -531 -1097
rect -493 -1131 -477 -1097
rect -419 -1131 -403 -1097
rect -365 -1131 -349 -1097
rect -291 -1131 -275 -1097
rect -237 -1131 -221 -1097
rect -163 -1131 -147 -1097
rect -109 -1131 -93 -1097
rect -35 -1131 -19 -1097
rect 19 -1131 35 -1097
rect 93 -1131 109 -1097
rect 147 -1131 163 -1097
rect 221 -1131 237 -1097
rect 275 -1131 291 -1097
rect 349 -1131 365 -1097
rect 403 -1131 419 -1097
rect 477 -1131 493 -1097
rect 531 -1131 547 -1097
rect 605 -1131 621 -1097
rect 659 -1131 675 -1097
rect 733 -1131 749 -1097
rect 787 -1131 803 -1097
rect 861 -1131 877 -1097
rect 915 -1131 931 -1097
rect -1091 -1199 -1057 -1137
rect 1057 -1199 1091 -1137
rect -1091 -1233 -995 -1199
rect 995 -1233 1091 -1199
<< viali >>
rect -915 1097 -877 1131
rect -787 1097 -749 1131
rect -659 1097 -621 1131
rect -531 1097 -493 1131
rect -403 1097 -365 1131
rect -275 1097 -237 1131
rect -147 1097 -109 1131
rect -19 1097 19 1131
rect 109 1097 147 1131
rect 237 1097 275 1131
rect 365 1097 403 1131
rect 493 1097 531 1131
rect 621 1097 659 1131
rect 749 1097 787 1131
rect 877 1097 915 1131
rect -977 -1038 -943 1038
rect -849 -1038 -815 1038
rect -721 -1038 -687 1038
rect -593 -1038 -559 1038
rect -465 -1038 -431 1038
rect -337 -1038 -303 1038
rect -209 -1038 -175 1038
rect -81 -1038 -47 1038
rect 47 -1038 81 1038
rect 175 -1038 209 1038
rect 303 -1038 337 1038
rect 431 -1038 465 1038
rect 559 -1038 593 1038
rect 687 -1038 721 1038
rect 815 -1038 849 1038
rect 943 -1038 977 1038
rect -915 -1131 -877 -1097
rect -787 -1131 -749 -1097
rect -659 -1131 -621 -1097
rect -531 -1131 -493 -1097
rect -403 -1131 -365 -1097
rect -275 -1131 -237 -1097
rect -147 -1131 -109 -1097
rect -19 -1131 19 -1097
rect 109 -1131 147 -1097
rect 237 -1131 275 -1097
rect 365 -1131 403 -1097
rect 493 -1131 531 -1097
rect 621 -1131 659 -1097
rect 749 -1131 787 -1097
rect 877 -1131 915 -1097
<< metal1 >>
rect -927 1131 -865 1137
rect -927 1097 -915 1131
rect -877 1097 -865 1131
rect -927 1091 -865 1097
rect -799 1131 -737 1137
rect -799 1097 -787 1131
rect -749 1097 -737 1131
rect -799 1091 -737 1097
rect -671 1131 -609 1137
rect -671 1097 -659 1131
rect -621 1097 -609 1131
rect -671 1091 -609 1097
rect -543 1131 -481 1137
rect -543 1097 -531 1131
rect -493 1097 -481 1131
rect -543 1091 -481 1097
rect -415 1131 -353 1137
rect -415 1097 -403 1131
rect -365 1097 -353 1131
rect -415 1091 -353 1097
rect -287 1131 -225 1137
rect -287 1097 -275 1131
rect -237 1097 -225 1131
rect -287 1091 -225 1097
rect -159 1131 -97 1137
rect -159 1097 -147 1131
rect -109 1097 -97 1131
rect -159 1091 -97 1097
rect -31 1131 31 1137
rect -31 1097 -19 1131
rect 19 1097 31 1131
rect -31 1091 31 1097
rect 97 1131 159 1137
rect 97 1097 109 1131
rect 147 1097 159 1131
rect 97 1091 159 1097
rect 225 1131 287 1137
rect 225 1097 237 1131
rect 275 1097 287 1131
rect 225 1091 287 1097
rect 353 1131 415 1137
rect 353 1097 365 1131
rect 403 1097 415 1131
rect 353 1091 415 1097
rect 481 1131 543 1137
rect 481 1097 493 1131
rect 531 1097 543 1131
rect 481 1091 543 1097
rect 609 1131 671 1137
rect 609 1097 621 1131
rect 659 1097 671 1131
rect 609 1091 671 1097
rect 737 1131 799 1137
rect 737 1097 749 1131
rect 787 1097 799 1131
rect 737 1091 799 1097
rect 865 1131 927 1137
rect 865 1097 877 1131
rect 915 1097 927 1131
rect 865 1091 927 1097
rect -983 1038 -937 1050
rect -983 -1038 -977 1038
rect -943 -1038 -937 1038
rect -983 -1050 -937 -1038
rect -855 1038 -809 1050
rect -855 -1038 -849 1038
rect -815 -1038 -809 1038
rect -855 -1050 -809 -1038
rect -727 1038 -681 1050
rect -727 -1038 -721 1038
rect -687 -1038 -681 1038
rect -727 -1050 -681 -1038
rect -599 1038 -553 1050
rect -599 -1038 -593 1038
rect -559 -1038 -553 1038
rect -599 -1050 -553 -1038
rect -471 1038 -425 1050
rect -471 -1038 -465 1038
rect -431 -1038 -425 1038
rect -471 -1050 -425 -1038
rect -343 1038 -297 1050
rect -343 -1038 -337 1038
rect -303 -1038 -297 1038
rect -343 -1050 -297 -1038
rect -215 1038 -169 1050
rect -215 -1038 -209 1038
rect -175 -1038 -169 1038
rect -215 -1050 -169 -1038
rect -87 1038 -41 1050
rect -87 -1038 -81 1038
rect -47 -1038 -41 1038
rect -87 -1050 -41 -1038
rect 41 1038 87 1050
rect 41 -1038 47 1038
rect 81 -1038 87 1038
rect 41 -1050 87 -1038
rect 169 1038 215 1050
rect 169 -1038 175 1038
rect 209 -1038 215 1038
rect 169 -1050 215 -1038
rect 297 1038 343 1050
rect 297 -1038 303 1038
rect 337 -1038 343 1038
rect 297 -1050 343 -1038
rect 425 1038 471 1050
rect 425 -1038 431 1038
rect 465 -1038 471 1038
rect 425 -1050 471 -1038
rect 553 1038 599 1050
rect 553 -1038 559 1038
rect 593 -1038 599 1038
rect 553 -1050 599 -1038
rect 681 1038 727 1050
rect 681 -1038 687 1038
rect 721 -1038 727 1038
rect 681 -1050 727 -1038
rect 809 1038 855 1050
rect 809 -1038 815 1038
rect 849 -1038 855 1038
rect 809 -1050 855 -1038
rect 937 1038 983 1050
rect 937 -1038 943 1038
rect 977 -1038 983 1038
rect 937 -1050 983 -1038
rect -927 -1097 -865 -1091
rect -927 -1131 -915 -1097
rect -877 -1131 -865 -1097
rect -927 -1137 -865 -1131
rect -799 -1097 -737 -1091
rect -799 -1131 -787 -1097
rect -749 -1131 -737 -1097
rect -799 -1137 -737 -1131
rect -671 -1097 -609 -1091
rect -671 -1131 -659 -1097
rect -621 -1131 -609 -1097
rect -671 -1137 -609 -1131
rect -543 -1097 -481 -1091
rect -543 -1131 -531 -1097
rect -493 -1131 -481 -1097
rect -543 -1137 -481 -1131
rect -415 -1097 -353 -1091
rect -415 -1131 -403 -1097
rect -365 -1131 -353 -1097
rect -415 -1137 -353 -1131
rect -287 -1097 -225 -1091
rect -287 -1131 -275 -1097
rect -237 -1131 -225 -1097
rect -287 -1137 -225 -1131
rect -159 -1097 -97 -1091
rect -159 -1131 -147 -1097
rect -109 -1131 -97 -1097
rect -159 -1137 -97 -1131
rect -31 -1097 31 -1091
rect -31 -1131 -19 -1097
rect 19 -1131 31 -1097
rect -31 -1137 31 -1131
rect 97 -1097 159 -1091
rect 97 -1131 109 -1097
rect 147 -1131 159 -1097
rect 97 -1137 159 -1131
rect 225 -1097 287 -1091
rect 225 -1131 237 -1097
rect 275 -1131 287 -1097
rect 225 -1137 287 -1131
rect 353 -1097 415 -1091
rect 353 -1131 365 -1097
rect 403 -1131 415 -1097
rect 353 -1137 415 -1131
rect 481 -1097 543 -1091
rect 481 -1131 493 -1097
rect 531 -1131 543 -1097
rect 481 -1137 543 -1131
rect 609 -1097 671 -1091
rect 609 -1131 621 -1097
rect 659 -1131 671 -1097
rect 609 -1137 671 -1131
rect 737 -1097 799 -1091
rect 737 -1131 749 -1097
rect 787 -1131 799 -1097
rect 737 -1137 799 -1131
rect 865 -1097 927 -1091
rect 865 -1131 877 -1097
rect 915 -1131 927 -1097
rect 865 -1137 927 -1131
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1074 -1216 1074 1216
string parameters w 10.5 l 0.35 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
