magic
tech sky130A
magscale 1 2
timestamp 1623973798
<< nwell >>
rect -76 1856 48274 2870
rect -10 12 12851 1856
<< pwell >>
rect 16186 -14940 20257 -14839
rect 16186 -16005 20597 -14940
rect 16186 -16006 20628 -16005
rect 16186 -16853 20597 -16006
rect 16186 -16859 20257 -16853
rect 5066 -21156 10212 -19683
rect -49 -21425 48734 -21156
rect -54 -22020 48734 -21425
rect -64 -23588 48734 -22020
<< psubdiff >>
rect 16343 -15023 16746 -14999
rect 16343 -16574 16746 -16550
rect 20146 -15047 20549 -15023
rect 20146 -16598 20549 -16574
rect 26499 -19058 26523 -18504
rect 40693 -19058 40717 -18504
rect 277 -23223 301 -21906
rect 48300 -23223 48324 -21906
<< nsubdiff >>
rect 30 1922 54 2730
rect 47950 1922 47974 2730
<< psubdiffcont >>
rect 16343 -16550 16746 -15023
rect 20146 -16574 20549 -15047
rect 26523 -19058 40693 -18504
rect 301 -23223 48300 -21906
<< nsubdiffcont >>
rect 54 1922 47950 2730
<< locali >>
rect 38 1922 54 2730
rect 47950 1922 47966 2730
rect 16343 -15023 16746 -15007
rect 16343 -16566 16746 -16550
rect 20146 -15047 20549 -15031
rect 20146 -16590 20549 -16574
rect 26507 -19058 26523 -18504
rect 40693 -19058 40709 -18504
rect 285 -23223 301 -21906
rect 48300 -23223 48316 -21906
<< viali >>
rect 98 1922 47896 2730
rect 13282 1802 22371 1836
rect 25121 1802 34210 1836
rect 36971 1802 46060 1836
rect 22433 -4893 22467 1635
rect 25025 -4862 25059 1666
rect 34272 -4893 34306 1635
rect 36864 -4862 36898 1666
rect 46122 -5166 46156 1477
rect 13577 -5683 45774 -5649
rect 16343 -16499 16746 -15063
rect 20146 -16523 20549 -15087
rect 26545 -19058 40648 -18504
rect 329 -23223 47950 -21906
<< metal1 >>
rect 86 2730 47908 2736
rect 86 1922 98 2730
rect 47896 1922 47908 2730
rect 86 1916 47908 1922
rect 192 1854 47860 1916
rect 13194 1836 23370 1854
rect 13194 1802 13282 1836
rect 22371 1802 23370 1836
rect 13194 1792 23370 1802
rect 22348 1785 23370 1792
rect 24106 1836 47860 1854
rect 24106 1802 25121 1836
rect 34210 1802 36971 1836
rect 46060 1802 47860 1836
rect 24106 1785 47860 1802
rect 22348 1666 25128 1785
rect 22348 1635 25025 1666
rect 1133 58 1439 66
rect 1133 -32 1143 58
rect 1431 -32 1441 58
rect 1133 -42 1439 -32
rect 13062 -1197 13548 -1173
rect 13062 -1704 13095 -1197
rect 13341 -1704 13548 -1197
rect 13062 -1732 13548 -1704
rect 22348 -4893 22433 1635
rect 22467 -4862 25025 1635
rect 25059 -4862 25128 1666
rect 22467 -4893 25128 -4862
rect 22348 -5333 25128 -4893
rect 34186 1762 47860 1785
rect 34186 1666 37006 1762
rect 34186 1635 36864 1666
rect 34186 -4893 34272 1635
rect 34306 -4862 36864 1635
rect 36898 -3090 37006 1666
rect 46064 1477 47860 1762
rect 36898 -3655 36966 -3090
rect 36898 -4862 37006 -3655
rect 34306 -4893 37006 -4862
rect 34186 -5321 37006 -4893
rect 46064 -5166 46122 1477
rect 46156 -3090 47860 1477
rect 46156 -3655 46973 -3090
rect 46156 -5166 47860 -3655
rect 46064 -5321 47860 -5166
rect 34186 -5333 47860 -5321
rect 22348 -5341 47860 -5333
rect 13273 -5409 47860 -5341
rect 13270 -5455 47860 -5409
rect 13273 -5611 47860 -5455
rect 13273 -5649 18005 -5611
rect 18809 -5649 47860 -5611
rect 13273 -5683 13577 -5649
rect 45774 -5683 47860 -5649
rect 13273 -5727 18005 -5683
rect 13273 -6513 13311 -5727
rect 16294 -5925 18005 -5727
rect 17995 -6435 18005 -5925
rect 18809 -5897 47860 -5683
rect 18809 -5925 46087 -5897
rect 18809 -6435 18819 -5925
rect 22467 -6149 25128 -5925
rect 22467 -6213 25025 -6149
rect 46640 -6513 47860 -5897
rect 17939 -14859 18877 -14837
rect 17939 -15001 17963 -14859
rect 18854 -15001 18877 -14859
rect 17939 -15038 18877 -15001
rect 16327 -15063 16764 -15048
rect 16327 -16499 16343 -15063
rect 16746 -16499 16764 -15063
rect 17939 -15129 17963 -15038
rect 18199 -15042 18877 -15038
rect 18199 -15043 18582 -15042
rect 18199 -15123 18240 -15043
rect 18320 -15123 18349 -15043
rect 18429 -15123 18458 -15043
rect 18538 -15123 18582 -15043
rect 18199 -15129 18582 -15123
rect 17939 -15130 18582 -15129
rect 18864 -15130 18877 -15042
rect 17939 -15155 18877 -15130
rect 20130 -15087 20567 -15072
rect 5767 -19484 6638 -19456
rect 5767 -19672 5786 -19484
rect 6612 -19672 6638 -19484
rect 5767 -19698 6638 -19672
rect 5767 -19709 6645 -19698
rect 5767 -19805 5785 -19709
rect 6015 -19711 6645 -19709
rect 6015 -19805 6342 -19711
rect 5767 -19807 6342 -19805
rect 6634 -19807 6645 -19711
rect 5767 -19816 6645 -19807
rect 5767 -19817 6638 -19816
rect 5814 -19986 6548 -19817
rect 9052 -21766 9891 -21704
rect 16327 -21766 16764 -16499
rect 18001 -16325 18992 -16315
rect 18001 -16326 18390 -16325
rect 18001 -16386 18077 -16326
rect 18356 -16385 18390 -16326
rect 18450 -16385 18478 -16325
rect 18538 -16385 18566 -16325
rect 18626 -16326 18992 -16325
rect 18626 -16385 18656 -16326
rect 18356 -16386 18656 -16385
rect 18935 -16386 18992 -16326
rect 18001 -16423 18992 -16386
rect 18001 -16611 18039 -16423
rect 18965 -16611 18992 -16423
rect 18001 -16633 18992 -16611
rect 20130 -16523 20146 -15087
rect 20549 -16523 20567 -15087
rect 20130 -21766 20567 -16523
rect 26342 -18504 40891 -18439
rect 26342 -19058 26545 -18504
rect 40648 -19058 40891 -18504
rect 26342 -19111 40891 -19058
rect 26345 -21766 27017 -19111
rect 27646 -19495 27698 -19111
rect 27882 -19495 27934 -19111
rect 28118 -19495 28170 -19111
rect 28354 -19495 28406 -19111
rect 28590 -19495 28642 -19111
rect 28826 -19495 28878 -19111
rect 29062 -19495 29114 -19111
rect 29298 -19495 29350 -19111
rect 29534 -19495 29586 -19111
rect 29770 -19495 29822 -19111
rect 30006 -19495 30058 -19111
rect 30242 -19495 30294 -19111
rect 30478 -19495 30530 -19111
rect 30714 -19495 30766 -19111
rect 30950 -19495 31002 -19111
rect 31186 -19495 31238 -19111
rect 31422 -19495 31474 -19111
rect 31658 -19495 31710 -19111
rect 31894 -19495 31946 -19111
rect 32130 -19495 32182 -19111
rect 32366 -19495 32418 -19111
rect 32602 -19495 32654 -19111
rect 32838 -19495 32890 -19111
rect 33074 -19495 33126 -19111
rect 33310 -19495 33362 -19111
rect 33546 -19495 33598 -19111
rect 33782 -19495 33834 -19111
rect 34018 -19495 34070 -19111
rect 34254 -19495 34306 -19111
rect 34490 -19495 34542 -19111
rect 34726 -19495 34778 -19111
rect 34962 -19495 35014 -19111
rect 35198 -19495 35250 -19111
rect 35434 -19495 35486 -19111
rect 35670 -19495 35722 -19111
rect 35906 -19495 35958 -19111
rect 36142 -19495 36194 -19111
rect 36378 -19495 36430 -19111
rect 36614 -19495 36666 -19111
rect 36850 -19495 36902 -19111
rect 37086 -19495 37138 -19111
rect 37322 -19495 37374 -19111
rect 37558 -19495 37610 -19111
rect 37794 -19495 37846 -19111
rect 38030 -19495 38082 -19111
rect 38266 -19495 38318 -19111
rect 38502 -19495 38554 -19111
rect 38738 -19495 38790 -19111
rect 38974 -19495 39026 -19111
rect 39210 -19495 39262 -19111
rect 39446 -19495 39498 -19111
rect 27399 -20187 27606 -20166
rect 27393 -20828 27403 -20187
rect 27509 -20241 27606 -20187
rect 27509 -20301 27537 -20241
rect 27597 -20301 27607 -20241
rect 27509 -20687 27606 -20301
rect 27509 -20747 27538 -20687
rect 27598 -20747 27608 -20687
rect 27509 -20828 27606 -20747
rect 27399 -20845 27606 -20828
rect 27646 -21766 27698 -21491
rect 27882 -21766 27934 -21491
rect 28118 -21766 28170 -21491
rect 28354 -21766 28406 -21491
rect 28590 -21766 28642 -21491
rect 28826 -21766 28878 -21491
rect 29062 -21766 29114 -21491
rect 29298 -21766 29350 -21491
rect 29534 -21766 29586 -21491
rect 29770 -21766 29822 -21491
rect 30006 -21766 30058 -21491
rect 30242 -21766 30294 -21491
rect 30478 -21766 30530 -21491
rect 30714 -21766 30766 -21491
rect 30950 -21766 31002 -21491
rect 31186 -21766 31238 -21491
rect 31422 -21766 31474 -21491
rect 31658 -21766 31710 -21491
rect 31894 -21766 31946 -21491
rect 32130 -21766 32182 -21491
rect 32366 -21766 32418 -21491
rect 32602 -21766 32654 -21491
rect 32838 -21766 32890 -21491
rect 33074 -21766 33126 -21491
rect 33310 -21766 33362 -21491
rect 33546 -21766 33598 -21491
rect 33782 -21766 33834 -21491
rect 34018 -21766 34070 -21491
rect 34254 -21766 34306 -21491
rect 34490 -21766 34542 -21491
rect 34726 -21766 34778 -21491
rect 34962 -21766 35014 -21491
rect 35198 -21766 35250 -21491
rect 35434 -21766 35486 -21491
rect 35670 -21766 35722 -21491
rect 35906 -21766 35958 -21491
rect 36142 -21766 36194 -21491
rect 36378 -21766 36430 -21491
rect 36614 -21766 36666 -21491
rect 36850 -21766 36902 -21491
rect 37086 -21766 37138 -21491
rect 37322 -21766 37374 -21491
rect 37558 -21766 37610 -21491
rect 37794 -21766 37846 -21491
rect 38030 -21766 38082 -21491
rect 38266 -21766 38318 -21491
rect 38502 -21766 38554 -21491
rect 38738 -21766 38790 -21491
rect 38974 -21766 39026 -21491
rect 39210 -21766 39262 -21491
rect 39446 -21766 39498 -21491
rect 5754 -21767 39782 -21766
rect 5754 -21900 39799 -21767
rect 40219 -21900 40891 -19111
rect 317 -21906 47962 -21900
rect 317 -23223 329 -21906
rect 47950 -23223 47962 -21906
rect 317 -23229 47962 -23223
<< via1 >>
rect 1143 -32 1431 58
rect 13095 -1704 13341 -1197
rect 18005 -5649 18809 -5611
rect 18005 -5683 18809 -5649
rect 18005 -6435 18809 -5683
rect 17963 -15001 18854 -14859
rect 17963 -15129 18199 -15038
rect 18240 -15123 18320 -15043
rect 18349 -15123 18429 -15043
rect 18458 -15123 18538 -15043
rect 18582 -15130 18864 -15042
rect 5786 -19672 6612 -19484
rect 5785 -19805 6015 -19709
rect 6342 -19807 6634 -19711
rect 18077 -16386 18356 -16326
rect 18390 -16385 18450 -16325
rect 18478 -16385 18538 -16325
rect 18566 -16385 18626 -16325
rect 18656 -16386 18935 -16326
rect 18039 -16611 18965 -16423
rect 27403 -20828 27509 -20187
rect 27537 -20301 27597 -20241
rect 27538 -20747 27598 -20687
<< metal2 >>
rect 1143 58 1431 68
rect 1143 -42 1431 -32
rect 10445 54 10690 64
rect 10445 -30 10455 54
rect 10680 -30 10690 54
rect 7186 -153 8123 -152
rect 7174 -162 8123 -153
rect 7174 -223 7186 -162
rect 7387 -164 8123 -162
rect 7387 -223 7531 -164
rect 7174 -224 7531 -223
rect 7787 -165 8123 -164
rect 7787 -224 7909 -165
rect 8109 -224 8123 -165
rect 7174 -264 8123 -224
rect 7174 -379 7192 -264
rect 8096 -379 8123 -264
rect 7174 -2425 8123 -379
rect 10445 -1178 10690 -30
rect 10445 -1719 10454 -1178
rect 10680 -1719 10690 -1178
rect 10445 -1727 10690 -1719
rect 13062 -1197 13548 -1173
rect 13062 -1704 13095 -1197
rect 13341 -1704 13548 -1197
rect 10454 -1729 10680 -1727
rect 13062 -1732 13548 -1704
rect 932 -2440 1881 -2430
rect 932 -3363 937 -2440
rect 1854 -3363 1881 -2440
rect 932 -12357 1881 -3363
rect 8123 -3373 8124 -3227
rect 7174 -3383 8123 -3373
rect 17934 -5611 18885 -5565
rect 17934 -6435 18005 -5611
rect 18809 -6435 18885 -5611
rect 17934 -14859 18885 -6435
rect 17934 -15001 17963 -14859
rect 18854 -15001 18885 -14859
rect 17934 -15038 18885 -15001
rect 17934 -15129 17963 -15038
rect 18199 -15042 18885 -15038
rect 18199 -15043 18582 -15042
rect 18199 -15123 18240 -15043
rect 18320 -15123 18349 -15043
rect 18429 -15123 18458 -15043
rect 18538 -15123 18582 -15043
rect 18199 -15129 18582 -15123
rect 17934 -15130 18582 -15129
rect 18864 -15130 18885 -15042
rect 17934 -15158 18885 -15130
rect 17170 -15263 18236 -15253
rect 17170 -15338 18236 -15328
rect 18547 -15264 19613 -15254
rect 18547 -15339 19613 -15329
rect 18001 -16325 18992 -16315
rect 18001 -16326 18390 -16325
rect 18001 -16386 18077 -16326
rect 18356 -16385 18390 -16326
rect 18450 -16385 18478 -16325
rect 18538 -16385 18566 -16325
rect 18626 -16326 18992 -16325
rect 18626 -16385 18656 -16326
rect 18356 -16386 18656 -16385
rect 18935 -16386 18992 -16326
rect 18001 -16423 18992 -16386
rect 18001 -16611 18039 -16423
rect 18965 -16611 18992 -16423
rect 18001 -16633 18992 -16611
rect 8971 -19405 9938 -19402
rect 8959 -19412 9959 -19405
rect 5767 -19484 6638 -19456
rect 5767 -19672 5786 -19484
rect 6612 -19672 6638 -19484
rect 8959 -19553 8971 -19412
rect 9938 -19553 9959 -19412
rect 8959 -19560 9959 -19553
rect 8957 -19580 9959 -19560
rect 8957 -19582 9640 -19580
rect 8957 -19647 8968 -19582
rect 9310 -19646 9640 -19582
rect 9939 -19581 9959 -19580
rect 9939 -19646 9960 -19581
rect 9310 -19647 9960 -19646
rect 8957 -19654 9960 -19647
rect 8957 -19662 9959 -19654
rect 5767 -19709 6638 -19672
rect 5767 -19805 5785 -19709
rect 6015 -19710 6638 -19709
rect 6015 -19805 6047 -19710
rect 5767 -19813 6047 -19805
rect 6167 -19813 6196 -19710
rect 6316 -19711 6638 -19710
rect 6316 -19807 6342 -19711
rect 6634 -19807 6638 -19711
rect 6316 -19813 6638 -19807
rect 5767 -19817 6638 -19813
rect 6047 -19823 6167 -19817
rect 6196 -19818 6470 -19817
rect 6196 -19823 6316 -19818
rect 27403 -20187 27509 -20177
rect 27537 -20241 27597 -20231
rect 27537 -20311 27597 -20301
rect 27538 -20687 27598 -20677
rect 27538 -20757 27598 -20747
rect 27403 -20838 27509 -20828
<< via2 >>
rect 1143 -32 1431 58
rect 10455 -30 10680 54
rect 7186 -223 7387 -162
rect 7531 -224 7787 -164
rect 7909 -224 8109 -165
rect 7192 -379 8096 -264
rect 10454 -1719 10680 -1178
rect 13095 -1704 13341 -1197
rect 937 -3363 1854 -2440
rect 7174 -3373 8123 -2425
rect 17170 -15328 18236 -15263
rect 18547 -15329 19613 -15264
rect 18077 -16386 18356 -16326
rect 18390 -16385 18450 -16325
rect 18478 -16385 18538 -16325
rect 18566 -16385 18626 -16325
rect 18656 -16386 18935 -16326
rect 18039 -16611 18965 -16423
rect 5786 -19672 6612 -19484
rect 8971 -19553 9938 -19412
rect 8968 -19647 9310 -19582
rect 9640 -19646 9939 -19580
rect 5785 -19805 6015 -19709
rect 6047 -19813 6167 -19710
rect 6196 -19813 6316 -19710
rect 6342 -19807 6634 -19711
rect 27403 -20828 27509 -20187
rect 27537 -20301 27597 -20241
rect 27538 -20747 27598 -20687
<< metal3 >>
rect -759 58 10914 114
rect -759 -32 1143 58
rect 1431 54 10914 58
rect 1431 -30 10455 54
rect 10680 -30 10914 54
rect 1431 -32 10914 -30
rect -759 -87 10914 -32
rect 7175 -162 8119 -156
rect 7175 -223 7186 -162
rect 7387 -164 8119 -162
rect 7387 -223 7531 -164
rect 7175 -224 7531 -223
rect 7787 -165 8119 -164
rect 7787 -224 7909 -165
rect 8109 -224 8119 -165
rect 7175 -264 8119 -224
rect 7175 -379 7192 -264
rect 8096 -379 8119 -264
rect 7175 -389 8119 -379
rect 10445 -1173 13551 -1168
rect 10444 -1178 13551 -1173
rect 10444 -1719 10454 -1178
rect 10680 -1197 13551 -1178
rect 10680 -1704 13095 -1197
rect 13341 -1704 13551 -1197
rect 10680 -1719 13551 -1704
rect 10444 -1724 13551 -1719
rect 10445 -1730 13551 -1724
rect 7164 -2425 8133 -2420
rect 932 -2435 7174 -2425
rect 927 -2440 7174 -2435
rect 927 -3363 937 -2440
rect 1854 -3363 7174 -2440
rect 927 -3368 7174 -3363
rect 932 -3373 7174 -3368
rect 8123 -3373 8133 -2425
rect 7164 -3378 8133 -3373
rect 13809 -5221 45514 -5218
rect -1038 -6128 378 -5250
rect 8729 -6100 8739 -5289
rect 10205 -6100 10215 -5289
rect 13809 -5314 29210 -5221
rect 29200 -5318 29210 -5314
rect 30103 -5223 45514 -5221
rect 30103 -5313 41055 -5223
rect 41936 -5313 45514 -5223
rect 30103 -5314 45514 -5313
rect 30103 -5318 30113 -5314
rect 29211 -5352 30101 -5318
rect 29211 -5494 29228 -5352
rect 30090 -5494 30101 -5352
rect 29211 -5513 30101 -5494
rect 41047 -5368 41947 -5314
rect 41047 -5510 41061 -5368
rect 41923 -5510 41947 -5368
rect 41047 -5566 41947 -5510
rect 8742 -7584 8752 -6804
rect 10173 -7584 10183 -6804
rect 26886 -8740 27110 -8737
rect 19396 -14196 19879 -8774
rect 26789 -14196 27115 -8740
rect 34139 -14196 34481 -8772
rect 41497 -8779 41839 -8768
rect 41497 -14196 41840 -8779
rect 19396 -14674 41884 -14196
rect 19396 -15256 19879 -14674
rect 17182 -15258 19879 -15256
rect 17160 -15263 19879 -15258
rect 17160 -15328 17170 -15263
rect 18236 -15264 19879 -15263
rect 18236 -15328 18547 -15264
rect 17160 -15329 18547 -15328
rect 19613 -15329 19879 -15264
rect 17160 -15333 19879 -15329
rect 17182 -15336 19879 -15333
rect 18275 -15337 19296 -15336
rect 18001 -16395 18071 -16315
rect 18941 -16395 18992 -16315
rect 18001 -16423 18992 -16395
rect 8742 -17316 8752 -16536
rect 10173 -17316 10183 -16536
rect 18001 -16611 18039 -16423
rect 18965 -16611 18992 -16423
rect 18001 -16633 18992 -16611
rect -1038 -18870 378 -17992
rect 36485 -19136 37355 -19120
rect 29213 -19183 30088 -19175
rect 29213 -19297 29225 -19183
rect 30069 -19297 30088 -19183
rect 29213 -19337 30088 -19297
rect 36485 -19302 36509 -19136
rect 37324 -19302 37355 -19136
rect 36485 -19337 37355 -19302
rect 8959 -19412 9959 -19405
rect 29205 -19411 29215 -19337
rect 30085 -19411 30095 -19337
rect 36475 -19412 36485 -19337
rect 37357 -19412 37367 -19337
rect 5767 -19484 6638 -19456
rect 5767 -19672 5786 -19484
rect 6612 -19672 6638 -19484
rect 8959 -19553 8971 -19412
rect 9938 -19553 9959 -19412
rect 8959 -19555 9959 -19553
rect 8957 -19580 9959 -19555
rect 8957 -19582 9640 -19580
rect 8957 -19647 8968 -19582
rect 9310 -19646 9640 -19582
rect 9939 -19581 9959 -19580
rect 9939 -19646 9960 -19581
rect 9310 -19647 9960 -19646
rect 8957 -19654 9960 -19647
rect 8957 -19657 9959 -19654
rect 8959 -19658 9959 -19657
rect 5767 -19706 6638 -19672
rect 5767 -19709 6644 -19706
rect 5767 -19805 5785 -19709
rect 6015 -19710 6644 -19709
rect 6015 -19805 6047 -19710
rect 5767 -19813 6047 -19805
rect 6167 -19813 6196 -19710
rect 6316 -19711 6644 -19710
rect 6316 -19807 6342 -19711
rect 6634 -19720 6644 -19711
rect 6634 -19807 8629 -19720
rect 6316 -19813 8629 -19807
rect 5767 -19817 8629 -19813
rect 5770 -19847 8629 -19817
rect 18021 -20187 27610 -20165
rect 18021 -20196 27403 -20187
rect 18021 -20800 18046 -20196
rect 18964 -20800 27403 -20196
rect 18021 -20828 27403 -20800
rect 27509 -20241 27610 -20187
rect 27509 -20301 27537 -20241
rect 27597 -20301 27610 -20241
rect 27509 -20687 27610 -20301
rect 27509 -20747 27538 -20687
rect 27598 -20747 27610 -20687
rect 27509 -20828 27610 -20747
rect 18021 -20846 27610 -20828
<< via3 >>
rect 29210 -5318 30103 -5221
rect 41055 -5313 41936 -5223
rect 29228 -5494 30090 -5352
rect 41061 -5510 41923 -5368
rect 8752 -7584 10173 -6804
rect 18071 -16325 18941 -16315
rect 18071 -16326 18390 -16325
rect 18071 -16386 18077 -16326
rect 18077 -16386 18356 -16326
rect 18356 -16385 18390 -16326
rect 18390 -16385 18450 -16325
rect 18450 -16385 18478 -16325
rect 18478 -16385 18538 -16325
rect 18538 -16385 18566 -16325
rect 18566 -16385 18626 -16325
rect 18626 -16326 18941 -16325
rect 18626 -16385 18656 -16326
rect 18356 -16386 18656 -16385
rect 18656 -16386 18935 -16326
rect 18935 -16386 18941 -16326
rect 18071 -16395 18941 -16386
rect 8752 -17316 10173 -16536
rect 18039 -16611 18965 -16423
rect 29225 -19297 30069 -19183
rect 36509 -19302 37324 -19136
rect 29215 -19411 30085 -19337
rect 36485 -19412 37357 -19337
rect 5786 -19672 6612 -19484
rect 8971 -19553 9938 -19412
rect 8968 -19647 9310 -19582
rect 9640 -19646 9939 -19580
rect 5785 -19805 6015 -19709
rect 6047 -19813 6167 -19710
rect 6196 -19813 6316 -19710
rect 6342 -19807 6634 -19711
rect 18046 -20800 18964 -20196
<< metal4 >>
rect 29210 -5220 30110 -5215
rect 29209 -5221 30110 -5220
rect 29209 -5318 29210 -5221
rect 30103 -5318 30110 -5221
rect 29209 -5319 30110 -5318
rect 29210 -5352 30110 -5319
rect 29210 -5494 29228 -5352
rect 30090 -5494 30110 -5352
rect 5771 -6804 10240 -6762
rect 5771 -7584 8752 -6804
rect 10173 -7584 10240 -6804
rect 29210 -7578 30110 -5494
rect 41048 -5223 41948 -5218
rect 41048 -5313 41055 -5223
rect 41936 -5313 41948 -5223
rect 41048 -5368 41948 -5313
rect 41048 -5510 41061 -5368
rect 41923 -5510 41948 -5368
rect 41048 -7578 41948 -5510
rect 46430 -7578 51308 -7564
rect 21893 -7580 51308 -7578
rect 5771 -7644 10240 -7584
rect 5771 -19484 6638 -7644
rect 21868 -8451 51308 -7580
rect 21868 -15215 22741 -8451
rect 29217 -15215 30090 -8451
rect 36484 -15215 37359 -8451
rect 43714 -15215 44587 -8451
rect 50435 -15214 51308 -8451
rect 46215 -15215 51308 -15214
rect 21868 -16088 51308 -15215
rect 17999 -16315 19001 -16312
rect 17999 -16395 18071 -16315
rect 18941 -16395 19001 -16315
rect 17999 -16423 19001 -16395
rect 8698 -16536 10240 -16476
rect 8698 -17316 8752 -16536
rect 10173 -17316 10240 -16536
rect 8698 -17364 10240 -17316
rect 17999 -16611 18039 -16423
rect 18965 -16611 19001 -16423
rect 5771 -19672 5786 -19484
rect 6612 -19672 6638 -19484
rect 8958 -18660 9960 -17364
rect 17999 -18660 19001 -16611
rect 29217 -17657 30090 -16088
rect 8958 -19412 19001 -18660
rect 29213 -19183 30090 -17657
rect 29213 -19297 29225 -19183
rect 30069 -19297 30090 -19183
rect 29213 -19337 30090 -19297
rect 29213 -19411 29215 -19337
rect 30085 -19411 30090 -19337
rect 29213 -19412 30090 -19411
rect 36484 -19136 37359 -16088
rect 43714 -16102 44587 -16088
rect 36484 -19302 36509 -19136
rect 37324 -19302 37359 -19136
rect 36484 -19337 37359 -19302
rect 36484 -19412 36485 -19337
rect 37357 -19412 37359 -19337
rect 8958 -19553 8971 -19412
rect 9938 -19553 19001 -19412
rect 36484 -19413 37359 -19412
rect 8958 -19555 19001 -19553
rect 8957 -19580 19001 -19555
rect 8957 -19582 9640 -19580
rect 8957 -19647 8968 -19582
rect 9310 -19646 9640 -19582
rect 9939 -19646 19001 -19580
rect 9310 -19647 19001 -19646
rect 8957 -19657 19001 -19647
rect 8958 -19662 19001 -19657
rect 5771 -19709 6638 -19672
rect 5771 -19805 5785 -19709
rect 6015 -19710 6638 -19709
rect 6015 -19805 6047 -19710
rect 5771 -19813 6047 -19805
rect 6167 -19813 6196 -19710
rect 6316 -19711 6638 -19710
rect 6316 -19807 6342 -19711
rect 6634 -19807 6638 -19711
rect 6316 -19813 6638 -19807
rect 5771 -19818 6638 -19813
rect 17999 -20196 19001 -19662
rect 17999 -20800 18046 -20196
rect 18964 -20800 19001 -20196
rect 17999 -20848 19001 -20800
use M9  M9_0
timestamp 1615944125
transform 1 0 17118 0 1 -15250
box -546 -1326 3146 243
use M6  M6_0
timestamp 1615925795
transform 1 0 27643 0 1 -20881
box -637 -1175 12467 2068
use M4  M4_0
timestamp 1615949206
transform 1 0 3689 0 1 -21635
box 4940 -92 6345 2059
use M3  M3_0
timestamp 1615949206
transform 1 0 4004 0 1 -22431
box 1612 645 2738 2732
use sky130_fd_pr__cap_mim_m3_1_2674SJ  sky130_fd_pr__cap_mim_m3_1_2674SJ_3
timestamp 1616037006
transform -1 0 22324 0 1 -11269
box -2550 -2500 2549 2500
use sky130_fd_pr__cap_mim_m3_1_2674SJ  sky130_fd_pr__cap_mim_m3_1_2674SJ_0
timestamp 1616037006
transform -1 0 44296 0 1 -11271
box -2550 -2500 2549 2500
use sky130_fd_pr__cap_mim_m3_1_2674SJ  sky130_fd_pr__cap_mim_m3_1_2674SJ_1
timestamp 1616037006
transform -1 0 36931 0 1 -11271
box -2550 -2500 2549 2500
use sky130_fd_pr__cap_mim_m3_1_2674SJ  sky130_fd_pr__cap_mim_m3_1_2674SJ_2
timestamp 1616037006
transform -1 0 29566 0 1 -11229
box -2550 -2500 2549 2500
use M7  M7_0
timestamp 1623972813
transform 1 0 14034 0 1 -435
box -1784 -6078 34024 3239
use M8  M8_0
timestamp 1616023926
transform 1 0 182 0 1 156
box -182 -156 2368 2112
use M5_B  M5_B_0
timestamp 1616024728
transform 1 0 2653 0 1 156
box -104 -385 10001 2080
use M1_2  M1_2_0
timestamp 1616093313
transform 1 0 2173 0 1 -10801
box -1795 -8069 14571 5551
<< labels >>
rlabel nwell 155 1973 1445 2651 1 vdd
rlabel metal3 -750 -35 -572 63 1 iref
rlabel metal4 50484 -13534 51240 -9354 1 vout
rlabel pwell 440 -22991 1856 -22113 1 vss
rlabel metal3 -1038 -6128 378 -5250 1 vin_n
rlabel metal3 -1038 -18870 378 -17992 1 vin_p
<< end >>
