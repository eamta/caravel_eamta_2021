magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -557 222 -499 228
rect -365 222 -307 228
rect -173 222 -115 228
rect 19 222 77 228
rect 211 222 269 228
rect 403 222 461 228
rect 595 222 653 228
rect -557 188 -545 222
rect -365 188 -353 222
rect -173 188 -161 222
rect 19 188 31 222
rect 211 188 223 222
rect 403 188 415 222
rect 595 188 607 222
rect -557 182 -499 188
rect -365 182 -307 188
rect -173 182 -115 188
rect 19 182 77 188
rect 211 182 269 188
rect 403 182 461 188
rect 595 182 653 188
rect -653 -188 -595 -182
rect -461 -188 -403 -182
rect -269 -188 -211 -182
rect -77 -188 -19 -182
rect 115 -188 173 -182
rect 307 -188 365 -182
rect 499 -188 557 -182
rect -653 -222 -641 -188
rect -461 -222 -449 -188
rect -269 -222 -257 -188
rect -77 -222 -65 -188
rect 115 -222 127 -188
rect 307 -222 319 -188
rect 499 -222 511 -188
rect -653 -228 -595 -222
rect -461 -228 -403 -222
rect -269 -228 -211 -222
rect -77 -228 -19 -222
rect 115 -228 173 -222
rect 307 -228 365 -222
rect 499 -228 557 -222
<< pwell >>
rect -839 -360 839 360
<< nmos >>
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
<< ndiff >>
rect -701 138 -639 150
rect -701 -138 -689 138
rect -655 -138 -639 138
rect -701 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 701 150
rect 639 -138 655 138
rect 689 -138 701 138
rect 639 -150 701 -138
<< ndiffc >>
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
<< psubdiff >>
rect -803 290 -707 324
rect 707 290 803 324
rect -803 228 -769 290
rect 769 228 803 290
rect -803 -290 -769 -228
rect 769 -290 803 -228
rect -803 -324 -707 -290
rect 707 -324 803 -290
<< psubdiffcont >>
rect -707 290 707 324
rect -803 -228 -769 228
rect 769 -228 803 228
rect -707 -324 707 -290
<< poly >>
rect -561 222 -495 238
rect -561 188 -545 222
rect -511 188 -495 222
rect -639 150 -609 176
rect -561 172 -495 188
rect -369 222 -303 238
rect -369 188 -353 222
rect -319 188 -303 222
rect -543 150 -513 172
rect -447 150 -417 176
rect -369 172 -303 188
rect -177 222 -111 238
rect -177 188 -161 222
rect -127 188 -111 222
rect -351 150 -321 172
rect -255 150 -225 176
rect -177 172 -111 188
rect 15 222 81 238
rect 15 188 31 222
rect 65 188 81 222
rect -159 150 -129 172
rect -63 150 -33 176
rect 15 172 81 188
rect 207 222 273 238
rect 207 188 223 222
rect 257 188 273 222
rect 33 150 63 172
rect 129 150 159 176
rect 207 172 273 188
rect 399 222 465 238
rect 399 188 415 222
rect 449 188 465 222
rect 225 150 255 172
rect 321 150 351 176
rect 399 172 465 188
rect 591 222 657 238
rect 591 188 607 222
rect 641 188 657 222
rect 417 150 447 172
rect 513 150 543 176
rect 591 172 657 188
rect 609 150 639 172
rect -639 -172 -609 -150
rect -657 -188 -591 -172
rect -543 -176 -513 -150
rect -447 -172 -417 -150
rect -657 -222 -641 -188
rect -607 -222 -591 -188
rect -657 -238 -591 -222
rect -465 -188 -399 -172
rect -351 -176 -321 -150
rect -255 -172 -225 -150
rect -465 -222 -449 -188
rect -415 -222 -399 -188
rect -465 -238 -399 -222
rect -273 -188 -207 -172
rect -159 -176 -129 -150
rect -63 -172 -33 -150
rect -273 -222 -257 -188
rect -223 -222 -207 -188
rect -273 -238 -207 -222
rect -81 -188 -15 -172
rect 33 -176 63 -150
rect 129 -172 159 -150
rect -81 -222 -65 -188
rect -31 -222 -15 -188
rect -81 -238 -15 -222
rect 111 -188 177 -172
rect 225 -176 255 -150
rect 321 -172 351 -150
rect 111 -222 127 -188
rect 161 -222 177 -188
rect 111 -238 177 -222
rect 303 -188 369 -172
rect 417 -176 447 -150
rect 513 -172 543 -150
rect 303 -222 319 -188
rect 353 -222 369 -188
rect 303 -238 369 -222
rect 495 -188 561 -172
rect 609 -176 639 -150
rect 495 -222 511 -188
rect 545 -222 561 -188
rect 495 -238 561 -222
<< polycont >>
rect -545 188 -511 222
rect -353 188 -319 222
rect -161 188 -127 222
rect 31 188 65 222
rect 223 188 257 222
rect 415 188 449 222
rect 607 188 641 222
rect -641 -222 -607 -188
rect -449 -222 -415 -188
rect -257 -222 -223 -188
rect -65 -222 -31 -188
rect 127 -222 161 -188
rect 319 -222 353 -188
rect 511 -222 545 -188
<< locali >>
rect -803 290 -707 324
rect 707 290 803 324
rect -803 228 -769 290
rect 769 228 803 290
rect -561 188 -545 222
rect -511 188 -495 222
rect -369 188 -353 222
rect -319 188 -303 222
rect -177 188 -161 222
rect -127 188 -111 222
rect 15 188 31 222
rect 65 188 81 222
rect 207 188 223 222
rect 257 188 273 222
rect 399 188 415 222
rect 449 188 465 222
rect 591 188 607 222
rect 641 188 657 222
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect -657 -222 -641 -188
rect -607 -222 -591 -188
rect -465 -222 -449 -188
rect -415 -222 -399 -188
rect -273 -222 -257 -188
rect -223 -222 -207 -188
rect -81 -222 -65 -188
rect -31 -222 -15 -188
rect 111 -222 127 -188
rect 161 -222 177 -188
rect 303 -222 319 -188
rect 353 -222 369 -188
rect 495 -222 511 -188
rect 545 -222 561 -188
rect -803 -290 -769 -228
rect 769 -290 803 -228
rect -803 -324 -707 -290
rect 707 -324 803 -290
<< viali >>
rect -545 188 -511 222
rect -353 188 -319 222
rect -161 188 -127 222
rect 31 188 65 222
rect 223 188 257 222
rect 415 188 449 222
rect 607 188 641 222
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect -641 -222 -607 -188
rect -449 -222 -415 -188
rect -257 -222 -223 -188
rect -65 -222 -31 -188
rect 127 -222 161 -188
rect 319 -222 353 -188
rect 511 -222 545 -188
<< metal1 >>
rect -557 222 -499 228
rect -557 188 -545 222
rect -511 188 -499 222
rect -557 182 -499 188
rect -365 222 -307 228
rect -365 188 -353 222
rect -319 188 -307 222
rect -365 182 -307 188
rect -173 222 -115 228
rect -173 188 -161 222
rect -127 188 -115 222
rect -173 182 -115 188
rect 19 222 77 228
rect 19 188 31 222
rect 65 188 77 222
rect 19 182 77 188
rect 211 222 269 228
rect 211 188 223 222
rect 257 188 269 222
rect 211 182 269 188
rect 403 222 461 228
rect 403 188 415 222
rect 449 188 461 222
rect 403 182 461 188
rect 595 222 653 228
rect 595 188 607 222
rect 641 188 653 222
rect 595 182 653 188
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
rect -653 -188 -595 -182
rect -653 -222 -641 -188
rect -607 -222 -595 -188
rect -653 -228 -595 -222
rect -461 -188 -403 -182
rect -461 -222 -449 -188
rect -415 -222 -403 -188
rect -461 -228 -403 -222
rect -269 -188 -211 -182
rect -269 -222 -257 -188
rect -223 -222 -211 -188
rect -269 -228 -211 -222
rect -77 -188 -19 -182
rect -77 -222 -65 -188
rect -31 -222 -19 -188
rect -77 -228 -19 -222
rect 115 -188 173 -182
rect 115 -222 127 -188
rect 161 -222 173 -188
rect 115 -228 173 -222
rect 307 -188 365 -182
rect 307 -222 319 -188
rect 353 -222 365 -188
rect 307 -228 365 -222
rect 499 -188 557 -182
rect 499 -222 511 -188
rect 545 -222 557 -188
rect 499 -228 557 -222
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -786 -307 786 307
string parameters w 1.5 l 0.150 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
