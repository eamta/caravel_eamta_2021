magic
tech sky130A
magscale 1 2
timestamp 1623972813
<< nwell >>
rect -1784 -5513 34024 3239
<< pmos >>
rect 11495 740 11635 2140
rect 11693 740 11833 2140
rect 11891 740 12031 2140
rect 12089 740 12229 2140
rect 12287 740 12427 2140
rect 12485 740 12625 2140
rect 12683 740 12823 2140
rect 12881 740 13021 2140
rect 13079 740 13219 2140
rect 13277 740 13417 2140
rect 13475 740 13615 2140
rect 13673 740 13813 2140
rect 13871 740 14011 2140
rect 14069 740 14209 2140
rect 14267 740 14407 2140
rect 14465 740 14605 2140
rect 14663 740 14803 2140
rect 14861 740 15001 2140
rect 15059 740 15199 2140
rect 15257 740 15397 2140
rect 15455 740 15595 2140
rect 15653 740 15793 2140
rect 15851 740 15991 2140
rect 16049 740 16189 2140
rect 16247 740 16387 2140
rect 16445 740 16585 2140
rect 16643 740 16783 2140
rect 16841 740 16981 2140
rect 17039 740 17179 2140
rect 17237 740 17377 2140
rect 17435 740 17575 2140
rect 17633 740 17773 2140
rect 17831 740 17971 2140
rect 18029 740 18169 2140
rect 18227 740 18367 2140
rect 18425 740 18565 2140
rect 18623 740 18763 2140
rect 18821 740 18961 2140
rect 19019 740 19159 2140
rect 19217 740 19357 2140
rect 19415 740 19555 2140
rect 19613 740 19753 2140
rect 11495 -896 11635 504
rect 11693 -896 11833 504
rect 11891 -896 12031 504
rect 12089 -896 12229 504
rect 12287 -896 12427 504
rect 12485 -896 12625 504
rect 12683 -896 12823 504
rect 12881 -896 13021 504
rect 13079 -896 13219 504
rect 13277 -896 13417 504
rect 13475 -896 13615 504
rect 13673 -896 13813 504
rect 13871 -896 14011 504
rect 14069 -896 14209 504
rect 14267 -896 14407 504
rect 14465 -896 14605 504
rect 14663 -896 14803 504
rect 14861 -896 15001 504
rect 15059 -896 15199 504
rect 15257 -896 15397 504
rect 15455 -896 15595 504
rect 15653 -896 15793 504
rect 15851 -896 15991 504
rect 16049 -896 16189 504
rect 16247 -896 16387 504
rect 16445 -896 16585 504
rect 16643 -896 16783 504
rect 16841 -896 16981 504
rect 17039 -896 17179 504
rect 17237 -896 17377 504
rect 17435 -896 17575 504
rect 17633 -896 17773 504
rect 17831 -896 17971 504
rect 18029 -896 18169 504
rect 18227 -896 18367 504
rect 18425 -896 18565 504
rect 18623 -896 18763 504
rect 18821 -896 18961 504
rect 19019 -896 19159 504
rect 19217 -896 19357 504
rect 19415 -896 19555 504
rect 19613 -896 19753 504
rect 11495 -2532 11635 -1132
rect 11693 -2532 11833 -1132
rect 11891 -2532 12031 -1132
rect 12089 -2532 12229 -1132
rect 12287 -2532 12427 -1132
rect 12485 -2532 12625 -1132
rect 12683 -2532 12823 -1132
rect 12881 -2532 13021 -1132
rect 13079 -2532 13219 -1132
rect 13277 -2532 13417 -1132
rect 13475 -2532 13615 -1132
rect 13673 -2532 13813 -1132
rect 13871 -2532 14011 -1132
rect 14069 -2532 14209 -1132
rect 14267 -2532 14407 -1132
rect 14465 -2532 14605 -1132
rect 14663 -2532 14803 -1132
rect 14861 -2532 15001 -1132
rect 15059 -2532 15199 -1132
rect 15257 -2532 15397 -1132
rect 15455 -2532 15595 -1132
rect 15653 -2532 15793 -1132
rect 15851 -2532 15991 -1132
rect 16049 -2532 16189 -1132
rect 16247 -2532 16387 -1132
rect 16445 -2532 16585 -1132
rect 16643 -2532 16783 -1132
rect 16841 -2532 16981 -1132
rect 17039 -2532 17179 -1132
rect 17237 -2532 17377 -1132
rect 17435 -2532 17575 -1132
rect 17633 -2532 17773 -1132
rect 17831 -2532 17971 -1132
rect 18029 -2532 18169 -1132
rect 18227 -2532 18367 -1132
rect 18425 -2532 18565 -1132
rect 18623 -2532 18763 -1132
rect 18821 -2532 18961 -1132
rect 19019 -2532 19159 -1132
rect 19217 -2532 19357 -1132
rect 19415 -2532 19555 -1132
rect 19613 -2532 19753 -1132
rect 11495 -4733 11635 -3333
rect 11693 -4733 11833 -3333
rect 11891 -4733 12031 -3333
rect 12089 -4733 12229 -3333
rect 12287 -4733 12427 -3333
rect 12485 -4733 12625 -3333
rect 12683 -4733 12823 -3333
rect 12881 -4733 13021 -3333
rect 13079 -4733 13219 -3333
rect 13277 -4733 13417 -3333
rect 13475 -4733 13615 -3333
rect 13673 -4733 13813 -3333
rect 13871 -4733 14011 -3333
rect 14069 -4733 14209 -3333
rect 14267 -4733 14407 -3333
rect 14465 -4733 14605 -3333
rect 14663 -4733 14803 -3333
rect 14861 -4733 15001 -3333
rect 15059 -4733 15199 -3333
rect 15257 -4733 15397 -3333
rect 15455 -4733 15595 -3333
rect 15653 -4733 15793 -3333
rect 15851 -4733 15991 -3333
rect 16049 -4733 16189 -3333
rect 16247 -4733 16387 -3333
rect 16445 -4733 16585 -3333
rect 16643 -4733 16783 -3333
rect 16841 -4733 16981 -3333
rect 17039 -4733 17179 -3333
rect 17237 -4733 17377 -3333
rect 17435 -4733 17575 -3333
rect 17633 -4733 17773 -3333
rect 17831 -4733 17971 -3333
rect 18029 -4733 18169 -3333
rect 18227 -4733 18367 -3333
rect 18425 -4733 18565 -3333
rect 18623 -4733 18763 -3333
rect 18821 -4733 18961 -3333
rect 19019 -4733 19159 -3333
rect 19217 -4733 19357 -3333
rect 19415 -4733 19555 -3333
rect 19613 -4733 19753 -3333
rect 23345 740 23485 2140
rect 23543 740 23683 2140
rect 23741 740 23881 2140
rect 23939 740 24079 2140
rect 24137 740 24277 2140
rect 24335 740 24475 2140
rect 24533 740 24673 2140
rect 24731 740 24871 2140
rect 24929 740 25069 2140
rect 25127 740 25267 2140
rect 25325 740 25465 2140
rect 25523 740 25663 2140
rect 25721 740 25861 2140
rect 25919 740 26059 2140
rect 26117 740 26257 2140
rect 26315 740 26455 2140
rect 26513 740 26653 2140
rect 26711 740 26851 2140
rect 26909 740 27049 2140
rect 27107 740 27247 2140
rect 27305 740 27445 2140
rect 27503 740 27643 2140
rect 27701 740 27841 2140
rect 27899 740 28039 2140
rect 28097 740 28237 2140
rect 28295 740 28435 2140
rect 28493 740 28633 2140
rect 28691 740 28831 2140
rect 28889 740 29029 2140
rect 29087 740 29227 2140
rect 29285 740 29425 2140
rect 29483 740 29623 2140
rect 29681 740 29821 2140
rect 29879 740 30019 2140
rect 30077 740 30217 2140
rect 30275 740 30415 2140
rect 30473 740 30613 2140
rect 30671 740 30811 2140
rect 30869 740 31009 2140
rect 31067 740 31207 2140
rect 31265 740 31405 2140
rect 31463 740 31603 2140
rect 23345 -896 23485 504
rect 23543 -896 23683 504
rect 23741 -896 23881 504
rect 23939 -896 24079 504
rect 24137 -896 24277 504
rect 24335 -896 24475 504
rect 24533 -896 24673 504
rect 24731 -896 24871 504
rect 24929 -896 25069 504
rect 25127 -896 25267 504
rect 25325 -896 25465 504
rect 25523 -896 25663 504
rect 25721 -896 25861 504
rect 25919 -896 26059 504
rect 26117 -896 26257 504
rect 26315 -896 26455 504
rect 26513 -896 26653 504
rect 26711 -896 26851 504
rect 26909 -896 27049 504
rect 27107 -896 27247 504
rect 27305 -896 27445 504
rect 27503 -896 27643 504
rect 27701 -896 27841 504
rect 27899 -896 28039 504
rect 28097 -896 28237 504
rect 28295 -896 28435 504
rect 28493 -896 28633 504
rect 28691 -896 28831 504
rect 28889 -896 29029 504
rect 29087 -896 29227 504
rect 29285 -896 29425 504
rect 29483 -896 29623 504
rect 29681 -896 29821 504
rect 29879 -896 30019 504
rect 30077 -896 30217 504
rect 30275 -896 30415 504
rect 30473 -896 30613 504
rect 30671 -896 30811 504
rect 30869 -896 31009 504
rect 31067 -896 31207 504
rect 31265 -896 31405 504
rect 31463 -896 31603 504
rect 23345 -2532 23485 -1132
rect 23543 -2532 23683 -1132
rect 23741 -2532 23881 -1132
rect 23939 -2532 24079 -1132
rect 24137 -2532 24277 -1132
rect 24335 -2532 24475 -1132
rect 24533 -2532 24673 -1132
rect 24731 -2532 24871 -1132
rect 24929 -2532 25069 -1132
rect 25127 -2532 25267 -1132
rect 25325 -2532 25465 -1132
rect 25523 -2532 25663 -1132
rect 25721 -2532 25861 -1132
rect 25919 -2532 26059 -1132
rect 26117 -2532 26257 -1132
rect 26315 -2532 26455 -1132
rect 26513 -2532 26653 -1132
rect 26711 -2532 26851 -1132
rect 26909 -2532 27049 -1132
rect 27107 -2532 27247 -1132
rect 27305 -2532 27445 -1132
rect 27503 -2532 27643 -1132
rect 27701 -2532 27841 -1132
rect 27899 -2532 28039 -1132
rect 28097 -2532 28237 -1132
rect 28295 -2532 28435 -1132
rect 28493 -2532 28633 -1132
rect 28691 -2532 28831 -1132
rect 28889 -2532 29029 -1132
rect 29087 -2532 29227 -1132
rect 29285 -2532 29425 -1132
rect 29483 -2532 29623 -1132
rect 29681 -2532 29821 -1132
rect 29879 -2532 30019 -1132
rect 30077 -2532 30217 -1132
rect 30275 -2532 30415 -1132
rect 30473 -2532 30613 -1132
rect 30671 -2532 30811 -1132
rect 30869 -2532 31009 -1132
rect 31067 -2532 31207 -1132
rect 31265 -2532 31405 -1132
rect 31463 -2532 31603 -1132
rect 23345 -4733 23485 -3333
rect 23543 -4733 23683 -3333
rect 23741 -4733 23881 -3333
rect 23939 -4733 24079 -3333
rect 24137 -4733 24277 -3333
rect 24335 -4733 24475 -3333
rect 24533 -4733 24673 -3333
rect 24731 -4733 24871 -3333
rect 24929 -4733 25069 -3333
rect 25127 -4733 25267 -3333
rect 25325 -4733 25465 -3333
rect 25523 -4733 25663 -3333
rect 25721 -4733 25861 -3333
rect 25919 -4733 26059 -3333
rect 26117 -4733 26257 -3333
rect 26315 -4733 26455 -3333
rect 26513 -4733 26653 -3333
rect 26711 -4733 26851 -3333
rect 26909 -4733 27049 -3333
rect 27107 -4733 27247 -3333
rect 27305 -4733 27445 -3333
rect 27503 -4733 27643 -3333
rect 27701 -4733 27841 -3333
rect 27899 -4733 28039 -3333
rect 28097 -4733 28237 -3333
rect 28295 -4733 28435 -3333
rect 28493 -4733 28633 -3333
rect 28691 -4733 28831 -3333
rect 28889 -4733 29029 -3333
rect 29087 -4733 29227 -3333
rect 29285 -4733 29425 -3333
rect 29483 -4733 29623 -3333
rect 29681 -4733 29821 -3333
rect 29879 -4733 30019 -3333
rect 30077 -4733 30217 -3333
rect 30275 -4733 30415 -3333
rect 30473 -4733 30613 -3333
rect 30671 -4733 30811 -3333
rect 30869 -4733 31009 -3333
rect 31067 -4733 31207 -3333
rect 31265 -4733 31405 -3333
rect 31463 -4733 31603 -3333
<< pdiff >>
rect 11437 2128 11495 2140
rect 11437 752 11449 2128
rect 11483 752 11495 2128
rect 11437 740 11495 752
rect 11635 2128 11693 2140
rect 11635 752 11647 2128
rect 11681 752 11693 2128
rect 11635 740 11693 752
rect 11833 2128 11891 2140
rect 11833 752 11845 2128
rect 11879 752 11891 2128
rect 11833 740 11891 752
rect 12031 2128 12089 2140
rect 12031 752 12043 2128
rect 12077 752 12089 2128
rect 12031 740 12089 752
rect 12229 2128 12287 2140
rect 12229 752 12241 2128
rect 12275 752 12287 2128
rect 12229 740 12287 752
rect 12427 2128 12485 2140
rect 12427 752 12439 2128
rect 12473 752 12485 2128
rect 12427 740 12485 752
rect 12625 2128 12683 2140
rect 12625 752 12637 2128
rect 12671 752 12683 2128
rect 12625 740 12683 752
rect 12823 2128 12881 2140
rect 12823 752 12835 2128
rect 12869 752 12881 2128
rect 12823 740 12881 752
rect 13021 2128 13079 2140
rect 13021 752 13033 2128
rect 13067 752 13079 2128
rect 13021 740 13079 752
rect 13219 2128 13277 2140
rect 13219 752 13231 2128
rect 13265 752 13277 2128
rect 13219 740 13277 752
rect 13417 2128 13475 2140
rect 13417 752 13429 2128
rect 13463 752 13475 2128
rect 13417 740 13475 752
rect 13615 2128 13673 2140
rect 13615 752 13627 2128
rect 13661 752 13673 2128
rect 13615 740 13673 752
rect 13813 2128 13871 2140
rect 13813 752 13825 2128
rect 13859 752 13871 2128
rect 13813 740 13871 752
rect 14011 2128 14069 2140
rect 14011 752 14023 2128
rect 14057 752 14069 2128
rect 14011 740 14069 752
rect 14209 2128 14267 2140
rect 14209 752 14221 2128
rect 14255 752 14267 2128
rect 14209 740 14267 752
rect 14407 2128 14465 2140
rect 14407 752 14419 2128
rect 14453 752 14465 2128
rect 14407 740 14465 752
rect 14605 2128 14663 2140
rect 14605 752 14617 2128
rect 14651 752 14663 2128
rect 14605 740 14663 752
rect 14803 2128 14861 2140
rect 14803 752 14815 2128
rect 14849 752 14861 2128
rect 14803 740 14861 752
rect 15001 2128 15059 2140
rect 15001 752 15013 2128
rect 15047 752 15059 2128
rect 15001 740 15059 752
rect 15199 2128 15257 2140
rect 15199 752 15211 2128
rect 15245 752 15257 2128
rect 15199 740 15257 752
rect 15397 2128 15455 2140
rect 15397 752 15409 2128
rect 15443 752 15455 2128
rect 15397 740 15455 752
rect 15595 2128 15653 2140
rect 15595 752 15607 2128
rect 15641 752 15653 2128
rect 15595 740 15653 752
rect 15793 2128 15851 2140
rect 15793 752 15805 2128
rect 15839 752 15851 2128
rect 15793 740 15851 752
rect 15991 2128 16049 2140
rect 15991 752 16003 2128
rect 16037 752 16049 2128
rect 15991 740 16049 752
rect 16189 2128 16247 2140
rect 16189 752 16201 2128
rect 16235 752 16247 2128
rect 16189 740 16247 752
rect 16387 2128 16445 2140
rect 16387 752 16399 2128
rect 16433 752 16445 2128
rect 16387 740 16445 752
rect 16585 2128 16643 2140
rect 16585 752 16597 2128
rect 16631 752 16643 2128
rect 16585 740 16643 752
rect 16783 2128 16841 2140
rect 16783 752 16795 2128
rect 16829 752 16841 2128
rect 16783 740 16841 752
rect 16981 2128 17039 2140
rect 16981 752 16993 2128
rect 17027 752 17039 2128
rect 16981 740 17039 752
rect 17179 2128 17237 2140
rect 17179 752 17191 2128
rect 17225 752 17237 2128
rect 17179 740 17237 752
rect 17377 2128 17435 2140
rect 17377 752 17389 2128
rect 17423 752 17435 2128
rect 17377 740 17435 752
rect 17575 2128 17633 2140
rect 17575 752 17587 2128
rect 17621 752 17633 2128
rect 17575 740 17633 752
rect 17773 2128 17831 2140
rect 17773 752 17785 2128
rect 17819 752 17831 2128
rect 17773 740 17831 752
rect 17971 2128 18029 2140
rect 17971 752 17983 2128
rect 18017 752 18029 2128
rect 17971 740 18029 752
rect 18169 2128 18227 2140
rect 18169 752 18181 2128
rect 18215 752 18227 2128
rect 18169 740 18227 752
rect 18367 2128 18425 2140
rect 18367 752 18379 2128
rect 18413 752 18425 2128
rect 18367 740 18425 752
rect 18565 2128 18623 2140
rect 18565 752 18577 2128
rect 18611 752 18623 2128
rect 18565 740 18623 752
rect 18763 2128 18821 2140
rect 18763 752 18775 2128
rect 18809 752 18821 2128
rect 18763 740 18821 752
rect 18961 2128 19019 2140
rect 18961 752 18973 2128
rect 19007 752 19019 2128
rect 18961 740 19019 752
rect 19159 2128 19217 2140
rect 19159 752 19171 2128
rect 19205 752 19217 2128
rect 19159 740 19217 752
rect 19357 2128 19415 2140
rect 19357 752 19369 2128
rect 19403 752 19415 2128
rect 19357 740 19415 752
rect 19555 2128 19613 2140
rect 19555 752 19567 2128
rect 19601 752 19613 2128
rect 19555 740 19613 752
rect 19753 2128 19811 2140
rect 19753 752 19765 2128
rect 19799 752 19811 2128
rect 19753 740 19811 752
rect 11437 492 11495 504
rect 11437 -884 11449 492
rect 11483 -884 11495 492
rect 11437 -896 11495 -884
rect 11635 492 11693 504
rect 11635 -884 11647 492
rect 11681 -884 11693 492
rect 11635 -896 11693 -884
rect 11833 492 11891 504
rect 11833 -884 11845 492
rect 11879 -884 11891 492
rect 11833 -896 11891 -884
rect 12031 492 12089 504
rect 12031 -884 12043 492
rect 12077 -884 12089 492
rect 12031 -896 12089 -884
rect 12229 492 12287 504
rect 12229 -884 12241 492
rect 12275 -884 12287 492
rect 12229 -896 12287 -884
rect 12427 492 12485 504
rect 12427 -884 12439 492
rect 12473 -884 12485 492
rect 12427 -896 12485 -884
rect 12625 492 12683 504
rect 12625 -884 12637 492
rect 12671 -884 12683 492
rect 12625 -896 12683 -884
rect 12823 492 12881 504
rect 12823 -884 12835 492
rect 12869 -884 12881 492
rect 12823 -896 12881 -884
rect 13021 492 13079 504
rect 13021 -884 13033 492
rect 13067 -884 13079 492
rect 13021 -896 13079 -884
rect 13219 492 13277 504
rect 13219 -884 13231 492
rect 13265 -884 13277 492
rect 13219 -896 13277 -884
rect 13417 492 13475 504
rect 13417 -884 13429 492
rect 13463 -884 13475 492
rect 13417 -896 13475 -884
rect 13615 492 13673 504
rect 13615 -884 13627 492
rect 13661 -884 13673 492
rect 13615 -896 13673 -884
rect 13813 492 13871 504
rect 13813 -884 13825 492
rect 13859 -884 13871 492
rect 13813 -896 13871 -884
rect 14011 492 14069 504
rect 14011 -884 14023 492
rect 14057 -884 14069 492
rect 14011 -896 14069 -884
rect 14209 492 14267 504
rect 14209 -884 14221 492
rect 14255 -884 14267 492
rect 14209 -896 14267 -884
rect 14407 492 14465 504
rect 14407 -884 14419 492
rect 14453 -884 14465 492
rect 14407 -896 14465 -884
rect 14605 492 14663 504
rect 14605 -884 14617 492
rect 14651 -884 14663 492
rect 14605 -896 14663 -884
rect 14803 492 14861 504
rect 14803 -884 14815 492
rect 14849 -884 14861 492
rect 14803 -896 14861 -884
rect 15001 492 15059 504
rect 15001 -884 15013 492
rect 15047 -884 15059 492
rect 15001 -896 15059 -884
rect 15199 492 15257 504
rect 15199 -884 15211 492
rect 15245 -884 15257 492
rect 15199 -896 15257 -884
rect 15397 492 15455 504
rect 15397 -884 15409 492
rect 15443 -884 15455 492
rect 15397 -896 15455 -884
rect 15595 492 15653 504
rect 15595 -884 15607 492
rect 15641 -884 15653 492
rect 15595 -896 15653 -884
rect 15793 492 15851 504
rect 15793 -884 15805 492
rect 15839 -884 15851 492
rect 15793 -896 15851 -884
rect 15991 492 16049 504
rect 15991 -884 16003 492
rect 16037 -884 16049 492
rect 15991 -896 16049 -884
rect 16189 492 16247 504
rect 16189 -884 16201 492
rect 16235 -884 16247 492
rect 16189 -896 16247 -884
rect 16387 492 16445 504
rect 16387 -884 16399 492
rect 16433 -884 16445 492
rect 16387 -896 16445 -884
rect 16585 492 16643 504
rect 16585 -884 16597 492
rect 16631 -884 16643 492
rect 16585 -896 16643 -884
rect 16783 492 16841 504
rect 16783 -884 16795 492
rect 16829 -884 16841 492
rect 16783 -896 16841 -884
rect 16981 492 17039 504
rect 16981 -884 16993 492
rect 17027 -884 17039 492
rect 16981 -896 17039 -884
rect 17179 492 17237 504
rect 17179 -884 17191 492
rect 17225 -884 17237 492
rect 17179 -896 17237 -884
rect 17377 492 17435 504
rect 17377 -884 17389 492
rect 17423 -884 17435 492
rect 17377 -896 17435 -884
rect 17575 492 17633 504
rect 17575 -884 17587 492
rect 17621 -884 17633 492
rect 17575 -896 17633 -884
rect 17773 492 17831 504
rect 17773 -884 17785 492
rect 17819 -884 17831 492
rect 17773 -896 17831 -884
rect 17971 492 18029 504
rect 17971 -884 17983 492
rect 18017 -884 18029 492
rect 17971 -896 18029 -884
rect 18169 492 18227 504
rect 18169 -884 18181 492
rect 18215 -884 18227 492
rect 18169 -896 18227 -884
rect 18367 492 18425 504
rect 18367 -884 18379 492
rect 18413 -884 18425 492
rect 18367 -896 18425 -884
rect 18565 492 18623 504
rect 18565 -884 18577 492
rect 18611 -884 18623 492
rect 18565 -896 18623 -884
rect 18763 492 18821 504
rect 18763 -884 18775 492
rect 18809 -884 18821 492
rect 18763 -896 18821 -884
rect 18961 492 19019 504
rect 18961 -884 18973 492
rect 19007 -884 19019 492
rect 18961 -896 19019 -884
rect 19159 492 19217 504
rect 19159 -884 19171 492
rect 19205 -884 19217 492
rect 19159 -896 19217 -884
rect 19357 492 19415 504
rect 19357 -884 19369 492
rect 19403 -884 19415 492
rect 19357 -896 19415 -884
rect 19555 492 19613 504
rect 19555 -884 19567 492
rect 19601 -884 19613 492
rect 19555 -896 19613 -884
rect 19753 492 19811 504
rect 19753 -884 19765 492
rect 19799 -884 19811 492
rect 19753 -896 19811 -884
rect 11437 -1144 11495 -1132
rect 11437 -2520 11449 -1144
rect 11483 -2520 11495 -1144
rect 11437 -2532 11495 -2520
rect 11635 -1144 11693 -1132
rect 11635 -2520 11647 -1144
rect 11681 -2520 11693 -1144
rect 11635 -2532 11693 -2520
rect 11833 -1144 11891 -1132
rect 11833 -2520 11845 -1144
rect 11879 -2520 11891 -1144
rect 11833 -2532 11891 -2520
rect 12031 -1144 12089 -1132
rect 12031 -2520 12043 -1144
rect 12077 -2520 12089 -1144
rect 12031 -2532 12089 -2520
rect 12229 -1144 12287 -1132
rect 12229 -2520 12241 -1144
rect 12275 -2520 12287 -1144
rect 12229 -2532 12287 -2520
rect 12427 -1144 12485 -1132
rect 12427 -2520 12439 -1144
rect 12473 -2520 12485 -1144
rect 12427 -2532 12485 -2520
rect 12625 -1144 12683 -1132
rect 12625 -2520 12637 -1144
rect 12671 -2520 12683 -1144
rect 12625 -2532 12683 -2520
rect 12823 -1144 12881 -1132
rect 12823 -2520 12835 -1144
rect 12869 -2520 12881 -1144
rect 12823 -2532 12881 -2520
rect 13021 -1144 13079 -1132
rect 13021 -2520 13033 -1144
rect 13067 -2520 13079 -1144
rect 13021 -2532 13079 -2520
rect 13219 -1144 13277 -1132
rect 13219 -2520 13231 -1144
rect 13265 -2520 13277 -1144
rect 13219 -2532 13277 -2520
rect 13417 -1144 13475 -1132
rect 13417 -2520 13429 -1144
rect 13463 -2520 13475 -1144
rect 13417 -2532 13475 -2520
rect 13615 -1144 13673 -1132
rect 13615 -2520 13627 -1144
rect 13661 -2520 13673 -1144
rect 13615 -2532 13673 -2520
rect 13813 -1144 13871 -1132
rect 13813 -2520 13825 -1144
rect 13859 -2520 13871 -1144
rect 13813 -2532 13871 -2520
rect 14011 -1144 14069 -1132
rect 14011 -2520 14023 -1144
rect 14057 -2520 14069 -1144
rect 14011 -2532 14069 -2520
rect 14209 -1144 14267 -1132
rect 14209 -2520 14221 -1144
rect 14255 -2520 14267 -1144
rect 14209 -2532 14267 -2520
rect 14407 -1144 14465 -1132
rect 14407 -2520 14419 -1144
rect 14453 -2520 14465 -1144
rect 14407 -2532 14465 -2520
rect 14605 -1144 14663 -1132
rect 14605 -2520 14617 -1144
rect 14651 -2520 14663 -1144
rect 14605 -2532 14663 -2520
rect 14803 -1144 14861 -1132
rect 14803 -2520 14815 -1144
rect 14849 -2520 14861 -1144
rect 14803 -2532 14861 -2520
rect 15001 -1144 15059 -1132
rect 15001 -2520 15013 -1144
rect 15047 -2520 15059 -1144
rect 15001 -2532 15059 -2520
rect 15199 -1144 15257 -1132
rect 15199 -2520 15211 -1144
rect 15245 -2520 15257 -1144
rect 15199 -2532 15257 -2520
rect 15397 -1144 15455 -1132
rect 15397 -2520 15409 -1144
rect 15443 -2520 15455 -1144
rect 15397 -2532 15455 -2520
rect 15595 -1144 15653 -1132
rect 15595 -2520 15607 -1144
rect 15641 -2520 15653 -1144
rect 15595 -2532 15653 -2520
rect 15793 -1144 15851 -1132
rect 15793 -2520 15805 -1144
rect 15839 -2520 15851 -1144
rect 15793 -2532 15851 -2520
rect 15991 -1144 16049 -1132
rect 15991 -2520 16003 -1144
rect 16037 -2520 16049 -1144
rect 15991 -2532 16049 -2520
rect 16189 -1144 16247 -1132
rect 16189 -2520 16201 -1144
rect 16235 -2520 16247 -1144
rect 16189 -2532 16247 -2520
rect 16387 -1144 16445 -1132
rect 16387 -2520 16399 -1144
rect 16433 -2520 16445 -1144
rect 16387 -2532 16445 -2520
rect 16585 -1144 16643 -1132
rect 16585 -2520 16597 -1144
rect 16631 -2520 16643 -1144
rect 16585 -2532 16643 -2520
rect 16783 -1144 16841 -1132
rect 16783 -2520 16795 -1144
rect 16829 -2520 16841 -1144
rect 16783 -2532 16841 -2520
rect 16981 -1144 17039 -1132
rect 16981 -2520 16993 -1144
rect 17027 -2520 17039 -1144
rect 16981 -2532 17039 -2520
rect 17179 -1144 17237 -1132
rect 17179 -2520 17191 -1144
rect 17225 -2520 17237 -1144
rect 17179 -2532 17237 -2520
rect 17377 -1144 17435 -1132
rect 17377 -2520 17389 -1144
rect 17423 -2520 17435 -1144
rect 17377 -2532 17435 -2520
rect 17575 -1144 17633 -1132
rect 17575 -2520 17587 -1144
rect 17621 -2520 17633 -1144
rect 17575 -2532 17633 -2520
rect 17773 -1144 17831 -1132
rect 17773 -2520 17785 -1144
rect 17819 -2520 17831 -1144
rect 17773 -2532 17831 -2520
rect 17971 -1144 18029 -1132
rect 17971 -2520 17983 -1144
rect 18017 -2520 18029 -1144
rect 17971 -2532 18029 -2520
rect 18169 -1144 18227 -1132
rect 18169 -2520 18181 -1144
rect 18215 -2520 18227 -1144
rect 18169 -2532 18227 -2520
rect 18367 -1144 18425 -1132
rect 18367 -2520 18379 -1144
rect 18413 -2520 18425 -1144
rect 18367 -2532 18425 -2520
rect 18565 -1144 18623 -1132
rect 18565 -2520 18577 -1144
rect 18611 -2520 18623 -1144
rect 18565 -2532 18623 -2520
rect 18763 -1144 18821 -1132
rect 18763 -2520 18775 -1144
rect 18809 -2520 18821 -1144
rect 18763 -2532 18821 -2520
rect 18961 -1144 19019 -1132
rect 18961 -2520 18973 -1144
rect 19007 -2520 19019 -1144
rect 18961 -2532 19019 -2520
rect 19159 -1144 19217 -1132
rect 19159 -2520 19171 -1144
rect 19205 -2520 19217 -1144
rect 19159 -2532 19217 -2520
rect 19357 -1144 19415 -1132
rect 19357 -2520 19369 -1144
rect 19403 -2520 19415 -1144
rect 19357 -2532 19415 -2520
rect 19555 -1144 19613 -1132
rect 19555 -2520 19567 -1144
rect 19601 -2520 19613 -1144
rect 19555 -2532 19613 -2520
rect 19753 -1144 19811 -1132
rect 19753 -2520 19765 -1144
rect 19799 -2520 19811 -1144
rect 19753 -2532 19811 -2520
rect 11437 -3345 11495 -3333
rect 11437 -4721 11449 -3345
rect 11483 -4721 11495 -3345
rect 11437 -4733 11495 -4721
rect 11635 -3345 11693 -3333
rect 11635 -4721 11647 -3345
rect 11681 -4721 11693 -3345
rect 11635 -4733 11693 -4721
rect 11833 -3345 11891 -3333
rect 11833 -4721 11845 -3345
rect 11879 -4721 11891 -3345
rect 11833 -4733 11891 -4721
rect 12031 -3345 12089 -3333
rect 12031 -4721 12043 -3345
rect 12077 -4721 12089 -3345
rect 12031 -4733 12089 -4721
rect 12229 -3345 12287 -3333
rect 12229 -4721 12241 -3345
rect 12275 -4721 12287 -3345
rect 12229 -4733 12287 -4721
rect 12427 -3345 12485 -3333
rect 12427 -4721 12439 -3345
rect 12473 -4721 12485 -3345
rect 12427 -4733 12485 -4721
rect 12625 -3345 12683 -3333
rect 12625 -4721 12637 -3345
rect 12671 -4721 12683 -3345
rect 12625 -4733 12683 -4721
rect 12823 -3345 12881 -3333
rect 12823 -4721 12835 -3345
rect 12869 -4721 12881 -3345
rect 12823 -4733 12881 -4721
rect 13021 -3345 13079 -3333
rect 13021 -4721 13033 -3345
rect 13067 -4721 13079 -3345
rect 13021 -4733 13079 -4721
rect 13219 -3345 13277 -3333
rect 13219 -4721 13231 -3345
rect 13265 -4721 13277 -3345
rect 13219 -4733 13277 -4721
rect 13417 -3345 13475 -3333
rect 13417 -4721 13429 -3345
rect 13463 -4721 13475 -3345
rect 13417 -4733 13475 -4721
rect 13615 -3345 13673 -3333
rect 13615 -4721 13627 -3345
rect 13661 -4721 13673 -3345
rect 13615 -4733 13673 -4721
rect 13813 -3345 13871 -3333
rect 13813 -4721 13825 -3345
rect 13859 -4721 13871 -3345
rect 13813 -4733 13871 -4721
rect 14011 -3345 14069 -3333
rect 14011 -4721 14023 -3345
rect 14057 -4721 14069 -3345
rect 14011 -4733 14069 -4721
rect 14209 -3345 14267 -3333
rect 14209 -4721 14221 -3345
rect 14255 -4721 14267 -3345
rect 14209 -4733 14267 -4721
rect 14407 -3345 14465 -3333
rect 14407 -4721 14419 -3345
rect 14453 -4721 14465 -3345
rect 14407 -4733 14465 -4721
rect 14605 -3345 14663 -3333
rect 14605 -4721 14617 -3345
rect 14651 -4721 14663 -3345
rect 14605 -4733 14663 -4721
rect 14803 -3345 14861 -3333
rect 14803 -4721 14815 -3345
rect 14849 -4721 14861 -3345
rect 14803 -4733 14861 -4721
rect 15001 -3345 15059 -3333
rect 15001 -4721 15013 -3345
rect 15047 -4721 15059 -3345
rect 15001 -4733 15059 -4721
rect 15199 -3345 15257 -3333
rect 15199 -4721 15211 -3345
rect 15245 -4721 15257 -3345
rect 15199 -4733 15257 -4721
rect 15397 -3345 15455 -3333
rect 15397 -4721 15409 -3345
rect 15443 -4721 15455 -3345
rect 15397 -4733 15455 -4721
rect 15595 -3345 15653 -3333
rect 15595 -4721 15607 -3345
rect 15641 -4721 15653 -3345
rect 15595 -4733 15653 -4721
rect 15793 -3345 15851 -3333
rect 15793 -4721 15805 -3345
rect 15839 -4721 15851 -3345
rect 15793 -4733 15851 -4721
rect 15991 -3345 16049 -3333
rect 15991 -4721 16003 -3345
rect 16037 -4721 16049 -3345
rect 15991 -4733 16049 -4721
rect 16189 -3345 16247 -3333
rect 16189 -4721 16201 -3345
rect 16235 -4721 16247 -3345
rect 16189 -4733 16247 -4721
rect 16387 -3345 16445 -3333
rect 16387 -4721 16399 -3345
rect 16433 -4721 16445 -3345
rect 16387 -4733 16445 -4721
rect 16585 -3345 16643 -3333
rect 16585 -4721 16597 -3345
rect 16631 -4721 16643 -3345
rect 16585 -4733 16643 -4721
rect 16783 -3345 16841 -3333
rect 16783 -4721 16795 -3345
rect 16829 -4721 16841 -3345
rect 16783 -4733 16841 -4721
rect 16981 -3345 17039 -3333
rect 16981 -4721 16993 -3345
rect 17027 -4721 17039 -3345
rect 16981 -4733 17039 -4721
rect 17179 -3345 17237 -3333
rect 17179 -4721 17191 -3345
rect 17225 -4721 17237 -3345
rect 17179 -4733 17237 -4721
rect 17377 -3345 17435 -3333
rect 17377 -4721 17389 -3345
rect 17423 -4721 17435 -3345
rect 17377 -4733 17435 -4721
rect 17575 -3345 17633 -3333
rect 17575 -4721 17587 -3345
rect 17621 -4721 17633 -3345
rect 17575 -4733 17633 -4721
rect 17773 -3345 17831 -3333
rect 17773 -4721 17785 -3345
rect 17819 -4721 17831 -3345
rect 17773 -4733 17831 -4721
rect 17971 -3345 18029 -3333
rect 17971 -4721 17983 -3345
rect 18017 -4721 18029 -3345
rect 17971 -4733 18029 -4721
rect 18169 -3345 18227 -3333
rect 18169 -4721 18181 -3345
rect 18215 -4721 18227 -3345
rect 18169 -4733 18227 -4721
rect 18367 -3345 18425 -3333
rect 18367 -4721 18379 -3345
rect 18413 -4721 18425 -3345
rect 18367 -4733 18425 -4721
rect 18565 -3345 18623 -3333
rect 18565 -4721 18577 -3345
rect 18611 -4721 18623 -3345
rect 18565 -4733 18623 -4721
rect 18763 -3345 18821 -3333
rect 18763 -4721 18775 -3345
rect 18809 -4721 18821 -3345
rect 18763 -4733 18821 -4721
rect 18961 -3345 19019 -3333
rect 18961 -4721 18973 -3345
rect 19007 -4721 19019 -3345
rect 18961 -4733 19019 -4721
rect 19159 -3345 19217 -3333
rect 19159 -4721 19171 -3345
rect 19205 -4721 19217 -3345
rect 19159 -4733 19217 -4721
rect 19357 -3345 19415 -3333
rect 19357 -4721 19369 -3345
rect 19403 -4721 19415 -3345
rect 19357 -4733 19415 -4721
rect 19555 -3345 19613 -3333
rect 19555 -4721 19567 -3345
rect 19601 -4721 19613 -3345
rect 19555 -4733 19613 -4721
rect 19753 -3345 19811 -3333
rect 19753 -4721 19765 -3345
rect 19799 -4721 19811 -3345
rect 19753 -4733 19811 -4721
rect 23287 2128 23345 2140
rect 23287 752 23299 2128
rect 23333 752 23345 2128
rect 23287 740 23345 752
rect 23485 2128 23543 2140
rect 23485 752 23497 2128
rect 23531 752 23543 2128
rect 23485 740 23543 752
rect 23683 2128 23741 2140
rect 23683 752 23695 2128
rect 23729 752 23741 2128
rect 23683 740 23741 752
rect 23881 2128 23939 2140
rect 23881 752 23893 2128
rect 23927 752 23939 2128
rect 23881 740 23939 752
rect 24079 2128 24137 2140
rect 24079 752 24091 2128
rect 24125 752 24137 2128
rect 24079 740 24137 752
rect 24277 2128 24335 2140
rect 24277 752 24289 2128
rect 24323 752 24335 2128
rect 24277 740 24335 752
rect 24475 2128 24533 2140
rect 24475 752 24487 2128
rect 24521 752 24533 2128
rect 24475 740 24533 752
rect 24673 2128 24731 2140
rect 24673 752 24685 2128
rect 24719 752 24731 2128
rect 24673 740 24731 752
rect 24871 2128 24929 2140
rect 24871 752 24883 2128
rect 24917 752 24929 2128
rect 24871 740 24929 752
rect 25069 2128 25127 2140
rect 25069 752 25081 2128
rect 25115 752 25127 2128
rect 25069 740 25127 752
rect 25267 2128 25325 2140
rect 25267 752 25279 2128
rect 25313 752 25325 2128
rect 25267 740 25325 752
rect 25465 2128 25523 2140
rect 25465 752 25477 2128
rect 25511 752 25523 2128
rect 25465 740 25523 752
rect 25663 2128 25721 2140
rect 25663 752 25675 2128
rect 25709 752 25721 2128
rect 25663 740 25721 752
rect 25861 2128 25919 2140
rect 25861 752 25873 2128
rect 25907 752 25919 2128
rect 25861 740 25919 752
rect 26059 2128 26117 2140
rect 26059 752 26071 2128
rect 26105 752 26117 2128
rect 26059 740 26117 752
rect 26257 2128 26315 2140
rect 26257 752 26269 2128
rect 26303 752 26315 2128
rect 26257 740 26315 752
rect 26455 2128 26513 2140
rect 26455 752 26467 2128
rect 26501 752 26513 2128
rect 26455 740 26513 752
rect 26653 2128 26711 2140
rect 26653 752 26665 2128
rect 26699 752 26711 2128
rect 26653 740 26711 752
rect 26851 2128 26909 2140
rect 26851 752 26863 2128
rect 26897 752 26909 2128
rect 26851 740 26909 752
rect 27049 2128 27107 2140
rect 27049 752 27061 2128
rect 27095 752 27107 2128
rect 27049 740 27107 752
rect 27247 2128 27305 2140
rect 27247 752 27259 2128
rect 27293 752 27305 2128
rect 27247 740 27305 752
rect 27445 2128 27503 2140
rect 27445 752 27457 2128
rect 27491 752 27503 2128
rect 27445 740 27503 752
rect 27643 2128 27701 2140
rect 27643 752 27655 2128
rect 27689 752 27701 2128
rect 27643 740 27701 752
rect 27841 2128 27899 2140
rect 27841 752 27853 2128
rect 27887 752 27899 2128
rect 27841 740 27899 752
rect 28039 2128 28097 2140
rect 28039 752 28051 2128
rect 28085 752 28097 2128
rect 28039 740 28097 752
rect 28237 2128 28295 2140
rect 28237 752 28249 2128
rect 28283 752 28295 2128
rect 28237 740 28295 752
rect 28435 2128 28493 2140
rect 28435 752 28447 2128
rect 28481 752 28493 2128
rect 28435 740 28493 752
rect 28633 2128 28691 2140
rect 28633 752 28645 2128
rect 28679 752 28691 2128
rect 28633 740 28691 752
rect 28831 2128 28889 2140
rect 28831 752 28843 2128
rect 28877 752 28889 2128
rect 28831 740 28889 752
rect 29029 2128 29087 2140
rect 29029 752 29041 2128
rect 29075 752 29087 2128
rect 29029 740 29087 752
rect 29227 2128 29285 2140
rect 29227 752 29239 2128
rect 29273 752 29285 2128
rect 29227 740 29285 752
rect 29425 2128 29483 2140
rect 29425 752 29437 2128
rect 29471 752 29483 2128
rect 29425 740 29483 752
rect 29623 2128 29681 2140
rect 29623 752 29635 2128
rect 29669 752 29681 2128
rect 29623 740 29681 752
rect 29821 2128 29879 2140
rect 29821 752 29833 2128
rect 29867 752 29879 2128
rect 29821 740 29879 752
rect 30019 2128 30077 2140
rect 30019 752 30031 2128
rect 30065 752 30077 2128
rect 30019 740 30077 752
rect 30217 2128 30275 2140
rect 30217 752 30229 2128
rect 30263 752 30275 2128
rect 30217 740 30275 752
rect 30415 2128 30473 2140
rect 30415 752 30427 2128
rect 30461 752 30473 2128
rect 30415 740 30473 752
rect 30613 2128 30671 2140
rect 30613 752 30625 2128
rect 30659 752 30671 2128
rect 30613 740 30671 752
rect 30811 2128 30869 2140
rect 30811 752 30823 2128
rect 30857 752 30869 2128
rect 30811 740 30869 752
rect 31009 2128 31067 2140
rect 31009 752 31021 2128
rect 31055 752 31067 2128
rect 31009 740 31067 752
rect 31207 2128 31265 2140
rect 31207 752 31219 2128
rect 31253 752 31265 2128
rect 31207 740 31265 752
rect 31405 2128 31463 2140
rect 31405 752 31417 2128
rect 31451 752 31463 2128
rect 31405 740 31463 752
rect 31603 2128 31661 2140
rect 31603 752 31615 2128
rect 31649 752 31661 2128
rect 31603 740 31661 752
rect 23287 492 23345 504
rect 23287 -884 23299 492
rect 23333 -884 23345 492
rect 23287 -896 23345 -884
rect 23485 492 23543 504
rect 23485 -884 23497 492
rect 23531 -884 23543 492
rect 23485 -896 23543 -884
rect 23683 492 23741 504
rect 23683 -884 23695 492
rect 23729 -884 23741 492
rect 23683 -896 23741 -884
rect 23881 492 23939 504
rect 23881 -884 23893 492
rect 23927 -884 23939 492
rect 23881 -896 23939 -884
rect 24079 492 24137 504
rect 24079 -884 24091 492
rect 24125 -884 24137 492
rect 24079 -896 24137 -884
rect 24277 492 24335 504
rect 24277 -884 24289 492
rect 24323 -884 24335 492
rect 24277 -896 24335 -884
rect 24475 492 24533 504
rect 24475 -884 24487 492
rect 24521 -884 24533 492
rect 24475 -896 24533 -884
rect 24673 492 24731 504
rect 24673 -884 24685 492
rect 24719 -884 24731 492
rect 24673 -896 24731 -884
rect 24871 492 24929 504
rect 24871 -884 24883 492
rect 24917 -884 24929 492
rect 24871 -896 24929 -884
rect 25069 492 25127 504
rect 25069 -884 25081 492
rect 25115 -884 25127 492
rect 25069 -896 25127 -884
rect 25267 492 25325 504
rect 25267 -884 25279 492
rect 25313 -884 25325 492
rect 25267 -896 25325 -884
rect 25465 492 25523 504
rect 25465 -884 25477 492
rect 25511 -884 25523 492
rect 25465 -896 25523 -884
rect 25663 492 25721 504
rect 25663 -884 25675 492
rect 25709 -884 25721 492
rect 25663 -896 25721 -884
rect 25861 492 25919 504
rect 25861 -884 25873 492
rect 25907 -884 25919 492
rect 25861 -896 25919 -884
rect 26059 492 26117 504
rect 26059 -884 26071 492
rect 26105 -884 26117 492
rect 26059 -896 26117 -884
rect 26257 492 26315 504
rect 26257 -884 26269 492
rect 26303 -884 26315 492
rect 26257 -896 26315 -884
rect 26455 492 26513 504
rect 26455 -884 26467 492
rect 26501 -884 26513 492
rect 26455 -896 26513 -884
rect 26653 492 26711 504
rect 26653 -884 26665 492
rect 26699 -884 26711 492
rect 26653 -896 26711 -884
rect 26851 492 26909 504
rect 26851 -884 26863 492
rect 26897 -884 26909 492
rect 26851 -896 26909 -884
rect 27049 492 27107 504
rect 27049 -884 27061 492
rect 27095 -884 27107 492
rect 27049 -896 27107 -884
rect 27247 492 27305 504
rect 27247 -884 27259 492
rect 27293 -884 27305 492
rect 27247 -896 27305 -884
rect 27445 492 27503 504
rect 27445 -884 27457 492
rect 27491 -884 27503 492
rect 27445 -896 27503 -884
rect 27643 492 27701 504
rect 27643 -884 27655 492
rect 27689 -884 27701 492
rect 27643 -896 27701 -884
rect 27841 492 27899 504
rect 27841 -884 27853 492
rect 27887 -884 27899 492
rect 27841 -896 27899 -884
rect 28039 492 28097 504
rect 28039 -884 28051 492
rect 28085 -884 28097 492
rect 28039 -896 28097 -884
rect 28237 492 28295 504
rect 28237 -884 28249 492
rect 28283 -884 28295 492
rect 28237 -896 28295 -884
rect 28435 492 28493 504
rect 28435 -884 28447 492
rect 28481 -884 28493 492
rect 28435 -896 28493 -884
rect 28633 492 28691 504
rect 28633 -884 28645 492
rect 28679 -884 28691 492
rect 28633 -896 28691 -884
rect 28831 492 28889 504
rect 28831 -884 28843 492
rect 28877 -884 28889 492
rect 28831 -896 28889 -884
rect 29029 492 29087 504
rect 29029 -884 29041 492
rect 29075 -884 29087 492
rect 29029 -896 29087 -884
rect 29227 492 29285 504
rect 29227 -884 29239 492
rect 29273 -884 29285 492
rect 29227 -896 29285 -884
rect 29425 492 29483 504
rect 29425 -884 29437 492
rect 29471 -884 29483 492
rect 29425 -896 29483 -884
rect 29623 492 29681 504
rect 29623 -884 29635 492
rect 29669 -884 29681 492
rect 29623 -896 29681 -884
rect 29821 492 29879 504
rect 29821 -884 29833 492
rect 29867 -884 29879 492
rect 29821 -896 29879 -884
rect 30019 492 30077 504
rect 30019 -884 30031 492
rect 30065 -884 30077 492
rect 30019 -896 30077 -884
rect 30217 492 30275 504
rect 30217 -884 30229 492
rect 30263 -884 30275 492
rect 30217 -896 30275 -884
rect 30415 492 30473 504
rect 30415 -884 30427 492
rect 30461 -884 30473 492
rect 30415 -896 30473 -884
rect 30613 492 30671 504
rect 30613 -884 30625 492
rect 30659 -884 30671 492
rect 30613 -896 30671 -884
rect 30811 492 30869 504
rect 30811 -884 30823 492
rect 30857 -884 30869 492
rect 30811 -896 30869 -884
rect 31009 492 31067 504
rect 31009 -884 31021 492
rect 31055 -884 31067 492
rect 31009 -896 31067 -884
rect 31207 492 31265 504
rect 31207 -884 31219 492
rect 31253 -884 31265 492
rect 31207 -896 31265 -884
rect 31405 492 31463 504
rect 31405 -884 31417 492
rect 31451 -884 31463 492
rect 31405 -896 31463 -884
rect 31603 492 31661 504
rect 31603 -884 31615 492
rect 31649 -884 31661 492
rect 31603 -896 31661 -884
rect 23287 -1144 23345 -1132
rect 23287 -2520 23299 -1144
rect 23333 -2520 23345 -1144
rect 23287 -2532 23345 -2520
rect 23485 -1144 23543 -1132
rect 23485 -2520 23497 -1144
rect 23531 -2520 23543 -1144
rect 23485 -2532 23543 -2520
rect 23683 -1144 23741 -1132
rect 23683 -2520 23695 -1144
rect 23729 -2520 23741 -1144
rect 23683 -2532 23741 -2520
rect 23881 -1144 23939 -1132
rect 23881 -2520 23893 -1144
rect 23927 -2520 23939 -1144
rect 23881 -2532 23939 -2520
rect 24079 -1144 24137 -1132
rect 24079 -2520 24091 -1144
rect 24125 -2520 24137 -1144
rect 24079 -2532 24137 -2520
rect 24277 -1144 24335 -1132
rect 24277 -2520 24289 -1144
rect 24323 -2520 24335 -1144
rect 24277 -2532 24335 -2520
rect 24475 -1144 24533 -1132
rect 24475 -2520 24487 -1144
rect 24521 -2520 24533 -1144
rect 24475 -2532 24533 -2520
rect 24673 -1144 24731 -1132
rect 24673 -2520 24685 -1144
rect 24719 -2520 24731 -1144
rect 24673 -2532 24731 -2520
rect 24871 -1144 24929 -1132
rect 24871 -2520 24883 -1144
rect 24917 -2520 24929 -1144
rect 24871 -2532 24929 -2520
rect 25069 -1144 25127 -1132
rect 25069 -2520 25081 -1144
rect 25115 -2520 25127 -1144
rect 25069 -2532 25127 -2520
rect 25267 -1144 25325 -1132
rect 25267 -2520 25279 -1144
rect 25313 -2520 25325 -1144
rect 25267 -2532 25325 -2520
rect 25465 -1144 25523 -1132
rect 25465 -2520 25477 -1144
rect 25511 -2520 25523 -1144
rect 25465 -2532 25523 -2520
rect 25663 -1144 25721 -1132
rect 25663 -2520 25675 -1144
rect 25709 -2520 25721 -1144
rect 25663 -2532 25721 -2520
rect 25861 -1144 25919 -1132
rect 25861 -2520 25873 -1144
rect 25907 -2520 25919 -1144
rect 25861 -2532 25919 -2520
rect 26059 -1144 26117 -1132
rect 26059 -2520 26071 -1144
rect 26105 -2520 26117 -1144
rect 26059 -2532 26117 -2520
rect 26257 -1144 26315 -1132
rect 26257 -2520 26269 -1144
rect 26303 -2520 26315 -1144
rect 26257 -2532 26315 -2520
rect 26455 -1144 26513 -1132
rect 26455 -2520 26467 -1144
rect 26501 -2520 26513 -1144
rect 26455 -2532 26513 -2520
rect 26653 -1144 26711 -1132
rect 26653 -2520 26665 -1144
rect 26699 -2520 26711 -1144
rect 26653 -2532 26711 -2520
rect 26851 -1144 26909 -1132
rect 26851 -2520 26863 -1144
rect 26897 -2520 26909 -1144
rect 26851 -2532 26909 -2520
rect 27049 -1144 27107 -1132
rect 27049 -2520 27061 -1144
rect 27095 -2520 27107 -1144
rect 27049 -2532 27107 -2520
rect 27247 -1144 27305 -1132
rect 27247 -2520 27259 -1144
rect 27293 -2520 27305 -1144
rect 27247 -2532 27305 -2520
rect 27445 -1144 27503 -1132
rect 27445 -2520 27457 -1144
rect 27491 -2520 27503 -1144
rect 27445 -2532 27503 -2520
rect 27643 -1144 27701 -1132
rect 27643 -2520 27655 -1144
rect 27689 -2520 27701 -1144
rect 27643 -2532 27701 -2520
rect 27841 -1144 27899 -1132
rect 27841 -2520 27853 -1144
rect 27887 -2520 27899 -1144
rect 27841 -2532 27899 -2520
rect 28039 -1144 28097 -1132
rect 28039 -2520 28051 -1144
rect 28085 -2520 28097 -1144
rect 28039 -2532 28097 -2520
rect 28237 -1144 28295 -1132
rect 28237 -2520 28249 -1144
rect 28283 -2520 28295 -1144
rect 28237 -2532 28295 -2520
rect 28435 -1144 28493 -1132
rect 28435 -2520 28447 -1144
rect 28481 -2520 28493 -1144
rect 28435 -2532 28493 -2520
rect 28633 -1144 28691 -1132
rect 28633 -2520 28645 -1144
rect 28679 -2520 28691 -1144
rect 28633 -2532 28691 -2520
rect 28831 -1144 28889 -1132
rect 28831 -2520 28843 -1144
rect 28877 -2520 28889 -1144
rect 28831 -2532 28889 -2520
rect 29029 -1144 29087 -1132
rect 29029 -2520 29041 -1144
rect 29075 -2520 29087 -1144
rect 29029 -2532 29087 -2520
rect 29227 -1144 29285 -1132
rect 29227 -2520 29239 -1144
rect 29273 -2520 29285 -1144
rect 29227 -2532 29285 -2520
rect 29425 -1144 29483 -1132
rect 29425 -2520 29437 -1144
rect 29471 -2520 29483 -1144
rect 29425 -2532 29483 -2520
rect 29623 -1144 29681 -1132
rect 29623 -2520 29635 -1144
rect 29669 -2520 29681 -1144
rect 29623 -2532 29681 -2520
rect 29821 -1144 29879 -1132
rect 29821 -2520 29833 -1144
rect 29867 -2520 29879 -1144
rect 29821 -2532 29879 -2520
rect 30019 -1144 30077 -1132
rect 30019 -2520 30031 -1144
rect 30065 -2520 30077 -1144
rect 30019 -2532 30077 -2520
rect 30217 -1144 30275 -1132
rect 30217 -2520 30229 -1144
rect 30263 -2520 30275 -1144
rect 30217 -2532 30275 -2520
rect 30415 -1144 30473 -1132
rect 30415 -2520 30427 -1144
rect 30461 -2520 30473 -1144
rect 30415 -2532 30473 -2520
rect 30613 -1144 30671 -1132
rect 30613 -2520 30625 -1144
rect 30659 -2520 30671 -1144
rect 30613 -2532 30671 -2520
rect 30811 -1144 30869 -1132
rect 30811 -2520 30823 -1144
rect 30857 -2520 30869 -1144
rect 30811 -2532 30869 -2520
rect 31009 -1144 31067 -1132
rect 31009 -2520 31021 -1144
rect 31055 -2520 31067 -1144
rect 31009 -2532 31067 -2520
rect 31207 -1144 31265 -1132
rect 31207 -2520 31219 -1144
rect 31253 -2520 31265 -1144
rect 31207 -2532 31265 -2520
rect 31405 -1144 31463 -1132
rect 31405 -2520 31417 -1144
rect 31451 -2520 31463 -1144
rect 31405 -2532 31463 -2520
rect 31603 -1144 31661 -1132
rect 31603 -2520 31615 -1144
rect 31649 -2520 31661 -1144
rect 31603 -2532 31661 -2520
rect 23287 -3345 23345 -3333
rect 23287 -4721 23299 -3345
rect 23333 -4721 23345 -3345
rect 23287 -4733 23345 -4721
rect 23485 -3345 23543 -3333
rect 23485 -4721 23497 -3345
rect 23531 -4721 23543 -3345
rect 23485 -4733 23543 -4721
rect 23683 -3345 23741 -3333
rect 23683 -4721 23695 -3345
rect 23729 -4721 23741 -3345
rect 23683 -4733 23741 -4721
rect 23881 -3345 23939 -3333
rect 23881 -4721 23893 -3345
rect 23927 -4721 23939 -3345
rect 23881 -4733 23939 -4721
rect 24079 -3345 24137 -3333
rect 24079 -4721 24091 -3345
rect 24125 -4721 24137 -3345
rect 24079 -4733 24137 -4721
rect 24277 -3345 24335 -3333
rect 24277 -4721 24289 -3345
rect 24323 -4721 24335 -3345
rect 24277 -4733 24335 -4721
rect 24475 -3345 24533 -3333
rect 24475 -4721 24487 -3345
rect 24521 -4721 24533 -3345
rect 24475 -4733 24533 -4721
rect 24673 -3345 24731 -3333
rect 24673 -4721 24685 -3345
rect 24719 -4721 24731 -3345
rect 24673 -4733 24731 -4721
rect 24871 -3345 24929 -3333
rect 24871 -4721 24883 -3345
rect 24917 -4721 24929 -3345
rect 24871 -4733 24929 -4721
rect 25069 -3345 25127 -3333
rect 25069 -4721 25081 -3345
rect 25115 -4721 25127 -3345
rect 25069 -4733 25127 -4721
rect 25267 -3345 25325 -3333
rect 25267 -4721 25279 -3345
rect 25313 -4721 25325 -3345
rect 25267 -4733 25325 -4721
rect 25465 -3345 25523 -3333
rect 25465 -4721 25477 -3345
rect 25511 -4721 25523 -3345
rect 25465 -4733 25523 -4721
rect 25663 -3345 25721 -3333
rect 25663 -4721 25675 -3345
rect 25709 -4721 25721 -3345
rect 25663 -4733 25721 -4721
rect 25861 -3345 25919 -3333
rect 25861 -4721 25873 -3345
rect 25907 -4721 25919 -3345
rect 25861 -4733 25919 -4721
rect 26059 -3345 26117 -3333
rect 26059 -4721 26071 -3345
rect 26105 -4721 26117 -3345
rect 26059 -4733 26117 -4721
rect 26257 -3345 26315 -3333
rect 26257 -4721 26269 -3345
rect 26303 -4721 26315 -3345
rect 26257 -4733 26315 -4721
rect 26455 -3345 26513 -3333
rect 26455 -4721 26467 -3345
rect 26501 -4721 26513 -3345
rect 26455 -4733 26513 -4721
rect 26653 -3345 26711 -3333
rect 26653 -4721 26665 -3345
rect 26699 -4721 26711 -3345
rect 26653 -4733 26711 -4721
rect 26851 -3345 26909 -3333
rect 26851 -4721 26863 -3345
rect 26897 -4721 26909 -3345
rect 26851 -4733 26909 -4721
rect 27049 -3345 27107 -3333
rect 27049 -4721 27061 -3345
rect 27095 -4721 27107 -3345
rect 27049 -4733 27107 -4721
rect 27247 -3345 27305 -3333
rect 27247 -4721 27259 -3345
rect 27293 -4721 27305 -3345
rect 27247 -4733 27305 -4721
rect 27445 -3345 27503 -3333
rect 27445 -4721 27457 -3345
rect 27491 -4721 27503 -3345
rect 27445 -4733 27503 -4721
rect 27643 -3345 27701 -3333
rect 27643 -4721 27655 -3345
rect 27689 -4721 27701 -3345
rect 27643 -4733 27701 -4721
rect 27841 -3345 27899 -3333
rect 27841 -4721 27853 -3345
rect 27887 -4721 27899 -3345
rect 27841 -4733 27899 -4721
rect 28039 -3345 28097 -3333
rect 28039 -4721 28051 -3345
rect 28085 -4721 28097 -3345
rect 28039 -4733 28097 -4721
rect 28237 -3345 28295 -3333
rect 28237 -4721 28249 -3345
rect 28283 -4721 28295 -3345
rect 28237 -4733 28295 -4721
rect 28435 -3345 28493 -3333
rect 28435 -4721 28447 -3345
rect 28481 -4721 28493 -3345
rect 28435 -4733 28493 -4721
rect 28633 -3345 28691 -3333
rect 28633 -4721 28645 -3345
rect 28679 -4721 28691 -3345
rect 28633 -4733 28691 -4721
rect 28831 -3345 28889 -3333
rect 28831 -4721 28843 -3345
rect 28877 -4721 28889 -3345
rect 28831 -4733 28889 -4721
rect 29029 -3345 29087 -3333
rect 29029 -4721 29041 -3345
rect 29075 -4721 29087 -3345
rect 29029 -4733 29087 -4721
rect 29227 -3345 29285 -3333
rect 29227 -4721 29239 -3345
rect 29273 -4721 29285 -3345
rect 29227 -4733 29285 -4721
rect 29425 -3345 29483 -3333
rect 29425 -4721 29437 -3345
rect 29471 -4721 29483 -3345
rect 29425 -4733 29483 -4721
rect 29623 -3345 29681 -3333
rect 29623 -4721 29635 -3345
rect 29669 -4721 29681 -3345
rect 29623 -4733 29681 -4721
rect 29821 -3345 29879 -3333
rect 29821 -4721 29833 -3345
rect 29867 -4721 29879 -3345
rect 29821 -4733 29879 -4721
rect 30019 -3345 30077 -3333
rect 30019 -4721 30031 -3345
rect 30065 -4721 30077 -3345
rect 30019 -4733 30077 -4721
rect 30217 -3345 30275 -3333
rect 30217 -4721 30229 -3345
rect 30263 -4721 30275 -3345
rect 30217 -4733 30275 -4721
rect 30415 -3345 30473 -3333
rect 30415 -4721 30427 -3345
rect 30461 -4721 30473 -3345
rect 30415 -4733 30473 -4721
rect 30613 -3345 30671 -3333
rect 30613 -4721 30625 -3345
rect 30659 -4721 30671 -3345
rect 30613 -4733 30671 -4721
rect 30811 -3345 30869 -3333
rect 30811 -4721 30823 -3345
rect 30857 -4721 30869 -3345
rect 30811 -4733 30869 -4721
rect 31009 -3345 31067 -3333
rect 31009 -4721 31021 -3345
rect 31055 -4721 31067 -3345
rect 31009 -4733 31067 -4721
rect 31207 -3345 31265 -3333
rect 31207 -4721 31219 -3345
rect 31253 -4721 31265 -3345
rect 31207 -4733 31265 -4721
rect 31405 -3345 31463 -3333
rect 31405 -4721 31417 -3345
rect 31451 -4721 31463 -3345
rect 31405 -4733 31463 -4721
rect 31603 -3345 31661 -3333
rect 31603 -4721 31615 -3345
rect 31649 -4721 31661 -3345
rect 31603 -4733 31661 -4721
<< pdiffc >>
rect 11449 752 11483 2128
rect 11647 752 11681 2128
rect 11845 752 11879 2128
rect 12043 752 12077 2128
rect 12241 752 12275 2128
rect 12439 752 12473 2128
rect 12637 752 12671 2128
rect 12835 752 12869 2128
rect 13033 752 13067 2128
rect 13231 752 13265 2128
rect 13429 752 13463 2128
rect 13627 752 13661 2128
rect 13825 752 13859 2128
rect 14023 752 14057 2128
rect 14221 752 14255 2128
rect 14419 752 14453 2128
rect 14617 752 14651 2128
rect 14815 752 14849 2128
rect 15013 752 15047 2128
rect 15211 752 15245 2128
rect 15409 752 15443 2128
rect 15607 752 15641 2128
rect 15805 752 15839 2128
rect 16003 752 16037 2128
rect 16201 752 16235 2128
rect 16399 752 16433 2128
rect 16597 752 16631 2128
rect 16795 752 16829 2128
rect 16993 752 17027 2128
rect 17191 752 17225 2128
rect 17389 752 17423 2128
rect 17587 752 17621 2128
rect 17785 752 17819 2128
rect 17983 752 18017 2128
rect 18181 752 18215 2128
rect 18379 752 18413 2128
rect 18577 752 18611 2128
rect 18775 752 18809 2128
rect 18973 752 19007 2128
rect 19171 752 19205 2128
rect 19369 752 19403 2128
rect 19567 752 19601 2128
rect 19765 752 19799 2128
rect 11449 -884 11483 492
rect 11647 -884 11681 492
rect 11845 -884 11879 492
rect 12043 -884 12077 492
rect 12241 -884 12275 492
rect 12439 -884 12473 492
rect 12637 -884 12671 492
rect 12835 -884 12869 492
rect 13033 -884 13067 492
rect 13231 -884 13265 492
rect 13429 -884 13463 492
rect 13627 -884 13661 492
rect 13825 -884 13859 492
rect 14023 -884 14057 492
rect 14221 -884 14255 492
rect 14419 -884 14453 492
rect 14617 -884 14651 492
rect 14815 -884 14849 492
rect 15013 -884 15047 492
rect 15211 -884 15245 492
rect 15409 -884 15443 492
rect 15607 -884 15641 492
rect 15805 -884 15839 492
rect 16003 -884 16037 492
rect 16201 -884 16235 492
rect 16399 -884 16433 492
rect 16597 -884 16631 492
rect 16795 -884 16829 492
rect 16993 -884 17027 492
rect 17191 -884 17225 492
rect 17389 -884 17423 492
rect 17587 -884 17621 492
rect 17785 -884 17819 492
rect 17983 -884 18017 492
rect 18181 -884 18215 492
rect 18379 -884 18413 492
rect 18577 -884 18611 492
rect 18775 -884 18809 492
rect 18973 -884 19007 492
rect 19171 -884 19205 492
rect 19369 -884 19403 492
rect 19567 -884 19601 492
rect 19765 -884 19799 492
rect 11449 -2520 11483 -1144
rect 11647 -2520 11681 -1144
rect 11845 -2520 11879 -1144
rect 12043 -2520 12077 -1144
rect 12241 -2520 12275 -1144
rect 12439 -2520 12473 -1144
rect 12637 -2520 12671 -1144
rect 12835 -2520 12869 -1144
rect 13033 -2520 13067 -1144
rect 13231 -2520 13265 -1144
rect 13429 -2520 13463 -1144
rect 13627 -2520 13661 -1144
rect 13825 -2520 13859 -1144
rect 14023 -2520 14057 -1144
rect 14221 -2520 14255 -1144
rect 14419 -2520 14453 -1144
rect 14617 -2520 14651 -1144
rect 14815 -2520 14849 -1144
rect 15013 -2520 15047 -1144
rect 15211 -2520 15245 -1144
rect 15409 -2520 15443 -1144
rect 15607 -2520 15641 -1144
rect 15805 -2520 15839 -1144
rect 16003 -2520 16037 -1144
rect 16201 -2520 16235 -1144
rect 16399 -2520 16433 -1144
rect 16597 -2520 16631 -1144
rect 16795 -2520 16829 -1144
rect 16993 -2520 17027 -1144
rect 17191 -2520 17225 -1144
rect 17389 -2520 17423 -1144
rect 17587 -2520 17621 -1144
rect 17785 -2520 17819 -1144
rect 17983 -2520 18017 -1144
rect 18181 -2520 18215 -1144
rect 18379 -2520 18413 -1144
rect 18577 -2520 18611 -1144
rect 18775 -2520 18809 -1144
rect 18973 -2520 19007 -1144
rect 19171 -2520 19205 -1144
rect 19369 -2520 19403 -1144
rect 19567 -2520 19601 -1144
rect 19765 -2520 19799 -1144
rect 11449 -4721 11483 -3345
rect 11647 -4721 11681 -3345
rect 11845 -4721 11879 -3345
rect 12043 -4721 12077 -3345
rect 12241 -4721 12275 -3345
rect 12439 -4721 12473 -3345
rect 12637 -4721 12671 -3345
rect 12835 -4721 12869 -3345
rect 13033 -4721 13067 -3345
rect 13231 -4721 13265 -3345
rect 13429 -4721 13463 -3345
rect 13627 -4721 13661 -3345
rect 13825 -4721 13859 -3345
rect 14023 -4721 14057 -3345
rect 14221 -4721 14255 -3345
rect 14419 -4721 14453 -3345
rect 14617 -4721 14651 -3345
rect 14815 -4721 14849 -3345
rect 15013 -4721 15047 -3345
rect 15211 -4721 15245 -3345
rect 15409 -4721 15443 -3345
rect 15607 -4721 15641 -3345
rect 15805 -4721 15839 -3345
rect 16003 -4721 16037 -3345
rect 16201 -4721 16235 -3345
rect 16399 -4721 16433 -3345
rect 16597 -4721 16631 -3345
rect 16795 -4721 16829 -3345
rect 16993 -4721 17027 -3345
rect 17191 -4721 17225 -3345
rect 17389 -4721 17423 -3345
rect 17587 -4721 17621 -3345
rect 17785 -4721 17819 -3345
rect 17983 -4721 18017 -3345
rect 18181 -4721 18215 -3345
rect 18379 -4721 18413 -3345
rect 18577 -4721 18611 -3345
rect 18775 -4721 18809 -3345
rect 18973 -4721 19007 -3345
rect 19171 -4721 19205 -3345
rect 19369 -4721 19403 -3345
rect 19567 -4721 19601 -3345
rect 19765 -4721 19799 -3345
rect 23299 752 23333 2128
rect 23497 752 23531 2128
rect 23695 752 23729 2128
rect 23893 752 23927 2128
rect 24091 752 24125 2128
rect 24289 752 24323 2128
rect 24487 752 24521 2128
rect 24685 752 24719 2128
rect 24883 752 24917 2128
rect 25081 752 25115 2128
rect 25279 752 25313 2128
rect 25477 752 25511 2128
rect 25675 752 25709 2128
rect 25873 752 25907 2128
rect 26071 752 26105 2128
rect 26269 752 26303 2128
rect 26467 752 26501 2128
rect 26665 752 26699 2128
rect 26863 752 26897 2128
rect 27061 752 27095 2128
rect 27259 752 27293 2128
rect 27457 752 27491 2128
rect 27655 752 27689 2128
rect 27853 752 27887 2128
rect 28051 752 28085 2128
rect 28249 752 28283 2128
rect 28447 752 28481 2128
rect 28645 752 28679 2128
rect 28843 752 28877 2128
rect 29041 752 29075 2128
rect 29239 752 29273 2128
rect 29437 752 29471 2128
rect 29635 752 29669 2128
rect 29833 752 29867 2128
rect 30031 752 30065 2128
rect 30229 752 30263 2128
rect 30427 752 30461 2128
rect 30625 752 30659 2128
rect 30823 752 30857 2128
rect 31021 752 31055 2128
rect 31219 752 31253 2128
rect 31417 752 31451 2128
rect 31615 752 31649 2128
rect 23299 -884 23333 492
rect 23497 -884 23531 492
rect 23695 -884 23729 492
rect 23893 -884 23927 492
rect 24091 -884 24125 492
rect 24289 -884 24323 492
rect 24487 -884 24521 492
rect 24685 -884 24719 492
rect 24883 -884 24917 492
rect 25081 -884 25115 492
rect 25279 -884 25313 492
rect 25477 -884 25511 492
rect 25675 -884 25709 492
rect 25873 -884 25907 492
rect 26071 -884 26105 492
rect 26269 -884 26303 492
rect 26467 -884 26501 492
rect 26665 -884 26699 492
rect 26863 -884 26897 492
rect 27061 -884 27095 492
rect 27259 -884 27293 492
rect 27457 -884 27491 492
rect 27655 -884 27689 492
rect 27853 -884 27887 492
rect 28051 -884 28085 492
rect 28249 -884 28283 492
rect 28447 -884 28481 492
rect 28645 -884 28679 492
rect 28843 -884 28877 492
rect 29041 -884 29075 492
rect 29239 -884 29273 492
rect 29437 -884 29471 492
rect 29635 -884 29669 492
rect 29833 -884 29867 492
rect 30031 -884 30065 492
rect 30229 -884 30263 492
rect 30427 -884 30461 492
rect 30625 -884 30659 492
rect 30823 -884 30857 492
rect 31021 -884 31055 492
rect 31219 -884 31253 492
rect 31417 -884 31451 492
rect 31615 -884 31649 492
rect 23299 -2520 23333 -1144
rect 23497 -2520 23531 -1144
rect 23695 -2520 23729 -1144
rect 23893 -2520 23927 -1144
rect 24091 -2520 24125 -1144
rect 24289 -2520 24323 -1144
rect 24487 -2520 24521 -1144
rect 24685 -2520 24719 -1144
rect 24883 -2520 24917 -1144
rect 25081 -2520 25115 -1144
rect 25279 -2520 25313 -1144
rect 25477 -2520 25511 -1144
rect 25675 -2520 25709 -1144
rect 25873 -2520 25907 -1144
rect 26071 -2520 26105 -1144
rect 26269 -2520 26303 -1144
rect 26467 -2520 26501 -1144
rect 26665 -2520 26699 -1144
rect 26863 -2520 26897 -1144
rect 27061 -2520 27095 -1144
rect 27259 -2520 27293 -1144
rect 27457 -2520 27491 -1144
rect 27655 -2520 27689 -1144
rect 27853 -2520 27887 -1144
rect 28051 -2520 28085 -1144
rect 28249 -2520 28283 -1144
rect 28447 -2520 28481 -1144
rect 28645 -2520 28679 -1144
rect 28843 -2520 28877 -1144
rect 29041 -2520 29075 -1144
rect 29239 -2520 29273 -1144
rect 29437 -2520 29471 -1144
rect 29635 -2520 29669 -1144
rect 29833 -2520 29867 -1144
rect 30031 -2520 30065 -1144
rect 30229 -2520 30263 -1144
rect 30427 -2520 30461 -1144
rect 30625 -2520 30659 -1144
rect 30823 -2520 30857 -1144
rect 31021 -2520 31055 -1144
rect 31219 -2520 31253 -1144
rect 31417 -2520 31451 -1144
rect 31615 -2520 31649 -1144
rect 23299 -4721 23333 -3345
rect 23497 -4721 23531 -3345
rect 23695 -4721 23729 -3345
rect 23893 -4721 23927 -3345
rect 24091 -4721 24125 -3345
rect 24289 -4721 24323 -3345
rect 24487 -4721 24521 -3345
rect 24685 -4721 24719 -3345
rect 24883 -4721 24917 -3345
rect 25081 -4721 25115 -3345
rect 25279 -4721 25313 -3345
rect 25477 -4721 25511 -3345
rect 25675 -4721 25709 -3345
rect 25873 -4721 25907 -3345
rect 26071 -4721 26105 -3345
rect 26269 -4721 26303 -3345
rect 26467 -4721 26501 -3345
rect 26665 -4721 26699 -3345
rect 26863 -4721 26897 -3345
rect 27061 -4721 27095 -3345
rect 27259 -4721 27293 -3345
rect 27457 -4721 27491 -3345
rect 27655 -4721 27689 -3345
rect 27853 -4721 27887 -3345
rect 28051 -4721 28085 -3345
rect 28249 -4721 28283 -3345
rect 28447 -4721 28481 -3345
rect 28645 -4721 28679 -3345
rect 28843 -4721 28877 -3345
rect 29041 -4721 29075 -3345
rect 29239 -4721 29273 -3345
rect 29437 -4721 29471 -3345
rect 29635 -4721 29669 -3345
rect 29833 -4721 29867 -3345
rect 30031 -4721 30065 -3345
rect 30229 -4721 30263 -3345
rect 30427 -4721 30461 -3345
rect 30625 -4721 30659 -3345
rect 30823 -4721 30857 -3345
rect 31021 -4721 31055 -3345
rect 31219 -4721 31253 -3345
rect 31417 -4721 31451 -3345
rect 31615 -4721 31649 -3345
<< nsubdiff >>
rect -848 2237 -752 2271
rect 8337 2237 8433 2271
rect -848 2175 -814 2237
rect 8399 2070 8433 2237
rect -814 -3034 -347 -2933
rect 7917 -3034 8399 -2933
rect -848 -5214 -814 -4353
rect 10991 2237 11087 2271
rect 20176 2237 20272 2271
rect 10991 2101 11025 2237
rect 8433 -3034 10991 -2933
rect 8399 -5214 8433 -4458
rect 20238 2070 20272 2237
rect 11025 -3034 11492 -2933
rect 19756 -3034 20238 -2933
rect 10991 -5214 11025 -4427
rect 22830 2237 22937 2271
rect 32026 2237 32122 2271
rect 22830 2101 22864 2237
rect 20272 -3034 22830 -2933
rect 20238 -5214 20272 -4458
rect 32088 1912 32122 2237
rect 22864 -3034 23342 -2933
rect 31606 -3034 32088 -2933
rect 22864 -4415 22875 -4353
rect 22830 -5214 22864 -4427
rect 32088 -5214 32122 -4731
rect -848 -5248 -457 -5214
rect 31740 -5248 32122 -5214
<< nsubdiffcont >>
rect -752 2237 8337 2271
rect -848 -4353 -814 2175
rect -347 -3034 7917 -2933
rect 8399 -4458 8433 2070
rect 11087 2237 20176 2271
rect 10991 -4427 11025 2101
rect 11492 -3034 19756 -2933
rect 20238 -4458 20272 2070
rect 22937 2237 32026 2271
rect 22830 -4427 22864 2101
rect 23342 -3034 31606 -2933
rect 32088 -4731 32122 1912
rect -457 -5248 31740 -5214
<< poly >>
rect 11495 2140 11635 2166
rect 11693 2140 11833 2166
rect 11891 2140 12031 2166
rect 12089 2140 12229 2166
rect 12287 2140 12427 2166
rect 12485 2140 12625 2166
rect 12683 2140 12823 2166
rect 12881 2140 13021 2166
rect 13079 2140 13219 2166
rect 13277 2140 13417 2166
rect 13475 2140 13615 2166
rect 13673 2140 13813 2166
rect 13871 2140 14011 2166
rect 14069 2140 14209 2166
rect 14267 2140 14407 2166
rect 14465 2140 14605 2166
rect 14663 2140 14803 2166
rect 14861 2140 15001 2166
rect 15059 2140 15199 2166
rect 15257 2140 15397 2166
rect 15455 2140 15595 2166
rect 15653 2140 15793 2166
rect 15851 2140 15991 2166
rect 16049 2140 16189 2166
rect 16247 2140 16387 2166
rect 16445 2140 16585 2166
rect 16643 2140 16783 2166
rect 16841 2140 16981 2166
rect 17039 2140 17179 2166
rect 17237 2140 17377 2166
rect 17435 2140 17575 2166
rect 17633 2140 17773 2166
rect 17831 2140 17971 2166
rect 18029 2140 18169 2166
rect 18227 2140 18367 2166
rect 18425 2140 18565 2166
rect 18623 2140 18763 2166
rect 18821 2140 18961 2166
rect 19019 2140 19159 2166
rect 19217 2140 19357 2166
rect 19415 2140 19555 2166
rect 19613 2140 19753 2166
rect 11495 693 11635 740
rect 11495 659 11511 693
rect 11619 659 11635 693
rect 11495 643 11635 659
rect 11693 693 11833 740
rect 11693 659 11709 693
rect 11817 659 11833 693
rect 11693 643 11833 659
rect 11891 693 12031 740
rect 11891 659 11907 693
rect 12015 659 12031 693
rect 11891 643 12031 659
rect 12089 693 12229 740
rect 12089 659 12105 693
rect 12213 659 12229 693
rect 12089 643 12229 659
rect 12287 693 12427 740
rect 12287 659 12303 693
rect 12411 659 12427 693
rect 12287 643 12427 659
rect 12485 693 12625 740
rect 12485 659 12501 693
rect 12609 659 12625 693
rect 12485 643 12625 659
rect 12683 693 12823 740
rect 12683 659 12699 693
rect 12807 659 12823 693
rect 12683 643 12823 659
rect 12881 693 13021 740
rect 12881 659 12897 693
rect 13005 659 13021 693
rect 12881 643 13021 659
rect 13079 693 13219 740
rect 13079 659 13095 693
rect 13203 659 13219 693
rect 13079 643 13219 659
rect 13277 693 13417 740
rect 13277 659 13293 693
rect 13401 659 13417 693
rect 13277 643 13417 659
rect 13475 693 13615 740
rect 13475 659 13491 693
rect 13599 659 13615 693
rect 13475 643 13615 659
rect 13673 693 13813 740
rect 13673 659 13689 693
rect 13797 659 13813 693
rect 13673 643 13813 659
rect 13871 693 14011 740
rect 13871 659 13887 693
rect 13995 659 14011 693
rect 13871 643 14011 659
rect 14069 693 14209 740
rect 14069 659 14085 693
rect 14193 659 14209 693
rect 14069 643 14209 659
rect 14267 693 14407 740
rect 14267 659 14283 693
rect 14391 659 14407 693
rect 14267 643 14407 659
rect 14465 693 14605 740
rect 14465 659 14481 693
rect 14589 659 14605 693
rect 14465 643 14605 659
rect 14663 693 14803 740
rect 14663 659 14679 693
rect 14787 659 14803 693
rect 14663 643 14803 659
rect 14861 693 15001 740
rect 14861 659 14877 693
rect 14985 659 15001 693
rect 14861 643 15001 659
rect 15059 693 15199 740
rect 15059 659 15075 693
rect 15183 659 15199 693
rect 15059 643 15199 659
rect 15257 693 15397 740
rect 15257 659 15273 693
rect 15381 659 15397 693
rect 15257 643 15397 659
rect 15455 693 15595 740
rect 15455 659 15471 693
rect 15579 659 15595 693
rect 15455 643 15595 659
rect 15653 693 15793 740
rect 15653 659 15669 693
rect 15777 659 15793 693
rect 15653 643 15793 659
rect 15851 693 15991 740
rect 15851 659 15867 693
rect 15975 659 15991 693
rect 15851 643 15991 659
rect 16049 693 16189 740
rect 16049 659 16065 693
rect 16173 659 16189 693
rect 16049 643 16189 659
rect 16247 693 16387 740
rect 16247 659 16263 693
rect 16371 659 16387 693
rect 16247 643 16387 659
rect 16445 693 16585 740
rect 16445 659 16461 693
rect 16569 659 16585 693
rect 16445 643 16585 659
rect 16643 693 16783 740
rect 16643 659 16659 693
rect 16767 659 16783 693
rect 16643 643 16783 659
rect 16841 693 16981 740
rect 16841 659 16857 693
rect 16965 659 16981 693
rect 16841 643 16981 659
rect 17039 693 17179 740
rect 17039 659 17055 693
rect 17163 659 17179 693
rect 17039 643 17179 659
rect 17237 693 17377 740
rect 17237 659 17253 693
rect 17361 659 17377 693
rect 17237 643 17377 659
rect 17435 693 17575 740
rect 17435 659 17451 693
rect 17559 659 17575 693
rect 17435 643 17575 659
rect 17633 693 17773 740
rect 17633 659 17649 693
rect 17757 659 17773 693
rect 17633 643 17773 659
rect 17831 693 17971 740
rect 17831 659 17847 693
rect 17955 659 17971 693
rect 17831 643 17971 659
rect 18029 693 18169 740
rect 18029 659 18045 693
rect 18153 659 18169 693
rect 18029 643 18169 659
rect 18227 693 18367 740
rect 18227 659 18243 693
rect 18351 659 18367 693
rect 18227 643 18367 659
rect 18425 693 18565 740
rect 18425 659 18441 693
rect 18549 659 18565 693
rect 18425 643 18565 659
rect 18623 693 18763 740
rect 18623 659 18639 693
rect 18747 659 18763 693
rect 18623 643 18763 659
rect 18821 693 18961 740
rect 18821 659 18837 693
rect 18945 659 18961 693
rect 18821 643 18961 659
rect 19019 693 19159 740
rect 19019 659 19035 693
rect 19143 659 19159 693
rect 19019 643 19159 659
rect 19217 693 19357 740
rect 19217 659 19233 693
rect 19341 659 19357 693
rect 19217 643 19357 659
rect 19415 693 19555 740
rect 19415 659 19431 693
rect 19539 659 19555 693
rect 19415 643 19555 659
rect 19613 693 19753 740
rect 19613 659 19629 693
rect 19737 659 19753 693
rect 19613 643 19753 659
rect 11495 585 11635 601
rect 11495 551 11511 585
rect 11619 551 11635 585
rect 11495 504 11635 551
rect 11693 585 11833 601
rect 11693 551 11709 585
rect 11817 551 11833 585
rect 11693 504 11833 551
rect 11891 585 12031 601
rect 11891 551 11907 585
rect 12015 551 12031 585
rect 11891 504 12031 551
rect 12089 585 12229 601
rect 12089 551 12105 585
rect 12213 551 12229 585
rect 12089 504 12229 551
rect 12287 585 12427 601
rect 12287 551 12303 585
rect 12411 551 12427 585
rect 12287 504 12427 551
rect 12485 585 12625 601
rect 12485 551 12501 585
rect 12609 551 12625 585
rect 12485 504 12625 551
rect 12683 585 12823 601
rect 12683 551 12699 585
rect 12807 551 12823 585
rect 12683 504 12823 551
rect 12881 585 13021 601
rect 12881 551 12897 585
rect 13005 551 13021 585
rect 12881 504 13021 551
rect 13079 585 13219 601
rect 13079 551 13095 585
rect 13203 551 13219 585
rect 13079 504 13219 551
rect 13277 585 13417 601
rect 13277 551 13293 585
rect 13401 551 13417 585
rect 13277 504 13417 551
rect 13475 585 13615 601
rect 13475 551 13491 585
rect 13599 551 13615 585
rect 13475 504 13615 551
rect 13673 585 13813 601
rect 13673 551 13689 585
rect 13797 551 13813 585
rect 13673 504 13813 551
rect 13871 585 14011 601
rect 13871 551 13887 585
rect 13995 551 14011 585
rect 13871 504 14011 551
rect 14069 585 14209 601
rect 14069 551 14085 585
rect 14193 551 14209 585
rect 14069 504 14209 551
rect 14267 585 14407 601
rect 14267 551 14283 585
rect 14391 551 14407 585
rect 14267 504 14407 551
rect 14465 585 14605 601
rect 14465 551 14481 585
rect 14589 551 14605 585
rect 14465 504 14605 551
rect 14663 585 14803 601
rect 14663 551 14679 585
rect 14787 551 14803 585
rect 14663 504 14803 551
rect 14861 585 15001 601
rect 14861 551 14877 585
rect 14985 551 15001 585
rect 14861 504 15001 551
rect 15059 585 15199 601
rect 15059 551 15075 585
rect 15183 551 15199 585
rect 15059 504 15199 551
rect 15257 585 15397 601
rect 15257 551 15273 585
rect 15381 551 15397 585
rect 15257 504 15397 551
rect 15455 585 15595 601
rect 15455 551 15471 585
rect 15579 551 15595 585
rect 15455 504 15595 551
rect 15653 585 15793 601
rect 15653 551 15669 585
rect 15777 551 15793 585
rect 15653 504 15793 551
rect 15851 585 15991 601
rect 15851 551 15867 585
rect 15975 551 15991 585
rect 15851 504 15991 551
rect 16049 585 16189 601
rect 16049 551 16065 585
rect 16173 551 16189 585
rect 16049 504 16189 551
rect 16247 585 16387 601
rect 16247 551 16263 585
rect 16371 551 16387 585
rect 16247 504 16387 551
rect 16445 585 16585 601
rect 16445 551 16461 585
rect 16569 551 16585 585
rect 16445 504 16585 551
rect 16643 585 16783 601
rect 16643 551 16659 585
rect 16767 551 16783 585
rect 16643 504 16783 551
rect 16841 585 16981 601
rect 16841 551 16857 585
rect 16965 551 16981 585
rect 16841 504 16981 551
rect 17039 585 17179 601
rect 17039 551 17055 585
rect 17163 551 17179 585
rect 17039 504 17179 551
rect 17237 585 17377 601
rect 17237 551 17253 585
rect 17361 551 17377 585
rect 17237 504 17377 551
rect 17435 585 17575 601
rect 17435 551 17451 585
rect 17559 551 17575 585
rect 17435 504 17575 551
rect 17633 585 17773 601
rect 17633 551 17649 585
rect 17757 551 17773 585
rect 17633 504 17773 551
rect 17831 585 17971 601
rect 17831 551 17847 585
rect 17955 551 17971 585
rect 17831 504 17971 551
rect 18029 585 18169 601
rect 18029 551 18045 585
rect 18153 551 18169 585
rect 18029 504 18169 551
rect 18227 585 18367 601
rect 18227 551 18243 585
rect 18351 551 18367 585
rect 18227 504 18367 551
rect 18425 585 18565 601
rect 18425 551 18441 585
rect 18549 551 18565 585
rect 18425 504 18565 551
rect 18623 585 18763 601
rect 18623 551 18639 585
rect 18747 551 18763 585
rect 18623 504 18763 551
rect 18821 585 18961 601
rect 18821 551 18837 585
rect 18945 551 18961 585
rect 18821 504 18961 551
rect 19019 585 19159 601
rect 19019 551 19035 585
rect 19143 551 19159 585
rect 19019 504 19159 551
rect 19217 585 19357 601
rect 19217 551 19233 585
rect 19341 551 19357 585
rect 19217 504 19357 551
rect 19415 585 19555 601
rect 19415 551 19431 585
rect 19539 551 19555 585
rect 19415 504 19555 551
rect 19613 585 19753 601
rect 19613 551 19629 585
rect 19737 551 19753 585
rect 19613 504 19753 551
rect 11495 -943 11635 -896
rect 11495 -977 11511 -943
rect 11619 -977 11635 -943
rect 11495 -993 11635 -977
rect 11693 -943 11833 -896
rect 11693 -977 11709 -943
rect 11817 -977 11833 -943
rect 11693 -993 11833 -977
rect 11891 -943 12031 -896
rect 11891 -977 11907 -943
rect 12015 -977 12031 -943
rect 11891 -993 12031 -977
rect 12089 -943 12229 -896
rect 12089 -977 12105 -943
rect 12213 -977 12229 -943
rect 12089 -993 12229 -977
rect 12287 -943 12427 -896
rect 12287 -977 12303 -943
rect 12411 -977 12427 -943
rect 12287 -993 12427 -977
rect 12485 -943 12625 -896
rect 12485 -977 12501 -943
rect 12609 -977 12625 -943
rect 12485 -993 12625 -977
rect 12683 -943 12823 -896
rect 12683 -977 12699 -943
rect 12807 -977 12823 -943
rect 12683 -993 12823 -977
rect 12881 -943 13021 -896
rect 12881 -977 12897 -943
rect 13005 -977 13021 -943
rect 12881 -993 13021 -977
rect 13079 -943 13219 -896
rect 13079 -977 13095 -943
rect 13203 -977 13219 -943
rect 13079 -993 13219 -977
rect 13277 -943 13417 -896
rect 13277 -977 13293 -943
rect 13401 -977 13417 -943
rect 13277 -993 13417 -977
rect 13475 -943 13615 -896
rect 13475 -977 13491 -943
rect 13599 -977 13615 -943
rect 13475 -993 13615 -977
rect 13673 -943 13813 -896
rect 13673 -977 13689 -943
rect 13797 -977 13813 -943
rect 13673 -993 13813 -977
rect 13871 -943 14011 -896
rect 13871 -977 13887 -943
rect 13995 -977 14011 -943
rect 13871 -993 14011 -977
rect 14069 -943 14209 -896
rect 14069 -977 14085 -943
rect 14193 -977 14209 -943
rect 14069 -993 14209 -977
rect 14267 -943 14407 -896
rect 14267 -977 14283 -943
rect 14391 -977 14407 -943
rect 14267 -993 14407 -977
rect 14465 -943 14605 -896
rect 14465 -977 14481 -943
rect 14589 -977 14605 -943
rect 14465 -993 14605 -977
rect 14663 -943 14803 -896
rect 14663 -977 14679 -943
rect 14787 -977 14803 -943
rect 14663 -993 14803 -977
rect 14861 -943 15001 -896
rect 14861 -977 14877 -943
rect 14985 -977 15001 -943
rect 14861 -993 15001 -977
rect 15059 -943 15199 -896
rect 15059 -977 15075 -943
rect 15183 -977 15199 -943
rect 15059 -993 15199 -977
rect 15257 -943 15397 -896
rect 15257 -977 15273 -943
rect 15381 -977 15397 -943
rect 15257 -993 15397 -977
rect 15455 -943 15595 -896
rect 15455 -977 15471 -943
rect 15579 -977 15595 -943
rect 15455 -993 15595 -977
rect 15653 -943 15793 -896
rect 15653 -977 15669 -943
rect 15777 -977 15793 -943
rect 15653 -993 15793 -977
rect 15851 -943 15991 -896
rect 15851 -977 15867 -943
rect 15975 -977 15991 -943
rect 15851 -993 15991 -977
rect 16049 -943 16189 -896
rect 16049 -977 16065 -943
rect 16173 -977 16189 -943
rect 16049 -993 16189 -977
rect 16247 -943 16387 -896
rect 16247 -977 16263 -943
rect 16371 -977 16387 -943
rect 16247 -993 16387 -977
rect 16445 -943 16585 -896
rect 16445 -977 16461 -943
rect 16569 -977 16585 -943
rect 16445 -993 16585 -977
rect 16643 -943 16783 -896
rect 16643 -977 16659 -943
rect 16767 -977 16783 -943
rect 16643 -993 16783 -977
rect 16841 -943 16981 -896
rect 16841 -977 16857 -943
rect 16965 -977 16981 -943
rect 16841 -993 16981 -977
rect 17039 -943 17179 -896
rect 17039 -977 17055 -943
rect 17163 -977 17179 -943
rect 17039 -993 17179 -977
rect 17237 -943 17377 -896
rect 17237 -977 17253 -943
rect 17361 -977 17377 -943
rect 17237 -993 17377 -977
rect 17435 -943 17575 -896
rect 17435 -977 17451 -943
rect 17559 -977 17575 -943
rect 17435 -993 17575 -977
rect 17633 -943 17773 -896
rect 17633 -977 17649 -943
rect 17757 -977 17773 -943
rect 17633 -993 17773 -977
rect 17831 -943 17971 -896
rect 17831 -977 17847 -943
rect 17955 -977 17971 -943
rect 17831 -993 17971 -977
rect 18029 -943 18169 -896
rect 18029 -977 18045 -943
rect 18153 -977 18169 -943
rect 18029 -993 18169 -977
rect 18227 -943 18367 -896
rect 18227 -977 18243 -943
rect 18351 -977 18367 -943
rect 18227 -993 18367 -977
rect 18425 -943 18565 -896
rect 18425 -977 18441 -943
rect 18549 -977 18565 -943
rect 18425 -993 18565 -977
rect 18623 -943 18763 -896
rect 18623 -977 18639 -943
rect 18747 -977 18763 -943
rect 18623 -993 18763 -977
rect 18821 -943 18961 -896
rect 18821 -977 18837 -943
rect 18945 -977 18961 -943
rect 18821 -993 18961 -977
rect 19019 -943 19159 -896
rect 19019 -977 19035 -943
rect 19143 -977 19159 -943
rect 19019 -993 19159 -977
rect 19217 -943 19357 -896
rect 19217 -977 19233 -943
rect 19341 -977 19357 -943
rect 19217 -993 19357 -977
rect 19415 -943 19555 -896
rect 19415 -977 19431 -943
rect 19539 -977 19555 -943
rect 19415 -993 19555 -977
rect 19613 -943 19753 -896
rect 19613 -977 19629 -943
rect 19737 -977 19753 -943
rect 19613 -993 19753 -977
rect 11495 -1051 11635 -1035
rect 11495 -1085 11511 -1051
rect 11619 -1085 11635 -1051
rect 11495 -1132 11635 -1085
rect 11693 -1051 11833 -1035
rect 11693 -1085 11709 -1051
rect 11817 -1085 11833 -1051
rect 11693 -1132 11833 -1085
rect 11891 -1051 12031 -1035
rect 11891 -1085 11907 -1051
rect 12015 -1085 12031 -1051
rect 11891 -1132 12031 -1085
rect 12089 -1051 12229 -1035
rect 12089 -1085 12105 -1051
rect 12213 -1085 12229 -1051
rect 12089 -1132 12229 -1085
rect 12287 -1051 12427 -1035
rect 12287 -1085 12303 -1051
rect 12411 -1085 12427 -1051
rect 12287 -1132 12427 -1085
rect 12485 -1051 12625 -1035
rect 12485 -1085 12501 -1051
rect 12609 -1085 12625 -1051
rect 12485 -1132 12625 -1085
rect 12683 -1051 12823 -1035
rect 12683 -1085 12699 -1051
rect 12807 -1085 12823 -1051
rect 12683 -1132 12823 -1085
rect 12881 -1051 13021 -1035
rect 12881 -1085 12897 -1051
rect 13005 -1085 13021 -1051
rect 12881 -1132 13021 -1085
rect 13079 -1051 13219 -1035
rect 13079 -1085 13095 -1051
rect 13203 -1085 13219 -1051
rect 13079 -1132 13219 -1085
rect 13277 -1051 13417 -1035
rect 13277 -1085 13293 -1051
rect 13401 -1085 13417 -1051
rect 13277 -1132 13417 -1085
rect 13475 -1051 13615 -1035
rect 13475 -1085 13491 -1051
rect 13599 -1085 13615 -1051
rect 13475 -1132 13615 -1085
rect 13673 -1051 13813 -1035
rect 13673 -1085 13689 -1051
rect 13797 -1085 13813 -1051
rect 13673 -1132 13813 -1085
rect 13871 -1051 14011 -1035
rect 13871 -1085 13887 -1051
rect 13995 -1085 14011 -1051
rect 13871 -1132 14011 -1085
rect 14069 -1051 14209 -1035
rect 14069 -1085 14085 -1051
rect 14193 -1085 14209 -1051
rect 14069 -1132 14209 -1085
rect 14267 -1051 14407 -1035
rect 14267 -1085 14283 -1051
rect 14391 -1085 14407 -1051
rect 14267 -1132 14407 -1085
rect 14465 -1051 14605 -1035
rect 14465 -1085 14481 -1051
rect 14589 -1085 14605 -1051
rect 14465 -1132 14605 -1085
rect 14663 -1051 14803 -1035
rect 14663 -1085 14679 -1051
rect 14787 -1085 14803 -1051
rect 14663 -1132 14803 -1085
rect 14861 -1051 15001 -1035
rect 14861 -1085 14877 -1051
rect 14985 -1085 15001 -1051
rect 14861 -1132 15001 -1085
rect 15059 -1051 15199 -1035
rect 15059 -1085 15075 -1051
rect 15183 -1085 15199 -1051
rect 15059 -1132 15199 -1085
rect 15257 -1051 15397 -1035
rect 15257 -1085 15273 -1051
rect 15381 -1085 15397 -1051
rect 15257 -1132 15397 -1085
rect 15455 -1051 15595 -1035
rect 15455 -1085 15471 -1051
rect 15579 -1085 15595 -1051
rect 15455 -1132 15595 -1085
rect 15653 -1051 15793 -1035
rect 15653 -1085 15669 -1051
rect 15777 -1085 15793 -1051
rect 15653 -1132 15793 -1085
rect 15851 -1051 15991 -1035
rect 15851 -1085 15867 -1051
rect 15975 -1085 15991 -1051
rect 15851 -1132 15991 -1085
rect 16049 -1051 16189 -1035
rect 16049 -1085 16065 -1051
rect 16173 -1085 16189 -1051
rect 16049 -1132 16189 -1085
rect 16247 -1051 16387 -1035
rect 16247 -1085 16263 -1051
rect 16371 -1085 16387 -1051
rect 16247 -1132 16387 -1085
rect 16445 -1051 16585 -1035
rect 16445 -1085 16461 -1051
rect 16569 -1085 16585 -1051
rect 16445 -1132 16585 -1085
rect 16643 -1051 16783 -1035
rect 16643 -1085 16659 -1051
rect 16767 -1085 16783 -1051
rect 16643 -1132 16783 -1085
rect 16841 -1051 16981 -1035
rect 16841 -1085 16857 -1051
rect 16965 -1085 16981 -1051
rect 16841 -1132 16981 -1085
rect 17039 -1051 17179 -1035
rect 17039 -1085 17055 -1051
rect 17163 -1085 17179 -1051
rect 17039 -1132 17179 -1085
rect 17237 -1051 17377 -1035
rect 17237 -1085 17253 -1051
rect 17361 -1085 17377 -1051
rect 17237 -1132 17377 -1085
rect 17435 -1051 17575 -1035
rect 17435 -1085 17451 -1051
rect 17559 -1085 17575 -1051
rect 17435 -1132 17575 -1085
rect 17633 -1051 17773 -1035
rect 17633 -1085 17649 -1051
rect 17757 -1085 17773 -1051
rect 17633 -1132 17773 -1085
rect 17831 -1051 17971 -1035
rect 17831 -1085 17847 -1051
rect 17955 -1085 17971 -1051
rect 17831 -1132 17971 -1085
rect 18029 -1051 18169 -1035
rect 18029 -1085 18045 -1051
rect 18153 -1085 18169 -1051
rect 18029 -1132 18169 -1085
rect 18227 -1051 18367 -1035
rect 18227 -1085 18243 -1051
rect 18351 -1085 18367 -1051
rect 18227 -1132 18367 -1085
rect 18425 -1051 18565 -1035
rect 18425 -1085 18441 -1051
rect 18549 -1085 18565 -1051
rect 18425 -1132 18565 -1085
rect 18623 -1051 18763 -1035
rect 18623 -1085 18639 -1051
rect 18747 -1085 18763 -1051
rect 18623 -1132 18763 -1085
rect 18821 -1051 18961 -1035
rect 18821 -1085 18837 -1051
rect 18945 -1085 18961 -1051
rect 18821 -1132 18961 -1085
rect 19019 -1051 19159 -1035
rect 19019 -1085 19035 -1051
rect 19143 -1085 19159 -1051
rect 19019 -1132 19159 -1085
rect 19217 -1051 19357 -1035
rect 19217 -1085 19233 -1051
rect 19341 -1085 19357 -1051
rect 19217 -1132 19357 -1085
rect 19415 -1051 19555 -1035
rect 19415 -1085 19431 -1051
rect 19539 -1085 19555 -1051
rect 19415 -1132 19555 -1085
rect 19613 -1051 19753 -1035
rect 19613 -1085 19629 -1051
rect 19737 -1085 19753 -1051
rect 19613 -1132 19753 -1085
rect 11495 -2579 11635 -2532
rect 11495 -2613 11511 -2579
rect 11619 -2613 11635 -2579
rect 11495 -2629 11635 -2613
rect 11693 -2579 11833 -2532
rect 11693 -2613 11709 -2579
rect 11817 -2613 11833 -2579
rect 11693 -2629 11833 -2613
rect 11891 -2579 12031 -2532
rect 11891 -2613 11907 -2579
rect 12015 -2613 12031 -2579
rect 11891 -2629 12031 -2613
rect 12089 -2579 12229 -2532
rect 12089 -2613 12105 -2579
rect 12213 -2613 12229 -2579
rect 12089 -2629 12229 -2613
rect 12287 -2579 12427 -2532
rect 12287 -2613 12303 -2579
rect 12411 -2613 12427 -2579
rect 12287 -2629 12427 -2613
rect 12485 -2579 12625 -2532
rect 12485 -2613 12501 -2579
rect 12609 -2613 12625 -2579
rect 12485 -2629 12625 -2613
rect 12683 -2579 12823 -2532
rect 12683 -2613 12699 -2579
rect 12807 -2613 12823 -2579
rect 12683 -2629 12823 -2613
rect 12881 -2579 13021 -2532
rect 12881 -2613 12897 -2579
rect 13005 -2613 13021 -2579
rect 12881 -2629 13021 -2613
rect 13079 -2579 13219 -2532
rect 13079 -2613 13095 -2579
rect 13203 -2613 13219 -2579
rect 13079 -2629 13219 -2613
rect 13277 -2579 13417 -2532
rect 13277 -2613 13293 -2579
rect 13401 -2613 13417 -2579
rect 13277 -2629 13417 -2613
rect 13475 -2579 13615 -2532
rect 13475 -2613 13491 -2579
rect 13599 -2613 13615 -2579
rect 13475 -2629 13615 -2613
rect 13673 -2579 13813 -2532
rect 13673 -2613 13689 -2579
rect 13797 -2613 13813 -2579
rect 13673 -2629 13813 -2613
rect 13871 -2579 14011 -2532
rect 13871 -2613 13887 -2579
rect 13995 -2613 14011 -2579
rect 13871 -2629 14011 -2613
rect 14069 -2579 14209 -2532
rect 14069 -2613 14085 -2579
rect 14193 -2613 14209 -2579
rect 14069 -2629 14209 -2613
rect 14267 -2579 14407 -2532
rect 14267 -2613 14283 -2579
rect 14391 -2613 14407 -2579
rect 14267 -2629 14407 -2613
rect 14465 -2579 14605 -2532
rect 14465 -2613 14481 -2579
rect 14589 -2613 14605 -2579
rect 14465 -2629 14605 -2613
rect 14663 -2579 14803 -2532
rect 14663 -2613 14679 -2579
rect 14787 -2613 14803 -2579
rect 14663 -2629 14803 -2613
rect 14861 -2579 15001 -2532
rect 14861 -2613 14877 -2579
rect 14985 -2613 15001 -2579
rect 14861 -2629 15001 -2613
rect 15059 -2579 15199 -2532
rect 15059 -2613 15075 -2579
rect 15183 -2613 15199 -2579
rect 15059 -2629 15199 -2613
rect 15257 -2579 15397 -2532
rect 15257 -2613 15273 -2579
rect 15381 -2613 15397 -2579
rect 15257 -2629 15397 -2613
rect 15455 -2579 15595 -2532
rect 15455 -2613 15471 -2579
rect 15579 -2613 15595 -2579
rect 15455 -2629 15595 -2613
rect 15653 -2579 15793 -2532
rect 15653 -2613 15669 -2579
rect 15777 -2613 15793 -2579
rect 15653 -2629 15793 -2613
rect 15851 -2579 15991 -2532
rect 15851 -2613 15867 -2579
rect 15975 -2613 15991 -2579
rect 15851 -2629 15991 -2613
rect 16049 -2579 16189 -2532
rect 16049 -2613 16065 -2579
rect 16173 -2613 16189 -2579
rect 16049 -2629 16189 -2613
rect 16247 -2579 16387 -2532
rect 16247 -2613 16263 -2579
rect 16371 -2613 16387 -2579
rect 16247 -2629 16387 -2613
rect 16445 -2579 16585 -2532
rect 16445 -2613 16461 -2579
rect 16569 -2613 16585 -2579
rect 16445 -2629 16585 -2613
rect 16643 -2579 16783 -2532
rect 16643 -2613 16659 -2579
rect 16767 -2613 16783 -2579
rect 16643 -2629 16783 -2613
rect 16841 -2579 16981 -2532
rect 16841 -2613 16857 -2579
rect 16965 -2613 16981 -2579
rect 16841 -2629 16981 -2613
rect 17039 -2579 17179 -2532
rect 17039 -2613 17055 -2579
rect 17163 -2613 17179 -2579
rect 17039 -2629 17179 -2613
rect 17237 -2579 17377 -2532
rect 17237 -2613 17253 -2579
rect 17361 -2613 17377 -2579
rect 17237 -2629 17377 -2613
rect 17435 -2579 17575 -2532
rect 17435 -2613 17451 -2579
rect 17559 -2613 17575 -2579
rect 17435 -2629 17575 -2613
rect 17633 -2579 17773 -2532
rect 17633 -2613 17649 -2579
rect 17757 -2613 17773 -2579
rect 17633 -2629 17773 -2613
rect 17831 -2579 17971 -2532
rect 17831 -2613 17847 -2579
rect 17955 -2613 17971 -2579
rect 17831 -2629 17971 -2613
rect 18029 -2579 18169 -2532
rect 18029 -2613 18045 -2579
rect 18153 -2613 18169 -2579
rect 18029 -2629 18169 -2613
rect 18227 -2579 18367 -2532
rect 18227 -2613 18243 -2579
rect 18351 -2613 18367 -2579
rect 18227 -2629 18367 -2613
rect 18425 -2579 18565 -2532
rect 18425 -2613 18441 -2579
rect 18549 -2613 18565 -2579
rect 18425 -2629 18565 -2613
rect 18623 -2579 18763 -2532
rect 18623 -2613 18639 -2579
rect 18747 -2613 18763 -2579
rect 18623 -2629 18763 -2613
rect 18821 -2579 18961 -2532
rect 18821 -2613 18837 -2579
rect 18945 -2613 18961 -2579
rect 18821 -2629 18961 -2613
rect 19019 -2579 19159 -2532
rect 19019 -2613 19035 -2579
rect 19143 -2613 19159 -2579
rect 19019 -2629 19159 -2613
rect 19217 -2579 19357 -2532
rect 19217 -2613 19233 -2579
rect 19341 -2613 19357 -2579
rect 19217 -2629 19357 -2613
rect 19415 -2579 19555 -2532
rect 19415 -2613 19431 -2579
rect 19539 -2613 19555 -2579
rect 19415 -2629 19555 -2613
rect 19613 -2579 19753 -2532
rect 19613 -2613 19629 -2579
rect 19737 -2613 19753 -2579
rect 19613 -2629 19753 -2613
rect 11495 -3252 11635 -3236
rect 11495 -3286 11511 -3252
rect 11619 -3286 11635 -3252
rect 11495 -3333 11635 -3286
rect 11693 -3252 11833 -3236
rect 11693 -3286 11709 -3252
rect 11817 -3286 11833 -3252
rect 11693 -3333 11833 -3286
rect 11891 -3252 12031 -3236
rect 11891 -3286 11907 -3252
rect 12015 -3286 12031 -3252
rect 11891 -3333 12031 -3286
rect 12089 -3252 12229 -3236
rect 12089 -3286 12105 -3252
rect 12213 -3286 12229 -3252
rect 12089 -3333 12229 -3286
rect 12287 -3252 12427 -3236
rect 12287 -3286 12303 -3252
rect 12411 -3286 12427 -3252
rect 12287 -3333 12427 -3286
rect 12485 -3252 12625 -3236
rect 12485 -3286 12501 -3252
rect 12609 -3286 12625 -3252
rect 12485 -3333 12625 -3286
rect 12683 -3252 12823 -3236
rect 12683 -3286 12699 -3252
rect 12807 -3286 12823 -3252
rect 12683 -3333 12823 -3286
rect 12881 -3252 13021 -3236
rect 12881 -3286 12897 -3252
rect 13005 -3286 13021 -3252
rect 12881 -3333 13021 -3286
rect 13079 -3252 13219 -3236
rect 13079 -3286 13095 -3252
rect 13203 -3286 13219 -3252
rect 13079 -3333 13219 -3286
rect 13277 -3252 13417 -3236
rect 13277 -3286 13293 -3252
rect 13401 -3286 13417 -3252
rect 13277 -3333 13417 -3286
rect 13475 -3252 13615 -3236
rect 13475 -3286 13491 -3252
rect 13599 -3286 13615 -3252
rect 13475 -3333 13615 -3286
rect 13673 -3252 13813 -3236
rect 13673 -3286 13689 -3252
rect 13797 -3286 13813 -3252
rect 13673 -3333 13813 -3286
rect 13871 -3252 14011 -3236
rect 13871 -3286 13887 -3252
rect 13995 -3286 14011 -3252
rect 13871 -3333 14011 -3286
rect 14069 -3252 14209 -3236
rect 14069 -3286 14085 -3252
rect 14193 -3286 14209 -3252
rect 14069 -3333 14209 -3286
rect 14267 -3252 14407 -3236
rect 14267 -3286 14283 -3252
rect 14391 -3286 14407 -3252
rect 14267 -3333 14407 -3286
rect 14465 -3252 14605 -3236
rect 14465 -3286 14481 -3252
rect 14589 -3286 14605 -3252
rect 14465 -3333 14605 -3286
rect 14663 -3252 14803 -3236
rect 14663 -3286 14679 -3252
rect 14787 -3286 14803 -3252
rect 14663 -3333 14803 -3286
rect 14861 -3252 15001 -3236
rect 14861 -3286 14877 -3252
rect 14985 -3286 15001 -3252
rect 14861 -3333 15001 -3286
rect 15059 -3252 15199 -3236
rect 15059 -3286 15075 -3252
rect 15183 -3286 15199 -3252
rect 15059 -3333 15199 -3286
rect 15257 -3252 15397 -3236
rect 15257 -3286 15273 -3252
rect 15381 -3286 15397 -3252
rect 15257 -3333 15397 -3286
rect 15455 -3252 15595 -3236
rect 15455 -3286 15471 -3252
rect 15579 -3286 15595 -3252
rect 15455 -3333 15595 -3286
rect 15653 -3252 15793 -3236
rect 15653 -3286 15669 -3252
rect 15777 -3286 15793 -3252
rect 15653 -3333 15793 -3286
rect 15851 -3252 15991 -3236
rect 15851 -3286 15867 -3252
rect 15975 -3286 15991 -3252
rect 15851 -3333 15991 -3286
rect 16049 -3252 16189 -3236
rect 16049 -3286 16065 -3252
rect 16173 -3286 16189 -3252
rect 16049 -3333 16189 -3286
rect 16247 -3252 16387 -3236
rect 16247 -3286 16263 -3252
rect 16371 -3286 16387 -3252
rect 16247 -3333 16387 -3286
rect 16445 -3252 16585 -3236
rect 16445 -3286 16461 -3252
rect 16569 -3286 16585 -3252
rect 16445 -3333 16585 -3286
rect 16643 -3252 16783 -3236
rect 16643 -3286 16659 -3252
rect 16767 -3286 16783 -3252
rect 16643 -3333 16783 -3286
rect 16841 -3252 16981 -3236
rect 16841 -3286 16857 -3252
rect 16965 -3286 16981 -3252
rect 16841 -3333 16981 -3286
rect 17039 -3252 17179 -3236
rect 17039 -3286 17055 -3252
rect 17163 -3286 17179 -3252
rect 17039 -3333 17179 -3286
rect 17237 -3252 17377 -3236
rect 17237 -3286 17253 -3252
rect 17361 -3286 17377 -3252
rect 17237 -3333 17377 -3286
rect 17435 -3252 17575 -3236
rect 17435 -3286 17451 -3252
rect 17559 -3286 17575 -3252
rect 17435 -3333 17575 -3286
rect 17633 -3252 17773 -3236
rect 17633 -3286 17649 -3252
rect 17757 -3286 17773 -3252
rect 17633 -3333 17773 -3286
rect 17831 -3252 17971 -3236
rect 17831 -3286 17847 -3252
rect 17955 -3286 17971 -3252
rect 17831 -3333 17971 -3286
rect 18029 -3252 18169 -3236
rect 18029 -3286 18045 -3252
rect 18153 -3286 18169 -3252
rect 18029 -3333 18169 -3286
rect 18227 -3252 18367 -3236
rect 18227 -3286 18243 -3252
rect 18351 -3286 18367 -3252
rect 18227 -3333 18367 -3286
rect 18425 -3252 18565 -3236
rect 18425 -3286 18441 -3252
rect 18549 -3286 18565 -3252
rect 18425 -3333 18565 -3286
rect 18623 -3252 18763 -3236
rect 18623 -3286 18639 -3252
rect 18747 -3286 18763 -3252
rect 18623 -3333 18763 -3286
rect 18821 -3252 18961 -3236
rect 18821 -3286 18837 -3252
rect 18945 -3286 18961 -3252
rect 18821 -3333 18961 -3286
rect 19019 -3252 19159 -3236
rect 19019 -3286 19035 -3252
rect 19143 -3286 19159 -3252
rect 19019 -3333 19159 -3286
rect 19217 -3252 19357 -3236
rect 19217 -3286 19233 -3252
rect 19341 -3286 19357 -3252
rect 19217 -3333 19357 -3286
rect 19415 -3252 19555 -3236
rect 19415 -3286 19431 -3252
rect 19539 -3286 19555 -3252
rect 19415 -3333 19555 -3286
rect 19613 -3252 19753 -3236
rect 19613 -3286 19629 -3252
rect 19737 -3286 19753 -3252
rect 19613 -3333 19753 -3286
rect 23345 2140 23485 2166
rect 23543 2140 23683 2166
rect 23741 2140 23881 2166
rect 23939 2140 24079 2166
rect 24137 2140 24277 2166
rect 24335 2140 24475 2166
rect 24533 2140 24673 2166
rect 24731 2140 24871 2166
rect 24929 2140 25069 2166
rect 25127 2140 25267 2166
rect 25325 2140 25465 2166
rect 25523 2140 25663 2166
rect 25721 2140 25861 2166
rect 25919 2140 26059 2166
rect 26117 2140 26257 2166
rect 26315 2140 26455 2166
rect 26513 2140 26653 2166
rect 26711 2140 26851 2166
rect 26909 2140 27049 2166
rect 27107 2140 27247 2166
rect 27305 2140 27445 2166
rect 27503 2140 27643 2166
rect 27701 2140 27841 2166
rect 27899 2140 28039 2166
rect 28097 2140 28237 2166
rect 28295 2140 28435 2166
rect 28493 2140 28633 2166
rect 28691 2140 28831 2166
rect 28889 2140 29029 2166
rect 29087 2140 29227 2166
rect 29285 2140 29425 2166
rect 29483 2140 29623 2166
rect 29681 2140 29821 2166
rect 29879 2140 30019 2166
rect 30077 2140 30217 2166
rect 30275 2140 30415 2166
rect 30473 2140 30613 2166
rect 30671 2140 30811 2166
rect 30869 2140 31009 2166
rect 31067 2140 31207 2166
rect 31265 2140 31405 2166
rect 31463 2140 31603 2166
rect 11495 -4759 11635 -4733
rect 11693 -4759 11833 -4733
rect 11891 -4759 12031 -4733
rect 12089 -4759 12229 -4733
rect 12287 -4759 12427 -4733
rect 12485 -4759 12625 -4733
rect 12683 -4759 12823 -4733
rect 12881 -4759 13021 -4733
rect 13079 -4759 13219 -4733
rect 13277 -4759 13417 -4733
rect 13475 -4759 13615 -4733
rect 13673 -4759 13813 -4733
rect 13871 -4759 14011 -4733
rect 14069 -4759 14209 -4733
rect 14267 -4759 14407 -4733
rect 14465 -4759 14605 -4733
rect 14663 -4759 14803 -4733
rect 14861 -4759 15001 -4733
rect 15059 -4759 15199 -4733
rect 15257 -4759 15397 -4733
rect 15455 -4759 15595 -4733
rect 15653 -4759 15793 -4733
rect 15851 -4759 15991 -4733
rect 16049 -4759 16189 -4733
rect 16247 -4759 16387 -4733
rect 16445 -4759 16585 -4733
rect 16643 -4759 16783 -4733
rect 16841 -4759 16981 -4733
rect 17039 -4759 17179 -4733
rect 17237 -4759 17377 -4733
rect 17435 -4759 17575 -4733
rect 17633 -4759 17773 -4733
rect 17831 -4759 17971 -4733
rect 18029 -4759 18169 -4733
rect 18227 -4759 18367 -4733
rect 18425 -4759 18565 -4733
rect 18623 -4759 18763 -4733
rect 18821 -4759 18961 -4733
rect 19019 -4759 19159 -4733
rect 19217 -4759 19357 -4733
rect 19415 -4759 19555 -4733
rect 19613 -4759 19753 -4733
rect 23345 693 23485 740
rect 23345 659 23361 693
rect 23469 659 23485 693
rect 23345 643 23485 659
rect 23543 693 23683 740
rect 23543 659 23559 693
rect 23667 659 23683 693
rect 23543 643 23683 659
rect 23741 693 23881 740
rect 23741 659 23757 693
rect 23865 659 23881 693
rect 23741 643 23881 659
rect 23939 693 24079 740
rect 23939 659 23955 693
rect 24063 659 24079 693
rect 23939 643 24079 659
rect 24137 693 24277 740
rect 24137 659 24153 693
rect 24261 659 24277 693
rect 24137 643 24277 659
rect 24335 693 24475 740
rect 24335 659 24351 693
rect 24459 659 24475 693
rect 24335 643 24475 659
rect 24533 693 24673 740
rect 24533 659 24549 693
rect 24657 659 24673 693
rect 24533 643 24673 659
rect 24731 693 24871 740
rect 24731 659 24747 693
rect 24855 659 24871 693
rect 24731 643 24871 659
rect 24929 693 25069 740
rect 24929 659 24945 693
rect 25053 659 25069 693
rect 24929 643 25069 659
rect 25127 693 25267 740
rect 25127 659 25143 693
rect 25251 659 25267 693
rect 25127 643 25267 659
rect 25325 693 25465 740
rect 25325 659 25341 693
rect 25449 659 25465 693
rect 25325 643 25465 659
rect 25523 693 25663 740
rect 25523 659 25539 693
rect 25647 659 25663 693
rect 25523 643 25663 659
rect 25721 693 25861 740
rect 25721 659 25737 693
rect 25845 659 25861 693
rect 25721 643 25861 659
rect 25919 693 26059 740
rect 25919 659 25935 693
rect 26043 659 26059 693
rect 25919 643 26059 659
rect 26117 693 26257 740
rect 26117 659 26133 693
rect 26241 659 26257 693
rect 26117 643 26257 659
rect 26315 693 26455 740
rect 26315 659 26331 693
rect 26439 659 26455 693
rect 26315 643 26455 659
rect 26513 693 26653 740
rect 26513 659 26529 693
rect 26637 659 26653 693
rect 26513 643 26653 659
rect 26711 693 26851 740
rect 26711 659 26727 693
rect 26835 659 26851 693
rect 26711 643 26851 659
rect 26909 693 27049 740
rect 26909 659 26925 693
rect 27033 659 27049 693
rect 26909 643 27049 659
rect 27107 693 27247 740
rect 27107 659 27123 693
rect 27231 659 27247 693
rect 27107 643 27247 659
rect 27305 693 27445 740
rect 27305 659 27321 693
rect 27429 659 27445 693
rect 27305 643 27445 659
rect 27503 693 27643 740
rect 27503 659 27519 693
rect 27627 659 27643 693
rect 27503 643 27643 659
rect 27701 693 27841 740
rect 27701 659 27717 693
rect 27825 659 27841 693
rect 27701 643 27841 659
rect 27899 693 28039 740
rect 27899 659 27915 693
rect 28023 659 28039 693
rect 27899 643 28039 659
rect 28097 693 28237 740
rect 28097 659 28113 693
rect 28221 659 28237 693
rect 28097 643 28237 659
rect 28295 693 28435 740
rect 28295 659 28311 693
rect 28419 659 28435 693
rect 28295 643 28435 659
rect 28493 693 28633 740
rect 28493 659 28509 693
rect 28617 659 28633 693
rect 28493 643 28633 659
rect 28691 693 28831 740
rect 28691 659 28707 693
rect 28815 659 28831 693
rect 28691 643 28831 659
rect 28889 693 29029 740
rect 28889 659 28905 693
rect 29013 659 29029 693
rect 28889 643 29029 659
rect 29087 693 29227 740
rect 29087 659 29103 693
rect 29211 659 29227 693
rect 29087 643 29227 659
rect 29285 693 29425 740
rect 29285 659 29301 693
rect 29409 659 29425 693
rect 29285 643 29425 659
rect 29483 693 29623 740
rect 29483 659 29499 693
rect 29607 659 29623 693
rect 29483 643 29623 659
rect 29681 693 29821 740
rect 29681 659 29697 693
rect 29805 659 29821 693
rect 29681 643 29821 659
rect 29879 693 30019 740
rect 29879 659 29895 693
rect 30003 659 30019 693
rect 29879 643 30019 659
rect 30077 693 30217 740
rect 30077 659 30093 693
rect 30201 659 30217 693
rect 30077 643 30217 659
rect 30275 693 30415 740
rect 30275 659 30291 693
rect 30399 659 30415 693
rect 30275 643 30415 659
rect 30473 693 30613 740
rect 30473 659 30489 693
rect 30597 659 30613 693
rect 30473 643 30613 659
rect 30671 693 30811 740
rect 30671 659 30687 693
rect 30795 659 30811 693
rect 30671 643 30811 659
rect 30869 693 31009 740
rect 30869 659 30885 693
rect 30993 659 31009 693
rect 30869 643 31009 659
rect 31067 693 31207 740
rect 31067 659 31083 693
rect 31191 659 31207 693
rect 31067 643 31207 659
rect 31265 693 31405 740
rect 31265 659 31281 693
rect 31389 659 31405 693
rect 31265 643 31405 659
rect 31463 693 31603 740
rect 31463 659 31479 693
rect 31587 659 31603 693
rect 31463 643 31603 659
rect 23345 585 23485 601
rect 23345 551 23361 585
rect 23469 551 23485 585
rect 23345 504 23485 551
rect 23543 585 23683 601
rect 23543 551 23559 585
rect 23667 551 23683 585
rect 23543 504 23683 551
rect 23741 585 23881 601
rect 23741 551 23757 585
rect 23865 551 23881 585
rect 23741 504 23881 551
rect 23939 585 24079 601
rect 23939 551 23955 585
rect 24063 551 24079 585
rect 23939 504 24079 551
rect 24137 585 24277 601
rect 24137 551 24153 585
rect 24261 551 24277 585
rect 24137 504 24277 551
rect 24335 585 24475 601
rect 24335 551 24351 585
rect 24459 551 24475 585
rect 24335 504 24475 551
rect 24533 585 24673 601
rect 24533 551 24549 585
rect 24657 551 24673 585
rect 24533 504 24673 551
rect 24731 585 24871 601
rect 24731 551 24747 585
rect 24855 551 24871 585
rect 24731 504 24871 551
rect 24929 585 25069 601
rect 24929 551 24945 585
rect 25053 551 25069 585
rect 24929 504 25069 551
rect 25127 585 25267 601
rect 25127 551 25143 585
rect 25251 551 25267 585
rect 25127 504 25267 551
rect 25325 585 25465 601
rect 25325 551 25341 585
rect 25449 551 25465 585
rect 25325 504 25465 551
rect 25523 585 25663 601
rect 25523 551 25539 585
rect 25647 551 25663 585
rect 25523 504 25663 551
rect 25721 585 25861 601
rect 25721 551 25737 585
rect 25845 551 25861 585
rect 25721 504 25861 551
rect 25919 585 26059 601
rect 25919 551 25935 585
rect 26043 551 26059 585
rect 25919 504 26059 551
rect 26117 585 26257 601
rect 26117 551 26133 585
rect 26241 551 26257 585
rect 26117 504 26257 551
rect 26315 585 26455 601
rect 26315 551 26331 585
rect 26439 551 26455 585
rect 26315 504 26455 551
rect 26513 585 26653 601
rect 26513 551 26529 585
rect 26637 551 26653 585
rect 26513 504 26653 551
rect 26711 585 26851 601
rect 26711 551 26727 585
rect 26835 551 26851 585
rect 26711 504 26851 551
rect 26909 585 27049 601
rect 26909 551 26925 585
rect 27033 551 27049 585
rect 26909 504 27049 551
rect 27107 585 27247 601
rect 27107 551 27123 585
rect 27231 551 27247 585
rect 27107 504 27247 551
rect 27305 585 27445 601
rect 27305 551 27321 585
rect 27429 551 27445 585
rect 27305 504 27445 551
rect 27503 585 27643 601
rect 27503 551 27519 585
rect 27627 551 27643 585
rect 27503 504 27643 551
rect 27701 585 27841 601
rect 27701 551 27717 585
rect 27825 551 27841 585
rect 27701 504 27841 551
rect 27899 585 28039 601
rect 27899 551 27915 585
rect 28023 551 28039 585
rect 27899 504 28039 551
rect 28097 585 28237 601
rect 28097 551 28113 585
rect 28221 551 28237 585
rect 28097 504 28237 551
rect 28295 585 28435 601
rect 28295 551 28311 585
rect 28419 551 28435 585
rect 28295 504 28435 551
rect 28493 585 28633 601
rect 28493 551 28509 585
rect 28617 551 28633 585
rect 28493 504 28633 551
rect 28691 585 28831 601
rect 28691 551 28707 585
rect 28815 551 28831 585
rect 28691 504 28831 551
rect 28889 585 29029 601
rect 28889 551 28905 585
rect 29013 551 29029 585
rect 28889 504 29029 551
rect 29087 585 29227 601
rect 29087 551 29103 585
rect 29211 551 29227 585
rect 29087 504 29227 551
rect 29285 585 29425 601
rect 29285 551 29301 585
rect 29409 551 29425 585
rect 29285 504 29425 551
rect 29483 585 29623 601
rect 29483 551 29499 585
rect 29607 551 29623 585
rect 29483 504 29623 551
rect 29681 585 29821 601
rect 29681 551 29697 585
rect 29805 551 29821 585
rect 29681 504 29821 551
rect 29879 585 30019 601
rect 29879 551 29895 585
rect 30003 551 30019 585
rect 29879 504 30019 551
rect 30077 585 30217 601
rect 30077 551 30093 585
rect 30201 551 30217 585
rect 30077 504 30217 551
rect 30275 585 30415 601
rect 30275 551 30291 585
rect 30399 551 30415 585
rect 30275 504 30415 551
rect 30473 585 30613 601
rect 30473 551 30489 585
rect 30597 551 30613 585
rect 30473 504 30613 551
rect 30671 585 30811 601
rect 30671 551 30687 585
rect 30795 551 30811 585
rect 30671 504 30811 551
rect 30869 585 31009 601
rect 30869 551 30885 585
rect 30993 551 31009 585
rect 30869 504 31009 551
rect 31067 585 31207 601
rect 31067 551 31083 585
rect 31191 551 31207 585
rect 31067 504 31207 551
rect 31265 585 31405 601
rect 31265 551 31281 585
rect 31389 551 31405 585
rect 31265 504 31405 551
rect 31463 585 31603 601
rect 31463 551 31479 585
rect 31587 551 31603 585
rect 31463 504 31603 551
rect 23345 -943 23485 -896
rect 23345 -977 23361 -943
rect 23469 -977 23485 -943
rect 23345 -993 23485 -977
rect 23543 -943 23683 -896
rect 23543 -977 23559 -943
rect 23667 -977 23683 -943
rect 23543 -993 23683 -977
rect 23741 -943 23881 -896
rect 23741 -977 23757 -943
rect 23865 -977 23881 -943
rect 23741 -993 23881 -977
rect 23939 -943 24079 -896
rect 23939 -977 23955 -943
rect 24063 -977 24079 -943
rect 23939 -993 24079 -977
rect 24137 -943 24277 -896
rect 24137 -977 24153 -943
rect 24261 -977 24277 -943
rect 24137 -993 24277 -977
rect 24335 -943 24475 -896
rect 24335 -977 24351 -943
rect 24459 -977 24475 -943
rect 24335 -993 24475 -977
rect 24533 -943 24673 -896
rect 24533 -977 24549 -943
rect 24657 -977 24673 -943
rect 24533 -993 24673 -977
rect 24731 -943 24871 -896
rect 24731 -977 24747 -943
rect 24855 -977 24871 -943
rect 24731 -993 24871 -977
rect 24929 -943 25069 -896
rect 24929 -977 24945 -943
rect 25053 -977 25069 -943
rect 24929 -993 25069 -977
rect 25127 -943 25267 -896
rect 25127 -977 25143 -943
rect 25251 -977 25267 -943
rect 25127 -993 25267 -977
rect 25325 -943 25465 -896
rect 25325 -977 25341 -943
rect 25449 -977 25465 -943
rect 25325 -993 25465 -977
rect 25523 -943 25663 -896
rect 25523 -977 25539 -943
rect 25647 -977 25663 -943
rect 25523 -993 25663 -977
rect 25721 -943 25861 -896
rect 25721 -977 25737 -943
rect 25845 -977 25861 -943
rect 25721 -993 25861 -977
rect 25919 -943 26059 -896
rect 25919 -977 25935 -943
rect 26043 -977 26059 -943
rect 25919 -993 26059 -977
rect 26117 -943 26257 -896
rect 26117 -977 26133 -943
rect 26241 -977 26257 -943
rect 26117 -993 26257 -977
rect 26315 -943 26455 -896
rect 26315 -977 26331 -943
rect 26439 -977 26455 -943
rect 26315 -993 26455 -977
rect 26513 -943 26653 -896
rect 26513 -977 26529 -943
rect 26637 -977 26653 -943
rect 26513 -993 26653 -977
rect 26711 -943 26851 -896
rect 26711 -977 26727 -943
rect 26835 -977 26851 -943
rect 26711 -993 26851 -977
rect 26909 -943 27049 -896
rect 26909 -977 26925 -943
rect 27033 -977 27049 -943
rect 26909 -993 27049 -977
rect 27107 -943 27247 -896
rect 27107 -977 27123 -943
rect 27231 -977 27247 -943
rect 27107 -993 27247 -977
rect 27305 -943 27445 -896
rect 27305 -977 27321 -943
rect 27429 -977 27445 -943
rect 27305 -993 27445 -977
rect 27503 -943 27643 -896
rect 27503 -977 27519 -943
rect 27627 -977 27643 -943
rect 27503 -993 27643 -977
rect 27701 -943 27841 -896
rect 27701 -977 27717 -943
rect 27825 -977 27841 -943
rect 27701 -993 27841 -977
rect 27899 -943 28039 -896
rect 27899 -977 27915 -943
rect 28023 -977 28039 -943
rect 27899 -993 28039 -977
rect 28097 -943 28237 -896
rect 28097 -977 28113 -943
rect 28221 -977 28237 -943
rect 28097 -993 28237 -977
rect 28295 -943 28435 -896
rect 28295 -977 28311 -943
rect 28419 -977 28435 -943
rect 28295 -993 28435 -977
rect 28493 -943 28633 -896
rect 28493 -977 28509 -943
rect 28617 -977 28633 -943
rect 28493 -993 28633 -977
rect 28691 -943 28831 -896
rect 28691 -977 28707 -943
rect 28815 -977 28831 -943
rect 28691 -993 28831 -977
rect 28889 -943 29029 -896
rect 28889 -977 28905 -943
rect 29013 -977 29029 -943
rect 28889 -993 29029 -977
rect 29087 -943 29227 -896
rect 29087 -977 29103 -943
rect 29211 -977 29227 -943
rect 29087 -993 29227 -977
rect 29285 -943 29425 -896
rect 29285 -977 29301 -943
rect 29409 -977 29425 -943
rect 29285 -993 29425 -977
rect 29483 -943 29623 -896
rect 29483 -977 29499 -943
rect 29607 -977 29623 -943
rect 29483 -993 29623 -977
rect 29681 -943 29821 -896
rect 29681 -977 29697 -943
rect 29805 -977 29821 -943
rect 29681 -993 29821 -977
rect 29879 -943 30019 -896
rect 29879 -977 29895 -943
rect 30003 -977 30019 -943
rect 29879 -993 30019 -977
rect 30077 -943 30217 -896
rect 30077 -977 30093 -943
rect 30201 -977 30217 -943
rect 30077 -993 30217 -977
rect 30275 -943 30415 -896
rect 30275 -977 30291 -943
rect 30399 -977 30415 -943
rect 30275 -993 30415 -977
rect 30473 -943 30613 -896
rect 30473 -977 30489 -943
rect 30597 -977 30613 -943
rect 30473 -993 30613 -977
rect 30671 -943 30811 -896
rect 30671 -977 30687 -943
rect 30795 -977 30811 -943
rect 30671 -993 30811 -977
rect 30869 -943 31009 -896
rect 30869 -977 30885 -943
rect 30993 -977 31009 -943
rect 30869 -993 31009 -977
rect 31067 -943 31207 -896
rect 31067 -977 31083 -943
rect 31191 -977 31207 -943
rect 31067 -993 31207 -977
rect 31265 -943 31405 -896
rect 31265 -977 31281 -943
rect 31389 -977 31405 -943
rect 31265 -993 31405 -977
rect 31463 -943 31603 -896
rect 31463 -977 31479 -943
rect 31587 -977 31603 -943
rect 31463 -993 31603 -977
rect 23345 -1051 23485 -1035
rect 23345 -1085 23361 -1051
rect 23469 -1085 23485 -1051
rect 23345 -1132 23485 -1085
rect 23543 -1051 23683 -1035
rect 23543 -1085 23559 -1051
rect 23667 -1085 23683 -1051
rect 23543 -1132 23683 -1085
rect 23741 -1051 23881 -1035
rect 23741 -1085 23757 -1051
rect 23865 -1085 23881 -1051
rect 23741 -1132 23881 -1085
rect 23939 -1051 24079 -1035
rect 23939 -1085 23955 -1051
rect 24063 -1085 24079 -1051
rect 23939 -1132 24079 -1085
rect 24137 -1051 24277 -1035
rect 24137 -1085 24153 -1051
rect 24261 -1085 24277 -1051
rect 24137 -1132 24277 -1085
rect 24335 -1051 24475 -1035
rect 24335 -1085 24351 -1051
rect 24459 -1085 24475 -1051
rect 24335 -1132 24475 -1085
rect 24533 -1051 24673 -1035
rect 24533 -1085 24549 -1051
rect 24657 -1085 24673 -1051
rect 24533 -1132 24673 -1085
rect 24731 -1051 24871 -1035
rect 24731 -1085 24747 -1051
rect 24855 -1085 24871 -1051
rect 24731 -1132 24871 -1085
rect 24929 -1051 25069 -1035
rect 24929 -1085 24945 -1051
rect 25053 -1085 25069 -1051
rect 24929 -1132 25069 -1085
rect 25127 -1051 25267 -1035
rect 25127 -1085 25143 -1051
rect 25251 -1085 25267 -1051
rect 25127 -1132 25267 -1085
rect 25325 -1051 25465 -1035
rect 25325 -1085 25341 -1051
rect 25449 -1085 25465 -1051
rect 25325 -1132 25465 -1085
rect 25523 -1051 25663 -1035
rect 25523 -1085 25539 -1051
rect 25647 -1085 25663 -1051
rect 25523 -1132 25663 -1085
rect 25721 -1051 25861 -1035
rect 25721 -1085 25737 -1051
rect 25845 -1085 25861 -1051
rect 25721 -1132 25861 -1085
rect 25919 -1051 26059 -1035
rect 25919 -1085 25935 -1051
rect 26043 -1085 26059 -1051
rect 25919 -1132 26059 -1085
rect 26117 -1051 26257 -1035
rect 26117 -1085 26133 -1051
rect 26241 -1085 26257 -1051
rect 26117 -1132 26257 -1085
rect 26315 -1051 26455 -1035
rect 26315 -1085 26331 -1051
rect 26439 -1085 26455 -1051
rect 26315 -1132 26455 -1085
rect 26513 -1051 26653 -1035
rect 26513 -1085 26529 -1051
rect 26637 -1085 26653 -1051
rect 26513 -1132 26653 -1085
rect 26711 -1051 26851 -1035
rect 26711 -1085 26727 -1051
rect 26835 -1085 26851 -1051
rect 26711 -1132 26851 -1085
rect 26909 -1051 27049 -1035
rect 26909 -1085 26925 -1051
rect 27033 -1085 27049 -1051
rect 26909 -1132 27049 -1085
rect 27107 -1051 27247 -1035
rect 27107 -1085 27123 -1051
rect 27231 -1085 27247 -1051
rect 27107 -1132 27247 -1085
rect 27305 -1051 27445 -1035
rect 27305 -1085 27321 -1051
rect 27429 -1085 27445 -1051
rect 27305 -1132 27445 -1085
rect 27503 -1051 27643 -1035
rect 27503 -1085 27519 -1051
rect 27627 -1085 27643 -1051
rect 27503 -1132 27643 -1085
rect 27701 -1051 27841 -1035
rect 27701 -1085 27717 -1051
rect 27825 -1085 27841 -1051
rect 27701 -1132 27841 -1085
rect 27899 -1051 28039 -1035
rect 27899 -1085 27915 -1051
rect 28023 -1085 28039 -1051
rect 27899 -1132 28039 -1085
rect 28097 -1051 28237 -1035
rect 28097 -1085 28113 -1051
rect 28221 -1085 28237 -1051
rect 28097 -1132 28237 -1085
rect 28295 -1051 28435 -1035
rect 28295 -1085 28311 -1051
rect 28419 -1085 28435 -1051
rect 28295 -1132 28435 -1085
rect 28493 -1051 28633 -1035
rect 28493 -1085 28509 -1051
rect 28617 -1085 28633 -1051
rect 28493 -1132 28633 -1085
rect 28691 -1051 28831 -1035
rect 28691 -1085 28707 -1051
rect 28815 -1085 28831 -1051
rect 28691 -1132 28831 -1085
rect 28889 -1051 29029 -1035
rect 28889 -1085 28905 -1051
rect 29013 -1085 29029 -1051
rect 28889 -1132 29029 -1085
rect 29087 -1051 29227 -1035
rect 29087 -1085 29103 -1051
rect 29211 -1085 29227 -1051
rect 29087 -1132 29227 -1085
rect 29285 -1051 29425 -1035
rect 29285 -1085 29301 -1051
rect 29409 -1085 29425 -1051
rect 29285 -1132 29425 -1085
rect 29483 -1051 29623 -1035
rect 29483 -1085 29499 -1051
rect 29607 -1085 29623 -1051
rect 29483 -1132 29623 -1085
rect 29681 -1051 29821 -1035
rect 29681 -1085 29697 -1051
rect 29805 -1085 29821 -1051
rect 29681 -1132 29821 -1085
rect 29879 -1051 30019 -1035
rect 29879 -1085 29895 -1051
rect 30003 -1085 30019 -1051
rect 29879 -1132 30019 -1085
rect 30077 -1051 30217 -1035
rect 30077 -1085 30093 -1051
rect 30201 -1085 30217 -1051
rect 30077 -1132 30217 -1085
rect 30275 -1051 30415 -1035
rect 30275 -1085 30291 -1051
rect 30399 -1085 30415 -1051
rect 30275 -1132 30415 -1085
rect 30473 -1051 30613 -1035
rect 30473 -1085 30489 -1051
rect 30597 -1085 30613 -1051
rect 30473 -1132 30613 -1085
rect 30671 -1051 30811 -1035
rect 30671 -1085 30687 -1051
rect 30795 -1085 30811 -1051
rect 30671 -1132 30811 -1085
rect 30869 -1051 31009 -1035
rect 30869 -1085 30885 -1051
rect 30993 -1085 31009 -1051
rect 30869 -1132 31009 -1085
rect 31067 -1051 31207 -1035
rect 31067 -1085 31083 -1051
rect 31191 -1085 31207 -1051
rect 31067 -1132 31207 -1085
rect 31265 -1051 31405 -1035
rect 31265 -1085 31281 -1051
rect 31389 -1085 31405 -1051
rect 31265 -1132 31405 -1085
rect 31463 -1051 31603 -1035
rect 31463 -1085 31479 -1051
rect 31587 -1085 31603 -1051
rect 31463 -1132 31603 -1085
rect 23345 -2579 23485 -2532
rect 23345 -2613 23361 -2579
rect 23469 -2613 23485 -2579
rect 23345 -2629 23485 -2613
rect 23543 -2579 23683 -2532
rect 23543 -2613 23559 -2579
rect 23667 -2613 23683 -2579
rect 23543 -2629 23683 -2613
rect 23741 -2579 23881 -2532
rect 23741 -2613 23757 -2579
rect 23865 -2613 23881 -2579
rect 23741 -2629 23881 -2613
rect 23939 -2579 24079 -2532
rect 23939 -2613 23955 -2579
rect 24063 -2613 24079 -2579
rect 23939 -2629 24079 -2613
rect 24137 -2579 24277 -2532
rect 24137 -2613 24153 -2579
rect 24261 -2613 24277 -2579
rect 24137 -2629 24277 -2613
rect 24335 -2579 24475 -2532
rect 24335 -2613 24351 -2579
rect 24459 -2613 24475 -2579
rect 24335 -2629 24475 -2613
rect 24533 -2579 24673 -2532
rect 24533 -2613 24549 -2579
rect 24657 -2613 24673 -2579
rect 24533 -2629 24673 -2613
rect 24731 -2579 24871 -2532
rect 24731 -2613 24747 -2579
rect 24855 -2613 24871 -2579
rect 24731 -2629 24871 -2613
rect 24929 -2579 25069 -2532
rect 24929 -2613 24945 -2579
rect 25053 -2613 25069 -2579
rect 24929 -2629 25069 -2613
rect 25127 -2579 25267 -2532
rect 25127 -2613 25143 -2579
rect 25251 -2613 25267 -2579
rect 25127 -2629 25267 -2613
rect 25325 -2579 25465 -2532
rect 25325 -2613 25341 -2579
rect 25449 -2613 25465 -2579
rect 25325 -2629 25465 -2613
rect 25523 -2579 25663 -2532
rect 25523 -2613 25539 -2579
rect 25647 -2613 25663 -2579
rect 25523 -2629 25663 -2613
rect 25721 -2579 25861 -2532
rect 25721 -2613 25737 -2579
rect 25845 -2613 25861 -2579
rect 25721 -2629 25861 -2613
rect 25919 -2579 26059 -2532
rect 25919 -2613 25935 -2579
rect 26043 -2613 26059 -2579
rect 25919 -2629 26059 -2613
rect 26117 -2579 26257 -2532
rect 26117 -2613 26133 -2579
rect 26241 -2613 26257 -2579
rect 26117 -2629 26257 -2613
rect 26315 -2579 26455 -2532
rect 26315 -2613 26331 -2579
rect 26439 -2613 26455 -2579
rect 26315 -2629 26455 -2613
rect 26513 -2579 26653 -2532
rect 26513 -2613 26529 -2579
rect 26637 -2613 26653 -2579
rect 26513 -2629 26653 -2613
rect 26711 -2579 26851 -2532
rect 26711 -2613 26727 -2579
rect 26835 -2613 26851 -2579
rect 26711 -2629 26851 -2613
rect 26909 -2579 27049 -2532
rect 26909 -2613 26925 -2579
rect 27033 -2613 27049 -2579
rect 26909 -2629 27049 -2613
rect 27107 -2579 27247 -2532
rect 27107 -2613 27123 -2579
rect 27231 -2613 27247 -2579
rect 27107 -2629 27247 -2613
rect 27305 -2579 27445 -2532
rect 27305 -2613 27321 -2579
rect 27429 -2613 27445 -2579
rect 27305 -2629 27445 -2613
rect 27503 -2579 27643 -2532
rect 27503 -2613 27519 -2579
rect 27627 -2613 27643 -2579
rect 27503 -2629 27643 -2613
rect 27701 -2579 27841 -2532
rect 27701 -2613 27717 -2579
rect 27825 -2613 27841 -2579
rect 27701 -2629 27841 -2613
rect 27899 -2579 28039 -2532
rect 27899 -2613 27915 -2579
rect 28023 -2613 28039 -2579
rect 27899 -2629 28039 -2613
rect 28097 -2579 28237 -2532
rect 28097 -2613 28113 -2579
rect 28221 -2613 28237 -2579
rect 28097 -2629 28237 -2613
rect 28295 -2579 28435 -2532
rect 28295 -2613 28311 -2579
rect 28419 -2613 28435 -2579
rect 28295 -2629 28435 -2613
rect 28493 -2579 28633 -2532
rect 28493 -2613 28509 -2579
rect 28617 -2613 28633 -2579
rect 28493 -2629 28633 -2613
rect 28691 -2579 28831 -2532
rect 28691 -2613 28707 -2579
rect 28815 -2613 28831 -2579
rect 28691 -2629 28831 -2613
rect 28889 -2579 29029 -2532
rect 28889 -2613 28905 -2579
rect 29013 -2613 29029 -2579
rect 28889 -2629 29029 -2613
rect 29087 -2579 29227 -2532
rect 29087 -2613 29103 -2579
rect 29211 -2613 29227 -2579
rect 29087 -2629 29227 -2613
rect 29285 -2579 29425 -2532
rect 29285 -2613 29301 -2579
rect 29409 -2613 29425 -2579
rect 29285 -2629 29425 -2613
rect 29483 -2579 29623 -2532
rect 29483 -2613 29499 -2579
rect 29607 -2613 29623 -2579
rect 29483 -2629 29623 -2613
rect 29681 -2579 29821 -2532
rect 29681 -2613 29697 -2579
rect 29805 -2613 29821 -2579
rect 29681 -2629 29821 -2613
rect 29879 -2579 30019 -2532
rect 29879 -2613 29895 -2579
rect 30003 -2613 30019 -2579
rect 29879 -2629 30019 -2613
rect 30077 -2579 30217 -2532
rect 30077 -2613 30093 -2579
rect 30201 -2613 30217 -2579
rect 30077 -2629 30217 -2613
rect 30275 -2579 30415 -2532
rect 30275 -2613 30291 -2579
rect 30399 -2613 30415 -2579
rect 30275 -2629 30415 -2613
rect 30473 -2579 30613 -2532
rect 30473 -2613 30489 -2579
rect 30597 -2613 30613 -2579
rect 30473 -2629 30613 -2613
rect 30671 -2579 30811 -2532
rect 30671 -2613 30687 -2579
rect 30795 -2613 30811 -2579
rect 30671 -2629 30811 -2613
rect 30869 -2579 31009 -2532
rect 30869 -2613 30885 -2579
rect 30993 -2613 31009 -2579
rect 30869 -2629 31009 -2613
rect 31067 -2579 31207 -2532
rect 31067 -2613 31083 -2579
rect 31191 -2613 31207 -2579
rect 31067 -2629 31207 -2613
rect 31265 -2579 31405 -2532
rect 31265 -2613 31281 -2579
rect 31389 -2613 31405 -2579
rect 31265 -2629 31405 -2613
rect 31463 -2579 31603 -2532
rect 31463 -2613 31479 -2579
rect 31587 -2613 31603 -2579
rect 31463 -2629 31603 -2613
rect 23345 -3252 23485 -3236
rect 23345 -3286 23361 -3252
rect 23469 -3286 23485 -3252
rect 23345 -3333 23485 -3286
rect 23543 -3252 23683 -3236
rect 23543 -3286 23559 -3252
rect 23667 -3286 23683 -3252
rect 23543 -3333 23683 -3286
rect 23741 -3252 23881 -3236
rect 23741 -3286 23757 -3252
rect 23865 -3286 23881 -3252
rect 23741 -3333 23881 -3286
rect 23939 -3252 24079 -3236
rect 23939 -3286 23955 -3252
rect 24063 -3286 24079 -3252
rect 23939 -3333 24079 -3286
rect 24137 -3252 24277 -3236
rect 24137 -3286 24153 -3252
rect 24261 -3286 24277 -3252
rect 24137 -3333 24277 -3286
rect 24335 -3252 24475 -3236
rect 24335 -3286 24351 -3252
rect 24459 -3286 24475 -3252
rect 24335 -3333 24475 -3286
rect 24533 -3252 24673 -3236
rect 24533 -3286 24549 -3252
rect 24657 -3286 24673 -3252
rect 24533 -3333 24673 -3286
rect 24731 -3252 24871 -3236
rect 24731 -3286 24747 -3252
rect 24855 -3286 24871 -3252
rect 24731 -3333 24871 -3286
rect 24929 -3252 25069 -3236
rect 24929 -3286 24945 -3252
rect 25053 -3286 25069 -3252
rect 24929 -3333 25069 -3286
rect 25127 -3252 25267 -3236
rect 25127 -3286 25143 -3252
rect 25251 -3286 25267 -3252
rect 25127 -3333 25267 -3286
rect 25325 -3252 25465 -3236
rect 25325 -3286 25341 -3252
rect 25449 -3286 25465 -3252
rect 25325 -3333 25465 -3286
rect 25523 -3252 25663 -3236
rect 25523 -3286 25539 -3252
rect 25647 -3286 25663 -3252
rect 25523 -3333 25663 -3286
rect 25721 -3252 25861 -3236
rect 25721 -3286 25737 -3252
rect 25845 -3286 25861 -3252
rect 25721 -3333 25861 -3286
rect 25919 -3252 26059 -3236
rect 25919 -3286 25935 -3252
rect 26043 -3286 26059 -3252
rect 25919 -3333 26059 -3286
rect 26117 -3252 26257 -3236
rect 26117 -3286 26133 -3252
rect 26241 -3286 26257 -3252
rect 26117 -3333 26257 -3286
rect 26315 -3252 26455 -3236
rect 26315 -3286 26331 -3252
rect 26439 -3286 26455 -3252
rect 26315 -3333 26455 -3286
rect 26513 -3252 26653 -3236
rect 26513 -3286 26529 -3252
rect 26637 -3286 26653 -3252
rect 26513 -3333 26653 -3286
rect 26711 -3252 26851 -3236
rect 26711 -3286 26727 -3252
rect 26835 -3286 26851 -3252
rect 26711 -3333 26851 -3286
rect 26909 -3252 27049 -3236
rect 26909 -3286 26925 -3252
rect 27033 -3286 27049 -3252
rect 26909 -3333 27049 -3286
rect 27107 -3252 27247 -3236
rect 27107 -3286 27123 -3252
rect 27231 -3286 27247 -3252
rect 27107 -3333 27247 -3286
rect 27305 -3252 27445 -3236
rect 27305 -3286 27321 -3252
rect 27429 -3286 27445 -3252
rect 27305 -3333 27445 -3286
rect 27503 -3252 27643 -3236
rect 27503 -3286 27519 -3252
rect 27627 -3286 27643 -3252
rect 27503 -3333 27643 -3286
rect 27701 -3252 27841 -3236
rect 27701 -3286 27717 -3252
rect 27825 -3286 27841 -3252
rect 27701 -3333 27841 -3286
rect 27899 -3252 28039 -3236
rect 27899 -3286 27915 -3252
rect 28023 -3286 28039 -3252
rect 27899 -3333 28039 -3286
rect 28097 -3252 28237 -3236
rect 28097 -3286 28113 -3252
rect 28221 -3286 28237 -3252
rect 28097 -3333 28237 -3286
rect 28295 -3252 28435 -3236
rect 28295 -3286 28311 -3252
rect 28419 -3286 28435 -3252
rect 28295 -3333 28435 -3286
rect 28493 -3252 28633 -3236
rect 28493 -3286 28509 -3252
rect 28617 -3286 28633 -3252
rect 28493 -3333 28633 -3286
rect 28691 -3252 28831 -3236
rect 28691 -3286 28707 -3252
rect 28815 -3286 28831 -3252
rect 28691 -3333 28831 -3286
rect 28889 -3252 29029 -3236
rect 28889 -3286 28905 -3252
rect 29013 -3286 29029 -3252
rect 28889 -3333 29029 -3286
rect 29087 -3252 29227 -3236
rect 29087 -3286 29103 -3252
rect 29211 -3286 29227 -3252
rect 29087 -3333 29227 -3286
rect 29285 -3252 29425 -3236
rect 29285 -3286 29301 -3252
rect 29409 -3286 29425 -3252
rect 29285 -3333 29425 -3286
rect 29483 -3252 29623 -3236
rect 29483 -3286 29499 -3252
rect 29607 -3286 29623 -3252
rect 29483 -3333 29623 -3286
rect 29681 -3252 29821 -3236
rect 29681 -3286 29697 -3252
rect 29805 -3286 29821 -3252
rect 29681 -3333 29821 -3286
rect 29879 -3252 30019 -3236
rect 29879 -3286 29895 -3252
rect 30003 -3286 30019 -3252
rect 29879 -3333 30019 -3286
rect 30077 -3252 30217 -3236
rect 30077 -3286 30093 -3252
rect 30201 -3286 30217 -3252
rect 30077 -3333 30217 -3286
rect 30275 -3252 30415 -3236
rect 30275 -3286 30291 -3252
rect 30399 -3286 30415 -3252
rect 30275 -3333 30415 -3286
rect 30473 -3252 30613 -3236
rect 30473 -3286 30489 -3252
rect 30597 -3286 30613 -3252
rect 30473 -3333 30613 -3286
rect 30671 -3252 30811 -3236
rect 30671 -3286 30687 -3252
rect 30795 -3286 30811 -3252
rect 30671 -3333 30811 -3286
rect 30869 -3252 31009 -3236
rect 30869 -3286 30885 -3252
rect 30993 -3286 31009 -3252
rect 30869 -3333 31009 -3286
rect 31067 -3252 31207 -3236
rect 31067 -3286 31083 -3252
rect 31191 -3286 31207 -3252
rect 31067 -3333 31207 -3286
rect 31265 -3252 31405 -3236
rect 31265 -3286 31281 -3252
rect 31389 -3286 31405 -3252
rect 31265 -3333 31405 -3286
rect 31463 -3252 31603 -3236
rect 31463 -3286 31479 -3252
rect 31587 -3286 31603 -3252
rect 31463 -3333 31603 -3286
rect 23345 -4759 23485 -4733
rect 23543 -4759 23683 -4733
rect 23741 -4759 23881 -4733
rect 23939 -4759 24079 -4733
rect 24137 -4759 24277 -4733
rect 24335 -4759 24475 -4733
rect 24533 -4759 24673 -4733
rect 24731 -4759 24871 -4733
rect 24929 -4759 25069 -4733
rect 25127 -4759 25267 -4733
rect 25325 -4759 25465 -4733
rect 25523 -4759 25663 -4733
rect 25721 -4759 25861 -4733
rect 25919 -4759 26059 -4733
rect 26117 -4759 26257 -4733
rect 26315 -4759 26455 -4733
rect 26513 -4759 26653 -4733
rect 26711 -4759 26851 -4733
rect 26909 -4759 27049 -4733
rect 27107 -4759 27247 -4733
rect 27305 -4759 27445 -4733
rect 27503 -4759 27643 -4733
rect 27701 -4759 27841 -4733
rect 27899 -4759 28039 -4733
rect 28097 -4759 28237 -4733
rect 28295 -4759 28435 -4733
rect 28493 -4759 28633 -4733
rect 28691 -4759 28831 -4733
rect 28889 -4759 29029 -4733
rect 29087 -4759 29227 -4733
rect 29285 -4759 29425 -4733
rect 29483 -4759 29623 -4733
rect 29681 -4759 29821 -4733
rect 29879 -4759 30019 -4733
rect 30077 -4759 30217 -4733
rect 30275 -4759 30415 -4733
rect 30473 -4759 30613 -4733
rect 30671 -4759 30811 -4733
rect 30869 -4759 31009 -4733
rect 31067 -4759 31207 -4733
rect 31265 -4759 31405 -4733
rect 31463 -4759 31603 -4733
<< polycont >>
rect 11511 659 11619 693
rect 11709 659 11817 693
rect 11907 659 12015 693
rect 12105 659 12213 693
rect 12303 659 12411 693
rect 12501 659 12609 693
rect 12699 659 12807 693
rect 12897 659 13005 693
rect 13095 659 13203 693
rect 13293 659 13401 693
rect 13491 659 13599 693
rect 13689 659 13797 693
rect 13887 659 13995 693
rect 14085 659 14193 693
rect 14283 659 14391 693
rect 14481 659 14589 693
rect 14679 659 14787 693
rect 14877 659 14985 693
rect 15075 659 15183 693
rect 15273 659 15381 693
rect 15471 659 15579 693
rect 15669 659 15777 693
rect 15867 659 15975 693
rect 16065 659 16173 693
rect 16263 659 16371 693
rect 16461 659 16569 693
rect 16659 659 16767 693
rect 16857 659 16965 693
rect 17055 659 17163 693
rect 17253 659 17361 693
rect 17451 659 17559 693
rect 17649 659 17757 693
rect 17847 659 17955 693
rect 18045 659 18153 693
rect 18243 659 18351 693
rect 18441 659 18549 693
rect 18639 659 18747 693
rect 18837 659 18945 693
rect 19035 659 19143 693
rect 19233 659 19341 693
rect 19431 659 19539 693
rect 19629 659 19737 693
rect 11511 551 11619 585
rect 11709 551 11817 585
rect 11907 551 12015 585
rect 12105 551 12213 585
rect 12303 551 12411 585
rect 12501 551 12609 585
rect 12699 551 12807 585
rect 12897 551 13005 585
rect 13095 551 13203 585
rect 13293 551 13401 585
rect 13491 551 13599 585
rect 13689 551 13797 585
rect 13887 551 13995 585
rect 14085 551 14193 585
rect 14283 551 14391 585
rect 14481 551 14589 585
rect 14679 551 14787 585
rect 14877 551 14985 585
rect 15075 551 15183 585
rect 15273 551 15381 585
rect 15471 551 15579 585
rect 15669 551 15777 585
rect 15867 551 15975 585
rect 16065 551 16173 585
rect 16263 551 16371 585
rect 16461 551 16569 585
rect 16659 551 16767 585
rect 16857 551 16965 585
rect 17055 551 17163 585
rect 17253 551 17361 585
rect 17451 551 17559 585
rect 17649 551 17757 585
rect 17847 551 17955 585
rect 18045 551 18153 585
rect 18243 551 18351 585
rect 18441 551 18549 585
rect 18639 551 18747 585
rect 18837 551 18945 585
rect 19035 551 19143 585
rect 19233 551 19341 585
rect 19431 551 19539 585
rect 19629 551 19737 585
rect 11511 -977 11619 -943
rect 11709 -977 11817 -943
rect 11907 -977 12015 -943
rect 12105 -977 12213 -943
rect 12303 -977 12411 -943
rect 12501 -977 12609 -943
rect 12699 -977 12807 -943
rect 12897 -977 13005 -943
rect 13095 -977 13203 -943
rect 13293 -977 13401 -943
rect 13491 -977 13599 -943
rect 13689 -977 13797 -943
rect 13887 -977 13995 -943
rect 14085 -977 14193 -943
rect 14283 -977 14391 -943
rect 14481 -977 14589 -943
rect 14679 -977 14787 -943
rect 14877 -977 14985 -943
rect 15075 -977 15183 -943
rect 15273 -977 15381 -943
rect 15471 -977 15579 -943
rect 15669 -977 15777 -943
rect 15867 -977 15975 -943
rect 16065 -977 16173 -943
rect 16263 -977 16371 -943
rect 16461 -977 16569 -943
rect 16659 -977 16767 -943
rect 16857 -977 16965 -943
rect 17055 -977 17163 -943
rect 17253 -977 17361 -943
rect 17451 -977 17559 -943
rect 17649 -977 17757 -943
rect 17847 -977 17955 -943
rect 18045 -977 18153 -943
rect 18243 -977 18351 -943
rect 18441 -977 18549 -943
rect 18639 -977 18747 -943
rect 18837 -977 18945 -943
rect 19035 -977 19143 -943
rect 19233 -977 19341 -943
rect 19431 -977 19539 -943
rect 19629 -977 19737 -943
rect 11511 -1085 11619 -1051
rect 11709 -1085 11817 -1051
rect 11907 -1085 12015 -1051
rect 12105 -1085 12213 -1051
rect 12303 -1085 12411 -1051
rect 12501 -1085 12609 -1051
rect 12699 -1085 12807 -1051
rect 12897 -1085 13005 -1051
rect 13095 -1085 13203 -1051
rect 13293 -1085 13401 -1051
rect 13491 -1085 13599 -1051
rect 13689 -1085 13797 -1051
rect 13887 -1085 13995 -1051
rect 14085 -1085 14193 -1051
rect 14283 -1085 14391 -1051
rect 14481 -1085 14589 -1051
rect 14679 -1085 14787 -1051
rect 14877 -1085 14985 -1051
rect 15075 -1085 15183 -1051
rect 15273 -1085 15381 -1051
rect 15471 -1085 15579 -1051
rect 15669 -1085 15777 -1051
rect 15867 -1085 15975 -1051
rect 16065 -1085 16173 -1051
rect 16263 -1085 16371 -1051
rect 16461 -1085 16569 -1051
rect 16659 -1085 16767 -1051
rect 16857 -1085 16965 -1051
rect 17055 -1085 17163 -1051
rect 17253 -1085 17361 -1051
rect 17451 -1085 17559 -1051
rect 17649 -1085 17757 -1051
rect 17847 -1085 17955 -1051
rect 18045 -1085 18153 -1051
rect 18243 -1085 18351 -1051
rect 18441 -1085 18549 -1051
rect 18639 -1085 18747 -1051
rect 18837 -1085 18945 -1051
rect 19035 -1085 19143 -1051
rect 19233 -1085 19341 -1051
rect 19431 -1085 19539 -1051
rect 19629 -1085 19737 -1051
rect 11511 -2613 11619 -2579
rect 11709 -2613 11817 -2579
rect 11907 -2613 12015 -2579
rect 12105 -2613 12213 -2579
rect 12303 -2613 12411 -2579
rect 12501 -2613 12609 -2579
rect 12699 -2613 12807 -2579
rect 12897 -2613 13005 -2579
rect 13095 -2613 13203 -2579
rect 13293 -2613 13401 -2579
rect 13491 -2613 13599 -2579
rect 13689 -2613 13797 -2579
rect 13887 -2613 13995 -2579
rect 14085 -2613 14193 -2579
rect 14283 -2613 14391 -2579
rect 14481 -2613 14589 -2579
rect 14679 -2613 14787 -2579
rect 14877 -2613 14985 -2579
rect 15075 -2613 15183 -2579
rect 15273 -2613 15381 -2579
rect 15471 -2613 15579 -2579
rect 15669 -2613 15777 -2579
rect 15867 -2613 15975 -2579
rect 16065 -2613 16173 -2579
rect 16263 -2613 16371 -2579
rect 16461 -2613 16569 -2579
rect 16659 -2613 16767 -2579
rect 16857 -2613 16965 -2579
rect 17055 -2613 17163 -2579
rect 17253 -2613 17361 -2579
rect 17451 -2613 17559 -2579
rect 17649 -2613 17757 -2579
rect 17847 -2613 17955 -2579
rect 18045 -2613 18153 -2579
rect 18243 -2613 18351 -2579
rect 18441 -2613 18549 -2579
rect 18639 -2613 18747 -2579
rect 18837 -2613 18945 -2579
rect 19035 -2613 19143 -2579
rect 19233 -2613 19341 -2579
rect 19431 -2613 19539 -2579
rect 19629 -2613 19737 -2579
rect 11511 -3286 11619 -3252
rect 11709 -3286 11817 -3252
rect 11907 -3286 12015 -3252
rect 12105 -3286 12213 -3252
rect 12303 -3286 12411 -3252
rect 12501 -3286 12609 -3252
rect 12699 -3286 12807 -3252
rect 12897 -3286 13005 -3252
rect 13095 -3286 13203 -3252
rect 13293 -3286 13401 -3252
rect 13491 -3286 13599 -3252
rect 13689 -3286 13797 -3252
rect 13887 -3286 13995 -3252
rect 14085 -3286 14193 -3252
rect 14283 -3286 14391 -3252
rect 14481 -3286 14589 -3252
rect 14679 -3286 14787 -3252
rect 14877 -3286 14985 -3252
rect 15075 -3286 15183 -3252
rect 15273 -3286 15381 -3252
rect 15471 -3286 15579 -3252
rect 15669 -3286 15777 -3252
rect 15867 -3286 15975 -3252
rect 16065 -3286 16173 -3252
rect 16263 -3286 16371 -3252
rect 16461 -3286 16569 -3252
rect 16659 -3286 16767 -3252
rect 16857 -3286 16965 -3252
rect 17055 -3286 17163 -3252
rect 17253 -3286 17361 -3252
rect 17451 -3286 17559 -3252
rect 17649 -3286 17757 -3252
rect 17847 -3286 17955 -3252
rect 18045 -3286 18153 -3252
rect 18243 -3286 18351 -3252
rect 18441 -3286 18549 -3252
rect 18639 -3286 18747 -3252
rect 18837 -3286 18945 -3252
rect 19035 -3286 19143 -3252
rect 19233 -3286 19341 -3252
rect 19431 -3286 19539 -3252
rect 19629 -3286 19737 -3252
rect 23361 659 23469 693
rect 23559 659 23667 693
rect 23757 659 23865 693
rect 23955 659 24063 693
rect 24153 659 24261 693
rect 24351 659 24459 693
rect 24549 659 24657 693
rect 24747 659 24855 693
rect 24945 659 25053 693
rect 25143 659 25251 693
rect 25341 659 25449 693
rect 25539 659 25647 693
rect 25737 659 25845 693
rect 25935 659 26043 693
rect 26133 659 26241 693
rect 26331 659 26439 693
rect 26529 659 26637 693
rect 26727 659 26835 693
rect 26925 659 27033 693
rect 27123 659 27231 693
rect 27321 659 27429 693
rect 27519 659 27627 693
rect 27717 659 27825 693
rect 27915 659 28023 693
rect 28113 659 28221 693
rect 28311 659 28419 693
rect 28509 659 28617 693
rect 28707 659 28815 693
rect 28905 659 29013 693
rect 29103 659 29211 693
rect 29301 659 29409 693
rect 29499 659 29607 693
rect 29697 659 29805 693
rect 29895 659 30003 693
rect 30093 659 30201 693
rect 30291 659 30399 693
rect 30489 659 30597 693
rect 30687 659 30795 693
rect 30885 659 30993 693
rect 31083 659 31191 693
rect 31281 659 31389 693
rect 31479 659 31587 693
rect 23361 551 23469 585
rect 23559 551 23667 585
rect 23757 551 23865 585
rect 23955 551 24063 585
rect 24153 551 24261 585
rect 24351 551 24459 585
rect 24549 551 24657 585
rect 24747 551 24855 585
rect 24945 551 25053 585
rect 25143 551 25251 585
rect 25341 551 25449 585
rect 25539 551 25647 585
rect 25737 551 25845 585
rect 25935 551 26043 585
rect 26133 551 26241 585
rect 26331 551 26439 585
rect 26529 551 26637 585
rect 26727 551 26835 585
rect 26925 551 27033 585
rect 27123 551 27231 585
rect 27321 551 27429 585
rect 27519 551 27627 585
rect 27717 551 27825 585
rect 27915 551 28023 585
rect 28113 551 28221 585
rect 28311 551 28419 585
rect 28509 551 28617 585
rect 28707 551 28815 585
rect 28905 551 29013 585
rect 29103 551 29211 585
rect 29301 551 29409 585
rect 29499 551 29607 585
rect 29697 551 29805 585
rect 29895 551 30003 585
rect 30093 551 30201 585
rect 30291 551 30399 585
rect 30489 551 30597 585
rect 30687 551 30795 585
rect 30885 551 30993 585
rect 31083 551 31191 585
rect 31281 551 31389 585
rect 31479 551 31587 585
rect 23361 -977 23469 -943
rect 23559 -977 23667 -943
rect 23757 -977 23865 -943
rect 23955 -977 24063 -943
rect 24153 -977 24261 -943
rect 24351 -977 24459 -943
rect 24549 -977 24657 -943
rect 24747 -977 24855 -943
rect 24945 -977 25053 -943
rect 25143 -977 25251 -943
rect 25341 -977 25449 -943
rect 25539 -977 25647 -943
rect 25737 -977 25845 -943
rect 25935 -977 26043 -943
rect 26133 -977 26241 -943
rect 26331 -977 26439 -943
rect 26529 -977 26637 -943
rect 26727 -977 26835 -943
rect 26925 -977 27033 -943
rect 27123 -977 27231 -943
rect 27321 -977 27429 -943
rect 27519 -977 27627 -943
rect 27717 -977 27825 -943
rect 27915 -977 28023 -943
rect 28113 -977 28221 -943
rect 28311 -977 28419 -943
rect 28509 -977 28617 -943
rect 28707 -977 28815 -943
rect 28905 -977 29013 -943
rect 29103 -977 29211 -943
rect 29301 -977 29409 -943
rect 29499 -977 29607 -943
rect 29697 -977 29805 -943
rect 29895 -977 30003 -943
rect 30093 -977 30201 -943
rect 30291 -977 30399 -943
rect 30489 -977 30597 -943
rect 30687 -977 30795 -943
rect 30885 -977 30993 -943
rect 31083 -977 31191 -943
rect 31281 -977 31389 -943
rect 31479 -977 31587 -943
rect 23361 -1085 23469 -1051
rect 23559 -1085 23667 -1051
rect 23757 -1085 23865 -1051
rect 23955 -1085 24063 -1051
rect 24153 -1085 24261 -1051
rect 24351 -1085 24459 -1051
rect 24549 -1085 24657 -1051
rect 24747 -1085 24855 -1051
rect 24945 -1085 25053 -1051
rect 25143 -1085 25251 -1051
rect 25341 -1085 25449 -1051
rect 25539 -1085 25647 -1051
rect 25737 -1085 25845 -1051
rect 25935 -1085 26043 -1051
rect 26133 -1085 26241 -1051
rect 26331 -1085 26439 -1051
rect 26529 -1085 26637 -1051
rect 26727 -1085 26835 -1051
rect 26925 -1085 27033 -1051
rect 27123 -1085 27231 -1051
rect 27321 -1085 27429 -1051
rect 27519 -1085 27627 -1051
rect 27717 -1085 27825 -1051
rect 27915 -1085 28023 -1051
rect 28113 -1085 28221 -1051
rect 28311 -1085 28419 -1051
rect 28509 -1085 28617 -1051
rect 28707 -1085 28815 -1051
rect 28905 -1085 29013 -1051
rect 29103 -1085 29211 -1051
rect 29301 -1085 29409 -1051
rect 29499 -1085 29607 -1051
rect 29697 -1085 29805 -1051
rect 29895 -1085 30003 -1051
rect 30093 -1085 30201 -1051
rect 30291 -1085 30399 -1051
rect 30489 -1085 30597 -1051
rect 30687 -1085 30795 -1051
rect 30885 -1085 30993 -1051
rect 31083 -1085 31191 -1051
rect 31281 -1085 31389 -1051
rect 31479 -1085 31587 -1051
rect 23361 -2613 23469 -2579
rect 23559 -2613 23667 -2579
rect 23757 -2613 23865 -2579
rect 23955 -2613 24063 -2579
rect 24153 -2613 24261 -2579
rect 24351 -2613 24459 -2579
rect 24549 -2613 24657 -2579
rect 24747 -2613 24855 -2579
rect 24945 -2613 25053 -2579
rect 25143 -2613 25251 -2579
rect 25341 -2613 25449 -2579
rect 25539 -2613 25647 -2579
rect 25737 -2613 25845 -2579
rect 25935 -2613 26043 -2579
rect 26133 -2613 26241 -2579
rect 26331 -2613 26439 -2579
rect 26529 -2613 26637 -2579
rect 26727 -2613 26835 -2579
rect 26925 -2613 27033 -2579
rect 27123 -2613 27231 -2579
rect 27321 -2613 27429 -2579
rect 27519 -2613 27627 -2579
rect 27717 -2613 27825 -2579
rect 27915 -2613 28023 -2579
rect 28113 -2613 28221 -2579
rect 28311 -2613 28419 -2579
rect 28509 -2613 28617 -2579
rect 28707 -2613 28815 -2579
rect 28905 -2613 29013 -2579
rect 29103 -2613 29211 -2579
rect 29301 -2613 29409 -2579
rect 29499 -2613 29607 -2579
rect 29697 -2613 29805 -2579
rect 29895 -2613 30003 -2579
rect 30093 -2613 30201 -2579
rect 30291 -2613 30399 -2579
rect 30489 -2613 30597 -2579
rect 30687 -2613 30795 -2579
rect 30885 -2613 30993 -2579
rect 31083 -2613 31191 -2579
rect 31281 -2613 31389 -2579
rect 31479 -2613 31587 -2579
rect 23361 -3286 23469 -3252
rect 23559 -3286 23667 -3252
rect 23757 -3286 23865 -3252
rect 23955 -3286 24063 -3252
rect 24153 -3286 24261 -3252
rect 24351 -3286 24459 -3252
rect 24549 -3286 24657 -3252
rect 24747 -3286 24855 -3252
rect 24945 -3286 25053 -3252
rect 25143 -3286 25251 -3252
rect 25341 -3286 25449 -3252
rect 25539 -3286 25647 -3252
rect 25737 -3286 25845 -3252
rect 25935 -3286 26043 -3252
rect 26133 -3286 26241 -3252
rect 26331 -3286 26439 -3252
rect 26529 -3286 26637 -3252
rect 26727 -3286 26835 -3252
rect 26925 -3286 27033 -3252
rect 27123 -3286 27231 -3252
rect 27321 -3286 27429 -3252
rect 27519 -3286 27627 -3252
rect 27717 -3286 27825 -3252
rect 27915 -3286 28023 -3252
rect 28113 -3286 28221 -3252
rect 28311 -3286 28419 -3252
rect 28509 -3286 28617 -3252
rect 28707 -3286 28815 -3252
rect 28905 -3286 29013 -3252
rect 29103 -3286 29211 -3252
rect 29301 -3286 29409 -3252
rect 29499 -3286 29607 -3252
rect 29697 -3286 29805 -3252
rect 29895 -3286 30003 -3252
rect 30093 -3286 30201 -3252
rect 30291 -3286 30399 -3252
rect 30489 -3286 30597 -3252
rect 30687 -3286 30795 -3252
rect 30885 -3286 30993 -3252
rect 31083 -3286 31191 -3252
rect 31281 -3286 31389 -3252
rect 31479 -3286 31587 -3252
<< locali >>
rect -848 2237 -752 2271
rect 8337 2237 8433 2271
rect -848 2175 -814 2237
rect 8399 2070 8433 2237
rect -814 -3034 -347 -2933
rect 7917 -3034 8399 -2933
rect -848 -5214 -814 -4353
rect 10991 2237 11087 2271
rect 20176 2237 20272 2271
rect 10991 2101 11025 2237
rect 8433 -3034 10991 -2933
rect 8399 -5214 8433 -4458
rect 11449 2128 11483 2144
rect 11449 736 11483 752
rect 11647 2128 11681 2144
rect 11647 736 11681 752
rect 11845 2128 11879 2144
rect 11845 736 11879 752
rect 12043 2128 12077 2144
rect 12043 736 12077 752
rect 12241 2128 12275 2144
rect 12241 736 12275 752
rect 12439 2128 12473 2144
rect 12439 736 12473 752
rect 12637 2128 12671 2144
rect 12637 736 12671 752
rect 12835 2128 12869 2144
rect 12835 736 12869 752
rect 13033 2128 13067 2144
rect 13033 736 13067 752
rect 13231 2128 13265 2144
rect 13231 736 13265 752
rect 13429 2128 13463 2144
rect 13429 736 13463 752
rect 13627 2128 13661 2144
rect 13627 736 13661 752
rect 13825 2128 13859 2144
rect 13825 736 13859 752
rect 14023 2128 14057 2144
rect 14023 736 14057 752
rect 14221 2128 14255 2144
rect 14221 736 14255 752
rect 14419 2128 14453 2144
rect 14419 736 14453 752
rect 14617 2128 14651 2144
rect 14617 736 14651 752
rect 14815 2128 14849 2144
rect 14815 736 14849 752
rect 15013 2128 15047 2144
rect 15013 736 15047 752
rect 15211 2128 15245 2144
rect 15211 736 15245 752
rect 15409 2128 15443 2144
rect 15409 736 15443 752
rect 15607 2128 15641 2144
rect 15607 736 15641 752
rect 15805 2128 15839 2144
rect 15805 736 15839 752
rect 16003 2128 16037 2144
rect 16003 736 16037 752
rect 16201 2128 16235 2144
rect 16201 736 16235 752
rect 16399 2128 16433 2144
rect 16399 736 16433 752
rect 16597 2128 16631 2144
rect 16597 736 16631 752
rect 16795 2128 16829 2144
rect 16795 736 16829 752
rect 16993 2128 17027 2144
rect 16993 736 17027 752
rect 17191 2128 17225 2144
rect 17191 736 17225 752
rect 17389 2128 17423 2144
rect 17389 736 17423 752
rect 17587 2128 17621 2144
rect 17587 736 17621 752
rect 17785 2128 17819 2144
rect 17785 736 17819 752
rect 17983 2128 18017 2144
rect 17983 736 18017 752
rect 18181 2128 18215 2144
rect 18181 736 18215 752
rect 18379 2128 18413 2144
rect 18379 736 18413 752
rect 18577 2128 18611 2144
rect 18577 736 18611 752
rect 18775 2128 18809 2144
rect 18775 736 18809 752
rect 18973 2128 19007 2144
rect 18973 736 19007 752
rect 19171 2128 19205 2144
rect 19171 736 19205 752
rect 19369 2128 19403 2144
rect 19369 736 19403 752
rect 19567 2128 19601 2144
rect 19567 736 19601 752
rect 19765 2128 19799 2144
rect 19765 736 19799 752
rect 20238 2070 20272 2237
rect 11495 659 11511 693
rect 11619 659 11635 693
rect 11693 659 11709 693
rect 11817 659 11833 693
rect 11891 659 11907 693
rect 12015 659 12031 693
rect 12089 659 12105 693
rect 12213 659 12229 693
rect 12287 659 12303 693
rect 12411 659 12427 693
rect 12485 659 12501 693
rect 12609 659 12625 693
rect 12683 659 12699 693
rect 12807 659 12823 693
rect 12881 659 12897 693
rect 13005 659 13021 693
rect 13079 659 13095 693
rect 13203 659 13219 693
rect 13277 659 13293 693
rect 13401 659 13417 693
rect 13475 659 13491 693
rect 13599 659 13615 693
rect 13673 659 13689 693
rect 13797 659 13813 693
rect 13871 659 13887 693
rect 13995 659 14011 693
rect 14069 659 14085 693
rect 14193 659 14209 693
rect 14267 659 14283 693
rect 14391 659 14407 693
rect 14465 659 14481 693
rect 14589 659 14605 693
rect 14663 659 14679 693
rect 14787 659 14803 693
rect 14861 659 14877 693
rect 14985 659 15001 693
rect 15059 659 15075 693
rect 15183 659 15199 693
rect 15257 659 15273 693
rect 15381 659 15397 693
rect 15455 659 15471 693
rect 15579 659 15595 693
rect 15653 659 15669 693
rect 15777 659 15793 693
rect 15851 659 15867 693
rect 15975 659 15991 693
rect 16049 659 16065 693
rect 16173 659 16189 693
rect 16247 659 16263 693
rect 16371 659 16387 693
rect 16445 659 16461 693
rect 16569 659 16585 693
rect 16643 659 16659 693
rect 16767 659 16783 693
rect 16841 659 16857 693
rect 16965 659 16981 693
rect 17039 659 17055 693
rect 17163 659 17179 693
rect 17237 659 17253 693
rect 17361 659 17377 693
rect 17435 659 17451 693
rect 17559 659 17575 693
rect 17633 659 17649 693
rect 17757 659 17773 693
rect 17831 659 17847 693
rect 17955 659 17971 693
rect 18029 659 18045 693
rect 18153 659 18169 693
rect 18227 659 18243 693
rect 18351 659 18367 693
rect 18425 659 18441 693
rect 18549 659 18565 693
rect 18623 659 18639 693
rect 18747 659 18763 693
rect 18821 659 18837 693
rect 18945 659 18961 693
rect 19019 659 19035 693
rect 19143 659 19159 693
rect 19217 659 19233 693
rect 19341 659 19357 693
rect 19415 659 19431 693
rect 19539 659 19555 693
rect 19613 659 19629 693
rect 19737 659 19753 693
rect 11495 551 11511 585
rect 11619 551 11635 585
rect 11693 551 11709 585
rect 11817 551 11833 585
rect 11891 551 11907 585
rect 12015 551 12031 585
rect 12089 551 12105 585
rect 12213 551 12229 585
rect 12287 551 12303 585
rect 12411 551 12427 585
rect 12485 551 12501 585
rect 12609 551 12625 585
rect 12683 551 12699 585
rect 12807 551 12823 585
rect 12881 551 12897 585
rect 13005 551 13021 585
rect 13079 551 13095 585
rect 13203 551 13219 585
rect 13277 551 13293 585
rect 13401 551 13417 585
rect 13475 551 13491 585
rect 13599 551 13615 585
rect 13673 551 13689 585
rect 13797 551 13813 585
rect 13871 551 13887 585
rect 13995 551 14011 585
rect 14069 551 14085 585
rect 14193 551 14209 585
rect 14267 551 14283 585
rect 14391 551 14407 585
rect 14465 551 14481 585
rect 14589 551 14605 585
rect 14663 551 14679 585
rect 14787 551 14803 585
rect 14861 551 14877 585
rect 14985 551 15001 585
rect 15059 551 15075 585
rect 15183 551 15199 585
rect 15257 551 15273 585
rect 15381 551 15397 585
rect 15455 551 15471 585
rect 15579 551 15595 585
rect 15653 551 15669 585
rect 15777 551 15793 585
rect 15851 551 15867 585
rect 15975 551 15991 585
rect 16049 551 16065 585
rect 16173 551 16189 585
rect 16247 551 16263 585
rect 16371 551 16387 585
rect 16445 551 16461 585
rect 16569 551 16585 585
rect 16643 551 16659 585
rect 16767 551 16783 585
rect 16841 551 16857 585
rect 16965 551 16981 585
rect 17039 551 17055 585
rect 17163 551 17179 585
rect 17237 551 17253 585
rect 17361 551 17377 585
rect 17435 551 17451 585
rect 17559 551 17575 585
rect 17633 551 17649 585
rect 17757 551 17773 585
rect 17831 551 17847 585
rect 17955 551 17971 585
rect 18029 551 18045 585
rect 18153 551 18169 585
rect 18227 551 18243 585
rect 18351 551 18367 585
rect 18425 551 18441 585
rect 18549 551 18565 585
rect 18623 551 18639 585
rect 18747 551 18763 585
rect 18821 551 18837 585
rect 18945 551 18961 585
rect 19019 551 19035 585
rect 19143 551 19159 585
rect 19217 551 19233 585
rect 19341 551 19357 585
rect 19415 551 19431 585
rect 19539 551 19555 585
rect 19613 551 19629 585
rect 19737 551 19753 585
rect 11449 492 11483 508
rect 11449 -900 11483 -884
rect 11647 492 11681 508
rect 11647 -900 11681 -884
rect 11845 492 11879 508
rect 11845 -900 11879 -884
rect 12043 492 12077 508
rect 12043 -900 12077 -884
rect 12241 492 12275 508
rect 12241 -900 12275 -884
rect 12439 492 12473 508
rect 12439 -900 12473 -884
rect 12637 492 12671 508
rect 12637 -900 12671 -884
rect 12835 492 12869 508
rect 12835 -900 12869 -884
rect 13033 492 13067 508
rect 13033 -900 13067 -884
rect 13231 492 13265 508
rect 13231 -900 13265 -884
rect 13429 492 13463 508
rect 13429 -900 13463 -884
rect 13627 492 13661 508
rect 13627 -900 13661 -884
rect 13825 492 13859 508
rect 13825 -900 13859 -884
rect 14023 492 14057 508
rect 14023 -900 14057 -884
rect 14221 492 14255 508
rect 14221 -900 14255 -884
rect 14419 492 14453 508
rect 14419 -900 14453 -884
rect 14617 492 14651 508
rect 14617 -900 14651 -884
rect 14815 492 14849 508
rect 14815 -900 14849 -884
rect 15013 492 15047 508
rect 15013 -900 15047 -884
rect 15211 492 15245 508
rect 15211 -900 15245 -884
rect 15409 492 15443 508
rect 15409 -900 15443 -884
rect 15607 492 15641 508
rect 15607 -900 15641 -884
rect 15805 492 15839 508
rect 15805 -900 15839 -884
rect 16003 492 16037 508
rect 16003 -900 16037 -884
rect 16201 492 16235 508
rect 16201 -900 16235 -884
rect 16399 492 16433 508
rect 16399 -900 16433 -884
rect 16597 492 16631 508
rect 16597 -900 16631 -884
rect 16795 492 16829 508
rect 16795 -900 16829 -884
rect 16993 492 17027 508
rect 16993 -900 17027 -884
rect 17191 492 17225 508
rect 17191 -900 17225 -884
rect 17389 492 17423 508
rect 17389 -900 17423 -884
rect 17587 492 17621 508
rect 17587 -900 17621 -884
rect 17785 492 17819 508
rect 17785 -900 17819 -884
rect 17983 492 18017 508
rect 17983 -900 18017 -884
rect 18181 492 18215 508
rect 18181 -900 18215 -884
rect 18379 492 18413 508
rect 18379 -900 18413 -884
rect 18577 492 18611 508
rect 18577 -900 18611 -884
rect 18775 492 18809 508
rect 18775 -900 18809 -884
rect 18973 492 19007 508
rect 18973 -900 19007 -884
rect 19171 492 19205 508
rect 19171 -900 19205 -884
rect 19369 492 19403 508
rect 19369 -900 19403 -884
rect 19567 492 19601 508
rect 19567 -900 19601 -884
rect 19765 492 19799 508
rect 19765 -900 19799 -884
rect 11495 -977 11511 -943
rect 11619 -977 11635 -943
rect 11693 -977 11709 -943
rect 11817 -977 11833 -943
rect 11891 -977 11907 -943
rect 12015 -977 12031 -943
rect 12089 -977 12105 -943
rect 12213 -977 12229 -943
rect 12287 -977 12303 -943
rect 12411 -977 12427 -943
rect 12485 -977 12501 -943
rect 12609 -977 12625 -943
rect 12683 -977 12699 -943
rect 12807 -977 12823 -943
rect 12881 -977 12897 -943
rect 13005 -977 13021 -943
rect 13079 -977 13095 -943
rect 13203 -977 13219 -943
rect 13277 -977 13293 -943
rect 13401 -977 13417 -943
rect 13475 -977 13491 -943
rect 13599 -977 13615 -943
rect 13673 -977 13689 -943
rect 13797 -977 13813 -943
rect 13871 -977 13887 -943
rect 13995 -977 14011 -943
rect 14069 -977 14085 -943
rect 14193 -977 14209 -943
rect 14267 -977 14283 -943
rect 14391 -977 14407 -943
rect 14465 -977 14481 -943
rect 14589 -977 14605 -943
rect 14663 -977 14679 -943
rect 14787 -977 14803 -943
rect 14861 -977 14877 -943
rect 14985 -977 15001 -943
rect 15059 -977 15075 -943
rect 15183 -977 15199 -943
rect 15257 -977 15273 -943
rect 15381 -977 15397 -943
rect 15455 -977 15471 -943
rect 15579 -977 15595 -943
rect 15653 -977 15669 -943
rect 15777 -977 15793 -943
rect 15851 -977 15867 -943
rect 15975 -977 15991 -943
rect 16049 -977 16065 -943
rect 16173 -977 16189 -943
rect 16247 -977 16263 -943
rect 16371 -977 16387 -943
rect 16445 -977 16461 -943
rect 16569 -977 16585 -943
rect 16643 -977 16659 -943
rect 16767 -977 16783 -943
rect 16841 -977 16857 -943
rect 16965 -977 16981 -943
rect 17039 -977 17055 -943
rect 17163 -977 17179 -943
rect 17237 -977 17253 -943
rect 17361 -977 17377 -943
rect 17435 -977 17451 -943
rect 17559 -977 17575 -943
rect 17633 -977 17649 -943
rect 17757 -977 17773 -943
rect 17831 -977 17847 -943
rect 17955 -977 17971 -943
rect 18029 -977 18045 -943
rect 18153 -977 18169 -943
rect 18227 -977 18243 -943
rect 18351 -977 18367 -943
rect 18425 -977 18441 -943
rect 18549 -977 18565 -943
rect 18623 -977 18639 -943
rect 18747 -977 18763 -943
rect 18821 -977 18837 -943
rect 18945 -977 18961 -943
rect 19019 -977 19035 -943
rect 19143 -977 19159 -943
rect 19217 -977 19233 -943
rect 19341 -977 19357 -943
rect 19415 -977 19431 -943
rect 19539 -977 19555 -943
rect 19613 -977 19629 -943
rect 19737 -977 19753 -943
rect 11495 -1085 11511 -1051
rect 11619 -1085 11635 -1051
rect 11693 -1085 11709 -1051
rect 11817 -1085 11833 -1051
rect 11891 -1085 11907 -1051
rect 12015 -1085 12031 -1051
rect 12089 -1085 12105 -1051
rect 12213 -1085 12229 -1051
rect 12287 -1085 12303 -1051
rect 12411 -1085 12427 -1051
rect 12485 -1085 12501 -1051
rect 12609 -1085 12625 -1051
rect 12683 -1085 12699 -1051
rect 12807 -1085 12823 -1051
rect 12881 -1085 12897 -1051
rect 13005 -1085 13021 -1051
rect 13079 -1085 13095 -1051
rect 13203 -1085 13219 -1051
rect 13277 -1085 13293 -1051
rect 13401 -1085 13417 -1051
rect 13475 -1085 13491 -1051
rect 13599 -1085 13615 -1051
rect 13673 -1085 13689 -1051
rect 13797 -1085 13813 -1051
rect 13871 -1085 13887 -1051
rect 13995 -1085 14011 -1051
rect 14069 -1085 14085 -1051
rect 14193 -1085 14209 -1051
rect 14267 -1085 14283 -1051
rect 14391 -1085 14407 -1051
rect 14465 -1085 14481 -1051
rect 14589 -1085 14605 -1051
rect 14663 -1085 14679 -1051
rect 14787 -1085 14803 -1051
rect 14861 -1085 14877 -1051
rect 14985 -1085 15001 -1051
rect 15059 -1085 15075 -1051
rect 15183 -1085 15199 -1051
rect 15257 -1085 15273 -1051
rect 15381 -1085 15397 -1051
rect 15455 -1085 15471 -1051
rect 15579 -1085 15595 -1051
rect 15653 -1085 15669 -1051
rect 15777 -1085 15793 -1051
rect 15851 -1085 15867 -1051
rect 15975 -1085 15991 -1051
rect 16049 -1085 16065 -1051
rect 16173 -1085 16189 -1051
rect 16247 -1085 16263 -1051
rect 16371 -1085 16387 -1051
rect 16445 -1085 16461 -1051
rect 16569 -1085 16585 -1051
rect 16643 -1085 16659 -1051
rect 16767 -1085 16783 -1051
rect 16841 -1085 16857 -1051
rect 16965 -1085 16981 -1051
rect 17039 -1085 17055 -1051
rect 17163 -1085 17179 -1051
rect 17237 -1085 17253 -1051
rect 17361 -1085 17377 -1051
rect 17435 -1085 17451 -1051
rect 17559 -1085 17575 -1051
rect 17633 -1085 17649 -1051
rect 17757 -1085 17773 -1051
rect 17831 -1085 17847 -1051
rect 17955 -1085 17971 -1051
rect 18029 -1085 18045 -1051
rect 18153 -1085 18169 -1051
rect 18227 -1085 18243 -1051
rect 18351 -1085 18367 -1051
rect 18425 -1085 18441 -1051
rect 18549 -1085 18565 -1051
rect 18623 -1085 18639 -1051
rect 18747 -1085 18763 -1051
rect 18821 -1085 18837 -1051
rect 18945 -1085 18961 -1051
rect 19019 -1085 19035 -1051
rect 19143 -1085 19159 -1051
rect 19217 -1085 19233 -1051
rect 19341 -1085 19357 -1051
rect 19415 -1085 19431 -1051
rect 19539 -1085 19555 -1051
rect 19613 -1085 19629 -1051
rect 19737 -1085 19753 -1051
rect 11449 -1144 11483 -1128
rect 11449 -2536 11483 -2520
rect 11647 -1144 11681 -1128
rect 11647 -2536 11681 -2520
rect 11845 -1144 11879 -1128
rect 11845 -2536 11879 -2520
rect 12043 -1144 12077 -1128
rect 12043 -2536 12077 -2520
rect 12241 -1144 12275 -1128
rect 12241 -2536 12275 -2520
rect 12439 -1144 12473 -1128
rect 12439 -2536 12473 -2520
rect 12637 -1144 12671 -1128
rect 12637 -2536 12671 -2520
rect 12835 -1144 12869 -1128
rect 12835 -2536 12869 -2520
rect 13033 -1144 13067 -1128
rect 13033 -2536 13067 -2520
rect 13231 -1144 13265 -1128
rect 13231 -2536 13265 -2520
rect 13429 -1144 13463 -1128
rect 13429 -2536 13463 -2520
rect 13627 -1144 13661 -1128
rect 13627 -2536 13661 -2520
rect 13825 -1144 13859 -1128
rect 13825 -2536 13859 -2520
rect 14023 -1144 14057 -1128
rect 14023 -2536 14057 -2520
rect 14221 -1144 14255 -1128
rect 14221 -2536 14255 -2520
rect 14419 -1144 14453 -1128
rect 14419 -2536 14453 -2520
rect 14617 -1144 14651 -1128
rect 14617 -2536 14651 -2520
rect 14815 -1144 14849 -1128
rect 14815 -2536 14849 -2520
rect 15013 -1144 15047 -1128
rect 15013 -2536 15047 -2520
rect 15211 -1144 15245 -1128
rect 15211 -2536 15245 -2520
rect 15409 -1144 15443 -1128
rect 15409 -2536 15443 -2520
rect 15607 -1144 15641 -1128
rect 15607 -2536 15641 -2520
rect 15805 -1144 15839 -1128
rect 15805 -2536 15839 -2520
rect 16003 -1144 16037 -1128
rect 16003 -2536 16037 -2520
rect 16201 -1144 16235 -1128
rect 16201 -2536 16235 -2520
rect 16399 -1144 16433 -1128
rect 16399 -2536 16433 -2520
rect 16597 -1144 16631 -1128
rect 16597 -2536 16631 -2520
rect 16795 -1144 16829 -1128
rect 16795 -2536 16829 -2520
rect 16993 -1144 17027 -1128
rect 16993 -2536 17027 -2520
rect 17191 -1144 17225 -1128
rect 17191 -2536 17225 -2520
rect 17389 -1144 17423 -1128
rect 17389 -2536 17423 -2520
rect 17587 -1144 17621 -1128
rect 17587 -2536 17621 -2520
rect 17785 -1144 17819 -1128
rect 17785 -2536 17819 -2520
rect 17983 -1144 18017 -1128
rect 17983 -2536 18017 -2520
rect 18181 -1144 18215 -1128
rect 18181 -2536 18215 -2520
rect 18379 -1144 18413 -1128
rect 18379 -2536 18413 -2520
rect 18577 -1144 18611 -1128
rect 18577 -2536 18611 -2520
rect 18775 -1144 18809 -1128
rect 18775 -2536 18809 -2520
rect 18973 -1144 19007 -1128
rect 18973 -2536 19007 -2520
rect 19171 -1144 19205 -1128
rect 19171 -2536 19205 -2520
rect 19369 -1144 19403 -1128
rect 19369 -2536 19403 -2520
rect 19567 -1144 19601 -1128
rect 19567 -2536 19601 -2520
rect 19765 -1144 19799 -1128
rect 19765 -2536 19799 -2520
rect 11495 -2613 11511 -2579
rect 11619 -2613 11635 -2579
rect 11693 -2613 11709 -2579
rect 11817 -2613 11833 -2579
rect 11891 -2613 11907 -2579
rect 12015 -2613 12031 -2579
rect 12089 -2613 12105 -2579
rect 12213 -2613 12229 -2579
rect 12287 -2613 12303 -2579
rect 12411 -2613 12427 -2579
rect 12485 -2613 12501 -2579
rect 12609 -2613 12625 -2579
rect 12683 -2613 12699 -2579
rect 12807 -2613 12823 -2579
rect 12881 -2613 12897 -2579
rect 13005 -2613 13021 -2579
rect 13079 -2613 13095 -2579
rect 13203 -2613 13219 -2579
rect 13277 -2613 13293 -2579
rect 13401 -2613 13417 -2579
rect 13475 -2613 13491 -2579
rect 13599 -2613 13615 -2579
rect 13673 -2613 13689 -2579
rect 13797 -2613 13813 -2579
rect 13871 -2613 13887 -2579
rect 13995 -2613 14011 -2579
rect 14069 -2613 14085 -2579
rect 14193 -2613 14209 -2579
rect 14267 -2613 14283 -2579
rect 14391 -2613 14407 -2579
rect 14465 -2613 14481 -2579
rect 14589 -2613 14605 -2579
rect 14663 -2613 14679 -2579
rect 14787 -2613 14803 -2579
rect 14861 -2613 14877 -2579
rect 14985 -2613 15001 -2579
rect 15059 -2613 15075 -2579
rect 15183 -2613 15199 -2579
rect 15257 -2613 15273 -2579
rect 15381 -2613 15397 -2579
rect 15455 -2613 15471 -2579
rect 15579 -2613 15595 -2579
rect 15653 -2613 15669 -2579
rect 15777 -2613 15793 -2579
rect 15851 -2613 15867 -2579
rect 15975 -2613 15991 -2579
rect 16049 -2613 16065 -2579
rect 16173 -2613 16189 -2579
rect 16247 -2613 16263 -2579
rect 16371 -2613 16387 -2579
rect 16445 -2613 16461 -2579
rect 16569 -2613 16585 -2579
rect 16643 -2613 16659 -2579
rect 16767 -2613 16783 -2579
rect 16841 -2613 16857 -2579
rect 16965 -2613 16981 -2579
rect 17039 -2613 17055 -2579
rect 17163 -2613 17179 -2579
rect 17237 -2613 17253 -2579
rect 17361 -2613 17377 -2579
rect 17435 -2613 17451 -2579
rect 17559 -2613 17575 -2579
rect 17633 -2613 17649 -2579
rect 17757 -2613 17773 -2579
rect 17831 -2613 17847 -2579
rect 17955 -2613 17971 -2579
rect 18029 -2613 18045 -2579
rect 18153 -2613 18169 -2579
rect 18227 -2613 18243 -2579
rect 18351 -2613 18367 -2579
rect 18425 -2613 18441 -2579
rect 18549 -2613 18565 -2579
rect 18623 -2613 18639 -2579
rect 18747 -2613 18763 -2579
rect 18821 -2613 18837 -2579
rect 18945 -2613 18961 -2579
rect 19019 -2613 19035 -2579
rect 19143 -2613 19159 -2579
rect 19217 -2613 19233 -2579
rect 19341 -2613 19357 -2579
rect 19415 -2613 19431 -2579
rect 19539 -2613 19555 -2579
rect 19613 -2613 19629 -2579
rect 19737 -2613 19753 -2579
rect 11025 -3034 11492 -2933
rect 19756 -3034 20238 -2933
rect 11495 -3286 11511 -3252
rect 11619 -3286 11635 -3252
rect 11693 -3286 11709 -3252
rect 11817 -3286 11833 -3252
rect 11891 -3286 11907 -3252
rect 12015 -3286 12031 -3252
rect 12089 -3286 12105 -3252
rect 12213 -3286 12229 -3252
rect 12287 -3286 12303 -3252
rect 12411 -3286 12427 -3252
rect 12485 -3286 12501 -3252
rect 12609 -3286 12625 -3252
rect 12683 -3286 12699 -3252
rect 12807 -3286 12823 -3252
rect 12881 -3286 12897 -3252
rect 13005 -3286 13021 -3252
rect 13079 -3286 13095 -3252
rect 13203 -3286 13219 -3252
rect 13277 -3286 13293 -3252
rect 13401 -3286 13417 -3252
rect 13475 -3286 13491 -3252
rect 13599 -3286 13615 -3252
rect 13673 -3286 13689 -3252
rect 13797 -3286 13813 -3252
rect 13871 -3286 13887 -3252
rect 13995 -3286 14011 -3252
rect 14069 -3286 14085 -3252
rect 14193 -3286 14209 -3252
rect 14267 -3286 14283 -3252
rect 14391 -3286 14407 -3252
rect 14465 -3286 14481 -3252
rect 14589 -3286 14605 -3252
rect 14663 -3286 14679 -3252
rect 14787 -3286 14803 -3252
rect 14861 -3286 14877 -3252
rect 14985 -3286 15001 -3252
rect 15059 -3286 15075 -3252
rect 15183 -3286 15199 -3252
rect 15257 -3286 15273 -3252
rect 15381 -3286 15397 -3252
rect 15455 -3286 15471 -3252
rect 15579 -3286 15595 -3252
rect 15653 -3286 15669 -3252
rect 15777 -3286 15793 -3252
rect 15851 -3286 15867 -3252
rect 15975 -3286 15991 -3252
rect 16049 -3286 16065 -3252
rect 16173 -3286 16189 -3252
rect 16247 -3286 16263 -3252
rect 16371 -3286 16387 -3252
rect 16445 -3286 16461 -3252
rect 16569 -3286 16585 -3252
rect 16643 -3286 16659 -3252
rect 16767 -3286 16783 -3252
rect 16841 -3286 16857 -3252
rect 16965 -3286 16981 -3252
rect 17039 -3286 17055 -3252
rect 17163 -3286 17179 -3252
rect 17237 -3286 17253 -3252
rect 17361 -3286 17377 -3252
rect 17435 -3286 17451 -3252
rect 17559 -3286 17575 -3252
rect 17633 -3286 17649 -3252
rect 17757 -3286 17773 -3252
rect 17831 -3286 17847 -3252
rect 17955 -3286 17971 -3252
rect 18029 -3286 18045 -3252
rect 18153 -3286 18169 -3252
rect 18227 -3286 18243 -3252
rect 18351 -3286 18367 -3252
rect 18425 -3286 18441 -3252
rect 18549 -3286 18565 -3252
rect 18623 -3286 18639 -3252
rect 18747 -3286 18763 -3252
rect 18821 -3286 18837 -3252
rect 18945 -3286 18961 -3252
rect 19019 -3286 19035 -3252
rect 19143 -3286 19159 -3252
rect 19217 -3286 19233 -3252
rect 19341 -3286 19357 -3252
rect 19415 -3286 19431 -3252
rect 19539 -3286 19555 -3252
rect 19613 -3286 19629 -3252
rect 19737 -3286 19753 -3252
rect 10991 -5214 11025 -4427
rect 11449 -3345 11483 -3329
rect 11449 -4737 11483 -4721
rect 11647 -3345 11681 -3329
rect 11647 -4737 11681 -4721
rect 11845 -3345 11879 -3329
rect 11845 -4737 11879 -4721
rect 12043 -3345 12077 -3329
rect 12043 -4737 12077 -4721
rect 12241 -3345 12275 -3329
rect 12241 -4737 12275 -4721
rect 12439 -3345 12473 -3329
rect 12439 -4737 12473 -4721
rect 12637 -3345 12671 -3329
rect 12637 -4737 12671 -4721
rect 12835 -3345 12869 -3329
rect 12835 -4737 12869 -4721
rect 13033 -3345 13067 -3329
rect 13033 -4737 13067 -4721
rect 13231 -3345 13265 -3329
rect 13231 -4737 13265 -4721
rect 13429 -3345 13463 -3329
rect 13429 -4737 13463 -4721
rect 13627 -3345 13661 -3329
rect 13627 -4737 13661 -4721
rect 13825 -3345 13859 -3329
rect 13825 -4737 13859 -4721
rect 14023 -3345 14057 -3329
rect 14023 -4737 14057 -4721
rect 14221 -3345 14255 -3329
rect 14221 -4737 14255 -4721
rect 14419 -3345 14453 -3329
rect 14419 -4737 14453 -4721
rect 14617 -3345 14651 -3329
rect 14617 -4737 14651 -4721
rect 14815 -3345 14849 -3329
rect 14815 -4737 14849 -4721
rect 15013 -3345 15047 -3329
rect 15013 -4737 15047 -4721
rect 15211 -3345 15245 -3329
rect 15211 -4737 15245 -4721
rect 15409 -3345 15443 -3329
rect 15409 -4737 15443 -4721
rect 15607 -3345 15641 -3329
rect 15607 -4737 15641 -4721
rect 15805 -3345 15839 -3329
rect 15805 -4737 15839 -4721
rect 16003 -3345 16037 -3329
rect 16003 -4737 16037 -4721
rect 16201 -3345 16235 -3329
rect 16201 -4737 16235 -4721
rect 16399 -3345 16433 -3329
rect 16399 -4737 16433 -4721
rect 16597 -3345 16631 -3329
rect 16597 -4737 16631 -4721
rect 16795 -3345 16829 -3329
rect 16795 -4737 16829 -4721
rect 16993 -3345 17027 -3329
rect 16993 -4737 17027 -4721
rect 17191 -3345 17225 -3329
rect 17191 -4737 17225 -4721
rect 17389 -3345 17423 -3329
rect 17389 -4737 17423 -4721
rect 17587 -3345 17621 -3329
rect 17587 -4737 17621 -4721
rect 17785 -3345 17819 -3329
rect 17785 -4737 17819 -4721
rect 17983 -3345 18017 -3329
rect 17983 -4737 18017 -4721
rect 18181 -3345 18215 -3329
rect 18181 -4737 18215 -4721
rect 18379 -3345 18413 -3329
rect 18379 -4737 18413 -4721
rect 18577 -3345 18611 -3329
rect 18577 -4737 18611 -4721
rect 18775 -3345 18809 -3329
rect 18775 -4737 18809 -4721
rect 18973 -3345 19007 -3329
rect 18973 -4737 19007 -4721
rect 19171 -3345 19205 -3329
rect 19171 -4737 19205 -4721
rect 19369 -3345 19403 -3329
rect 19369 -4737 19403 -4721
rect 19567 -3345 19601 -3329
rect 19567 -4737 19601 -4721
rect 19765 -3345 19799 -3329
rect 19765 -4737 19799 -4721
rect 22830 2237 22937 2271
rect 32026 2237 32122 2271
rect 22830 2101 22864 2237
rect 20272 -3034 22830 -2933
rect 20238 -5214 20272 -4458
rect 23299 2128 23333 2144
rect 23299 736 23333 752
rect 23497 2128 23531 2144
rect 23497 736 23531 752
rect 23695 2128 23729 2144
rect 23695 736 23729 752
rect 23893 2128 23927 2144
rect 23893 736 23927 752
rect 24091 2128 24125 2144
rect 24091 736 24125 752
rect 24289 2128 24323 2144
rect 24289 736 24323 752
rect 24487 2128 24521 2144
rect 24487 736 24521 752
rect 24685 2128 24719 2144
rect 24685 736 24719 752
rect 24883 2128 24917 2144
rect 24883 736 24917 752
rect 25081 2128 25115 2144
rect 25081 736 25115 752
rect 25279 2128 25313 2144
rect 25279 736 25313 752
rect 25477 2128 25511 2144
rect 25477 736 25511 752
rect 25675 2128 25709 2144
rect 25675 736 25709 752
rect 25873 2128 25907 2144
rect 25873 736 25907 752
rect 26071 2128 26105 2144
rect 26071 736 26105 752
rect 26269 2128 26303 2144
rect 26269 736 26303 752
rect 26467 2128 26501 2144
rect 26467 736 26501 752
rect 26665 2128 26699 2144
rect 26665 736 26699 752
rect 26863 2128 26897 2144
rect 26863 736 26897 752
rect 27061 2128 27095 2144
rect 27061 736 27095 752
rect 27259 2128 27293 2144
rect 27259 736 27293 752
rect 27457 2128 27491 2144
rect 27457 736 27491 752
rect 27655 2128 27689 2144
rect 27655 736 27689 752
rect 27853 2128 27887 2144
rect 27853 736 27887 752
rect 28051 2128 28085 2144
rect 28051 736 28085 752
rect 28249 2128 28283 2144
rect 28249 736 28283 752
rect 28447 2128 28481 2144
rect 28447 736 28481 752
rect 28645 2128 28679 2144
rect 28645 736 28679 752
rect 28843 2128 28877 2144
rect 28843 736 28877 752
rect 29041 2128 29075 2144
rect 29041 736 29075 752
rect 29239 2128 29273 2144
rect 29239 736 29273 752
rect 29437 2128 29471 2144
rect 29437 736 29471 752
rect 29635 2128 29669 2144
rect 29635 736 29669 752
rect 29833 2128 29867 2144
rect 29833 736 29867 752
rect 30031 2128 30065 2144
rect 30031 736 30065 752
rect 30229 2128 30263 2144
rect 30229 736 30263 752
rect 30427 2128 30461 2144
rect 30427 736 30461 752
rect 30625 2128 30659 2144
rect 30625 736 30659 752
rect 30823 2128 30857 2144
rect 30823 736 30857 752
rect 31021 2128 31055 2144
rect 31021 736 31055 752
rect 31219 2128 31253 2144
rect 31219 736 31253 752
rect 31417 2128 31451 2144
rect 31417 736 31451 752
rect 31615 2128 31649 2144
rect 31615 736 31649 752
rect 32088 1912 32122 2237
rect 23345 659 23361 693
rect 23469 659 23485 693
rect 23543 659 23559 693
rect 23667 659 23683 693
rect 23741 659 23757 693
rect 23865 659 23881 693
rect 23939 659 23955 693
rect 24063 659 24079 693
rect 24137 659 24153 693
rect 24261 659 24277 693
rect 24335 659 24351 693
rect 24459 659 24475 693
rect 24533 659 24549 693
rect 24657 659 24673 693
rect 24731 659 24747 693
rect 24855 659 24871 693
rect 24929 659 24945 693
rect 25053 659 25069 693
rect 25127 659 25143 693
rect 25251 659 25267 693
rect 25325 659 25341 693
rect 25449 659 25465 693
rect 25523 659 25539 693
rect 25647 659 25663 693
rect 25721 659 25737 693
rect 25845 659 25861 693
rect 25919 659 25935 693
rect 26043 659 26059 693
rect 26117 659 26133 693
rect 26241 659 26257 693
rect 26315 659 26331 693
rect 26439 659 26455 693
rect 26513 659 26529 693
rect 26637 659 26653 693
rect 26711 659 26727 693
rect 26835 659 26851 693
rect 26909 659 26925 693
rect 27033 659 27049 693
rect 27107 659 27123 693
rect 27231 659 27247 693
rect 27305 659 27321 693
rect 27429 659 27445 693
rect 27503 659 27519 693
rect 27627 659 27643 693
rect 27701 659 27717 693
rect 27825 659 27841 693
rect 27899 659 27915 693
rect 28023 659 28039 693
rect 28097 659 28113 693
rect 28221 659 28237 693
rect 28295 659 28311 693
rect 28419 659 28435 693
rect 28493 659 28509 693
rect 28617 659 28633 693
rect 28691 659 28707 693
rect 28815 659 28831 693
rect 28889 659 28905 693
rect 29013 659 29029 693
rect 29087 659 29103 693
rect 29211 659 29227 693
rect 29285 659 29301 693
rect 29409 659 29425 693
rect 29483 659 29499 693
rect 29607 659 29623 693
rect 29681 659 29697 693
rect 29805 659 29821 693
rect 29879 659 29895 693
rect 30003 659 30019 693
rect 30077 659 30093 693
rect 30201 659 30217 693
rect 30275 659 30291 693
rect 30399 659 30415 693
rect 30473 659 30489 693
rect 30597 659 30613 693
rect 30671 659 30687 693
rect 30795 659 30811 693
rect 30869 659 30885 693
rect 30993 659 31009 693
rect 31067 659 31083 693
rect 31191 659 31207 693
rect 31265 659 31281 693
rect 31389 659 31405 693
rect 31463 659 31479 693
rect 31587 659 31603 693
rect 23345 551 23361 585
rect 23469 551 23485 585
rect 23543 551 23559 585
rect 23667 551 23683 585
rect 23741 551 23757 585
rect 23865 551 23881 585
rect 23939 551 23955 585
rect 24063 551 24079 585
rect 24137 551 24153 585
rect 24261 551 24277 585
rect 24335 551 24351 585
rect 24459 551 24475 585
rect 24533 551 24549 585
rect 24657 551 24673 585
rect 24731 551 24747 585
rect 24855 551 24871 585
rect 24929 551 24945 585
rect 25053 551 25069 585
rect 25127 551 25143 585
rect 25251 551 25267 585
rect 25325 551 25341 585
rect 25449 551 25465 585
rect 25523 551 25539 585
rect 25647 551 25663 585
rect 25721 551 25737 585
rect 25845 551 25861 585
rect 25919 551 25935 585
rect 26043 551 26059 585
rect 26117 551 26133 585
rect 26241 551 26257 585
rect 26315 551 26331 585
rect 26439 551 26455 585
rect 26513 551 26529 585
rect 26637 551 26653 585
rect 26711 551 26727 585
rect 26835 551 26851 585
rect 26909 551 26925 585
rect 27033 551 27049 585
rect 27107 551 27123 585
rect 27231 551 27247 585
rect 27305 551 27321 585
rect 27429 551 27445 585
rect 27503 551 27519 585
rect 27627 551 27643 585
rect 27701 551 27717 585
rect 27825 551 27841 585
rect 27899 551 27915 585
rect 28023 551 28039 585
rect 28097 551 28113 585
rect 28221 551 28237 585
rect 28295 551 28311 585
rect 28419 551 28435 585
rect 28493 551 28509 585
rect 28617 551 28633 585
rect 28691 551 28707 585
rect 28815 551 28831 585
rect 28889 551 28905 585
rect 29013 551 29029 585
rect 29087 551 29103 585
rect 29211 551 29227 585
rect 29285 551 29301 585
rect 29409 551 29425 585
rect 29483 551 29499 585
rect 29607 551 29623 585
rect 29681 551 29697 585
rect 29805 551 29821 585
rect 29879 551 29895 585
rect 30003 551 30019 585
rect 30077 551 30093 585
rect 30201 551 30217 585
rect 30275 551 30291 585
rect 30399 551 30415 585
rect 30473 551 30489 585
rect 30597 551 30613 585
rect 30671 551 30687 585
rect 30795 551 30811 585
rect 30869 551 30885 585
rect 30993 551 31009 585
rect 31067 551 31083 585
rect 31191 551 31207 585
rect 31265 551 31281 585
rect 31389 551 31405 585
rect 31463 551 31479 585
rect 31587 551 31603 585
rect 23299 492 23333 508
rect 23299 -900 23333 -884
rect 23497 492 23531 508
rect 23497 -900 23531 -884
rect 23695 492 23729 508
rect 23695 -900 23729 -884
rect 23893 492 23927 508
rect 23893 -900 23927 -884
rect 24091 492 24125 508
rect 24091 -900 24125 -884
rect 24289 492 24323 508
rect 24289 -900 24323 -884
rect 24487 492 24521 508
rect 24487 -900 24521 -884
rect 24685 492 24719 508
rect 24685 -900 24719 -884
rect 24883 492 24917 508
rect 24883 -900 24917 -884
rect 25081 492 25115 508
rect 25081 -900 25115 -884
rect 25279 492 25313 508
rect 25279 -900 25313 -884
rect 25477 492 25511 508
rect 25477 -900 25511 -884
rect 25675 492 25709 508
rect 25675 -900 25709 -884
rect 25873 492 25907 508
rect 25873 -900 25907 -884
rect 26071 492 26105 508
rect 26071 -900 26105 -884
rect 26269 492 26303 508
rect 26269 -900 26303 -884
rect 26467 492 26501 508
rect 26467 -900 26501 -884
rect 26665 492 26699 508
rect 26665 -900 26699 -884
rect 26863 492 26897 508
rect 26863 -900 26897 -884
rect 27061 492 27095 508
rect 27061 -900 27095 -884
rect 27259 492 27293 508
rect 27259 -900 27293 -884
rect 27457 492 27491 508
rect 27457 -900 27491 -884
rect 27655 492 27689 508
rect 27655 -900 27689 -884
rect 27853 492 27887 508
rect 27853 -900 27887 -884
rect 28051 492 28085 508
rect 28051 -900 28085 -884
rect 28249 492 28283 508
rect 28249 -900 28283 -884
rect 28447 492 28481 508
rect 28447 -900 28481 -884
rect 28645 492 28679 508
rect 28645 -900 28679 -884
rect 28843 492 28877 508
rect 28843 -900 28877 -884
rect 29041 492 29075 508
rect 29041 -900 29075 -884
rect 29239 492 29273 508
rect 29239 -900 29273 -884
rect 29437 492 29471 508
rect 29437 -900 29471 -884
rect 29635 492 29669 508
rect 29635 -900 29669 -884
rect 29833 492 29867 508
rect 29833 -900 29867 -884
rect 30031 492 30065 508
rect 30031 -900 30065 -884
rect 30229 492 30263 508
rect 30229 -900 30263 -884
rect 30427 492 30461 508
rect 30427 -900 30461 -884
rect 30625 492 30659 508
rect 30625 -900 30659 -884
rect 30823 492 30857 508
rect 30823 -900 30857 -884
rect 31021 492 31055 508
rect 31021 -900 31055 -884
rect 31219 492 31253 508
rect 31219 -900 31253 -884
rect 31417 492 31451 508
rect 31417 -900 31451 -884
rect 31615 492 31649 508
rect 31615 -900 31649 -884
rect 23345 -977 23361 -943
rect 23469 -977 23485 -943
rect 23543 -977 23559 -943
rect 23667 -977 23683 -943
rect 23741 -977 23757 -943
rect 23865 -977 23881 -943
rect 23939 -977 23955 -943
rect 24063 -977 24079 -943
rect 24137 -977 24153 -943
rect 24261 -977 24277 -943
rect 24335 -977 24351 -943
rect 24459 -977 24475 -943
rect 24533 -977 24549 -943
rect 24657 -977 24673 -943
rect 24731 -977 24747 -943
rect 24855 -977 24871 -943
rect 24929 -977 24945 -943
rect 25053 -977 25069 -943
rect 25127 -977 25143 -943
rect 25251 -977 25267 -943
rect 25325 -977 25341 -943
rect 25449 -977 25465 -943
rect 25523 -977 25539 -943
rect 25647 -977 25663 -943
rect 25721 -977 25737 -943
rect 25845 -977 25861 -943
rect 25919 -977 25935 -943
rect 26043 -977 26059 -943
rect 26117 -977 26133 -943
rect 26241 -977 26257 -943
rect 26315 -977 26331 -943
rect 26439 -977 26455 -943
rect 26513 -977 26529 -943
rect 26637 -977 26653 -943
rect 26711 -977 26727 -943
rect 26835 -977 26851 -943
rect 26909 -977 26925 -943
rect 27033 -977 27049 -943
rect 27107 -977 27123 -943
rect 27231 -977 27247 -943
rect 27305 -977 27321 -943
rect 27429 -977 27445 -943
rect 27503 -977 27519 -943
rect 27627 -977 27643 -943
rect 27701 -977 27717 -943
rect 27825 -977 27841 -943
rect 27899 -977 27915 -943
rect 28023 -977 28039 -943
rect 28097 -977 28113 -943
rect 28221 -977 28237 -943
rect 28295 -977 28311 -943
rect 28419 -977 28435 -943
rect 28493 -977 28509 -943
rect 28617 -977 28633 -943
rect 28691 -977 28707 -943
rect 28815 -977 28831 -943
rect 28889 -977 28905 -943
rect 29013 -977 29029 -943
rect 29087 -977 29103 -943
rect 29211 -977 29227 -943
rect 29285 -977 29301 -943
rect 29409 -977 29425 -943
rect 29483 -977 29499 -943
rect 29607 -977 29623 -943
rect 29681 -977 29697 -943
rect 29805 -977 29821 -943
rect 29879 -977 29895 -943
rect 30003 -977 30019 -943
rect 30077 -977 30093 -943
rect 30201 -977 30217 -943
rect 30275 -977 30291 -943
rect 30399 -977 30415 -943
rect 30473 -977 30489 -943
rect 30597 -977 30613 -943
rect 30671 -977 30687 -943
rect 30795 -977 30811 -943
rect 30869 -977 30885 -943
rect 30993 -977 31009 -943
rect 31067 -977 31083 -943
rect 31191 -977 31207 -943
rect 31265 -977 31281 -943
rect 31389 -977 31405 -943
rect 31463 -977 31479 -943
rect 31587 -977 31603 -943
rect 23345 -1085 23361 -1051
rect 23469 -1085 23485 -1051
rect 23543 -1085 23559 -1051
rect 23667 -1085 23683 -1051
rect 23741 -1085 23757 -1051
rect 23865 -1085 23881 -1051
rect 23939 -1085 23955 -1051
rect 24063 -1085 24079 -1051
rect 24137 -1085 24153 -1051
rect 24261 -1085 24277 -1051
rect 24335 -1085 24351 -1051
rect 24459 -1085 24475 -1051
rect 24533 -1085 24549 -1051
rect 24657 -1085 24673 -1051
rect 24731 -1085 24747 -1051
rect 24855 -1085 24871 -1051
rect 24929 -1085 24945 -1051
rect 25053 -1085 25069 -1051
rect 25127 -1085 25143 -1051
rect 25251 -1085 25267 -1051
rect 25325 -1085 25341 -1051
rect 25449 -1085 25465 -1051
rect 25523 -1085 25539 -1051
rect 25647 -1085 25663 -1051
rect 25721 -1085 25737 -1051
rect 25845 -1085 25861 -1051
rect 25919 -1085 25935 -1051
rect 26043 -1085 26059 -1051
rect 26117 -1085 26133 -1051
rect 26241 -1085 26257 -1051
rect 26315 -1085 26331 -1051
rect 26439 -1085 26455 -1051
rect 26513 -1085 26529 -1051
rect 26637 -1085 26653 -1051
rect 26711 -1085 26727 -1051
rect 26835 -1085 26851 -1051
rect 26909 -1085 26925 -1051
rect 27033 -1085 27049 -1051
rect 27107 -1085 27123 -1051
rect 27231 -1085 27247 -1051
rect 27305 -1085 27321 -1051
rect 27429 -1085 27445 -1051
rect 27503 -1085 27519 -1051
rect 27627 -1085 27643 -1051
rect 27701 -1085 27717 -1051
rect 27825 -1085 27841 -1051
rect 27899 -1085 27915 -1051
rect 28023 -1085 28039 -1051
rect 28097 -1085 28113 -1051
rect 28221 -1085 28237 -1051
rect 28295 -1085 28311 -1051
rect 28419 -1085 28435 -1051
rect 28493 -1085 28509 -1051
rect 28617 -1085 28633 -1051
rect 28691 -1085 28707 -1051
rect 28815 -1085 28831 -1051
rect 28889 -1085 28905 -1051
rect 29013 -1085 29029 -1051
rect 29087 -1085 29103 -1051
rect 29211 -1085 29227 -1051
rect 29285 -1085 29301 -1051
rect 29409 -1085 29425 -1051
rect 29483 -1085 29499 -1051
rect 29607 -1085 29623 -1051
rect 29681 -1085 29697 -1051
rect 29805 -1085 29821 -1051
rect 29879 -1085 29895 -1051
rect 30003 -1085 30019 -1051
rect 30077 -1085 30093 -1051
rect 30201 -1085 30217 -1051
rect 30275 -1085 30291 -1051
rect 30399 -1085 30415 -1051
rect 30473 -1085 30489 -1051
rect 30597 -1085 30613 -1051
rect 30671 -1085 30687 -1051
rect 30795 -1085 30811 -1051
rect 30869 -1085 30885 -1051
rect 30993 -1085 31009 -1051
rect 31067 -1085 31083 -1051
rect 31191 -1085 31207 -1051
rect 31265 -1085 31281 -1051
rect 31389 -1085 31405 -1051
rect 31463 -1085 31479 -1051
rect 31587 -1085 31603 -1051
rect 23299 -1144 23333 -1128
rect 23299 -2536 23333 -2520
rect 23497 -1144 23531 -1128
rect 23497 -2536 23531 -2520
rect 23695 -1144 23729 -1128
rect 23695 -2536 23729 -2520
rect 23893 -1144 23927 -1128
rect 23893 -2536 23927 -2520
rect 24091 -1144 24125 -1128
rect 24091 -2536 24125 -2520
rect 24289 -1144 24323 -1128
rect 24289 -2536 24323 -2520
rect 24487 -1144 24521 -1128
rect 24487 -2536 24521 -2520
rect 24685 -1144 24719 -1128
rect 24685 -2536 24719 -2520
rect 24883 -1144 24917 -1128
rect 24883 -2536 24917 -2520
rect 25081 -1144 25115 -1128
rect 25081 -2536 25115 -2520
rect 25279 -1144 25313 -1128
rect 25279 -2536 25313 -2520
rect 25477 -1144 25511 -1128
rect 25477 -2536 25511 -2520
rect 25675 -1144 25709 -1128
rect 25675 -2536 25709 -2520
rect 25873 -1144 25907 -1128
rect 25873 -2536 25907 -2520
rect 26071 -1144 26105 -1128
rect 26071 -2536 26105 -2520
rect 26269 -1144 26303 -1128
rect 26269 -2536 26303 -2520
rect 26467 -1144 26501 -1128
rect 26467 -2536 26501 -2520
rect 26665 -1144 26699 -1128
rect 26665 -2536 26699 -2520
rect 26863 -1144 26897 -1128
rect 26863 -2536 26897 -2520
rect 27061 -1144 27095 -1128
rect 27061 -2536 27095 -2520
rect 27259 -1144 27293 -1128
rect 27259 -2536 27293 -2520
rect 27457 -1144 27491 -1128
rect 27457 -2536 27491 -2520
rect 27655 -1144 27689 -1128
rect 27655 -2536 27689 -2520
rect 27853 -1144 27887 -1128
rect 27853 -2536 27887 -2520
rect 28051 -1144 28085 -1128
rect 28051 -2536 28085 -2520
rect 28249 -1144 28283 -1128
rect 28249 -2536 28283 -2520
rect 28447 -1144 28481 -1128
rect 28447 -2536 28481 -2520
rect 28645 -1144 28679 -1128
rect 28645 -2536 28679 -2520
rect 28843 -1144 28877 -1128
rect 28843 -2536 28877 -2520
rect 29041 -1144 29075 -1128
rect 29041 -2536 29075 -2520
rect 29239 -1144 29273 -1128
rect 29239 -2536 29273 -2520
rect 29437 -1144 29471 -1128
rect 29437 -2536 29471 -2520
rect 29635 -1144 29669 -1128
rect 29635 -2536 29669 -2520
rect 29833 -1144 29867 -1128
rect 29833 -2536 29867 -2520
rect 30031 -1144 30065 -1128
rect 30031 -2536 30065 -2520
rect 30229 -1144 30263 -1128
rect 30229 -2536 30263 -2520
rect 30427 -1144 30461 -1128
rect 30427 -2536 30461 -2520
rect 30625 -1144 30659 -1128
rect 30625 -2536 30659 -2520
rect 30823 -1144 30857 -1128
rect 30823 -2536 30857 -2520
rect 31021 -1144 31055 -1128
rect 31021 -2536 31055 -2520
rect 31219 -1144 31253 -1128
rect 31219 -2536 31253 -2520
rect 31417 -1144 31451 -1128
rect 31417 -2536 31451 -2520
rect 31615 -1144 31649 -1128
rect 31615 -2536 31649 -2520
rect 23345 -2613 23361 -2579
rect 23469 -2613 23485 -2579
rect 23543 -2613 23559 -2579
rect 23667 -2613 23683 -2579
rect 23741 -2613 23757 -2579
rect 23865 -2613 23881 -2579
rect 23939 -2613 23955 -2579
rect 24063 -2613 24079 -2579
rect 24137 -2613 24153 -2579
rect 24261 -2613 24277 -2579
rect 24335 -2613 24351 -2579
rect 24459 -2613 24475 -2579
rect 24533 -2613 24549 -2579
rect 24657 -2613 24673 -2579
rect 24731 -2613 24747 -2579
rect 24855 -2613 24871 -2579
rect 24929 -2613 24945 -2579
rect 25053 -2613 25069 -2579
rect 25127 -2613 25143 -2579
rect 25251 -2613 25267 -2579
rect 25325 -2613 25341 -2579
rect 25449 -2613 25465 -2579
rect 25523 -2613 25539 -2579
rect 25647 -2613 25663 -2579
rect 25721 -2613 25737 -2579
rect 25845 -2613 25861 -2579
rect 25919 -2613 25935 -2579
rect 26043 -2613 26059 -2579
rect 26117 -2613 26133 -2579
rect 26241 -2613 26257 -2579
rect 26315 -2613 26331 -2579
rect 26439 -2613 26455 -2579
rect 26513 -2613 26529 -2579
rect 26637 -2613 26653 -2579
rect 26711 -2613 26727 -2579
rect 26835 -2613 26851 -2579
rect 26909 -2613 26925 -2579
rect 27033 -2613 27049 -2579
rect 27107 -2613 27123 -2579
rect 27231 -2613 27247 -2579
rect 27305 -2613 27321 -2579
rect 27429 -2613 27445 -2579
rect 27503 -2613 27519 -2579
rect 27627 -2613 27643 -2579
rect 27701 -2613 27717 -2579
rect 27825 -2613 27841 -2579
rect 27899 -2613 27915 -2579
rect 28023 -2613 28039 -2579
rect 28097 -2613 28113 -2579
rect 28221 -2613 28237 -2579
rect 28295 -2613 28311 -2579
rect 28419 -2613 28435 -2579
rect 28493 -2613 28509 -2579
rect 28617 -2613 28633 -2579
rect 28691 -2613 28707 -2579
rect 28815 -2613 28831 -2579
rect 28889 -2613 28905 -2579
rect 29013 -2613 29029 -2579
rect 29087 -2613 29103 -2579
rect 29211 -2613 29227 -2579
rect 29285 -2613 29301 -2579
rect 29409 -2613 29425 -2579
rect 29483 -2613 29499 -2579
rect 29607 -2613 29623 -2579
rect 29681 -2613 29697 -2579
rect 29805 -2613 29821 -2579
rect 29879 -2613 29895 -2579
rect 30003 -2613 30019 -2579
rect 30077 -2613 30093 -2579
rect 30201 -2613 30217 -2579
rect 30275 -2613 30291 -2579
rect 30399 -2613 30415 -2579
rect 30473 -2613 30489 -2579
rect 30597 -2613 30613 -2579
rect 30671 -2613 30687 -2579
rect 30795 -2613 30811 -2579
rect 30869 -2613 30885 -2579
rect 30993 -2613 31009 -2579
rect 31067 -2613 31083 -2579
rect 31191 -2613 31207 -2579
rect 31265 -2613 31281 -2579
rect 31389 -2613 31405 -2579
rect 31463 -2613 31479 -2579
rect 31587 -2613 31603 -2579
rect 22864 -3034 23342 -2933
rect 31606 -3034 32088 -2933
rect 23345 -3286 23361 -3252
rect 23469 -3286 23485 -3252
rect 23543 -3286 23559 -3252
rect 23667 -3286 23683 -3252
rect 23741 -3286 23757 -3252
rect 23865 -3286 23881 -3252
rect 23939 -3286 23955 -3252
rect 24063 -3286 24079 -3252
rect 24137 -3286 24153 -3252
rect 24261 -3286 24277 -3252
rect 24335 -3286 24351 -3252
rect 24459 -3286 24475 -3252
rect 24533 -3286 24549 -3252
rect 24657 -3286 24673 -3252
rect 24731 -3286 24747 -3252
rect 24855 -3286 24871 -3252
rect 24929 -3286 24945 -3252
rect 25053 -3286 25069 -3252
rect 25127 -3286 25143 -3252
rect 25251 -3286 25267 -3252
rect 25325 -3286 25341 -3252
rect 25449 -3286 25465 -3252
rect 25523 -3286 25539 -3252
rect 25647 -3286 25663 -3252
rect 25721 -3286 25737 -3252
rect 25845 -3286 25861 -3252
rect 25919 -3286 25935 -3252
rect 26043 -3286 26059 -3252
rect 26117 -3286 26133 -3252
rect 26241 -3286 26257 -3252
rect 26315 -3286 26331 -3252
rect 26439 -3286 26455 -3252
rect 26513 -3286 26529 -3252
rect 26637 -3286 26653 -3252
rect 26711 -3286 26727 -3252
rect 26835 -3286 26851 -3252
rect 26909 -3286 26925 -3252
rect 27033 -3286 27049 -3252
rect 27107 -3286 27123 -3252
rect 27231 -3286 27247 -3252
rect 27305 -3286 27321 -3252
rect 27429 -3286 27445 -3252
rect 27503 -3286 27519 -3252
rect 27627 -3286 27643 -3252
rect 27701 -3286 27717 -3252
rect 27825 -3286 27841 -3252
rect 27899 -3286 27915 -3252
rect 28023 -3286 28039 -3252
rect 28097 -3286 28113 -3252
rect 28221 -3286 28237 -3252
rect 28295 -3286 28311 -3252
rect 28419 -3286 28435 -3252
rect 28493 -3286 28509 -3252
rect 28617 -3286 28633 -3252
rect 28691 -3286 28707 -3252
rect 28815 -3286 28831 -3252
rect 28889 -3286 28905 -3252
rect 29013 -3286 29029 -3252
rect 29087 -3286 29103 -3252
rect 29211 -3286 29227 -3252
rect 29285 -3286 29301 -3252
rect 29409 -3286 29425 -3252
rect 29483 -3286 29499 -3252
rect 29607 -3286 29623 -3252
rect 29681 -3286 29697 -3252
rect 29805 -3286 29821 -3252
rect 29879 -3286 29895 -3252
rect 30003 -3286 30019 -3252
rect 30077 -3286 30093 -3252
rect 30201 -3286 30217 -3252
rect 30275 -3286 30291 -3252
rect 30399 -3286 30415 -3252
rect 30473 -3286 30489 -3252
rect 30597 -3286 30613 -3252
rect 30671 -3286 30687 -3252
rect 30795 -3286 30811 -3252
rect 30869 -3286 30885 -3252
rect 30993 -3286 31009 -3252
rect 31067 -3286 31083 -3252
rect 31191 -3286 31207 -3252
rect 31265 -3286 31281 -3252
rect 31389 -3286 31405 -3252
rect 31463 -3286 31479 -3252
rect 31587 -3286 31603 -3252
rect 23299 -3345 23333 -3329
rect 22864 -4415 22875 -4353
rect 22830 -5214 22864 -4427
rect 23299 -4737 23333 -4721
rect 23497 -3345 23531 -3329
rect 23497 -4737 23531 -4721
rect 23695 -3345 23729 -3329
rect 23695 -4737 23729 -4721
rect 23893 -3345 23927 -3329
rect 23893 -4737 23927 -4721
rect 24091 -3345 24125 -3329
rect 24091 -4737 24125 -4721
rect 24289 -3345 24323 -3329
rect 24289 -4737 24323 -4721
rect 24487 -3345 24521 -3329
rect 24487 -4737 24521 -4721
rect 24685 -3345 24719 -3329
rect 24685 -4737 24719 -4721
rect 24883 -3345 24917 -3329
rect 24883 -4737 24917 -4721
rect 25081 -3345 25115 -3329
rect 25081 -4737 25115 -4721
rect 25279 -3345 25313 -3329
rect 25279 -4737 25313 -4721
rect 25477 -3345 25511 -3329
rect 25477 -4737 25511 -4721
rect 25675 -3345 25709 -3329
rect 25675 -4737 25709 -4721
rect 25873 -3345 25907 -3329
rect 25873 -4737 25907 -4721
rect 26071 -3345 26105 -3329
rect 26071 -4737 26105 -4721
rect 26269 -3345 26303 -3329
rect 26269 -4737 26303 -4721
rect 26467 -3345 26501 -3329
rect 26467 -4737 26501 -4721
rect 26665 -3345 26699 -3329
rect 26665 -4737 26699 -4721
rect 26863 -3345 26897 -3329
rect 26863 -4737 26897 -4721
rect 27061 -3345 27095 -3329
rect 27061 -4737 27095 -4721
rect 27259 -3345 27293 -3329
rect 27259 -4737 27293 -4721
rect 27457 -3345 27491 -3329
rect 27457 -4737 27491 -4721
rect 27655 -3345 27689 -3329
rect 27655 -4737 27689 -4721
rect 27853 -3345 27887 -3329
rect 27853 -4737 27887 -4721
rect 28051 -3345 28085 -3329
rect 28051 -4737 28085 -4721
rect 28249 -3345 28283 -3329
rect 28249 -4737 28283 -4721
rect 28447 -3345 28481 -3329
rect 28447 -4737 28481 -4721
rect 28645 -3345 28679 -3329
rect 28645 -4737 28679 -4721
rect 28843 -3345 28877 -3329
rect 28843 -4737 28877 -4721
rect 29041 -3345 29075 -3329
rect 29041 -4737 29075 -4721
rect 29239 -3345 29273 -3329
rect 29239 -4737 29273 -4721
rect 29437 -3345 29471 -3329
rect 29437 -4737 29471 -4721
rect 29635 -3345 29669 -3329
rect 29635 -4737 29669 -4721
rect 29833 -3345 29867 -3329
rect 29833 -4737 29867 -4721
rect 30031 -3345 30065 -3329
rect 30031 -4737 30065 -4721
rect 30229 -3345 30263 -3329
rect 30229 -4737 30263 -4721
rect 30427 -3345 30461 -3329
rect 30427 -4737 30461 -4721
rect 30625 -3345 30659 -3329
rect 30625 -4737 30659 -4721
rect 30823 -3345 30857 -3329
rect 30823 -4737 30857 -4721
rect 31021 -3345 31055 -3329
rect 31021 -4737 31055 -4721
rect 31219 -3345 31253 -3329
rect 31219 -4737 31253 -4721
rect 31417 -3345 31451 -3329
rect 31417 -4737 31451 -4721
rect 31615 -3345 31649 -3329
rect 31615 -4737 31649 -4721
rect 32088 -5214 32122 -4731
rect -848 -5248 -457 -5214
rect 31740 -5248 32122 -5214
<< viali >>
rect 11449 752 11483 2128
rect 11647 752 11681 2128
rect 11845 752 11879 2128
rect 12043 752 12077 2128
rect 12241 752 12275 2128
rect 12439 752 12473 2128
rect 12637 752 12671 2128
rect 12835 752 12869 2128
rect 13033 752 13067 2128
rect 13231 752 13265 2128
rect 13429 752 13463 2128
rect 13627 752 13661 2128
rect 13825 752 13859 2128
rect 14023 752 14057 2128
rect 14221 752 14255 2128
rect 14419 752 14453 2128
rect 14617 752 14651 2128
rect 14815 752 14849 2128
rect 15013 752 15047 2128
rect 15211 752 15245 2128
rect 15409 752 15443 2128
rect 15607 752 15641 2128
rect 15805 752 15839 2128
rect 16003 752 16037 2128
rect 16201 752 16235 2128
rect 16399 752 16433 2128
rect 16597 752 16631 2128
rect 16795 752 16829 2128
rect 16993 752 17027 2128
rect 17191 752 17225 2128
rect 17389 752 17423 2128
rect 17587 752 17621 2128
rect 17785 752 17819 2128
rect 17983 752 18017 2128
rect 18181 752 18215 2128
rect 18379 752 18413 2128
rect 18577 752 18611 2128
rect 18775 752 18809 2128
rect 18973 752 19007 2128
rect 19171 752 19205 2128
rect 19369 752 19403 2128
rect 19567 752 19601 2128
rect 19765 752 19799 2128
rect 11511 659 11619 693
rect 11709 659 11817 693
rect 11907 659 12015 693
rect 12105 659 12213 693
rect 12303 659 12411 693
rect 12501 659 12609 693
rect 12699 659 12807 693
rect 12897 659 13005 693
rect 13095 659 13203 693
rect 13293 659 13401 693
rect 13491 659 13599 693
rect 13689 659 13797 693
rect 13887 659 13995 693
rect 14085 659 14193 693
rect 14283 659 14391 693
rect 14481 659 14589 693
rect 14679 659 14787 693
rect 14877 659 14985 693
rect 15075 659 15183 693
rect 15273 659 15381 693
rect 15471 659 15579 693
rect 15669 659 15777 693
rect 15867 659 15975 693
rect 16065 659 16173 693
rect 16263 659 16371 693
rect 16461 659 16569 693
rect 16659 659 16767 693
rect 16857 659 16965 693
rect 17055 659 17163 693
rect 17253 659 17361 693
rect 17451 659 17559 693
rect 17649 659 17757 693
rect 17847 659 17955 693
rect 18045 659 18153 693
rect 18243 659 18351 693
rect 18441 659 18549 693
rect 18639 659 18747 693
rect 18837 659 18945 693
rect 19035 659 19143 693
rect 19233 659 19341 693
rect 19431 659 19539 693
rect 19629 659 19737 693
rect 11511 551 11619 585
rect 11709 551 11817 585
rect 11907 551 12015 585
rect 12105 551 12213 585
rect 12303 551 12411 585
rect 12501 551 12609 585
rect 12699 551 12807 585
rect 12897 551 13005 585
rect 13095 551 13203 585
rect 13293 551 13401 585
rect 13491 551 13599 585
rect 13689 551 13797 585
rect 13887 551 13995 585
rect 14085 551 14193 585
rect 14283 551 14391 585
rect 14481 551 14589 585
rect 14679 551 14787 585
rect 14877 551 14985 585
rect 15075 551 15183 585
rect 15273 551 15381 585
rect 15471 551 15579 585
rect 15669 551 15777 585
rect 15867 551 15975 585
rect 16065 551 16173 585
rect 16263 551 16371 585
rect 16461 551 16569 585
rect 16659 551 16767 585
rect 16857 551 16965 585
rect 17055 551 17163 585
rect 17253 551 17361 585
rect 17451 551 17559 585
rect 17649 551 17757 585
rect 17847 551 17955 585
rect 18045 551 18153 585
rect 18243 551 18351 585
rect 18441 551 18549 585
rect 18639 551 18747 585
rect 18837 551 18945 585
rect 19035 551 19143 585
rect 19233 551 19341 585
rect 19431 551 19539 585
rect 19629 551 19737 585
rect 11449 -884 11483 492
rect 11647 -884 11681 492
rect 11845 -884 11879 492
rect 12043 -884 12077 492
rect 12241 -884 12275 492
rect 12439 -884 12473 492
rect 12637 -884 12671 492
rect 12835 -884 12869 492
rect 13033 -884 13067 492
rect 13231 -884 13265 492
rect 13429 -884 13463 492
rect 13627 -884 13661 492
rect 13825 -884 13859 492
rect 14023 -884 14057 492
rect 14221 -884 14255 492
rect 14419 -884 14453 492
rect 14617 -884 14651 492
rect 14815 -884 14849 492
rect 15013 -884 15047 492
rect 15211 -884 15245 492
rect 15409 -884 15443 492
rect 15607 -884 15641 492
rect 15805 -884 15839 492
rect 16003 -884 16037 492
rect 16201 -884 16235 492
rect 16399 -884 16433 492
rect 16597 -884 16631 492
rect 16795 -884 16829 492
rect 16993 -884 17027 492
rect 17191 -884 17225 492
rect 17389 -884 17423 492
rect 17587 -884 17621 492
rect 17785 -884 17819 492
rect 17983 -884 18017 492
rect 18181 -884 18215 492
rect 18379 -884 18413 492
rect 18577 -884 18611 492
rect 18775 -884 18809 492
rect 18973 -884 19007 492
rect 19171 -884 19205 492
rect 19369 -884 19403 492
rect 19567 -884 19601 492
rect 19765 -884 19799 492
rect 11511 -977 11619 -943
rect 11709 -977 11817 -943
rect 11907 -977 12015 -943
rect 12105 -977 12213 -943
rect 12303 -977 12411 -943
rect 12501 -977 12609 -943
rect 12699 -977 12807 -943
rect 12897 -977 13005 -943
rect 13095 -977 13203 -943
rect 13293 -977 13401 -943
rect 13491 -977 13599 -943
rect 13689 -977 13797 -943
rect 13887 -977 13995 -943
rect 14085 -977 14193 -943
rect 14283 -977 14391 -943
rect 14481 -977 14589 -943
rect 14679 -977 14787 -943
rect 14877 -977 14985 -943
rect 15075 -977 15183 -943
rect 15273 -977 15381 -943
rect 15471 -977 15579 -943
rect 15669 -977 15777 -943
rect 15867 -977 15975 -943
rect 16065 -977 16173 -943
rect 16263 -977 16371 -943
rect 16461 -977 16569 -943
rect 16659 -977 16767 -943
rect 16857 -977 16965 -943
rect 17055 -977 17163 -943
rect 17253 -977 17361 -943
rect 17451 -977 17559 -943
rect 17649 -977 17757 -943
rect 17847 -977 17955 -943
rect 18045 -977 18153 -943
rect 18243 -977 18351 -943
rect 18441 -977 18549 -943
rect 18639 -977 18747 -943
rect 18837 -977 18945 -943
rect 19035 -977 19143 -943
rect 19233 -977 19341 -943
rect 19431 -977 19539 -943
rect 19629 -977 19737 -943
rect 11511 -1085 11619 -1051
rect 11709 -1085 11817 -1051
rect 11907 -1085 12015 -1051
rect 12105 -1085 12213 -1051
rect 12303 -1085 12411 -1051
rect 12501 -1085 12609 -1051
rect 12699 -1085 12807 -1051
rect 12897 -1085 13005 -1051
rect 13095 -1085 13203 -1051
rect 13293 -1085 13401 -1051
rect 13491 -1085 13599 -1051
rect 13689 -1085 13797 -1051
rect 13887 -1085 13995 -1051
rect 14085 -1085 14193 -1051
rect 14283 -1085 14391 -1051
rect 14481 -1085 14589 -1051
rect 14679 -1085 14787 -1051
rect 14877 -1085 14985 -1051
rect 15075 -1085 15183 -1051
rect 15273 -1085 15381 -1051
rect 15471 -1085 15579 -1051
rect 15669 -1085 15777 -1051
rect 15867 -1085 15975 -1051
rect 16065 -1085 16173 -1051
rect 16263 -1085 16371 -1051
rect 16461 -1085 16569 -1051
rect 16659 -1085 16767 -1051
rect 16857 -1085 16965 -1051
rect 17055 -1085 17163 -1051
rect 17253 -1085 17361 -1051
rect 17451 -1085 17559 -1051
rect 17649 -1085 17757 -1051
rect 17847 -1085 17955 -1051
rect 18045 -1085 18153 -1051
rect 18243 -1085 18351 -1051
rect 18441 -1085 18549 -1051
rect 18639 -1085 18747 -1051
rect 18837 -1085 18945 -1051
rect 19035 -1085 19143 -1051
rect 19233 -1085 19341 -1051
rect 19431 -1085 19539 -1051
rect 19629 -1085 19737 -1051
rect 11449 -2520 11483 -1144
rect 11647 -2520 11681 -1144
rect 11845 -2520 11879 -1144
rect 12043 -2520 12077 -1144
rect 12241 -2520 12275 -1144
rect 12439 -2520 12473 -1144
rect 12637 -2520 12671 -1144
rect 12835 -2520 12869 -1144
rect 13033 -2520 13067 -1144
rect 13231 -2520 13265 -1144
rect 13429 -2520 13463 -1144
rect 13627 -2520 13661 -1144
rect 13825 -2520 13859 -1144
rect 14023 -2520 14057 -1144
rect 14221 -2520 14255 -1144
rect 14419 -2520 14453 -1144
rect 14617 -2520 14651 -1144
rect 14815 -2520 14849 -1144
rect 15013 -2520 15047 -1144
rect 15211 -2520 15245 -1144
rect 15409 -2520 15443 -1144
rect 15607 -2520 15641 -1144
rect 15805 -2520 15839 -1144
rect 16003 -2520 16037 -1144
rect 16201 -2520 16235 -1144
rect 16399 -2520 16433 -1144
rect 16597 -2520 16631 -1144
rect 16795 -2520 16829 -1144
rect 16993 -2520 17027 -1144
rect 17191 -2520 17225 -1144
rect 17389 -2520 17423 -1144
rect 17587 -2520 17621 -1144
rect 17785 -2520 17819 -1144
rect 17983 -2520 18017 -1144
rect 18181 -2520 18215 -1144
rect 18379 -2520 18413 -1144
rect 18577 -2520 18611 -1144
rect 18775 -2520 18809 -1144
rect 18973 -2520 19007 -1144
rect 19171 -2520 19205 -1144
rect 19369 -2520 19403 -1144
rect 19567 -2520 19601 -1144
rect 19765 -2520 19799 -1144
rect 11511 -2613 11619 -2579
rect 11709 -2613 11817 -2579
rect 11907 -2613 12015 -2579
rect 12105 -2613 12213 -2579
rect 12303 -2613 12411 -2579
rect 12501 -2613 12609 -2579
rect 12699 -2613 12807 -2579
rect 12897 -2613 13005 -2579
rect 13095 -2613 13203 -2579
rect 13293 -2613 13401 -2579
rect 13491 -2613 13599 -2579
rect 13689 -2613 13797 -2579
rect 13887 -2613 13995 -2579
rect 14085 -2613 14193 -2579
rect 14283 -2613 14391 -2579
rect 14481 -2613 14589 -2579
rect 14679 -2613 14787 -2579
rect 14877 -2613 14985 -2579
rect 15075 -2613 15183 -2579
rect 15273 -2613 15381 -2579
rect 15471 -2613 15579 -2579
rect 15669 -2613 15777 -2579
rect 15867 -2613 15975 -2579
rect 16065 -2613 16173 -2579
rect 16263 -2613 16371 -2579
rect 16461 -2613 16569 -2579
rect 16659 -2613 16767 -2579
rect 16857 -2613 16965 -2579
rect 17055 -2613 17163 -2579
rect 17253 -2613 17361 -2579
rect 17451 -2613 17559 -2579
rect 17649 -2613 17757 -2579
rect 17847 -2613 17955 -2579
rect 18045 -2613 18153 -2579
rect 18243 -2613 18351 -2579
rect 18441 -2613 18549 -2579
rect 18639 -2613 18747 -2579
rect 18837 -2613 18945 -2579
rect 19035 -2613 19143 -2579
rect 19233 -2613 19341 -2579
rect 19431 -2613 19539 -2579
rect 19629 -2613 19737 -2579
rect 11511 -3286 11619 -3252
rect 11709 -3286 11817 -3252
rect 11907 -3286 12015 -3252
rect 12105 -3286 12213 -3252
rect 12303 -3286 12411 -3252
rect 12501 -3286 12609 -3252
rect 12699 -3286 12807 -3252
rect 12897 -3286 13005 -3252
rect 13095 -3286 13203 -3252
rect 13293 -3286 13401 -3252
rect 13491 -3286 13599 -3252
rect 13689 -3286 13797 -3252
rect 13887 -3286 13995 -3252
rect 14085 -3286 14193 -3252
rect 14283 -3286 14391 -3252
rect 14481 -3286 14589 -3252
rect 14679 -3286 14787 -3252
rect 14877 -3286 14985 -3252
rect 15075 -3286 15183 -3252
rect 15273 -3286 15381 -3252
rect 15471 -3286 15579 -3252
rect 15669 -3286 15777 -3252
rect 15867 -3286 15975 -3252
rect 16065 -3286 16173 -3252
rect 16263 -3286 16371 -3252
rect 16461 -3286 16569 -3252
rect 16659 -3286 16767 -3252
rect 16857 -3286 16965 -3252
rect 17055 -3286 17163 -3252
rect 17253 -3286 17361 -3252
rect 17451 -3286 17559 -3252
rect 17649 -3286 17757 -3252
rect 17847 -3286 17955 -3252
rect 18045 -3286 18153 -3252
rect 18243 -3286 18351 -3252
rect 18441 -3286 18549 -3252
rect 18639 -3286 18747 -3252
rect 18837 -3286 18945 -3252
rect 19035 -3286 19143 -3252
rect 19233 -3286 19341 -3252
rect 19431 -3286 19539 -3252
rect 19629 -3286 19737 -3252
rect 11449 -4721 11483 -3345
rect 11647 -4721 11681 -3345
rect 11845 -4721 11879 -3345
rect 12043 -4721 12077 -3345
rect 12241 -4721 12275 -3345
rect 12439 -4721 12473 -3345
rect 12637 -4721 12671 -3345
rect 12835 -4721 12869 -3345
rect 13033 -4721 13067 -3345
rect 13231 -4721 13265 -3345
rect 13429 -4721 13463 -3345
rect 13627 -4721 13661 -3345
rect 13825 -4721 13859 -3345
rect 14023 -4721 14057 -3345
rect 14221 -4721 14255 -3345
rect 14419 -4721 14453 -3345
rect 14617 -4721 14651 -3345
rect 14815 -4721 14849 -3345
rect 15013 -4721 15047 -3345
rect 15211 -4721 15245 -3345
rect 15409 -4721 15443 -3345
rect 15607 -4721 15641 -3345
rect 15805 -4721 15839 -3345
rect 16003 -4721 16037 -3345
rect 16201 -4721 16235 -3345
rect 16399 -4721 16433 -3345
rect 16597 -4721 16631 -3345
rect 16795 -4721 16829 -3345
rect 16993 -4721 17027 -3345
rect 17191 -4721 17225 -3345
rect 17389 -4721 17423 -3345
rect 17587 -4721 17621 -3345
rect 17785 -4721 17819 -3345
rect 17983 -4721 18017 -3345
rect 18181 -4721 18215 -3345
rect 18379 -4721 18413 -3345
rect 18577 -4721 18611 -3345
rect 18775 -4721 18809 -3345
rect 18973 -4721 19007 -3345
rect 19171 -4721 19205 -3345
rect 19369 -4721 19403 -3345
rect 19567 -4721 19601 -3345
rect 19765 -4721 19799 -3345
rect 23299 752 23333 2128
rect 23497 752 23531 2128
rect 23695 752 23729 2128
rect 23893 752 23927 2128
rect 24091 752 24125 2128
rect 24289 752 24323 2128
rect 24487 752 24521 2128
rect 24685 752 24719 2128
rect 24883 752 24917 2128
rect 25081 752 25115 2128
rect 25279 752 25313 2128
rect 25477 752 25511 2128
rect 25675 752 25709 2128
rect 25873 752 25907 2128
rect 26071 752 26105 2128
rect 26269 752 26303 2128
rect 26467 752 26501 2128
rect 26665 752 26699 2128
rect 26863 752 26897 2128
rect 27061 752 27095 2128
rect 27259 752 27293 2128
rect 27457 752 27491 2128
rect 27655 752 27689 2128
rect 27853 752 27887 2128
rect 28051 752 28085 2128
rect 28249 752 28283 2128
rect 28447 752 28481 2128
rect 28645 752 28679 2128
rect 28843 752 28877 2128
rect 29041 752 29075 2128
rect 29239 752 29273 2128
rect 29437 752 29471 2128
rect 29635 752 29669 2128
rect 29833 752 29867 2128
rect 30031 752 30065 2128
rect 30229 752 30263 2128
rect 30427 752 30461 2128
rect 30625 752 30659 2128
rect 30823 752 30857 2128
rect 31021 752 31055 2128
rect 31219 752 31253 2128
rect 31417 752 31451 2128
rect 31615 752 31649 2128
rect 23361 659 23469 693
rect 23559 659 23667 693
rect 23757 659 23865 693
rect 23955 659 24063 693
rect 24153 659 24261 693
rect 24351 659 24459 693
rect 24549 659 24657 693
rect 24747 659 24855 693
rect 24945 659 25053 693
rect 25143 659 25251 693
rect 25341 659 25449 693
rect 25539 659 25647 693
rect 25737 659 25845 693
rect 25935 659 26043 693
rect 26133 659 26241 693
rect 26331 659 26439 693
rect 26529 659 26637 693
rect 26727 659 26835 693
rect 26925 659 27033 693
rect 27123 659 27231 693
rect 27321 659 27429 693
rect 27519 659 27627 693
rect 27717 659 27825 693
rect 27915 659 28023 693
rect 28113 659 28221 693
rect 28311 659 28419 693
rect 28509 659 28617 693
rect 28707 659 28815 693
rect 28905 659 29013 693
rect 29103 659 29211 693
rect 29301 659 29409 693
rect 29499 659 29607 693
rect 29697 659 29805 693
rect 29895 659 30003 693
rect 30093 659 30201 693
rect 30291 659 30399 693
rect 30489 659 30597 693
rect 30687 659 30795 693
rect 30885 659 30993 693
rect 31083 659 31191 693
rect 31281 659 31389 693
rect 31479 659 31587 693
rect 23361 551 23469 585
rect 23559 551 23667 585
rect 23757 551 23865 585
rect 23955 551 24063 585
rect 24153 551 24261 585
rect 24351 551 24459 585
rect 24549 551 24657 585
rect 24747 551 24855 585
rect 24945 551 25053 585
rect 25143 551 25251 585
rect 25341 551 25449 585
rect 25539 551 25647 585
rect 25737 551 25845 585
rect 25935 551 26043 585
rect 26133 551 26241 585
rect 26331 551 26439 585
rect 26529 551 26637 585
rect 26727 551 26835 585
rect 26925 551 27033 585
rect 27123 551 27231 585
rect 27321 551 27429 585
rect 27519 551 27627 585
rect 27717 551 27825 585
rect 27915 551 28023 585
rect 28113 551 28221 585
rect 28311 551 28419 585
rect 28509 551 28617 585
rect 28707 551 28815 585
rect 28905 551 29013 585
rect 29103 551 29211 585
rect 29301 551 29409 585
rect 29499 551 29607 585
rect 29697 551 29805 585
rect 29895 551 30003 585
rect 30093 551 30201 585
rect 30291 551 30399 585
rect 30489 551 30597 585
rect 30687 551 30795 585
rect 30885 551 30993 585
rect 31083 551 31191 585
rect 31281 551 31389 585
rect 31479 551 31587 585
rect 23299 -884 23333 492
rect 23497 -884 23531 492
rect 23695 -884 23729 492
rect 23893 -884 23927 492
rect 24091 -884 24125 492
rect 24289 -884 24323 492
rect 24487 -884 24521 492
rect 24685 -884 24719 492
rect 24883 -884 24917 492
rect 25081 -884 25115 492
rect 25279 -884 25313 492
rect 25477 -884 25511 492
rect 25675 -884 25709 492
rect 25873 -884 25907 492
rect 26071 -884 26105 492
rect 26269 -884 26303 492
rect 26467 -884 26501 492
rect 26665 -884 26699 492
rect 26863 -884 26897 492
rect 27061 -884 27095 492
rect 27259 -884 27293 492
rect 27457 -884 27491 492
rect 27655 -884 27689 492
rect 27853 -884 27887 492
rect 28051 -884 28085 492
rect 28249 -884 28283 492
rect 28447 -884 28481 492
rect 28645 -884 28679 492
rect 28843 -884 28877 492
rect 29041 -884 29075 492
rect 29239 -884 29273 492
rect 29437 -884 29471 492
rect 29635 -884 29669 492
rect 29833 -884 29867 492
rect 30031 -884 30065 492
rect 30229 -884 30263 492
rect 30427 -884 30461 492
rect 30625 -884 30659 492
rect 30823 -884 30857 492
rect 31021 -884 31055 492
rect 31219 -884 31253 492
rect 31417 -884 31451 492
rect 31615 -884 31649 492
rect 23361 -977 23469 -943
rect 23559 -977 23667 -943
rect 23757 -977 23865 -943
rect 23955 -977 24063 -943
rect 24153 -977 24261 -943
rect 24351 -977 24459 -943
rect 24549 -977 24657 -943
rect 24747 -977 24855 -943
rect 24945 -977 25053 -943
rect 25143 -977 25251 -943
rect 25341 -977 25449 -943
rect 25539 -977 25647 -943
rect 25737 -977 25845 -943
rect 25935 -977 26043 -943
rect 26133 -977 26241 -943
rect 26331 -977 26439 -943
rect 26529 -977 26637 -943
rect 26727 -977 26835 -943
rect 26925 -977 27033 -943
rect 27123 -977 27231 -943
rect 27321 -977 27429 -943
rect 27519 -977 27627 -943
rect 27717 -977 27825 -943
rect 27915 -977 28023 -943
rect 28113 -977 28221 -943
rect 28311 -977 28419 -943
rect 28509 -977 28617 -943
rect 28707 -977 28815 -943
rect 28905 -977 29013 -943
rect 29103 -977 29211 -943
rect 29301 -977 29409 -943
rect 29499 -977 29607 -943
rect 29697 -977 29805 -943
rect 29895 -977 30003 -943
rect 30093 -977 30201 -943
rect 30291 -977 30399 -943
rect 30489 -977 30597 -943
rect 30687 -977 30795 -943
rect 30885 -977 30993 -943
rect 31083 -977 31191 -943
rect 31281 -977 31389 -943
rect 31479 -977 31587 -943
rect 23361 -1085 23469 -1051
rect 23559 -1085 23667 -1051
rect 23757 -1085 23865 -1051
rect 23955 -1085 24063 -1051
rect 24153 -1085 24261 -1051
rect 24351 -1085 24459 -1051
rect 24549 -1085 24657 -1051
rect 24747 -1085 24855 -1051
rect 24945 -1085 25053 -1051
rect 25143 -1085 25251 -1051
rect 25341 -1085 25449 -1051
rect 25539 -1085 25647 -1051
rect 25737 -1085 25845 -1051
rect 25935 -1085 26043 -1051
rect 26133 -1085 26241 -1051
rect 26331 -1085 26439 -1051
rect 26529 -1085 26637 -1051
rect 26727 -1085 26835 -1051
rect 26925 -1085 27033 -1051
rect 27123 -1085 27231 -1051
rect 27321 -1085 27429 -1051
rect 27519 -1085 27627 -1051
rect 27717 -1085 27825 -1051
rect 27915 -1085 28023 -1051
rect 28113 -1085 28221 -1051
rect 28311 -1085 28419 -1051
rect 28509 -1085 28617 -1051
rect 28707 -1085 28815 -1051
rect 28905 -1085 29013 -1051
rect 29103 -1085 29211 -1051
rect 29301 -1085 29409 -1051
rect 29499 -1085 29607 -1051
rect 29697 -1085 29805 -1051
rect 29895 -1085 30003 -1051
rect 30093 -1085 30201 -1051
rect 30291 -1085 30399 -1051
rect 30489 -1085 30597 -1051
rect 30687 -1085 30795 -1051
rect 30885 -1085 30993 -1051
rect 31083 -1085 31191 -1051
rect 31281 -1085 31389 -1051
rect 31479 -1085 31587 -1051
rect 23299 -2520 23333 -1144
rect 23497 -2520 23531 -1144
rect 23695 -2520 23729 -1144
rect 23893 -2520 23927 -1144
rect 24091 -2520 24125 -1144
rect 24289 -2520 24323 -1144
rect 24487 -2520 24521 -1144
rect 24685 -2520 24719 -1144
rect 24883 -2520 24917 -1144
rect 25081 -2520 25115 -1144
rect 25279 -2520 25313 -1144
rect 25477 -2520 25511 -1144
rect 25675 -2520 25709 -1144
rect 25873 -2520 25907 -1144
rect 26071 -2520 26105 -1144
rect 26269 -2520 26303 -1144
rect 26467 -2520 26501 -1144
rect 26665 -2520 26699 -1144
rect 26863 -2520 26897 -1144
rect 27061 -2520 27095 -1144
rect 27259 -2520 27293 -1144
rect 27457 -2520 27491 -1144
rect 27655 -2520 27689 -1144
rect 27853 -2520 27887 -1144
rect 28051 -2520 28085 -1144
rect 28249 -2520 28283 -1144
rect 28447 -2520 28481 -1144
rect 28645 -2520 28679 -1144
rect 28843 -2520 28877 -1144
rect 29041 -2520 29075 -1144
rect 29239 -2520 29273 -1144
rect 29437 -2520 29471 -1144
rect 29635 -2520 29669 -1144
rect 29833 -2520 29867 -1144
rect 30031 -2520 30065 -1144
rect 30229 -2520 30263 -1144
rect 30427 -2520 30461 -1144
rect 30625 -2520 30659 -1144
rect 30823 -2520 30857 -1144
rect 31021 -2520 31055 -1144
rect 31219 -2520 31253 -1144
rect 31417 -2520 31451 -1144
rect 31615 -2520 31649 -1144
rect 23361 -2613 23469 -2579
rect 23559 -2613 23667 -2579
rect 23757 -2613 23865 -2579
rect 23955 -2613 24063 -2579
rect 24153 -2613 24261 -2579
rect 24351 -2613 24459 -2579
rect 24549 -2613 24657 -2579
rect 24747 -2613 24855 -2579
rect 24945 -2613 25053 -2579
rect 25143 -2613 25251 -2579
rect 25341 -2613 25449 -2579
rect 25539 -2613 25647 -2579
rect 25737 -2613 25845 -2579
rect 25935 -2613 26043 -2579
rect 26133 -2613 26241 -2579
rect 26331 -2613 26439 -2579
rect 26529 -2613 26637 -2579
rect 26727 -2613 26835 -2579
rect 26925 -2613 27033 -2579
rect 27123 -2613 27231 -2579
rect 27321 -2613 27429 -2579
rect 27519 -2613 27627 -2579
rect 27717 -2613 27825 -2579
rect 27915 -2613 28023 -2579
rect 28113 -2613 28221 -2579
rect 28311 -2613 28419 -2579
rect 28509 -2613 28617 -2579
rect 28707 -2613 28815 -2579
rect 28905 -2613 29013 -2579
rect 29103 -2613 29211 -2579
rect 29301 -2613 29409 -2579
rect 29499 -2613 29607 -2579
rect 29697 -2613 29805 -2579
rect 29895 -2613 30003 -2579
rect 30093 -2613 30201 -2579
rect 30291 -2613 30399 -2579
rect 30489 -2613 30597 -2579
rect 30687 -2613 30795 -2579
rect 30885 -2613 30993 -2579
rect 31083 -2613 31191 -2579
rect 31281 -2613 31389 -2579
rect 31479 -2613 31587 -2579
rect 23361 -3286 23469 -3252
rect 23559 -3286 23667 -3252
rect 23757 -3286 23865 -3252
rect 23955 -3286 24063 -3252
rect 24153 -3286 24261 -3252
rect 24351 -3286 24459 -3252
rect 24549 -3286 24657 -3252
rect 24747 -3286 24855 -3252
rect 24945 -3286 25053 -3252
rect 25143 -3286 25251 -3252
rect 25341 -3286 25449 -3252
rect 25539 -3286 25647 -3252
rect 25737 -3286 25845 -3252
rect 25935 -3286 26043 -3252
rect 26133 -3286 26241 -3252
rect 26331 -3286 26439 -3252
rect 26529 -3286 26637 -3252
rect 26727 -3286 26835 -3252
rect 26925 -3286 27033 -3252
rect 27123 -3286 27231 -3252
rect 27321 -3286 27429 -3252
rect 27519 -3286 27627 -3252
rect 27717 -3286 27825 -3252
rect 27915 -3286 28023 -3252
rect 28113 -3286 28221 -3252
rect 28311 -3286 28419 -3252
rect 28509 -3286 28617 -3252
rect 28707 -3286 28815 -3252
rect 28905 -3286 29013 -3252
rect 29103 -3286 29211 -3252
rect 29301 -3286 29409 -3252
rect 29499 -3286 29607 -3252
rect 29697 -3286 29805 -3252
rect 29895 -3286 30003 -3252
rect 30093 -3286 30201 -3252
rect 30291 -3286 30399 -3252
rect 30489 -3286 30597 -3252
rect 30687 -3286 30795 -3252
rect 30885 -3286 30993 -3252
rect 31083 -3286 31191 -3252
rect 31281 -3286 31389 -3252
rect 31479 -3286 31587 -3252
rect 23299 -4721 23333 -3345
rect 23497 -4721 23531 -3345
rect 23695 -4721 23729 -3345
rect 23893 -4721 23927 -3345
rect 24091 -4721 24125 -3345
rect 24289 -4721 24323 -3345
rect 24487 -4721 24521 -3345
rect 24685 -4721 24719 -3345
rect 24883 -4721 24917 -3345
rect 25081 -4721 25115 -3345
rect 25279 -4721 25313 -3345
rect 25477 -4721 25511 -3345
rect 25675 -4721 25709 -3345
rect 25873 -4721 25907 -3345
rect 26071 -4721 26105 -3345
rect 26269 -4721 26303 -3345
rect 26467 -4721 26501 -3345
rect 26665 -4721 26699 -3345
rect 26863 -4721 26897 -3345
rect 27061 -4721 27095 -3345
rect 27259 -4721 27293 -3345
rect 27457 -4721 27491 -3345
rect 27655 -4721 27689 -3345
rect 27853 -4721 27887 -3345
rect 28051 -4721 28085 -3345
rect 28249 -4721 28283 -3345
rect 28447 -4721 28481 -3345
rect 28645 -4721 28679 -3345
rect 28843 -4721 28877 -3345
rect 29041 -4721 29075 -3345
rect 29239 -4721 29273 -3345
rect 29437 -4721 29471 -3345
rect 29635 -4721 29669 -3345
rect 29833 -4721 29867 -3345
rect 30031 -4721 30065 -3345
rect 30229 -4721 30263 -3345
rect 30427 -4721 30461 -3345
rect 30625 -4721 30659 -3345
rect 30823 -4721 30857 -3345
rect 31021 -4721 31055 -3345
rect 31219 -4721 31253 -3345
rect 31417 -4721 31451 -3345
rect 31615 -4721 31649 -3345
<< metal1 >>
rect -396 2128 -350 2327
rect 0 2128 46 2327
rect 396 2128 442 2327
rect 792 2128 838 2327
rect 1188 2128 1234 2327
rect 1584 2128 1630 2327
rect 1980 2128 2026 2327
rect 2376 2128 2422 2327
rect 2772 2128 2818 2327
rect 3168 2128 3214 2327
rect 3564 2128 3610 2327
rect 3960 2128 4006 2327
rect 4356 2128 4402 2327
rect 4752 2128 4798 2327
rect 5148 2128 5194 2327
rect 5544 2128 5590 2327
rect 5940 2128 5986 2327
rect 6336 2128 6382 2327
rect 6732 2128 6778 2327
rect 7128 2128 7174 2327
rect 7524 2128 7570 2327
rect 7920 2129 7966 2327
rect -409 752 -399 2128
rect -347 752 -337 2128
rect -211 752 -201 2128
rect -149 752 -139 2128
rect -13 752 -3 2128
rect 49 752 59 2128
rect 185 752 195 2128
rect 247 752 257 2128
rect 383 752 393 2128
rect 445 752 455 2128
rect 581 752 591 2128
rect 643 752 653 2128
rect 779 752 789 2128
rect 841 752 851 2128
rect 977 752 987 2128
rect 1039 752 1049 2128
rect 1175 752 1185 2128
rect 1237 752 1247 2128
rect 1373 752 1383 2128
rect 1435 752 1445 2128
rect 1571 752 1581 2128
rect 1633 752 1643 2128
rect 1769 752 1779 2128
rect 1831 752 1841 2128
rect 1967 752 1977 2128
rect 2029 752 2039 2128
rect 2165 752 2175 2128
rect 2227 752 2237 2128
rect 2363 752 2373 2128
rect 2425 752 2435 2128
rect 2561 752 2571 2128
rect 2623 752 2633 2128
rect 2759 752 2769 2128
rect 2821 752 2831 2128
rect 2957 752 2967 2128
rect 3019 752 3029 2128
rect 3155 752 3165 2128
rect 3217 752 3227 2128
rect 3353 752 3363 2128
rect 3415 752 3425 2128
rect 3551 752 3561 2128
rect 3613 752 3623 2128
rect 3749 752 3759 2128
rect 3811 752 3821 2128
rect 3947 752 3957 2128
rect 4009 752 4019 2128
rect 4145 752 4155 2128
rect 4207 752 4217 2128
rect 4343 752 4353 2128
rect 4405 752 4415 2128
rect 4541 752 4551 2128
rect 4603 752 4613 2128
rect 4739 752 4749 2128
rect 4801 752 4811 2128
rect 4937 752 4947 2128
rect 4999 752 5009 2128
rect 5135 752 5145 2128
rect 5197 752 5207 2128
rect 5333 752 5343 2128
rect 5395 752 5405 2128
rect 5531 752 5541 2128
rect 5593 752 5603 2128
rect 5729 752 5739 2128
rect 5791 752 5801 2128
rect 5927 752 5937 2128
rect 5989 752 5999 2128
rect 6125 752 6135 2128
rect 6187 752 6197 2128
rect 6323 752 6333 2128
rect 6385 752 6395 2128
rect 6521 752 6531 2128
rect 6583 752 6593 2128
rect 6719 752 6729 2128
rect 6781 752 6791 2128
rect 6917 752 6927 2128
rect 6979 752 6989 2128
rect 7115 752 7125 2128
rect 7177 752 7187 2128
rect 7313 752 7323 2128
rect 7375 752 7385 2128
rect 7511 752 7521 2128
rect 7573 752 7583 2128
rect 7709 752 7719 2128
rect 7771 752 7781 2128
rect 7907 753 7917 2129
rect 7969 753 7979 2129
rect -637 545 8207 699
rect -637 -743 -483 545
rect -637 -877 -627 -743
rect -493 -877 -483 -743
rect -637 -937 -483 -877
rect -409 -884 -399 492
rect -347 -884 -337 492
rect -211 -884 -201 492
rect -149 -884 -139 492
rect -13 -884 -3 492
rect 49 -884 59 492
rect 185 -884 195 492
rect 247 -884 257 492
rect 383 -884 393 492
rect 445 -884 455 492
rect 581 -884 591 492
rect 643 -884 653 492
rect 779 -884 789 492
rect 841 -884 851 492
rect 977 -884 987 492
rect 1039 -884 1049 492
rect 1175 -884 1185 492
rect 1237 -884 1247 492
rect 1373 -884 1383 492
rect 1435 -884 1445 492
rect 1571 -884 1581 492
rect 1633 -884 1643 492
rect 1769 -884 1779 492
rect 1831 -884 1841 492
rect 1967 -884 1977 492
rect 2029 -884 2039 492
rect 2165 -884 2175 492
rect 2227 -884 2237 492
rect 2363 -884 2373 492
rect 2425 -884 2435 492
rect 2561 -884 2571 492
rect 2623 -884 2633 492
rect 2759 -884 2769 492
rect 2821 -884 2831 492
rect 2957 -884 2967 492
rect 3019 -884 3029 492
rect 3155 -884 3165 492
rect 3217 -884 3227 492
rect 3353 -884 3363 492
rect 3415 -884 3425 492
rect 3551 -884 3561 492
rect 3613 -884 3623 492
rect 3749 -884 3759 492
rect 3811 -884 3821 492
rect 3947 -884 3957 492
rect 4009 -884 4019 492
rect 4145 -884 4155 492
rect 4207 -884 4217 492
rect 4343 -884 4353 492
rect 4405 -884 4415 492
rect 4541 -884 4551 492
rect 4603 -884 4613 492
rect 4739 -884 4749 492
rect 4801 -884 4811 492
rect 4937 -884 4947 492
rect 4999 -884 5009 492
rect 5135 -884 5145 492
rect 5197 -884 5207 492
rect 5333 -884 5343 492
rect 5395 -884 5405 492
rect 5531 -884 5541 492
rect 5593 -884 5603 492
rect 5729 -884 5739 492
rect 5791 -884 5801 492
rect 5927 -884 5937 492
rect 5989 -884 5999 492
rect 6125 -884 6135 492
rect 6187 -884 6197 492
rect 6323 -884 6333 492
rect 6385 -884 6395 492
rect 6521 -884 6531 492
rect 6583 -884 6593 492
rect 6719 -884 6729 492
rect 6781 -884 6791 492
rect 6917 -884 6927 492
rect 6979 -884 6989 492
rect 7115 -884 7125 492
rect 7177 -884 7187 492
rect 7313 -884 7323 492
rect 7375 -884 7385 492
rect 7511 -884 7521 492
rect 7573 -884 7583 492
rect 7709 -884 7719 492
rect 7771 -884 7781 492
rect 7907 -883 7917 493
rect 7969 -883 7979 493
rect 8053 -743 8207 545
rect 8053 -877 8063 -743
rect 8197 -877 8207 -743
rect 8053 -937 8207 -877
rect -637 -947 8207 -937
rect -637 -1081 -627 -947
rect -493 -1081 8063 -947
rect 8197 -1081 8207 -947
rect -637 -1091 8207 -1081
rect -637 -1151 -483 -1091
rect -637 -1285 -627 -1151
rect -493 -1285 -483 -1151
rect -637 -2573 -483 -1285
rect -409 -2520 -399 -1144
rect -347 -2520 -337 -1144
rect -211 -2520 -201 -1144
rect -149 -2520 -139 -1144
rect -13 -2520 -3 -1144
rect 49 -2520 59 -1144
rect 185 -2520 195 -1144
rect 247 -2520 257 -1144
rect 383 -2520 393 -1144
rect 445 -2520 455 -1144
rect 581 -2520 591 -1144
rect 643 -2520 653 -1144
rect 779 -2520 789 -1144
rect 841 -2520 851 -1144
rect 977 -2520 987 -1144
rect 1039 -2520 1049 -1144
rect 1175 -2520 1185 -1144
rect 1237 -2520 1247 -1144
rect 1373 -2520 1383 -1144
rect 1435 -2520 1445 -1144
rect 1571 -2520 1581 -1144
rect 1633 -2520 1643 -1144
rect 1769 -2520 1779 -1144
rect 1831 -2520 1841 -1144
rect 1967 -2520 1977 -1144
rect 2029 -2520 2039 -1144
rect 2165 -2520 2175 -1144
rect 2227 -2520 2237 -1144
rect 2363 -2520 2373 -1144
rect 2425 -2520 2435 -1144
rect 2561 -2520 2571 -1144
rect 2623 -2520 2633 -1144
rect 2759 -2520 2769 -1144
rect 2821 -2520 2831 -1144
rect 2957 -2520 2967 -1144
rect 3019 -2520 3029 -1144
rect 3155 -2520 3165 -1144
rect 3217 -2520 3227 -1144
rect 3353 -2520 3363 -1144
rect 3415 -2520 3425 -1144
rect 3551 -2520 3561 -1144
rect 3613 -2520 3623 -1144
rect 3749 -2520 3759 -1144
rect 3811 -2520 3821 -1144
rect 3947 -2520 3957 -1144
rect 4009 -2520 4019 -1144
rect 4145 -2520 4155 -1144
rect 4207 -2520 4217 -1144
rect 4343 -2520 4353 -1144
rect 4405 -2520 4415 -1144
rect 4541 -2520 4551 -1144
rect 4603 -2520 4613 -1144
rect 4739 -2520 4749 -1144
rect 4801 -2520 4811 -1144
rect 4937 -2520 4947 -1144
rect 4999 -2520 5009 -1144
rect 5135 -2520 5145 -1144
rect 5197 -2520 5207 -1144
rect 5333 -2520 5343 -1144
rect 5395 -2520 5405 -1144
rect 5531 -2520 5541 -1144
rect 5593 -2520 5603 -1144
rect 5729 -2520 5739 -1144
rect 5791 -2520 5801 -1144
rect 5927 -2520 5937 -1144
rect 5989 -2520 5999 -1144
rect 6125 -2520 6135 -1144
rect 6187 -2520 6197 -1144
rect 6323 -2520 6333 -1144
rect 6385 -2520 6395 -1144
rect 6521 -2520 6531 -1144
rect 6583 -2520 6593 -1144
rect 6719 -2520 6729 -1144
rect 6781 -2520 6791 -1144
rect 6917 -2520 6927 -1144
rect 6979 -2520 6989 -1144
rect 7115 -2520 7125 -1144
rect 7177 -2520 7187 -1144
rect 7313 -2520 7323 -1144
rect 7375 -2520 7385 -1144
rect 7511 -2520 7521 -1144
rect 7573 -2520 7583 -1144
rect 7709 -2520 7719 -1144
rect 7771 -2520 7781 -1144
rect 7907 -2519 7917 -1143
rect 7969 -2519 7979 -1143
rect 8053 -1151 8207 -1091
rect 8053 -1285 8063 -1151
rect 8197 -1285 8207 -1151
rect 8053 -2573 8207 -1285
rect -637 -2643 8207 -2573
rect -637 -3208 -483 -2643
rect 8053 -3208 8207 -2643
rect -637 -3292 8207 -3208
rect -409 -4721 -399 -3345
rect -347 -4721 -337 -3345
rect -211 -4721 -201 -3345
rect -149 -4721 -139 -3345
rect -13 -4721 -3 -3345
rect 49 -4721 59 -3345
rect 185 -4721 195 -3345
rect 247 -4721 257 -3345
rect 383 -4721 393 -3345
rect 445 -4721 455 -3345
rect 581 -4721 591 -3345
rect 643 -4721 653 -3345
rect 779 -4721 789 -3345
rect 841 -4721 851 -3345
rect 977 -4721 987 -3345
rect 1039 -4721 1049 -3345
rect 1175 -4721 1185 -3345
rect 1237 -4721 1247 -3345
rect 1373 -4721 1383 -3345
rect 1435 -4721 1445 -3345
rect 1571 -4721 1581 -3345
rect 1633 -4721 1643 -3345
rect 1769 -4721 1779 -3345
rect 1831 -4721 1841 -3345
rect 1967 -4721 1977 -3345
rect 2029 -4721 2039 -3345
rect 2165 -4721 2175 -3345
rect 2227 -4721 2237 -3345
rect 2363 -4721 2373 -3345
rect 2425 -4721 2435 -3345
rect 2561 -4721 2571 -3345
rect 2623 -4721 2633 -3345
rect 2759 -4721 2769 -3345
rect 2821 -4721 2831 -3345
rect 2957 -4721 2967 -3345
rect 3019 -4721 3029 -3345
rect 3155 -4721 3165 -3345
rect 3217 -4721 3227 -3345
rect 3353 -4721 3363 -3345
rect 3415 -4721 3425 -3345
rect 3551 -4721 3561 -3345
rect 3613 -4721 3623 -3345
rect 3749 -4721 3759 -3345
rect 3811 -4721 3821 -3345
rect 3947 -4721 3957 -3345
rect 4009 -4721 4019 -3345
rect 4145 -4721 4155 -3345
rect 4207 -4721 4217 -3345
rect 4343 -4721 4353 -3345
rect 4405 -4721 4415 -3345
rect 4541 -4721 4551 -3345
rect 4603 -4721 4613 -3345
rect 4739 -4721 4749 -3345
rect 4801 -4721 4811 -3345
rect 4937 -4721 4947 -3345
rect 4999 -4721 5009 -3345
rect 5135 -4721 5145 -3345
rect 5197 -4721 5207 -3345
rect 5333 -4721 5343 -3345
rect 5395 -4721 5405 -3345
rect 5531 -4721 5541 -3345
rect 5593 -4721 5603 -3345
rect 5729 -4721 5739 -3345
rect 5791 -4721 5801 -3345
rect 5927 -4721 5937 -3345
rect 5989 -4721 5999 -3345
rect 6125 -4721 6135 -3345
rect 6187 -4721 6197 -3345
rect 6323 -4721 6333 -3345
rect 6385 -4721 6395 -3345
rect 6521 -4721 6531 -3345
rect 6583 -4721 6593 -3345
rect 6719 -4721 6729 -3345
rect 6781 -4721 6791 -3345
rect 6917 -4721 6927 -3345
rect 6979 -4721 6989 -3345
rect 7115 -4721 7125 -3345
rect 7177 -4721 7187 -3345
rect 7313 -4721 7323 -3345
rect 7375 -4721 7385 -3345
rect 7511 -4721 7521 -3345
rect 7573 -4721 7583 -3345
rect 7709 -4721 7719 -3345
rect 7771 -4721 7781 -3345
rect 7907 -4720 7917 -3344
rect 7969 -4720 7979 -3344
rect -396 -5127 -350 -4721
rect 0 -5127 46 -4721
rect 396 -5127 442 -4721
rect 792 -5127 838 -4721
rect 1188 -5127 1234 -4721
rect 1584 -5127 1630 -4721
rect 1980 -5127 2026 -4721
rect 2376 -5127 2422 -4721
rect 2772 -5127 2818 -4721
rect 3168 -5127 3214 -4721
rect 3564 -5127 3610 -4721
rect 3960 -5127 4006 -4721
rect 4356 -5127 4402 -4721
rect 4752 -5127 4798 -4721
rect 5148 -5127 5194 -4721
rect 5544 -5127 5590 -4721
rect 5940 -5127 5986 -4721
rect 6336 -5127 6382 -4721
rect 6732 -5127 6778 -4721
rect 7128 -5127 7174 -4721
rect 7524 -5127 7570 -4721
rect 7920 -5127 7966 -4721
rect 9137 -5127 10357 2327
rect 11443 2128 11489 2327
rect 11641 2128 11687 2140
rect 11839 2128 11885 2327
rect 12037 2128 12083 2140
rect 12235 2128 12281 2327
rect 12433 2128 12479 2140
rect 12631 2128 12677 2327
rect 12829 2128 12875 2140
rect 13027 2128 13073 2327
rect 13225 2128 13271 2140
rect 13423 2128 13469 2327
rect 13621 2128 13667 2140
rect 13819 2128 13865 2327
rect 14017 2128 14063 2140
rect 14215 2128 14261 2327
rect 14413 2128 14459 2140
rect 14611 2128 14657 2327
rect 14809 2128 14855 2140
rect 15007 2128 15053 2327
rect 15205 2128 15251 2140
rect 15403 2128 15449 2327
rect 15601 2128 15647 2140
rect 15799 2128 15845 2327
rect 15997 2128 16043 2140
rect 16195 2128 16241 2327
rect 16393 2128 16439 2140
rect 16591 2128 16637 2327
rect 16789 2128 16835 2140
rect 16987 2128 17033 2327
rect 17185 2128 17231 2140
rect 17383 2128 17429 2327
rect 17581 2128 17627 2140
rect 17779 2128 17825 2327
rect 17977 2128 18023 2140
rect 18175 2128 18221 2327
rect 18373 2128 18419 2140
rect 18571 2128 18617 2327
rect 18769 2128 18815 2140
rect 18967 2128 19013 2327
rect 19165 2128 19211 2140
rect 19363 2128 19409 2327
rect 19561 2128 19607 2140
rect 19759 2129 19805 2327
rect 11430 752 11440 2128
rect 11492 752 11502 2128
rect 11628 752 11638 2128
rect 11690 752 11700 2128
rect 11826 752 11836 2128
rect 11888 752 11898 2128
rect 12024 752 12034 2128
rect 12086 752 12096 2128
rect 12222 752 12232 2128
rect 12284 752 12294 2128
rect 12420 752 12430 2128
rect 12482 752 12492 2128
rect 12618 752 12628 2128
rect 12680 752 12690 2128
rect 12816 752 12826 2128
rect 12878 752 12888 2128
rect 13014 752 13024 2128
rect 13076 752 13086 2128
rect 13212 752 13222 2128
rect 13274 752 13284 2128
rect 13410 752 13420 2128
rect 13472 752 13482 2128
rect 13608 752 13618 2128
rect 13670 752 13680 2128
rect 13806 752 13816 2128
rect 13868 752 13878 2128
rect 14004 752 14014 2128
rect 14066 752 14076 2128
rect 14202 752 14212 2128
rect 14264 752 14274 2128
rect 14400 752 14410 2128
rect 14462 752 14472 2128
rect 14598 752 14608 2128
rect 14660 752 14670 2128
rect 14796 752 14806 2128
rect 14858 752 14868 2128
rect 14994 752 15004 2128
rect 15056 752 15066 2128
rect 15192 752 15202 2128
rect 15254 752 15264 2128
rect 15390 752 15400 2128
rect 15452 752 15462 2128
rect 15588 752 15598 2128
rect 15650 752 15660 2128
rect 15786 752 15796 2128
rect 15848 752 15858 2128
rect 15984 752 15994 2128
rect 16046 752 16056 2128
rect 16182 752 16192 2128
rect 16244 752 16254 2128
rect 16380 752 16390 2128
rect 16442 752 16452 2128
rect 16578 752 16588 2128
rect 16640 752 16650 2128
rect 16776 752 16786 2128
rect 16838 752 16848 2128
rect 16974 752 16984 2128
rect 17036 752 17046 2128
rect 17172 752 17182 2128
rect 17234 752 17244 2128
rect 17370 752 17380 2128
rect 17432 752 17442 2128
rect 17568 752 17578 2128
rect 17630 752 17640 2128
rect 17766 752 17776 2128
rect 17828 752 17838 2128
rect 17964 752 17974 2128
rect 18026 752 18036 2128
rect 18162 752 18172 2128
rect 18224 752 18234 2128
rect 18360 752 18370 2128
rect 18422 752 18432 2128
rect 18558 752 18568 2128
rect 18620 752 18630 2128
rect 18756 752 18766 2128
rect 18818 752 18828 2128
rect 18954 752 18964 2128
rect 19016 752 19026 2128
rect 19152 752 19162 2128
rect 19214 752 19224 2128
rect 19350 752 19360 2128
rect 19412 752 19422 2128
rect 19548 752 19558 2128
rect 19610 752 19620 2128
rect 19746 753 19756 2129
rect 19808 753 19818 2129
rect 19759 752 19765 753
rect 19799 752 19805 753
rect 11443 740 11489 752
rect 11641 740 11687 752
rect 11839 740 11885 752
rect 12037 740 12083 752
rect 12235 740 12281 752
rect 12433 740 12479 752
rect 12631 740 12677 752
rect 12829 740 12875 752
rect 13027 740 13073 752
rect 13225 740 13271 752
rect 13423 740 13469 752
rect 13621 740 13667 752
rect 13819 740 13865 752
rect 14017 740 14063 752
rect 14215 740 14261 752
rect 14413 740 14459 752
rect 14611 740 14657 752
rect 14809 740 14855 752
rect 15007 740 15053 752
rect 15205 740 15251 752
rect 15403 740 15449 752
rect 15601 740 15647 752
rect 15799 740 15845 752
rect 15997 740 16043 752
rect 16195 740 16241 752
rect 16393 740 16439 752
rect 16591 740 16637 752
rect 16789 740 16835 752
rect 16987 740 17033 752
rect 17185 740 17231 752
rect 17383 740 17429 752
rect 17581 740 17627 752
rect 17779 740 17825 752
rect 17977 740 18023 752
rect 18175 740 18221 752
rect 18373 740 18419 752
rect 18571 740 18617 752
rect 18769 740 18815 752
rect 18967 740 19013 752
rect 19165 740 19211 752
rect 19363 740 19409 752
rect 19561 740 19607 752
rect 19759 740 19805 752
rect 11202 693 20046 699
rect 11202 659 11511 693
rect 11619 659 11709 693
rect 11817 659 11907 693
rect 12015 659 12105 693
rect 12213 659 12303 693
rect 12411 659 12501 693
rect 12609 659 12699 693
rect 12807 659 12897 693
rect 13005 659 13095 693
rect 13203 659 13293 693
rect 13401 659 13491 693
rect 13599 659 13689 693
rect 13797 659 13887 693
rect 13995 659 14085 693
rect 14193 659 14283 693
rect 14391 659 14481 693
rect 14589 659 14679 693
rect 14787 659 14877 693
rect 14985 659 15075 693
rect 15183 659 15273 693
rect 15381 659 15471 693
rect 15579 659 15669 693
rect 15777 659 15867 693
rect 15975 659 16065 693
rect 16173 659 16263 693
rect 16371 659 16461 693
rect 16569 659 16659 693
rect 16767 659 16857 693
rect 16965 659 17055 693
rect 17163 659 17253 693
rect 17361 659 17451 693
rect 17559 659 17649 693
rect 17757 659 17847 693
rect 17955 659 18045 693
rect 18153 659 18243 693
rect 18351 659 18441 693
rect 18549 659 18639 693
rect 18747 659 18837 693
rect 18945 659 19035 693
rect 19143 659 19233 693
rect 19341 659 19431 693
rect 19539 659 19629 693
rect 19737 659 20046 693
rect 11202 585 20046 659
rect 11202 551 11511 585
rect 11619 551 11709 585
rect 11817 551 11907 585
rect 12015 551 12105 585
rect 12213 551 12303 585
rect 12411 551 12501 585
rect 12609 551 12699 585
rect 12807 551 12897 585
rect 13005 551 13095 585
rect 13203 551 13293 585
rect 13401 551 13491 585
rect 13599 551 13689 585
rect 13797 551 13887 585
rect 13995 551 14085 585
rect 14193 551 14283 585
rect 14391 551 14481 585
rect 14589 551 14679 585
rect 14787 551 14877 585
rect 14985 551 15075 585
rect 15183 551 15273 585
rect 15381 551 15471 585
rect 15579 551 15669 585
rect 15777 551 15867 585
rect 15975 551 16065 585
rect 16173 551 16263 585
rect 16371 551 16461 585
rect 16569 551 16659 585
rect 16767 551 16857 585
rect 16965 551 17055 585
rect 17163 551 17253 585
rect 17361 551 17451 585
rect 17559 551 17649 585
rect 17757 551 17847 585
rect 17955 551 18045 585
rect 18153 551 18243 585
rect 18351 551 18441 585
rect 18549 551 18639 585
rect 18747 551 18837 585
rect 18945 551 19035 585
rect 19143 551 19233 585
rect 19341 551 19431 585
rect 19539 551 19629 585
rect 19737 551 20046 585
rect 11202 545 20046 551
rect 11202 -743 11356 545
rect 11443 492 11489 504
rect 11641 492 11687 504
rect 11839 492 11885 504
rect 12037 492 12083 504
rect 12235 492 12281 504
rect 12433 492 12479 504
rect 12631 492 12677 504
rect 12829 492 12875 504
rect 13027 492 13073 504
rect 13225 492 13271 504
rect 13423 492 13469 504
rect 13621 492 13667 504
rect 13819 492 13865 504
rect 14017 492 14063 504
rect 14215 492 14261 504
rect 14413 492 14459 504
rect 14611 492 14657 504
rect 14809 492 14855 504
rect 15007 492 15053 504
rect 15205 492 15251 504
rect 15403 492 15449 504
rect 15601 492 15647 504
rect 15799 492 15845 504
rect 15997 492 16043 504
rect 16195 492 16241 504
rect 16393 492 16439 504
rect 16591 492 16637 504
rect 16789 492 16835 504
rect 16987 492 17033 504
rect 17185 492 17231 504
rect 17383 492 17429 504
rect 17581 492 17627 504
rect 17779 492 17825 504
rect 17977 492 18023 504
rect 18175 492 18221 504
rect 18373 492 18419 504
rect 18571 492 18617 504
rect 18769 492 18815 504
rect 18967 492 19013 504
rect 19165 492 19211 504
rect 19363 492 19409 504
rect 19561 492 19607 504
rect 19759 493 19805 504
rect 11202 -877 11212 -743
rect 11346 -877 11356 -743
rect 11202 -937 11356 -877
rect 11430 -884 11440 492
rect 11492 -884 11502 492
rect 11628 -884 11638 492
rect 11690 -884 11700 492
rect 11826 -884 11836 492
rect 11888 -884 11898 492
rect 12024 -884 12034 492
rect 12086 -884 12096 492
rect 12222 -884 12232 492
rect 12284 -884 12294 492
rect 12420 -884 12430 492
rect 12482 -884 12492 492
rect 12618 -884 12628 492
rect 12680 -884 12690 492
rect 12816 -884 12826 492
rect 12878 -884 12888 492
rect 13014 -884 13024 492
rect 13076 -884 13086 492
rect 13212 -884 13222 492
rect 13274 -884 13284 492
rect 13410 -884 13420 492
rect 13472 -884 13482 492
rect 13608 -884 13618 492
rect 13670 -884 13680 492
rect 13806 -884 13816 492
rect 13868 -884 13878 492
rect 14004 -884 14014 492
rect 14066 -884 14076 492
rect 14202 -884 14212 492
rect 14264 -884 14274 492
rect 14400 -884 14410 492
rect 14462 -884 14472 492
rect 14598 -884 14608 492
rect 14660 -884 14670 492
rect 14796 -884 14806 492
rect 14858 -884 14868 492
rect 14994 -884 15004 492
rect 15056 -884 15066 492
rect 15192 -884 15202 492
rect 15254 -884 15264 492
rect 15390 -884 15400 492
rect 15452 -884 15462 492
rect 15588 -884 15598 492
rect 15650 -884 15660 492
rect 15786 -884 15796 492
rect 15848 -884 15858 492
rect 15984 -884 15994 492
rect 16046 -884 16056 492
rect 16182 -884 16192 492
rect 16244 -884 16254 492
rect 16380 -884 16390 492
rect 16442 -884 16452 492
rect 16578 -884 16588 492
rect 16640 -884 16650 492
rect 16776 -884 16786 492
rect 16838 -884 16848 492
rect 16974 -884 16984 492
rect 17036 -884 17046 492
rect 17172 -884 17182 492
rect 17234 -884 17244 492
rect 17370 -884 17380 492
rect 17432 -884 17442 492
rect 17568 -884 17578 492
rect 17630 -884 17640 492
rect 17766 -884 17776 492
rect 17828 -884 17838 492
rect 17964 -884 17974 492
rect 18026 -884 18036 492
rect 18162 -884 18172 492
rect 18224 -884 18234 492
rect 18360 -884 18370 492
rect 18422 -884 18432 492
rect 18558 -884 18568 492
rect 18620 -884 18630 492
rect 18756 -884 18766 492
rect 18818 -884 18828 492
rect 18954 -884 18964 492
rect 19016 -884 19026 492
rect 19152 -884 19162 492
rect 19214 -884 19224 492
rect 19350 -884 19360 492
rect 19412 -884 19422 492
rect 19548 -884 19558 492
rect 19610 -884 19620 492
rect 19746 -883 19756 493
rect 19808 -883 19818 493
rect 19892 -743 20046 545
rect 19892 -877 19902 -743
rect 20036 -877 20046 -743
rect 19759 -884 19765 -883
rect 19799 -884 19805 -883
rect 11443 -896 11489 -884
rect 11641 -896 11687 -884
rect 11839 -896 11885 -884
rect 12037 -896 12083 -884
rect 12235 -896 12281 -884
rect 12433 -896 12479 -884
rect 12631 -896 12677 -884
rect 12829 -896 12875 -884
rect 13027 -896 13073 -884
rect 13225 -896 13271 -884
rect 13423 -896 13469 -884
rect 13621 -896 13667 -884
rect 13819 -896 13865 -884
rect 14017 -896 14063 -884
rect 14215 -896 14261 -884
rect 14413 -896 14459 -884
rect 14611 -896 14657 -884
rect 14809 -896 14855 -884
rect 15007 -896 15053 -884
rect 15205 -896 15251 -884
rect 15403 -896 15449 -884
rect 15601 -896 15647 -884
rect 15799 -896 15845 -884
rect 15997 -896 16043 -884
rect 16195 -896 16241 -884
rect 16393 -896 16439 -884
rect 16591 -896 16637 -884
rect 16789 -896 16835 -884
rect 16987 -896 17033 -884
rect 17185 -896 17231 -884
rect 17383 -896 17429 -884
rect 17581 -896 17627 -884
rect 17779 -896 17825 -884
rect 17977 -896 18023 -884
rect 18175 -896 18221 -884
rect 18373 -896 18419 -884
rect 18571 -896 18617 -884
rect 18769 -896 18815 -884
rect 18967 -896 19013 -884
rect 19165 -896 19211 -884
rect 19363 -896 19409 -884
rect 19561 -896 19607 -884
rect 19759 -896 19805 -884
rect 19892 -937 20046 -877
rect 11202 -943 20046 -937
rect 11202 -947 11511 -943
rect 11202 -1081 11212 -947
rect 11346 -977 11511 -947
rect 11619 -977 11709 -943
rect 11817 -977 11907 -943
rect 12015 -977 12105 -943
rect 12213 -977 12303 -943
rect 12411 -977 12501 -943
rect 12609 -977 12699 -943
rect 12807 -977 12897 -943
rect 13005 -977 13095 -943
rect 13203 -977 13293 -943
rect 13401 -977 13491 -943
rect 13599 -977 13689 -943
rect 13797 -977 13887 -943
rect 13995 -977 14085 -943
rect 14193 -977 14283 -943
rect 14391 -977 14481 -943
rect 14589 -977 14679 -943
rect 14787 -977 14877 -943
rect 14985 -977 15075 -943
rect 15183 -977 15273 -943
rect 15381 -977 15471 -943
rect 15579 -977 15669 -943
rect 15777 -977 15867 -943
rect 15975 -977 16065 -943
rect 16173 -977 16263 -943
rect 16371 -977 16461 -943
rect 16569 -977 16659 -943
rect 16767 -977 16857 -943
rect 16965 -977 17055 -943
rect 17163 -977 17253 -943
rect 17361 -977 17451 -943
rect 17559 -977 17649 -943
rect 17757 -977 17847 -943
rect 17955 -977 18045 -943
rect 18153 -977 18243 -943
rect 18351 -977 18441 -943
rect 18549 -977 18639 -943
rect 18747 -977 18837 -943
rect 18945 -977 19035 -943
rect 19143 -977 19233 -943
rect 19341 -977 19431 -943
rect 19539 -977 19629 -943
rect 19737 -947 20046 -943
rect 19737 -977 19902 -947
rect 11346 -1051 19902 -977
rect 11346 -1081 11511 -1051
rect 11202 -1085 11511 -1081
rect 11619 -1085 11709 -1051
rect 11817 -1085 11907 -1051
rect 12015 -1085 12105 -1051
rect 12213 -1085 12303 -1051
rect 12411 -1085 12501 -1051
rect 12609 -1085 12699 -1051
rect 12807 -1085 12897 -1051
rect 13005 -1085 13095 -1051
rect 13203 -1085 13293 -1051
rect 13401 -1085 13491 -1051
rect 13599 -1085 13689 -1051
rect 13797 -1085 13887 -1051
rect 13995 -1085 14085 -1051
rect 14193 -1085 14283 -1051
rect 14391 -1085 14481 -1051
rect 14589 -1085 14679 -1051
rect 14787 -1085 14877 -1051
rect 14985 -1085 15075 -1051
rect 15183 -1085 15273 -1051
rect 15381 -1085 15471 -1051
rect 15579 -1085 15669 -1051
rect 15777 -1085 15867 -1051
rect 15975 -1085 16065 -1051
rect 16173 -1085 16263 -1051
rect 16371 -1085 16461 -1051
rect 16569 -1085 16659 -1051
rect 16767 -1085 16857 -1051
rect 16965 -1085 17055 -1051
rect 17163 -1085 17253 -1051
rect 17361 -1085 17451 -1051
rect 17559 -1085 17649 -1051
rect 17757 -1085 17847 -1051
rect 17955 -1085 18045 -1051
rect 18153 -1085 18243 -1051
rect 18351 -1085 18441 -1051
rect 18549 -1085 18639 -1051
rect 18747 -1085 18837 -1051
rect 18945 -1085 19035 -1051
rect 19143 -1085 19233 -1051
rect 19341 -1085 19431 -1051
rect 19539 -1085 19629 -1051
rect 19737 -1081 19902 -1051
rect 20036 -1081 20046 -947
rect 19737 -1085 20046 -1081
rect 11202 -1091 20046 -1085
rect 11202 -1151 11356 -1091
rect 11443 -1144 11489 -1132
rect 11641 -1144 11687 -1132
rect 11839 -1144 11885 -1132
rect 12037 -1144 12083 -1132
rect 12235 -1144 12281 -1132
rect 12433 -1144 12479 -1132
rect 12631 -1144 12677 -1132
rect 12829 -1144 12875 -1132
rect 13027 -1144 13073 -1132
rect 13225 -1144 13271 -1132
rect 13423 -1144 13469 -1132
rect 13621 -1144 13667 -1132
rect 13819 -1144 13865 -1132
rect 14017 -1144 14063 -1132
rect 14215 -1144 14261 -1132
rect 14413 -1144 14459 -1132
rect 14611 -1144 14657 -1132
rect 14809 -1144 14855 -1132
rect 15007 -1144 15053 -1132
rect 15205 -1144 15251 -1132
rect 15403 -1144 15449 -1132
rect 15601 -1144 15647 -1132
rect 15799 -1144 15845 -1132
rect 15997 -1144 16043 -1132
rect 16195 -1144 16241 -1132
rect 16393 -1144 16439 -1132
rect 16591 -1144 16637 -1132
rect 16789 -1144 16835 -1132
rect 16987 -1144 17033 -1132
rect 17185 -1144 17231 -1132
rect 17383 -1144 17429 -1132
rect 17581 -1144 17627 -1132
rect 17779 -1144 17825 -1132
rect 17977 -1144 18023 -1132
rect 18175 -1144 18221 -1132
rect 18373 -1144 18419 -1132
rect 18571 -1144 18617 -1132
rect 18769 -1144 18815 -1132
rect 18967 -1144 19013 -1132
rect 19165 -1144 19211 -1132
rect 19363 -1144 19409 -1132
rect 19561 -1144 19607 -1132
rect 19759 -1143 19805 -1132
rect 11202 -1285 11212 -1151
rect 11346 -1285 11356 -1151
rect 11202 -2573 11356 -1285
rect 11430 -2520 11440 -1144
rect 11492 -2520 11502 -1144
rect 11628 -2520 11638 -1144
rect 11690 -2520 11700 -1144
rect 11826 -2520 11836 -1144
rect 11888 -2520 11898 -1144
rect 12024 -2520 12034 -1144
rect 12086 -2520 12096 -1144
rect 12222 -2520 12232 -1144
rect 12284 -2520 12294 -1144
rect 12420 -2520 12430 -1144
rect 12482 -2520 12492 -1144
rect 12618 -2520 12628 -1144
rect 12680 -2520 12690 -1144
rect 12816 -2520 12826 -1144
rect 12878 -2520 12888 -1144
rect 13014 -2520 13024 -1144
rect 13076 -2520 13086 -1144
rect 13212 -2520 13222 -1144
rect 13274 -2520 13284 -1144
rect 13410 -2520 13420 -1144
rect 13472 -2520 13482 -1144
rect 13608 -2520 13618 -1144
rect 13670 -2520 13680 -1144
rect 13806 -2520 13816 -1144
rect 13868 -2520 13878 -1144
rect 14004 -2520 14014 -1144
rect 14066 -2520 14076 -1144
rect 14202 -2520 14212 -1144
rect 14264 -2520 14274 -1144
rect 14400 -2520 14410 -1144
rect 14462 -2520 14472 -1144
rect 14598 -2520 14608 -1144
rect 14660 -2520 14670 -1144
rect 14796 -2520 14806 -1144
rect 14858 -2520 14868 -1144
rect 14994 -2520 15004 -1144
rect 15056 -2520 15066 -1144
rect 15192 -2520 15202 -1144
rect 15254 -2520 15264 -1144
rect 15390 -2520 15400 -1144
rect 15452 -2520 15462 -1144
rect 15588 -2520 15598 -1144
rect 15650 -2520 15660 -1144
rect 15786 -2520 15796 -1144
rect 15848 -2520 15858 -1144
rect 15984 -2520 15994 -1144
rect 16046 -2520 16056 -1144
rect 16182 -2520 16192 -1144
rect 16244 -2520 16254 -1144
rect 16380 -2520 16390 -1144
rect 16442 -2520 16452 -1144
rect 16578 -2520 16588 -1144
rect 16640 -2520 16650 -1144
rect 16776 -2520 16786 -1144
rect 16838 -2520 16848 -1144
rect 16974 -2520 16984 -1144
rect 17036 -2520 17046 -1144
rect 17172 -2520 17182 -1144
rect 17234 -2520 17244 -1144
rect 17370 -2520 17380 -1144
rect 17432 -2520 17442 -1144
rect 17568 -2520 17578 -1144
rect 17630 -2520 17640 -1144
rect 17766 -2520 17776 -1144
rect 17828 -2520 17838 -1144
rect 17964 -2520 17974 -1144
rect 18026 -2520 18036 -1144
rect 18162 -2520 18172 -1144
rect 18224 -2520 18234 -1144
rect 18360 -2520 18370 -1144
rect 18422 -2520 18432 -1144
rect 18558 -2520 18568 -1144
rect 18620 -2520 18630 -1144
rect 18756 -2520 18766 -1144
rect 18818 -2520 18828 -1144
rect 18954 -2520 18964 -1144
rect 19016 -2520 19026 -1144
rect 19152 -2520 19162 -1144
rect 19214 -2520 19224 -1144
rect 19350 -2520 19360 -1144
rect 19412 -2520 19422 -1144
rect 19548 -2520 19558 -1144
rect 19610 -2520 19620 -1144
rect 19746 -2519 19756 -1143
rect 19808 -2519 19818 -1143
rect 19892 -1151 20046 -1091
rect 19892 -1285 19902 -1151
rect 20036 -1285 20046 -1151
rect 19759 -2520 19765 -2519
rect 19799 -2520 19805 -2519
rect 11443 -2532 11489 -2520
rect 11641 -2532 11687 -2520
rect 11839 -2532 11885 -2520
rect 12037 -2532 12083 -2520
rect 12235 -2532 12281 -2520
rect 12433 -2532 12479 -2520
rect 12631 -2532 12677 -2520
rect 12829 -2532 12875 -2520
rect 13027 -2532 13073 -2520
rect 13225 -2532 13271 -2520
rect 13423 -2532 13469 -2520
rect 13621 -2532 13667 -2520
rect 13819 -2532 13865 -2520
rect 14017 -2532 14063 -2520
rect 14215 -2532 14261 -2520
rect 14413 -2532 14459 -2520
rect 14611 -2532 14657 -2520
rect 14809 -2532 14855 -2520
rect 15007 -2532 15053 -2520
rect 15205 -2532 15251 -2520
rect 15403 -2532 15449 -2520
rect 15601 -2532 15647 -2520
rect 15799 -2532 15845 -2520
rect 15997 -2532 16043 -2520
rect 16195 -2532 16241 -2520
rect 16393 -2532 16439 -2520
rect 16591 -2532 16637 -2520
rect 16789 -2532 16835 -2520
rect 16987 -2532 17033 -2520
rect 17185 -2532 17231 -2520
rect 17383 -2532 17429 -2520
rect 17581 -2532 17627 -2520
rect 17779 -2532 17825 -2520
rect 17977 -2532 18023 -2520
rect 18175 -2532 18221 -2520
rect 18373 -2532 18419 -2520
rect 18571 -2532 18617 -2520
rect 18769 -2532 18815 -2520
rect 18967 -2532 19013 -2520
rect 19165 -2532 19211 -2520
rect 19363 -2532 19409 -2520
rect 19561 -2532 19607 -2520
rect 19759 -2532 19805 -2520
rect 19892 -2573 20046 -1285
rect 11202 -2579 20046 -2573
rect 11202 -2613 11511 -2579
rect 11619 -2613 11709 -2579
rect 11817 -2613 11907 -2579
rect 12015 -2613 12105 -2579
rect 12213 -2613 12303 -2579
rect 12411 -2613 12501 -2579
rect 12609 -2613 12699 -2579
rect 12807 -2613 12897 -2579
rect 13005 -2613 13095 -2579
rect 13203 -2613 13293 -2579
rect 13401 -2613 13491 -2579
rect 13599 -2613 13689 -2579
rect 13797 -2613 13887 -2579
rect 13995 -2613 14085 -2579
rect 14193 -2613 14283 -2579
rect 14391 -2613 14481 -2579
rect 14589 -2613 14679 -2579
rect 14787 -2613 14877 -2579
rect 14985 -2613 15075 -2579
rect 15183 -2613 15273 -2579
rect 15381 -2613 15471 -2579
rect 15579 -2613 15669 -2579
rect 15777 -2613 15867 -2579
rect 15975 -2613 16065 -2579
rect 16173 -2613 16263 -2579
rect 16371 -2613 16461 -2579
rect 16569 -2613 16659 -2579
rect 16767 -2613 16857 -2579
rect 16965 -2613 17055 -2579
rect 17163 -2613 17253 -2579
rect 17361 -2613 17451 -2579
rect 17559 -2613 17649 -2579
rect 17757 -2613 17847 -2579
rect 17955 -2613 18045 -2579
rect 18153 -2613 18243 -2579
rect 18351 -2613 18441 -2579
rect 18549 -2613 18639 -2579
rect 18747 -2613 18837 -2579
rect 18945 -2613 19035 -2579
rect 19143 -2613 19233 -2579
rect 19341 -2613 19431 -2579
rect 19539 -2613 19629 -2579
rect 19737 -2613 20046 -2579
rect 11202 -2643 20046 -2613
rect 11202 -3208 11356 -2643
rect 19892 -3208 20046 -2643
rect 11202 -3252 20046 -3208
rect 11202 -3286 11511 -3252
rect 11619 -3286 11709 -3252
rect 11817 -3286 11907 -3252
rect 12015 -3286 12105 -3252
rect 12213 -3286 12303 -3252
rect 12411 -3286 12501 -3252
rect 12609 -3286 12699 -3252
rect 12807 -3286 12897 -3252
rect 13005 -3286 13095 -3252
rect 13203 -3286 13293 -3252
rect 13401 -3286 13491 -3252
rect 13599 -3286 13689 -3252
rect 13797 -3286 13887 -3252
rect 13995 -3286 14085 -3252
rect 14193 -3286 14283 -3252
rect 14391 -3286 14481 -3252
rect 14589 -3286 14679 -3252
rect 14787 -3286 14877 -3252
rect 14985 -3286 15075 -3252
rect 15183 -3286 15273 -3252
rect 15381 -3286 15471 -3252
rect 15579 -3286 15669 -3252
rect 15777 -3286 15867 -3252
rect 15975 -3286 16065 -3252
rect 16173 -3286 16263 -3252
rect 16371 -3286 16461 -3252
rect 16569 -3286 16659 -3252
rect 16767 -3286 16857 -3252
rect 16965 -3286 17055 -3252
rect 17163 -3286 17253 -3252
rect 17361 -3286 17451 -3252
rect 17559 -3286 17649 -3252
rect 17757 -3286 17847 -3252
rect 17955 -3286 18045 -3252
rect 18153 -3286 18243 -3252
rect 18351 -3286 18441 -3252
rect 18549 -3286 18639 -3252
rect 18747 -3286 18837 -3252
rect 18945 -3286 19035 -3252
rect 19143 -3286 19233 -3252
rect 19341 -3286 19431 -3252
rect 19539 -3286 19629 -3252
rect 19737 -3286 20046 -3252
rect 11202 -3292 20046 -3286
rect 11443 -3345 11489 -3333
rect 11641 -3345 11687 -3333
rect 11839 -3345 11885 -3333
rect 12037 -3345 12083 -3333
rect 12235 -3345 12281 -3333
rect 12433 -3345 12479 -3333
rect 12631 -3345 12677 -3333
rect 12829 -3345 12875 -3333
rect 13027 -3345 13073 -3333
rect 13225 -3345 13271 -3333
rect 13423 -3345 13469 -3333
rect 13621 -3345 13667 -3333
rect 13819 -3345 13865 -3333
rect 14017 -3345 14063 -3333
rect 14215 -3345 14261 -3333
rect 14413 -3345 14459 -3333
rect 14611 -3345 14657 -3333
rect 14809 -3345 14855 -3333
rect 15007 -3345 15053 -3333
rect 15205 -3345 15251 -3333
rect 15403 -3345 15449 -3333
rect 15601 -3345 15647 -3333
rect 15799 -3345 15845 -3333
rect 15997 -3345 16043 -3333
rect 16195 -3345 16241 -3333
rect 16393 -3345 16439 -3333
rect 16591 -3345 16637 -3333
rect 16789 -3345 16835 -3333
rect 16987 -3345 17033 -3333
rect 17185 -3345 17231 -3333
rect 17383 -3345 17429 -3333
rect 17581 -3345 17627 -3333
rect 17779 -3345 17825 -3333
rect 17977 -3345 18023 -3333
rect 18175 -3345 18221 -3333
rect 18373 -3345 18419 -3333
rect 18571 -3345 18617 -3333
rect 18769 -3345 18815 -3333
rect 18967 -3345 19013 -3333
rect 19165 -3345 19211 -3333
rect 19363 -3345 19409 -3333
rect 19561 -3345 19607 -3333
rect 19759 -3344 19805 -3333
rect 11430 -4721 11440 -3345
rect 11492 -4721 11502 -3345
rect 11628 -4721 11638 -3345
rect 11690 -4721 11700 -3345
rect 11826 -4721 11836 -3345
rect 11888 -4721 11898 -3345
rect 12024 -4721 12034 -3345
rect 12086 -4721 12096 -3345
rect 12222 -4721 12232 -3345
rect 12284 -4721 12294 -3345
rect 12420 -4721 12430 -3345
rect 12482 -4721 12492 -3345
rect 12618 -4721 12628 -3345
rect 12680 -4721 12690 -3345
rect 12816 -4721 12826 -3345
rect 12878 -4721 12888 -3345
rect 13014 -4721 13024 -3345
rect 13076 -4721 13086 -3345
rect 13212 -4721 13222 -3345
rect 13274 -4721 13284 -3345
rect 13410 -4721 13420 -3345
rect 13472 -4721 13482 -3345
rect 13608 -4721 13618 -3345
rect 13670 -4721 13680 -3345
rect 13806 -4721 13816 -3345
rect 13868 -4721 13878 -3345
rect 14004 -4721 14014 -3345
rect 14066 -4721 14076 -3345
rect 14202 -4721 14212 -3345
rect 14264 -4721 14274 -3345
rect 14400 -4721 14410 -3345
rect 14462 -4721 14472 -3345
rect 14598 -4721 14608 -3345
rect 14660 -4721 14670 -3345
rect 14796 -4721 14806 -3345
rect 14858 -4721 14868 -3345
rect 14994 -4721 15004 -3345
rect 15056 -4721 15066 -3345
rect 15192 -4721 15202 -3345
rect 15254 -4721 15264 -3345
rect 15390 -4721 15400 -3345
rect 15452 -4721 15462 -3345
rect 15588 -4721 15598 -3345
rect 15650 -4721 15660 -3345
rect 15786 -4721 15796 -3345
rect 15848 -4721 15858 -3345
rect 15984 -4721 15994 -3345
rect 16046 -4721 16056 -3345
rect 16182 -4721 16192 -3345
rect 16244 -4721 16254 -3345
rect 16380 -4721 16390 -3345
rect 16442 -4721 16452 -3345
rect 16578 -4721 16588 -3345
rect 16640 -4721 16650 -3345
rect 16776 -4721 16786 -3345
rect 16838 -4721 16848 -3345
rect 16974 -4721 16984 -3345
rect 17036 -4721 17046 -3345
rect 17172 -4721 17182 -3345
rect 17234 -4721 17244 -3345
rect 17370 -4721 17380 -3345
rect 17432 -4721 17442 -3345
rect 17568 -4721 17578 -3345
rect 17630 -4721 17640 -3345
rect 17766 -4721 17776 -3345
rect 17828 -4721 17838 -3345
rect 17964 -4721 17974 -3345
rect 18026 -4721 18036 -3345
rect 18162 -4721 18172 -3345
rect 18224 -4721 18234 -3345
rect 18360 -4721 18370 -3345
rect 18422 -4721 18432 -3345
rect 18558 -4721 18568 -3345
rect 18620 -4721 18630 -3345
rect 18756 -4721 18766 -3345
rect 18818 -4721 18828 -3345
rect 18954 -4721 18964 -3345
rect 19016 -4721 19026 -3345
rect 19152 -4721 19162 -3345
rect 19214 -4721 19224 -3345
rect 19350 -4721 19360 -3345
rect 19412 -4721 19422 -3345
rect 19548 -4721 19558 -3345
rect 19610 -4721 19620 -3345
rect 19746 -4720 19756 -3344
rect 19808 -4720 19818 -3344
rect 19759 -4721 19765 -4720
rect 19799 -4721 19805 -4720
rect 11443 -5127 11489 -4721
rect 11641 -4733 11687 -4721
rect 11839 -5127 11885 -4721
rect 12037 -4733 12083 -4721
rect 12235 -5127 12281 -4721
rect 12433 -4733 12479 -4721
rect 12631 -5127 12677 -4721
rect 12829 -4733 12875 -4721
rect 13027 -5127 13073 -4721
rect 13225 -4733 13271 -4721
rect 13423 -5127 13469 -4721
rect 13621 -4733 13667 -4721
rect 13819 -5127 13865 -4721
rect 14017 -4733 14063 -4721
rect 14215 -5127 14261 -4721
rect 14413 -4733 14459 -4721
rect 14611 -5127 14657 -4721
rect 14809 -4733 14855 -4721
rect 15007 -5127 15053 -4721
rect 15205 -4733 15251 -4721
rect 15403 -5127 15449 -4721
rect 15601 -4733 15647 -4721
rect 15799 -5127 15845 -4721
rect 15997 -4733 16043 -4721
rect 16195 -5127 16241 -4721
rect 16393 -4733 16439 -4721
rect 16591 -5127 16637 -4721
rect 16789 -4733 16835 -4721
rect 16987 -5127 17033 -4721
rect 17185 -4733 17231 -4721
rect 17383 -5127 17429 -4721
rect 17581 -4733 17627 -4721
rect 17779 -5127 17825 -4721
rect 17977 -4733 18023 -4721
rect 18175 -5127 18221 -4721
rect 18373 -4733 18419 -4721
rect 18571 -5127 18617 -4721
rect 18769 -4733 18815 -4721
rect 18967 -5127 19013 -4721
rect 19165 -4733 19211 -4721
rect 19363 -5127 19409 -4721
rect 19561 -4733 19607 -4721
rect 19759 -5127 19805 -4721
rect 20976 -5127 22196 2237
rect 23293 2128 23339 2327
rect 23491 2128 23537 2140
rect 23689 2128 23735 2327
rect 23887 2128 23933 2140
rect 24085 2128 24131 2327
rect 24283 2128 24329 2140
rect 24481 2128 24527 2327
rect 24679 2128 24725 2140
rect 24877 2128 24923 2327
rect 25075 2128 25121 2140
rect 25273 2128 25319 2327
rect 25471 2128 25517 2140
rect 25669 2128 25715 2327
rect 25867 2128 25913 2140
rect 26065 2128 26111 2327
rect 26263 2128 26309 2140
rect 26461 2128 26507 2327
rect 26659 2128 26705 2140
rect 26857 2128 26903 2327
rect 27055 2128 27101 2140
rect 27253 2128 27299 2327
rect 27451 2128 27497 2140
rect 27649 2128 27695 2327
rect 27847 2128 27893 2140
rect 28045 2128 28091 2327
rect 28243 2128 28289 2140
rect 28441 2128 28487 2327
rect 28639 2128 28685 2140
rect 28837 2128 28883 2327
rect 29035 2128 29081 2140
rect 29233 2128 29279 2327
rect 29431 2128 29477 2140
rect 29629 2128 29675 2327
rect 29827 2128 29873 2140
rect 30025 2128 30071 2327
rect 30223 2128 30269 2140
rect 30421 2128 30467 2327
rect 30619 2128 30665 2140
rect 30817 2128 30863 2327
rect 31015 2128 31061 2140
rect 31213 2128 31259 2327
rect 31411 2128 31457 2140
rect 31609 2129 31655 2327
rect 23280 752 23290 2128
rect 23342 752 23352 2128
rect 23478 752 23488 2128
rect 23540 752 23550 2128
rect 23676 752 23686 2128
rect 23738 752 23748 2128
rect 23874 752 23884 2128
rect 23936 752 23946 2128
rect 24072 752 24082 2128
rect 24134 752 24144 2128
rect 24270 752 24280 2128
rect 24332 752 24342 2128
rect 24468 752 24478 2128
rect 24530 752 24540 2128
rect 24666 752 24676 2128
rect 24728 752 24738 2128
rect 24864 752 24874 2128
rect 24926 752 24936 2128
rect 25062 752 25072 2128
rect 25124 752 25134 2128
rect 25260 752 25270 2128
rect 25322 752 25332 2128
rect 25458 752 25468 2128
rect 25520 752 25530 2128
rect 25656 752 25666 2128
rect 25718 752 25728 2128
rect 25854 752 25864 2128
rect 25916 752 25926 2128
rect 26052 752 26062 2128
rect 26114 752 26124 2128
rect 26250 752 26260 2128
rect 26312 752 26322 2128
rect 26448 752 26458 2128
rect 26510 752 26520 2128
rect 26646 752 26656 2128
rect 26708 752 26718 2128
rect 26844 752 26854 2128
rect 26906 752 26916 2128
rect 27042 752 27052 2128
rect 27104 752 27114 2128
rect 27240 752 27250 2128
rect 27302 752 27312 2128
rect 27438 752 27448 2128
rect 27500 752 27510 2128
rect 27636 752 27646 2128
rect 27698 752 27708 2128
rect 27834 752 27844 2128
rect 27896 752 27906 2128
rect 28032 752 28042 2128
rect 28094 752 28104 2128
rect 28230 752 28240 2128
rect 28292 752 28302 2128
rect 28428 752 28438 2128
rect 28490 752 28500 2128
rect 28626 752 28636 2128
rect 28688 752 28698 2128
rect 28824 752 28834 2128
rect 28886 752 28896 2128
rect 29022 752 29032 2128
rect 29084 752 29094 2128
rect 29220 752 29230 2128
rect 29282 752 29292 2128
rect 29418 752 29428 2128
rect 29480 752 29490 2128
rect 29616 752 29626 2128
rect 29678 752 29688 2128
rect 29814 752 29824 2128
rect 29876 752 29886 2128
rect 30012 752 30022 2128
rect 30074 752 30084 2128
rect 30210 752 30220 2128
rect 30272 752 30282 2128
rect 30408 752 30418 2128
rect 30470 752 30480 2128
rect 30606 752 30616 2128
rect 30668 752 30678 2128
rect 30804 752 30814 2128
rect 30866 752 30876 2128
rect 31002 752 31012 2128
rect 31064 752 31074 2128
rect 31200 752 31210 2128
rect 31262 752 31272 2128
rect 31398 752 31408 2128
rect 31460 752 31470 2128
rect 31596 753 31606 2129
rect 31658 753 31668 2129
rect 31609 752 31615 753
rect 31649 752 31655 753
rect 23293 740 23339 752
rect 23491 740 23537 752
rect 23689 740 23735 752
rect 23887 740 23933 752
rect 24085 740 24131 752
rect 24283 740 24329 752
rect 24481 740 24527 752
rect 24679 740 24725 752
rect 24877 740 24923 752
rect 25075 740 25121 752
rect 25273 740 25319 752
rect 25471 740 25517 752
rect 25669 740 25715 752
rect 25867 740 25913 752
rect 26065 740 26111 752
rect 26263 740 26309 752
rect 26461 740 26507 752
rect 26659 740 26705 752
rect 26857 740 26903 752
rect 27055 740 27101 752
rect 27253 740 27299 752
rect 27451 740 27497 752
rect 27649 740 27695 752
rect 27847 740 27893 752
rect 28045 740 28091 752
rect 28243 740 28289 752
rect 28441 740 28487 752
rect 28639 740 28685 752
rect 28837 740 28883 752
rect 29035 740 29081 752
rect 29233 740 29279 752
rect 29431 740 29477 752
rect 29629 740 29675 752
rect 29827 740 29873 752
rect 30025 740 30071 752
rect 30223 740 30269 752
rect 30421 740 30467 752
rect 30619 740 30665 752
rect 30817 740 30863 752
rect 31015 740 31061 752
rect 31213 740 31259 752
rect 31411 740 31457 752
rect 31609 740 31655 752
rect 23052 693 31896 699
rect 23052 659 23361 693
rect 23469 659 23559 693
rect 23667 659 23757 693
rect 23865 659 23955 693
rect 24063 659 24153 693
rect 24261 659 24351 693
rect 24459 659 24549 693
rect 24657 659 24747 693
rect 24855 659 24945 693
rect 25053 659 25143 693
rect 25251 659 25341 693
rect 25449 659 25539 693
rect 25647 659 25737 693
rect 25845 659 25935 693
rect 26043 659 26133 693
rect 26241 659 26331 693
rect 26439 659 26529 693
rect 26637 659 26727 693
rect 26835 659 26925 693
rect 27033 659 27123 693
rect 27231 659 27321 693
rect 27429 659 27519 693
rect 27627 659 27717 693
rect 27825 659 27915 693
rect 28023 659 28113 693
rect 28221 659 28311 693
rect 28419 659 28509 693
rect 28617 659 28707 693
rect 28815 659 28905 693
rect 29013 659 29103 693
rect 29211 659 29301 693
rect 29409 659 29499 693
rect 29607 659 29697 693
rect 29805 659 29895 693
rect 30003 659 30093 693
rect 30201 659 30291 693
rect 30399 659 30489 693
rect 30597 659 30687 693
rect 30795 659 30885 693
rect 30993 659 31083 693
rect 31191 659 31281 693
rect 31389 659 31479 693
rect 31587 659 31896 693
rect 23052 585 31896 659
rect 23052 551 23361 585
rect 23469 551 23559 585
rect 23667 551 23757 585
rect 23865 551 23955 585
rect 24063 551 24153 585
rect 24261 551 24351 585
rect 24459 551 24549 585
rect 24657 551 24747 585
rect 24855 551 24945 585
rect 25053 551 25143 585
rect 25251 551 25341 585
rect 25449 551 25539 585
rect 25647 551 25737 585
rect 25845 551 25935 585
rect 26043 551 26133 585
rect 26241 551 26331 585
rect 26439 551 26529 585
rect 26637 551 26727 585
rect 26835 551 26925 585
rect 27033 551 27123 585
rect 27231 551 27321 585
rect 27429 551 27519 585
rect 27627 551 27717 585
rect 27825 551 27915 585
rect 28023 551 28113 585
rect 28221 551 28311 585
rect 28419 551 28509 585
rect 28617 551 28707 585
rect 28815 551 28905 585
rect 29013 551 29103 585
rect 29211 551 29301 585
rect 29409 551 29499 585
rect 29607 551 29697 585
rect 29805 551 29895 585
rect 30003 551 30093 585
rect 30201 551 30291 585
rect 30399 551 30489 585
rect 30597 551 30687 585
rect 30795 551 30885 585
rect 30993 551 31083 585
rect 31191 551 31281 585
rect 31389 551 31479 585
rect 31587 551 31896 585
rect 23052 545 31896 551
rect 23052 -743 23206 545
rect 23293 492 23339 504
rect 23491 492 23537 504
rect 23689 492 23735 504
rect 23887 492 23933 504
rect 24085 492 24131 504
rect 24283 492 24329 504
rect 24481 492 24527 504
rect 24679 492 24725 504
rect 24877 492 24923 504
rect 25075 492 25121 504
rect 25273 492 25319 504
rect 25471 492 25517 504
rect 25669 492 25715 504
rect 25867 492 25913 504
rect 26065 492 26111 504
rect 26263 492 26309 504
rect 26461 492 26507 504
rect 26659 492 26705 504
rect 26857 492 26903 504
rect 27055 492 27101 504
rect 27253 492 27299 504
rect 27451 492 27497 504
rect 27649 492 27695 504
rect 27847 492 27893 504
rect 28045 492 28091 504
rect 28243 492 28289 504
rect 28441 492 28487 504
rect 28639 492 28685 504
rect 28837 492 28883 504
rect 29035 492 29081 504
rect 29233 492 29279 504
rect 29431 492 29477 504
rect 29629 492 29675 504
rect 29827 492 29873 504
rect 30025 492 30071 504
rect 30223 492 30269 504
rect 30421 492 30467 504
rect 30619 492 30665 504
rect 30817 492 30863 504
rect 31015 492 31061 504
rect 31213 492 31259 504
rect 31411 492 31457 504
rect 31609 493 31655 504
rect 23052 -877 23062 -743
rect 23196 -877 23206 -743
rect 23052 -937 23206 -877
rect 23280 -884 23290 492
rect 23342 -884 23352 492
rect 23478 -884 23488 492
rect 23540 -884 23550 492
rect 23676 -884 23686 492
rect 23738 -884 23748 492
rect 23874 -884 23884 492
rect 23936 -884 23946 492
rect 24072 -884 24082 492
rect 24134 -884 24144 492
rect 24270 -884 24280 492
rect 24332 -884 24342 492
rect 24468 -884 24478 492
rect 24530 -884 24540 492
rect 24666 -884 24676 492
rect 24728 -884 24738 492
rect 24864 -884 24874 492
rect 24926 -884 24936 492
rect 25062 -884 25072 492
rect 25124 -884 25134 492
rect 25260 -884 25270 492
rect 25322 -884 25332 492
rect 25458 -884 25468 492
rect 25520 -884 25530 492
rect 25656 -884 25666 492
rect 25718 -884 25728 492
rect 25854 -884 25864 492
rect 25916 -884 25926 492
rect 26052 -884 26062 492
rect 26114 -884 26124 492
rect 26250 -884 26260 492
rect 26312 -884 26322 492
rect 26448 -884 26458 492
rect 26510 -884 26520 492
rect 26646 -884 26656 492
rect 26708 -884 26718 492
rect 26844 -884 26854 492
rect 26906 -884 26916 492
rect 27042 -884 27052 492
rect 27104 -884 27114 492
rect 27240 -884 27250 492
rect 27302 -884 27312 492
rect 27438 -884 27448 492
rect 27500 -884 27510 492
rect 27636 -884 27646 492
rect 27698 -884 27708 492
rect 27834 -884 27844 492
rect 27896 -884 27906 492
rect 28032 -884 28042 492
rect 28094 -884 28104 492
rect 28230 -884 28240 492
rect 28292 -884 28302 492
rect 28428 -884 28438 492
rect 28490 -884 28500 492
rect 28626 -884 28636 492
rect 28688 -884 28698 492
rect 28824 -884 28834 492
rect 28886 -884 28896 492
rect 29022 -884 29032 492
rect 29084 -884 29094 492
rect 29220 -884 29230 492
rect 29282 -884 29292 492
rect 29418 -884 29428 492
rect 29480 -884 29490 492
rect 29616 -884 29626 492
rect 29678 -884 29688 492
rect 29814 -884 29824 492
rect 29876 -884 29886 492
rect 30012 -884 30022 492
rect 30074 -884 30084 492
rect 30210 -884 30220 492
rect 30272 -884 30282 492
rect 30408 -884 30418 492
rect 30470 -884 30480 492
rect 30606 -884 30616 492
rect 30668 -884 30678 492
rect 30804 -884 30814 492
rect 30866 -884 30876 492
rect 31002 -884 31012 492
rect 31064 -884 31074 492
rect 31200 -884 31210 492
rect 31262 -884 31272 492
rect 31398 -884 31408 492
rect 31460 -884 31470 492
rect 31596 -883 31606 493
rect 31658 -883 31668 493
rect 31609 -884 31615 -883
rect 31649 -884 31655 -883
rect 23293 -896 23339 -884
rect 23491 -896 23537 -884
rect 23689 -896 23735 -884
rect 23887 -896 23933 -884
rect 24085 -896 24131 -884
rect 24283 -896 24329 -884
rect 24481 -896 24527 -884
rect 24679 -896 24725 -884
rect 24877 -896 24923 -884
rect 25075 -896 25121 -884
rect 25273 -896 25319 -884
rect 25471 -896 25517 -884
rect 25669 -896 25715 -884
rect 25867 -896 25913 -884
rect 26065 -896 26111 -884
rect 26263 -896 26309 -884
rect 26461 -896 26507 -884
rect 26659 -896 26705 -884
rect 26857 -896 26903 -884
rect 27055 -896 27101 -884
rect 27253 -896 27299 -884
rect 27451 -896 27497 -884
rect 27649 -896 27695 -884
rect 27847 -896 27893 -884
rect 28045 -896 28091 -884
rect 28243 -896 28289 -884
rect 28441 -896 28487 -884
rect 28639 -896 28685 -884
rect 28837 -896 28883 -884
rect 29035 -896 29081 -884
rect 29233 -896 29279 -884
rect 29431 -896 29477 -884
rect 29629 -896 29675 -884
rect 29827 -896 29873 -884
rect 30025 -896 30071 -884
rect 30223 -896 30269 -884
rect 30421 -896 30467 -884
rect 30619 -896 30665 -884
rect 30817 -896 30863 -884
rect 31015 -896 31061 -884
rect 31213 -896 31259 -884
rect 31411 -896 31457 -884
rect 31609 -896 31655 -884
rect 31742 -937 31896 545
rect 23052 -943 31896 -937
rect 23052 -947 23361 -943
rect 23052 -1081 23062 -947
rect 23196 -977 23361 -947
rect 23469 -977 23559 -943
rect 23667 -977 23757 -943
rect 23865 -977 23955 -943
rect 24063 -977 24153 -943
rect 24261 -977 24351 -943
rect 24459 -977 24549 -943
rect 24657 -977 24747 -943
rect 24855 -977 24945 -943
rect 25053 -977 25143 -943
rect 25251 -977 25341 -943
rect 25449 -977 25539 -943
rect 25647 -977 25737 -943
rect 25845 -977 25935 -943
rect 26043 -977 26133 -943
rect 26241 -977 26331 -943
rect 26439 -977 26529 -943
rect 26637 -977 26727 -943
rect 26835 -977 26925 -943
rect 27033 -977 27123 -943
rect 27231 -977 27321 -943
rect 27429 -977 27519 -943
rect 27627 -977 27717 -943
rect 27825 -977 27915 -943
rect 28023 -977 28113 -943
rect 28221 -977 28311 -943
rect 28419 -977 28509 -943
rect 28617 -977 28707 -943
rect 28815 -977 28905 -943
rect 29013 -977 29103 -943
rect 29211 -977 29301 -943
rect 29409 -977 29499 -943
rect 29607 -977 29697 -943
rect 29805 -977 29895 -943
rect 30003 -977 30093 -943
rect 30201 -977 30291 -943
rect 30399 -977 30489 -943
rect 30597 -977 30687 -943
rect 30795 -977 30885 -943
rect 30993 -977 31083 -943
rect 31191 -977 31281 -943
rect 31389 -977 31479 -943
rect 31587 -977 31896 -943
rect 23196 -1051 31896 -977
rect 23196 -1081 23361 -1051
rect 23052 -1085 23361 -1081
rect 23469 -1085 23559 -1051
rect 23667 -1085 23757 -1051
rect 23865 -1085 23955 -1051
rect 24063 -1085 24153 -1051
rect 24261 -1085 24351 -1051
rect 24459 -1085 24549 -1051
rect 24657 -1085 24747 -1051
rect 24855 -1085 24945 -1051
rect 25053 -1085 25143 -1051
rect 25251 -1085 25341 -1051
rect 25449 -1085 25539 -1051
rect 25647 -1085 25737 -1051
rect 25845 -1085 25935 -1051
rect 26043 -1085 26133 -1051
rect 26241 -1085 26331 -1051
rect 26439 -1085 26529 -1051
rect 26637 -1085 26727 -1051
rect 26835 -1085 26925 -1051
rect 27033 -1085 27123 -1051
rect 27231 -1085 27321 -1051
rect 27429 -1085 27519 -1051
rect 27627 -1085 27717 -1051
rect 27825 -1085 27915 -1051
rect 28023 -1085 28113 -1051
rect 28221 -1085 28311 -1051
rect 28419 -1085 28509 -1051
rect 28617 -1085 28707 -1051
rect 28815 -1085 28905 -1051
rect 29013 -1085 29103 -1051
rect 29211 -1085 29301 -1051
rect 29409 -1085 29499 -1051
rect 29607 -1085 29697 -1051
rect 29805 -1085 29895 -1051
rect 30003 -1085 30093 -1051
rect 30201 -1085 30291 -1051
rect 30399 -1085 30489 -1051
rect 30597 -1085 30687 -1051
rect 30795 -1085 30885 -1051
rect 30993 -1085 31083 -1051
rect 31191 -1085 31281 -1051
rect 31389 -1085 31479 -1051
rect 31587 -1085 31896 -1051
rect 23052 -1091 31896 -1085
rect 23052 -1151 23206 -1091
rect 23293 -1144 23339 -1132
rect 23491 -1144 23537 -1132
rect 23689 -1144 23735 -1132
rect 23887 -1144 23933 -1132
rect 24085 -1144 24131 -1132
rect 24283 -1144 24329 -1132
rect 24481 -1144 24527 -1132
rect 24679 -1144 24725 -1132
rect 24877 -1144 24923 -1132
rect 25075 -1144 25121 -1132
rect 25273 -1144 25319 -1132
rect 25471 -1144 25517 -1132
rect 25669 -1144 25715 -1132
rect 25867 -1144 25913 -1132
rect 26065 -1144 26111 -1132
rect 26263 -1144 26309 -1132
rect 26461 -1144 26507 -1132
rect 26659 -1144 26705 -1132
rect 26857 -1144 26903 -1132
rect 27055 -1144 27101 -1132
rect 27253 -1144 27299 -1132
rect 27451 -1144 27497 -1132
rect 27649 -1144 27695 -1132
rect 27847 -1144 27893 -1132
rect 28045 -1144 28091 -1132
rect 28243 -1144 28289 -1132
rect 28441 -1144 28487 -1132
rect 28639 -1144 28685 -1132
rect 28837 -1144 28883 -1132
rect 29035 -1144 29081 -1132
rect 29233 -1144 29279 -1132
rect 29431 -1144 29477 -1132
rect 29629 -1144 29675 -1132
rect 29827 -1144 29873 -1132
rect 30025 -1144 30071 -1132
rect 30223 -1144 30269 -1132
rect 30421 -1144 30467 -1132
rect 30619 -1144 30665 -1132
rect 30817 -1144 30863 -1132
rect 31015 -1144 31061 -1132
rect 31213 -1144 31259 -1132
rect 31411 -1144 31457 -1132
rect 31609 -1143 31655 -1132
rect 23052 -1285 23062 -1151
rect 23196 -1285 23206 -1151
rect 23052 -2573 23206 -1285
rect 23280 -2520 23290 -1144
rect 23342 -2520 23352 -1144
rect 23478 -2520 23488 -1144
rect 23540 -2520 23550 -1144
rect 23676 -2520 23686 -1144
rect 23738 -2520 23748 -1144
rect 23874 -2520 23884 -1144
rect 23936 -2520 23946 -1144
rect 24072 -2520 24082 -1144
rect 24134 -2520 24144 -1144
rect 24270 -2520 24280 -1144
rect 24332 -2520 24342 -1144
rect 24468 -2520 24478 -1144
rect 24530 -2520 24540 -1144
rect 24666 -2520 24676 -1144
rect 24728 -2520 24738 -1144
rect 24864 -2520 24874 -1144
rect 24926 -2520 24936 -1144
rect 25062 -2520 25072 -1144
rect 25124 -2520 25134 -1144
rect 25260 -2520 25270 -1144
rect 25322 -2520 25332 -1144
rect 25458 -2520 25468 -1144
rect 25520 -2520 25530 -1144
rect 25656 -2520 25666 -1144
rect 25718 -2520 25728 -1144
rect 25854 -2520 25864 -1144
rect 25916 -2520 25926 -1144
rect 26052 -2520 26062 -1144
rect 26114 -2520 26124 -1144
rect 26250 -2520 26260 -1144
rect 26312 -2520 26322 -1144
rect 26448 -2520 26458 -1144
rect 26510 -2520 26520 -1144
rect 26646 -2520 26656 -1144
rect 26708 -2520 26718 -1144
rect 26844 -2520 26854 -1144
rect 26906 -2520 26916 -1144
rect 27042 -2520 27052 -1144
rect 27104 -2520 27114 -1144
rect 27240 -2520 27250 -1144
rect 27302 -2520 27312 -1144
rect 27438 -2520 27448 -1144
rect 27500 -2520 27510 -1144
rect 27636 -2520 27646 -1144
rect 27698 -2520 27708 -1144
rect 27834 -2520 27844 -1144
rect 27896 -2520 27906 -1144
rect 28032 -2520 28042 -1144
rect 28094 -2520 28104 -1144
rect 28230 -2520 28240 -1144
rect 28292 -2520 28302 -1144
rect 28428 -2520 28438 -1144
rect 28490 -2520 28500 -1144
rect 28626 -2520 28636 -1144
rect 28688 -2520 28698 -1144
rect 28824 -2520 28834 -1144
rect 28886 -2520 28896 -1144
rect 29022 -2520 29032 -1144
rect 29084 -2520 29094 -1144
rect 29220 -2520 29230 -1144
rect 29282 -2520 29292 -1144
rect 29418 -2520 29428 -1144
rect 29480 -2520 29490 -1144
rect 29616 -2520 29626 -1144
rect 29678 -2520 29688 -1144
rect 29814 -2520 29824 -1144
rect 29876 -2520 29886 -1144
rect 30012 -2520 30022 -1144
rect 30074 -2520 30084 -1144
rect 30210 -2520 30220 -1144
rect 30272 -2520 30282 -1144
rect 30408 -2520 30418 -1144
rect 30470 -2520 30480 -1144
rect 30606 -2520 30616 -1144
rect 30668 -2520 30678 -1144
rect 30804 -2520 30814 -1144
rect 30866 -2520 30876 -1144
rect 31002 -2520 31012 -1144
rect 31064 -2520 31074 -1144
rect 31200 -2520 31210 -1144
rect 31262 -2520 31272 -1144
rect 31398 -2520 31408 -1144
rect 31460 -2520 31470 -1144
rect 31596 -2519 31606 -1143
rect 31658 -2519 31668 -1143
rect 31609 -2520 31615 -2519
rect 31649 -2520 31655 -2519
rect 23293 -2532 23339 -2520
rect 23491 -2532 23537 -2520
rect 23689 -2532 23735 -2520
rect 23887 -2532 23933 -2520
rect 24085 -2532 24131 -2520
rect 24283 -2532 24329 -2520
rect 24481 -2532 24527 -2520
rect 24679 -2532 24725 -2520
rect 24877 -2532 24923 -2520
rect 25075 -2532 25121 -2520
rect 25273 -2532 25319 -2520
rect 25471 -2532 25517 -2520
rect 25669 -2532 25715 -2520
rect 25867 -2532 25913 -2520
rect 26065 -2532 26111 -2520
rect 26263 -2532 26309 -2520
rect 26461 -2532 26507 -2520
rect 26659 -2532 26705 -2520
rect 26857 -2532 26903 -2520
rect 27055 -2532 27101 -2520
rect 27253 -2532 27299 -2520
rect 27451 -2532 27497 -2520
rect 27649 -2532 27695 -2520
rect 27847 -2532 27893 -2520
rect 28045 -2532 28091 -2520
rect 28243 -2532 28289 -2520
rect 28441 -2532 28487 -2520
rect 28639 -2532 28685 -2520
rect 28837 -2532 28883 -2520
rect 29035 -2532 29081 -2520
rect 29233 -2532 29279 -2520
rect 29431 -2532 29477 -2520
rect 29629 -2532 29675 -2520
rect 29827 -2532 29873 -2520
rect 30025 -2532 30071 -2520
rect 30223 -2532 30269 -2520
rect 30421 -2532 30467 -2520
rect 30619 -2532 30665 -2520
rect 30817 -2532 30863 -2520
rect 31015 -2532 31061 -2520
rect 31213 -2532 31259 -2520
rect 31411 -2532 31457 -2520
rect 31609 -2532 31655 -2520
rect 31742 -2573 31896 -1091
rect 23052 -2579 31896 -2573
rect 23052 -2613 23361 -2579
rect 23469 -2613 23559 -2579
rect 23667 -2613 23757 -2579
rect 23865 -2613 23955 -2579
rect 24063 -2613 24153 -2579
rect 24261 -2613 24351 -2579
rect 24459 -2613 24549 -2579
rect 24657 -2613 24747 -2579
rect 24855 -2613 24945 -2579
rect 25053 -2613 25143 -2579
rect 25251 -2613 25341 -2579
rect 25449 -2613 25539 -2579
rect 25647 -2613 25737 -2579
rect 25845 -2613 25935 -2579
rect 26043 -2613 26133 -2579
rect 26241 -2613 26331 -2579
rect 26439 -2613 26529 -2579
rect 26637 -2613 26727 -2579
rect 26835 -2613 26925 -2579
rect 27033 -2613 27123 -2579
rect 27231 -2613 27321 -2579
rect 27429 -2613 27519 -2579
rect 27627 -2613 27717 -2579
rect 27825 -2613 27915 -2579
rect 28023 -2613 28113 -2579
rect 28221 -2613 28311 -2579
rect 28419 -2613 28509 -2579
rect 28617 -2613 28707 -2579
rect 28815 -2613 28905 -2579
rect 29013 -2613 29103 -2579
rect 29211 -2613 29301 -2579
rect 29409 -2613 29499 -2579
rect 29607 -2613 29697 -2579
rect 29805 -2613 29895 -2579
rect 30003 -2613 30093 -2579
rect 30201 -2613 30291 -2579
rect 30399 -2613 30489 -2579
rect 30597 -2613 30687 -2579
rect 30795 -2613 30885 -2579
rect 30993 -2613 31083 -2579
rect 31191 -2613 31281 -2579
rect 31389 -2613 31479 -2579
rect 31587 -2613 31896 -2579
rect 23052 -2643 31896 -2613
rect 23052 -3208 23206 -2643
rect 31742 -3208 31896 -2643
rect 23052 -3252 31896 -3208
rect 23052 -3286 23361 -3252
rect 23469 -3286 23559 -3252
rect 23667 -3286 23757 -3252
rect 23865 -3286 23955 -3252
rect 24063 -3286 24153 -3252
rect 24261 -3286 24351 -3252
rect 24459 -3286 24549 -3252
rect 24657 -3286 24747 -3252
rect 24855 -3286 24945 -3252
rect 25053 -3286 25143 -3252
rect 25251 -3286 25341 -3252
rect 25449 -3286 25539 -3252
rect 25647 -3286 25737 -3252
rect 25845 -3286 25935 -3252
rect 26043 -3286 26133 -3252
rect 26241 -3286 26331 -3252
rect 26439 -3286 26529 -3252
rect 26637 -3286 26727 -3252
rect 26835 -3286 26925 -3252
rect 27033 -3286 27123 -3252
rect 27231 -3286 27321 -3252
rect 27429 -3286 27519 -3252
rect 27627 -3286 27717 -3252
rect 27825 -3286 27915 -3252
rect 28023 -3286 28113 -3252
rect 28221 -3286 28311 -3252
rect 28419 -3286 28509 -3252
rect 28617 -3286 28707 -3252
rect 28815 -3286 28905 -3252
rect 29013 -3286 29103 -3252
rect 29211 -3286 29301 -3252
rect 29409 -3286 29499 -3252
rect 29607 -3286 29697 -3252
rect 29805 -3286 29895 -3252
rect 30003 -3286 30093 -3252
rect 30201 -3286 30291 -3252
rect 30399 -3286 30489 -3252
rect 30597 -3286 30687 -3252
rect 30795 -3286 30885 -3252
rect 30993 -3286 31083 -3252
rect 31191 -3286 31281 -3252
rect 31389 -3286 31479 -3252
rect 31587 -3286 31896 -3252
rect 23052 -3292 31896 -3286
rect 23293 -3345 23339 -3333
rect 23491 -3345 23537 -3333
rect 23689 -3345 23735 -3333
rect 23887 -3345 23933 -3333
rect 24085 -3345 24131 -3333
rect 24283 -3345 24329 -3333
rect 24481 -3345 24527 -3333
rect 24679 -3345 24725 -3333
rect 24877 -3345 24923 -3333
rect 25075 -3345 25121 -3333
rect 25273 -3345 25319 -3333
rect 25471 -3345 25517 -3333
rect 25669 -3345 25715 -3333
rect 25867 -3345 25913 -3333
rect 26065 -3345 26111 -3333
rect 26263 -3345 26309 -3333
rect 26461 -3345 26507 -3333
rect 26659 -3345 26705 -3333
rect 26857 -3345 26903 -3333
rect 27055 -3345 27101 -3333
rect 27253 -3345 27299 -3333
rect 27451 -3345 27497 -3333
rect 27649 -3345 27695 -3333
rect 27847 -3345 27893 -3333
rect 28045 -3345 28091 -3333
rect 28243 -3345 28289 -3333
rect 28441 -3345 28487 -3333
rect 28639 -3345 28685 -3333
rect 28837 -3345 28883 -3333
rect 29035 -3345 29081 -3333
rect 29233 -3345 29279 -3333
rect 29431 -3345 29477 -3333
rect 29629 -3345 29675 -3333
rect 29827 -3345 29873 -3333
rect 30025 -3345 30071 -3333
rect 30223 -3345 30269 -3333
rect 30421 -3345 30467 -3333
rect 30619 -3345 30665 -3333
rect 30817 -3345 30863 -3333
rect 31015 -3345 31061 -3333
rect 31213 -3345 31259 -3333
rect 31411 -3345 31457 -3333
rect 31609 -3344 31655 -3333
rect 23280 -4721 23290 -3345
rect 23342 -4721 23352 -3345
rect 23478 -4721 23488 -3345
rect 23540 -4721 23550 -3345
rect 23676 -4721 23686 -3345
rect 23738 -4721 23748 -3345
rect 23874 -4721 23884 -3345
rect 23936 -4721 23946 -3345
rect 24072 -4721 24082 -3345
rect 24134 -4721 24144 -3345
rect 24270 -4721 24280 -3345
rect 24332 -4721 24342 -3345
rect 24468 -4721 24478 -3345
rect 24530 -4721 24540 -3345
rect 24666 -4721 24676 -3345
rect 24728 -4721 24738 -3345
rect 24864 -4721 24874 -3345
rect 24926 -4721 24936 -3345
rect 25062 -4721 25072 -3345
rect 25124 -4721 25134 -3345
rect 25260 -4721 25270 -3345
rect 25322 -4721 25332 -3345
rect 25458 -4721 25468 -3345
rect 25520 -4721 25530 -3345
rect 25656 -4721 25666 -3345
rect 25718 -4721 25728 -3345
rect 25854 -4721 25864 -3345
rect 25916 -4721 25926 -3345
rect 26052 -4721 26062 -3345
rect 26114 -4721 26124 -3345
rect 26250 -4721 26260 -3345
rect 26312 -4721 26322 -3345
rect 26448 -4721 26458 -3345
rect 26510 -4721 26520 -3345
rect 26646 -4721 26656 -3345
rect 26708 -4721 26718 -3345
rect 26844 -4721 26854 -3345
rect 26906 -4721 26916 -3345
rect 27042 -4721 27052 -3345
rect 27104 -4721 27114 -3345
rect 27240 -4721 27250 -3345
rect 27302 -4721 27312 -3345
rect 27438 -4721 27448 -3345
rect 27500 -4721 27510 -3345
rect 27636 -4721 27646 -3345
rect 27698 -4721 27708 -3345
rect 27834 -4721 27844 -3345
rect 27896 -4721 27906 -3345
rect 28032 -4721 28042 -3345
rect 28094 -4721 28104 -3345
rect 28230 -4721 28240 -3345
rect 28292 -4721 28302 -3345
rect 28428 -4721 28438 -3345
rect 28490 -4721 28500 -3345
rect 28626 -4721 28636 -3345
rect 28688 -4721 28698 -3345
rect 28824 -4721 28834 -3345
rect 28886 -4721 28896 -3345
rect 29022 -4721 29032 -3345
rect 29084 -4721 29094 -3345
rect 29220 -4721 29230 -3345
rect 29282 -4721 29292 -3345
rect 29418 -4721 29428 -3345
rect 29480 -4721 29490 -3345
rect 29616 -4721 29626 -3345
rect 29678 -4721 29688 -3345
rect 29814 -4721 29824 -3345
rect 29876 -4721 29886 -3345
rect 30012 -4721 30022 -3345
rect 30074 -4721 30084 -3345
rect 30210 -4721 30220 -3345
rect 30272 -4721 30282 -3345
rect 30408 -4721 30418 -3345
rect 30470 -4721 30480 -3345
rect 30606 -4721 30616 -3345
rect 30668 -4721 30678 -3345
rect 30804 -4721 30814 -3345
rect 30866 -4721 30876 -3345
rect 31002 -4721 31012 -3345
rect 31064 -4721 31074 -3345
rect 31200 -4721 31210 -3345
rect 31262 -4721 31272 -3345
rect 31398 -4721 31408 -3345
rect 31460 -4721 31470 -3345
rect 31596 -4720 31606 -3344
rect 31658 -4720 31668 -3344
rect 31609 -4721 31615 -4720
rect 31649 -4721 31655 -4720
rect 23293 -5127 23339 -4721
rect 23491 -4733 23537 -4721
rect 23689 -5127 23735 -4721
rect 23887 -4733 23933 -4721
rect 24085 -5127 24131 -4721
rect 24283 -4733 24329 -4721
rect 24481 -5127 24527 -4721
rect 24679 -4733 24725 -4721
rect 24877 -5127 24923 -4721
rect 25075 -4733 25121 -4721
rect 25273 -5127 25319 -4721
rect 25471 -4733 25517 -4721
rect 25669 -5127 25715 -4721
rect 25867 -4733 25913 -4721
rect 26065 -5127 26111 -4721
rect 26263 -4733 26309 -4721
rect 26461 -5127 26507 -4721
rect 26659 -4733 26705 -4721
rect 26857 -5127 26903 -4721
rect 27055 -4733 27101 -4721
rect 27253 -5127 27299 -4721
rect 27451 -4733 27497 -4721
rect 27649 -5127 27695 -4721
rect 27847 -4733 27893 -4721
rect 28045 -5127 28091 -4721
rect 28243 -4733 28289 -4721
rect 28441 -5127 28487 -4721
rect 28639 -4733 28685 -4721
rect 28837 -5127 28883 -4721
rect 29035 -4733 29081 -4721
rect 29233 -5127 29279 -4721
rect 29431 -4733 29477 -4721
rect 29629 -5127 29675 -4721
rect 29827 -4733 29873 -4721
rect 30025 -5127 30071 -4721
rect 30223 -4733 30269 -4721
rect 30421 -5127 30467 -4721
rect 30619 -4733 30665 -4721
rect 30817 -5127 30863 -4721
rect 31015 -4733 31061 -4721
rect 31213 -5127 31259 -4721
rect 31411 -4733 31457 -4721
rect 31609 -5127 31655 -4721
rect 32606 -5127 33826 2327
rect -753 -6078 33826 -5127
<< via1 >>
rect -399 752 -347 2128
rect -201 752 -149 2128
rect -3 752 49 2128
rect 195 752 247 2128
rect 393 752 445 2128
rect 591 752 643 2128
rect 789 752 841 2128
rect 987 752 1039 2128
rect 1185 752 1237 2128
rect 1383 752 1435 2128
rect 1581 752 1633 2128
rect 1779 752 1831 2128
rect 1977 752 2029 2128
rect 2175 752 2227 2128
rect 2373 752 2425 2128
rect 2571 752 2623 2128
rect 2769 752 2821 2128
rect 2967 752 3019 2128
rect 3165 752 3217 2128
rect 3363 752 3415 2128
rect 3561 752 3613 2128
rect 3759 752 3811 2128
rect 3957 752 4009 2128
rect 4155 752 4207 2128
rect 4353 752 4405 2128
rect 4551 752 4603 2128
rect 4749 752 4801 2128
rect 4947 752 4999 2128
rect 5145 752 5197 2128
rect 5343 752 5395 2128
rect 5541 752 5593 2128
rect 5739 752 5791 2128
rect 5937 752 5989 2128
rect 6135 752 6187 2128
rect 6333 752 6385 2128
rect 6531 752 6583 2128
rect 6729 752 6781 2128
rect 6927 752 6979 2128
rect 7125 752 7177 2128
rect 7323 752 7375 2128
rect 7521 752 7573 2128
rect 7719 752 7771 2128
rect 7917 753 7969 2129
rect -627 -877 -493 -743
rect -399 -884 -347 492
rect -201 -884 -149 492
rect -3 -884 49 492
rect 195 -884 247 492
rect 393 -884 445 492
rect 591 -884 643 492
rect 789 -884 841 492
rect 987 -884 1039 492
rect 1185 -884 1237 492
rect 1383 -884 1435 492
rect 1581 -884 1633 492
rect 1779 -884 1831 492
rect 1977 -884 2029 492
rect 2175 -884 2227 492
rect 2373 -884 2425 492
rect 2571 -884 2623 492
rect 2769 -884 2821 492
rect 2967 -884 3019 492
rect 3165 -884 3217 492
rect 3363 -884 3415 492
rect 3561 -884 3613 492
rect 3759 -884 3811 492
rect 3957 -884 4009 492
rect 4155 -884 4207 492
rect 4353 -884 4405 492
rect 4551 -884 4603 492
rect 4749 -884 4801 492
rect 4947 -884 4999 492
rect 5145 -884 5197 492
rect 5343 -884 5395 492
rect 5541 -884 5593 492
rect 5739 -884 5791 492
rect 5937 -884 5989 492
rect 6135 -884 6187 492
rect 6333 -884 6385 492
rect 6531 -884 6583 492
rect 6729 -884 6781 492
rect 6927 -884 6979 492
rect 7125 -884 7177 492
rect 7323 -884 7375 492
rect 7521 -884 7573 492
rect 7719 -884 7771 492
rect 7917 -883 7969 493
rect 8063 -877 8197 -743
rect -627 -1081 -493 -947
rect 8063 -1081 8197 -947
rect -627 -1285 -493 -1151
rect -399 -2520 -347 -1144
rect -201 -2520 -149 -1144
rect -3 -2520 49 -1144
rect 195 -2520 247 -1144
rect 393 -2520 445 -1144
rect 591 -2520 643 -1144
rect 789 -2520 841 -1144
rect 987 -2520 1039 -1144
rect 1185 -2520 1237 -1144
rect 1383 -2520 1435 -1144
rect 1581 -2520 1633 -1144
rect 1779 -2520 1831 -1144
rect 1977 -2520 2029 -1144
rect 2175 -2520 2227 -1144
rect 2373 -2520 2425 -1144
rect 2571 -2520 2623 -1144
rect 2769 -2520 2821 -1144
rect 2967 -2520 3019 -1144
rect 3165 -2520 3217 -1144
rect 3363 -2520 3415 -1144
rect 3561 -2520 3613 -1144
rect 3759 -2520 3811 -1144
rect 3957 -2520 4009 -1144
rect 4155 -2520 4207 -1144
rect 4353 -2520 4405 -1144
rect 4551 -2520 4603 -1144
rect 4749 -2520 4801 -1144
rect 4947 -2520 4999 -1144
rect 5145 -2520 5197 -1144
rect 5343 -2520 5395 -1144
rect 5541 -2520 5593 -1144
rect 5739 -2520 5791 -1144
rect 5937 -2520 5989 -1144
rect 6135 -2520 6187 -1144
rect 6333 -2520 6385 -1144
rect 6531 -2520 6583 -1144
rect 6729 -2520 6781 -1144
rect 6927 -2520 6979 -1144
rect 7125 -2520 7177 -1144
rect 7323 -2520 7375 -1144
rect 7521 -2520 7573 -1144
rect 7719 -2520 7771 -1144
rect 7917 -2519 7969 -1143
rect 8063 -1285 8197 -1151
rect -399 -4721 -347 -3345
rect -201 -4721 -149 -3345
rect -3 -4721 49 -3345
rect 195 -4721 247 -3345
rect 393 -4721 445 -3345
rect 591 -4721 643 -3345
rect 789 -4721 841 -3345
rect 987 -4721 1039 -3345
rect 1185 -4721 1237 -3345
rect 1383 -4721 1435 -3345
rect 1581 -4721 1633 -3345
rect 1779 -4721 1831 -3345
rect 1977 -4721 2029 -3345
rect 2175 -4721 2227 -3345
rect 2373 -4721 2425 -3345
rect 2571 -4721 2623 -3345
rect 2769 -4721 2821 -3345
rect 2967 -4721 3019 -3345
rect 3165 -4721 3217 -3345
rect 3363 -4721 3415 -3345
rect 3561 -4721 3613 -3345
rect 3759 -4721 3811 -3345
rect 3957 -4721 4009 -3345
rect 4155 -4721 4207 -3345
rect 4353 -4721 4405 -3345
rect 4551 -4721 4603 -3345
rect 4749 -4721 4801 -3345
rect 4947 -4721 4999 -3345
rect 5145 -4721 5197 -3345
rect 5343 -4721 5395 -3345
rect 5541 -4721 5593 -3345
rect 5739 -4721 5791 -3345
rect 5937 -4721 5989 -3345
rect 6135 -4721 6187 -3345
rect 6333 -4721 6385 -3345
rect 6531 -4721 6583 -3345
rect 6729 -4721 6781 -3345
rect 6927 -4721 6979 -3345
rect 7125 -4721 7177 -3345
rect 7323 -4721 7375 -3345
rect 7521 -4721 7573 -3345
rect 7719 -4721 7771 -3345
rect 7917 -4720 7969 -3344
rect 11440 752 11449 2128
rect 11449 752 11483 2128
rect 11483 752 11492 2128
rect 11638 752 11647 2128
rect 11647 752 11681 2128
rect 11681 752 11690 2128
rect 11836 752 11845 2128
rect 11845 752 11879 2128
rect 11879 752 11888 2128
rect 12034 752 12043 2128
rect 12043 752 12077 2128
rect 12077 752 12086 2128
rect 12232 752 12241 2128
rect 12241 752 12275 2128
rect 12275 752 12284 2128
rect 12430 752 12439 2128
rect 12439 752 12473 2128
rect 12473 752 12482 2128
rect 12628 752 12637 2128
rect 12637 752 12671 2128
rect 12671 752 12680 2128
rect 12826 752 12835 2128
rect 12835 752 12869 2128
rect 12869 752 12878 2128
rect 13024 752 13033 2128
rect 13033 752 13067 2128
rect 13067 752 13076 2128
rect 13222 752 13231 2128
rect 13231 752 13265 2128
rect 13265 752 13274 2128
rect 13420 752 13429 2128
rect 13429 752 13463 2128
rect 13463 752 13472 2128
rect 13618 752 13627 2128
rect 13627 752 13661 2128
rect 13661 752 13670 2128
rect 13816 752 13825 2128
rect 13825 752 13859 2128
rect 13859 752 13868 2128
rect 14014 752 14023 2128
rect 14023 752 14057 2128
rect 14057 752 14066 2128
rect 14212 752 14221 2128
rect 14221 752 14255 2128
rect 14255 752 14264 2128
rect 14410 752 14419 2128
rect 14419 752 14453 2128
rect 14453 752 14462 2128
rect 14608 752 14617 2128
rect 14617 752 14651 2128
rect 14651 752 14660 2128
rect 14806 752 14815 2128
rect 14815 752 14849 2128
rect 14849 752 14858 2128
rect 15004 752 15013 2128
rect 15013 752 15047 2128
rect 15047 752 15056 2128
rect 15202 752 15211 2128
rect 15211 752 15245 2128
rect 15245 752 15254 2128
rect 15400 752 15409 2128
rect 15409 752 15443 2128
rect 15443 752 15452 2128
rect 15598 752 15607 2128
rect 15607 752 15641 2128
rect 15641 752 15650 2128
rect 15796 752 15805 2128
rect 15805 752 15839 2128
rect 15839 752 15848 2128
rect 15994 752 16003 2128
rect 16003 752 16037 2128
rect 16037 752 16046 2128
rect 16192 752 16201 2128
rect 16201 752 16235 2128
rect 16235 752 16244 2128
rect 16390 752 16399 2128
rect 16399 752 16433 2128
rect 16433 752 16442 2128
rect 16588 752 16597 2128
rect 16597 752 16631 2128
rect 16631 752 16640 2128
rect 16786 752 16795 2128
rect 16795 752 16829 2128
rect 16829 752 16838 2128
rect 16984 752 16993 2128
rect 16993 752 17027 2128
rect 17027 752 17036 2128
rect 17182 752 17191 2128
rect 17191 752 17225 2128
rect 17225 752 17234 2128
rect 17380 752 17389 2128
rect 17389 752 17423 2128
rect 17423 752 17432 2128
rect 17578 752 17587 2128
rect 17587 752 17621 2128
rect 17621 752 17630 2128
rect 17776 752 17785 2128
rect 17785 752 17819 2128
rect 17819 752 17828 2128
rect 17974 752 17983 2128
rect 17983 752 18017 2128
rect 18017 752 18026 2128
rect 18172 752 18181 2128
rect 18181 752 18215 2128
rect 18215 752 18224 2128
rect 18370 752 18379 2128
rect 18379 752 18413 2128
rect 18413 752 18422 2128
rect 18568 752 18577 2128
rect 18577 752 18611 2128
rect 18611 752 18620 2128
rect 18766 752 18775 2128
rect 18775 752 18809 2128
rect 18809 752 18818 2128
rect 18964 752 18973 2128
rect 18973 752 19007 2128
rect 19007 752 19016 2128
rect 19162 752 19171 2128
rect 19171 752 19205 2128
rect 19205 752 19214 2128
rect 19360 752 19369 2128
rect 19369 752 19403 2128
rect 19403 752 19412 2128
rect 19558 752 19567 2128
rect 19567 752 19601 2128
rect 19601 752 19610 2128
rect 19756 2128 19808 2129
rect 19756 753 19765 2128
rect 19765 753 19799 2128
rect 19799 753 19808 2128
rect 11212 -877 11346 -743
rect 11440 -884 11449 492
rect 11449 -884 11483 492
rect 11483 -884 11492 492
rect 11638 -884 11647 492
rect 11647 -884 11681 492
rect 11681 -884 11690 492
rect 11836 -884 11845 492
rect 11845 -884 11879 492
rect 11879 -884 11888 492
rect 12034 -884 12043 492
rect 12043 -884 12077 492
rect 12077 -884 12086 492
rect 12232 -884 12241 492
rect 12241 -884 12275 492
rect 12275 -884 12284 492
rect 12430 -884 12439 492
rect 12439 -884 12473 492
rect 12473 -884 12482 492
rect 12628 -884 12637 492
rect 12637 -884 12671 492
rect 12671 -884 12680 492
rect 12826 -884 12835 492
rect 12835 -884 12869 492
rect 12869 -884 12878 492
rect 13024 -884 13033 492
rect 13033 -884 13067 492
rect 13067 -884 13076 492
rect 13222 -884 13231 492
rect 13231 -884 13265 492
rect 13265 -884 13274 492
rect 13420 -884 13429 492
rect 13429 -884 13463 492
rect 13463 -884 13472 492
rect 13618 -884 13627 492
rect 13627 -884 13661 492
rect 13661 -884 13670 492
rect 13816 -884 13825 492
rect 13825 -884 13859 492
rect 13859 -884 13868 492
rect 14014 -884 14023 492
rect 14023 -884 14057 492
rect 14057 -884 14066 492
rect 14212 -884 14221 492
rect 14221 -884 14255 492
rect 14255 -884 14264 492
rect 14410 -884 14419 492
rect 14419 -884 14453 492
rect 14453 -884 14462 492
rect 14608 -884 14617 492
rect 14617 -884 14651 492
rect 14651 -884 14660 492
rect 14806 -884 14815 492
rect 14815 -884 14849 492
rect 14849 -884 14858 492
rect 15004 -884 15013 492
rect 15013 -884 15047 492
rect 15047 -884 15056 492
rect 15202 -884 15211 492
rect 15211 -884 15245 492
rect 15245 -884 15254 492
rect 15400 -884 15409 492
rect 15409 -884 15443 492
rect 15443 -884 15452 492
rect 15598 -884 15607 492
rect 15607 -884 15641 492
rect 15641 -884 15650 492
rect 15796 -884 15805 492
rect 15805 -884 15839 492
rect 15839 -884 15848 492
rect 15994 -884 16003 492
rect 16003 -884 16037 492
rect 16037 -884 16046 492
rect 16192 -884 16201 492
rect 16201 -884 16235 492
rect 16235 -884 16244 492
rect 16390 -884 16399 492
rect 16399 -884 16433 492
rect 16433 -884 16442 492
rect 16588 -884 16597 492
rect 16597 -884 16631 492
rect 16631 -884 16640 492
rect 16786 -884 16795 492
rect 16795 -884 16829 492
rect 16829 -884 16838 492
rect 16984 -884 16993 492
rect 16993 -884 17027 492
rect 17027 -884 17036 492
rect 17182 -884 17191 492
rect 17191 -884 17225 492
rect 17225 -884 17234 492
rect 17380 -884 17389 492
rect 17389 -884 17423 492
rect 17423 -884 17432 492
rect 17578 -884 17587 492
rect 17587 -884 17621 492
rect 17621 -884 17630 492
rect 17776 -884 17785 492
rect 17785 -884 17819 492
rect 17819 -884 17828 492
rect 17974 -884 17983 492
rect 17983 -884 18017 492
rect 18017 -884 18026 492
rect 18172 -884 18181 492
rect 18181 -884 18215 492
rect 18215 -884 18224 492
rect 18370 -884 18379 492
rect 18379 -884 18413 492
rect 18413 -884 18422 492
rect 18568 -884 18577 492
rect 18577 -884 18611 492
rect 18611 -884 18620 492
rect 18766 -884 18775 492
rect 18775 -884 18809 492
rect 18809 -884 18818 492
rect 18964 -884 18973 492
rect 18973 -884 19007 492
rect 19007 -884 19016 492
rect 19162 -884 19171 492
rect 19171 -884 19205 492
rect 19205 -884 19214 492
rect 19360 -884 19369 492
rect 19369 -884 19403 492
rect 19403 -884 19412 492
rect 19558 -884 19567 492
rect 19567 -884 19601 492
rect 19601 -884 19610 492
rect 19756 492 19808 493
rect 19756 -883 19765 492
rect 19765 -883 19799 492
rect 19799 -883 19808 492
rect 19902 -877 20036 -743
rect 11212 -1081 11346 -947
rect 19902 -1081 20036 -947
rect 11212 -1285 11346 -1151
rect 11440 -2520 11449 -1144
rect 11449 -2520 11483 -1144
rect 11483 -2520 11492 -1144
rect 11638 -2520 11647 -1144
rect 11647 -2520 11681 -1144
rect 11681 -2520 11690 -1144
rect 11836 -2520 11845 -1144
rect 11845 -2520 11879 -1144
rect 11879 -2520 11888 -1144
rect 12034 -2520 12043 -1144
rect 12043 -2520 12077 -1144
rect 12077 -2520 12086 -1144
rect 12232 -2520 12241 -1144
rect 12241 -2520 12275 -1144
rect 12275 -2520 12284 -1144
rect 12430 -2520 12439 -1144
rect 12439 -2520 12473 -1144
rect 12473 -2520 12482 -1144
rect 12628 -2520 12637 -1144
rect 12637 -2520 12671 -1144
rect 12671 -2520 12680 -1144
rect 12826 -2520 12835 -1144
rect 12835 -2520 12869 -1144
rect 12869 -2520 12878 -1144
rect 13024 -2520 13033 -1144
rect 13033 -2520 13067 -1144
rect 13067 -2520 13076 -1144
rect 13222 -2520 13231 -1144
rect 13231 -2520 13265 -1144
rect 13265 -2520 13274 -1144
rect 13420 -2520 13429 -1144
rect 13429 -2520 13463 -1144
rect 13463 -2520 13472 -1144
rect 13618 -2520 13627 -1144
rect 13627 -2520 13661 -1144
rect 13661 -2520 13670 -1144
rect 13816 -2520 13825 -1144
rect 13825 -2520 13859 -1144
rect 13859 -2520 13868 -1144
rect 14014 -2520 14023 -1144
rect 14023 -2520 14057 -1144
rect 14057 -2520 14066 -1144
rect 14212 -2520 14221 -1144
rect 14221 -2520 14255 -1144
rect 14255 -2520 14264 -1144
rect 14410 -2520 14419 -1144
rect 14419 -2520 14453 -1144
rect 14453 -2520 14462 -1144
rect 14608 -2520 14617 -1144
rect 14617 -2520 14651 -1144
rect 14651 -2520 14660 -1144
rect 14806 -2520 14815 -1144
rect 14815 -2520 14849 -1144
rect 14849 -2520 14858 -1144
rect 15004 -2520 15013 -1144
rect 15013 -2520 15047 -1144
rect 15047 -2520 15056 -1144
rect 15202 -2520 15211 -1144
rect 15211 -2520 15245 -1144
rect 15245 -2520 15254 -1144
rect 15400 -2520 15409 -1144
rect 15409 -2520 15443 -1144
rect 15443 -2520 15452 -1144
rect 15598 -2520 15607 -1144
rect 15607 -2520 15641 -1144
rect 15641 -2520 15650 -1144
rect 15796 -2520 15805 -1144
rect 15805 -2520 15839 -1144
rect 15839 -2520 15848 -1144
rect 15994 -2520 16003 -1144
rect 16003 -2520 16037 -1144
rect 16037 -2520 16046 -1144
rect 16192 -2520 16201 -1144
rect 16201 -2520 16235 -1144
rect 16235 -2520 16244 -1144
rect 16390 -2520 16399 -1144
rect 16399 -2520 16433 -1144
rect 16433 -2520 16442 -1144
rect 16588 -2520 16597 -1144
rect 16597 -2520 16631 -1144
rect 16631 -2520 16640 -1144
rect 16786 -2520 16795 -1144
rect 16795 -2520 16829 -1144
rect 16829 -2520 16838 -1144
rect 16984 -2520 16993 -1144
rect 16993 -2520 17027 -1144
rect 17027 -2520 17036 -1144
rect 17182 -2520 17191 -1144
rect 17191 -2520 17225 -1144
rect 17225 -2520 17234 -1144
rect 17380 -2520 17389 -1144
rect 17389 -2520 17423 -1144
rect 17423 -2520 17432 -1144
rect 17578 -2520 17587 -1144
rect 17587 -2520 17621 -1144
rect 17621 -2520 17630 -1144
rect 17776 -2520 17785 -1144
rect 17785 -2520 17819 -1144
rect 17819 -2520 17828 -1144
rect 17974 -2520 17983 -1144
rect 17983 -2520 18017 -1144
rect 18017 -2520 18026 -1144
rect 18172 -2520 18181 -1144
rect 18181 -2520 18215 -1144
rect 18215 -2520 18224 -1144
rect 18370 -2520 18379 -1144
rect 18379 -2520 18413 -1144
rect 18413 -2520 18422 -1144
rect 18568 -2520 18577 -1144
rect 18577 -2520 18611 -1144
rect 18611 -2520 18620 -1144
rect 18766 -2520 18775 -1144
rect 18775 -2520 18809 -1144
rect 18809 -2520 18818 -1144
rect 18964 -2520 18973 -1144
rect 18973 -2520 19007 -1144
rect 19007 -2520 19016 -1144
rect 19162 -2520 19171 -1144
rect 19171 -2520 19205 -1144
rect 19205 -2520 19214 -1144
rect 19360 -2520 19369 -1144
rect 19369 -2520 19403 -1144
rect 19403 -2520 19412 -1144
rect 19558 -2520 19567 -1144
rect 19567 -2520 19601 -1144
rect 19601 -2520 19610 -1144
rect 19756 -1144 19808 -1143
rect 19756 -2519 19765 -1144
rect 19765 -2519 19799 -1144
rect 19799 -2519 19808 -1144
rect 19902 -1285 20036 -1151
rect 11440 -4721 11449 -3345
rect 11449 -4721 11483 -3345
rect 11483 -4721 11492 -3345
rect 11638 -4721 11647 -3345
rect 11647 -4721 11681 -3345
rect 11681 -4721 11690 -3345
rect 11836 -4721 11845 -3345
rect 11845 -4721 11879 -3345
rect 11879 -4721 11888 -3345
rect 12034 -4721 12043 -3345
rect 12043 -4721 12077 -3345
rect 12077 -4721 12086 -3345
rect 12232 -4721 12241 -3345
rect 12241 -4721 12275 -3345
rect 12275 -4721 12284 -3345
rect 12430 -4721 12439 -3345
rect 12439 -4721 12473 -3345
rect 12473 -4721 12482 -3345
rect 12628 -4721 12637 -3345
rect 12637 -4721 12671 -3345
rect 12671 -4721 12680 -3345
rect 12826 -4721 12835 -3345
rect 12835 -4721 12869 -3345
rect 12869 -4721 12878 -3345
rect 13024 -4721 13033 -3345
rect 13033 -4721 13067 -3345
rect 13067 -4721 13076 -3345
rect 13222 -4721 13231 -3345
rect 13231 -4721 13265 -3345
rect 13265 -4721 13274 -3345
rect 13420 -4721 13429 -3345
rect 13429 -4721 13463 -3345
rect 13463 -4721 13472 -3345
rect 13618 -4721 13627 -3345
rect 13627 -4721 13661 -3345
rect 13661 -4721 13670 -3345
rect 13816 -4721 13825 -3345
rect 13825 -4721 13859 -3345
rect 13859 -4721 13868 -3345
rect 14014 -4721 14023 -3345
rect 14023 -4721 14057 -3345
rect 14057 -4721 14066 -3345
rect 14212 -4721 14221 -3345
rect 14221 -4721 14255 -3345
rect 14255 -4721 14264 -3345
rect 14410 -4721 14419 -3345
rect 14419 -4721 14453 -3345
rect 14453 -4721 14462 -3345
rect 14608 -4721 14617 -3345
rect 14617 -4721 14651 -3345
rect 14651 -4721 14660 -3345
rect 14806 -4721 14815 -3345
rect 14815 -4721 14849 -3345
rect 14849 -4721 14858 -3345
rect 15004 -4721 15013 -3345
rect 15013 -4721 15047 -3345
rect 15047 -4721 15056 -3345
rect 15202 -4721 15211 -3345
rect 15211 -4721 15245 -3345
rect 15245 -4721 15254 -3345
rect 15400 -4721 15409 -3345
rect 15409 -4721 15443 -3345
rect 15443 -4721 15452 -3345
rect 15598 -4721 15607 -3345
rect 15607 -4721 15641 -3345
rect 15641 -4721 15650 -3345
rect 15796 -4721 15805 -3345
rect 15805 -4721 15839 -3345
rect 15839 -4721 15848 -3345
rect 15994 -4721 16003 -3345
rect 16003 -4721 16037 -3345
rect 16037 -4721 16046 -3345
rect 16192 -4721 16201 -3345
rect 16201 -4721 16235 -3345
rect 16235 -4721 16244 -3345
rect 16390 -4721 16399 -3345
rect 16399 -4721 16433 -3345
rect 16433 -4721 16442 -3345
rect 16588 -4721 16597 -3345
rect 16597 -4721 16631 -3345
rect 16631 -4721 16640 -3345
rect 16786 -4721 16795 -3345
rect 16795 -4721 16829 -3345
rect 16829 -4721 16838 -3345
rect 16984 -4721 16993 -3345
rect 16993 -4721 17027 -3345
rect 17027 -4721 17036 -3345
rect 17182 -4721 17191 -3345
rect 17191 -4721 17225 -3345
rect 17225 -4721 17234 -3345
rect 17380 -4721 17389 -3345
rect 17389 -4721 17423 -3345
rect 17423 -4721 17432 -3345
rect 17578 -4721 17587 -3345
rect 17587 -4721 17621 -3345
rect 17621 -4721 17630 -3345
rect 17776 -4721 17785 -3345
rect 17785 -4721 17819 -3345
rect 17819 -4721 17828 -3345
rect 17974 -4721 17983 -3345
rect 17983 -4721 18017 -3345
rect 18017 -4721 18026 -3345
rect 18172 -4721 18181 -3345
rect 18181 -4721 18215 -3345
rect 18215 -4721 18224 -3345
rect 18370 -4721 18379 -3345
rect 18379 -4721 18413 -3345
rect 18413 -4721 18422 -3345
rect 18568 -4721 18577 -3345
rect 18577 -4721 18611 -3345
rect 18611 -4721 18620 -3345
rect 18766 -4721 18775 -3345
rect 18775 -4721 18809 -3345
rect 18809 -4721 18818 -3345
rect 18964 -4721 18973 -3345
rect 18973 -4721 19007 -3345
rect 19007 -4721 19016 -3345
rect 19162 -4721 19171 -3345
rect 19171 -4721 19205 -3345
rect 19205 -4721 19214 -3345
rect 19360 -4721 19369 -3345
rect 19369 -4721 19403 -3345
rect 19403 -4721 19412 -3345
rect 19558 -4721 19567 -3345
rect 19567 -4721 19601 -3345
rect 19601 -4721 19610 -3345
rect 19756 -3345 19808 -3344
rect 19756 -4720 19765 -3345
rect 19765 -4720 19799 -3345
rect 19799 -4720 19808 -3345
rect 23290 752 23299 2128
rect 23299 752 23333 2128
rect 23333 752 23342 2128
rect 23488 752 23497 2128
rect 23497 752 23531 2128
rect 23531 752 23540 2128
rect 23686 752 23695 2128
rect 23695 752 23729 2128
rect 23729 752 23738 2128
rect 23884 752 23893 2128
rect 23893 752 23927 2128
rect 23927 752 23936 2128
rect 24082 752 24091 2128
rect 24091 752 24125 2128
rect 24125 752 24134 2128
rect 24280 752 24289 2128
rect 24289 752 24323 2128
rect 24323 752 24332 2128
rect 24478 752 24487 2128
rect 24487 752 24521 2128
rect 24521 752 24530 2128
rect 24676 752 24685 2128
rect 24685 752 24719 2128
rect 24719 752 24728 2128
rect 24874 752 24883 2128
rect 24883 752 24917 2128
rect 24917 752 24926 2128
rect 25072 752 25081 2128
rect 25081 752 25115 2128
rect 25115 752 25124 2128
rect 25270 752 25279 2128
rect 25279 752 25313 2128
rect 25313 752 25322 2128
rect 25468 752 25477 2128
rect 25477 752 25511 2128
rect 25511 752 25520 2128
rect 25666 752 25675 2128
rect 25675 752 25709 2128
rect 25709 752 25718 2128
rect 25864 752 25873 2128
rect 25873 752 25907 2128
rect 25907 752 25916 2128
rect 26062 752 26071 2128
rect 26071 752 26105 2128
rect 26105 752 26114 2128
rect 26260 752 26269 2128
rect 26269 752 26303 2128
rect 26303 752 26312 2128
rect 26458 752 26467 2128
rect 26467 752 26501 2128
rect 26501 752 26510 2128
rect 26656 752 26665 2128
rect 26665 752 26699 2128
rect 26699 752 26708 2128
rect 26854 752 26863 2128
rect 26863 752 26897 2128
rect 26897 752 26906 2128
rect 27052 752 27061 2128
rect 27061 752 27095 2128
rect 27095 752 27104 2128
rect 27250 752 27259 2128
rect 27259 752 27293 2128
rect 27293 752 27302 2128
rect 27448 752 27457 2128
rect 27457 752 27491 2128
rect 27491 752 27500 2128
rect 27646 752 27655 2128
rect 27655 752 27689 2128
rect 27689 752 27698 2128
rect 27844 752 27853 2128
rect 27853 752 27887 2128
rect 27887 752 27896 2128
rect 28042 752 28051 2128
rect 28051 752 28085 2128
rect 28085 752 28094 2128
rect 28240 752 28249 2128
rect 28249 752 28283 2128
rect 28283 752 28292 2128
rect 28438 752 28447 2128
rect 28447 752 28481 2128
rect 28481 752 28490 2128
rect 28636 752 28645 2128
rect 28645 752 28679 2128
rect 28679 752 28688 2128
rect 28834 752 28843 2128
rect 28843 752 28877 2128
rect 28877 752 28886 2128
rect 29032 752 29041 2128
rect 29041 752 29075 2128
rect 29075 752 29084 2128
rect 29230 752 29239 2128
rect 29239 752 29273 2128
rect 29273 752 29282 2128
rect 29428 752 29437 2128
rect 29437 752 29471 2128
rect 29471 752 29480 2128
rect 29626 752 29635 2128
rect 29635 752 29669 2128
rect 29669 752 29678 2128
rect 29824 752 29833 2128
rect 29833 752 29867 2128
rect 29867 752 29876 2128
rect 30022 752 30031 2128
rect 30031 752 30065 2128
rect 30065 752 30074 2128
rect 30220 752 30229 2128
rect 30229 752 30263 2128
rect 30263 752 30272 2128
rect 30418 752 30427 2128
rect 30427 752 30461 2128
rect 30461 752 30470 2128
rect 30616 752 30625 2128
rect 30625 752 30659 2128
rect 30659 752 30668 2128
rect 30814 752 30823 2128
rect 30823 752 30857 2128
rect 30857 752 30866 2128
rect 31012 752 31021 2128
rect 31021 752 31055 2128
rect 31055 752 31064 2128
rect 31210 752 31219 2128
rect 31219 752 31253 2128
rect 31253 752 31262 2128
rect 31408 752 31417 2128
rect 31417 752 31451 2128
rect 31451 752 31460 2128
rect 31606 2128 31658 2129
rect 31606 753 31615 2128
rect 31615 753 31649 2128
rect 31649 753 31658 2128
rect 23062 -877 23196 -743
rect 23290 -884 23299 492
rect 23299 -884 23333 492
rect 23333 -884 23342 492
rect 23488 -884 23497 492
rect 23497 -884 23531 492
rect 23531 -884 23540 492
rect 23686 -884 23695 492
rect 23695 -884 23729 492
rect 23729 -884 23738 492
rect 23884 -884 23893 492
rect 23893 -884 23927 492
rect 23927 -884 23936 492
rect 24082 -884 24091 492
rect 24091 -884 24125 492
rect 24125 -884 24134 492
rect 24280 -884 24289 492
rect 24289 -884 24323 492
rect 24323 -884 24332 492
rect 24478 -884 24487 492
rect 24487 -884 24521 492
rect 24521 -884 24530 492
rect 24676 -884 24685 492
rect 24685 -884 24719 492
rect 24719 -884 24728 492
rect 24874 -884 24883 492
rect 24883 -884 24917 492
rect 24917 -884 24926 492
rect 25072 -884 25081 492
rect 25081 -884 25115 492
rect 25115 -884 25124 492
rect 25270 -884 25279 492
rect 25279 -884 25313 492
rect 25313 -884 25322 492
rect 25468 -884 25477 492
rect 25477 -884 25511 492
rect 25511 -884 25520 492
rect 25666 -884 25675 492
rect 25675 -884 25709 492
rect 25709 -884 25718 492
rect 25864 -884 25873 492
rect 25873 -884 25907 492
rect 25907 -884 25916 492
rect 26062 -884 26071 492
rect 26071 -884 26105 492
rect 26105 -884 26114 492
rect 26260 -884 26269 492
rect 26269 -884 26303 492
rect 26303 -884 26312 492
rect 26458 -884 26467 492
rect 26467 -884 26501 492
rect 26501 -884 26510 492
rect 26656 -884 26665 492
rect 26665 -884 26699 492
rect 26699 -884 26708 492
rect 26854 -884 26863 492
rect 26863 -884 26897 492
rect 26897 -884 26906 492
rect 27052 -884 27061 492
rect 27061 -884 27095 492
rect 27095 -884 27104 492
rect 27250 -884 27259 492
rect 27259 -884 27293 492
rect 27293 -884 27302 492
rect 27448 -884 27457 492
rect 27457 -884 27491 492
rect 27491 -884 27500 492
rect 27646 -884 27655 492
rect 27655 -884 27689 492
rect 27689 -884 27698 492
rect 27844 -884 27853 492
rect 27853 -884 27887 492
rect 27887 -884 27896 492
rect 28042 -884 28051 492
rect 28051 -884 28085 492
rect 28085 -884 28094 492
rect 28240 -884 28249 492
rect 28249 -884 28283 492
rect 28283 -884 28292 492
rect 28438 -884 28447 492
rect 28447 -884 28481 492
rect 28481 -884 28490 492
rect 28636 -884 28645 492
rect 28645 -884 28679 492
rect 28679 -884 28688 492
rect 28834 -884 28843 492
rect 28843 -884 28877 492
rect 28877 -884 28886 492
rect 29032 -884 29041 492
rect 29041 -884 29075 492
rect 29075 -884 29084 492
rect 29230 -884 29239 492
rect 29239 -884 29273 492
rect 29273 -884 29282 492
rect 29428 -884 29437 492
rect 29437 -884 29471 492
rect 29471 -884 29480 492
rect 29626 -884 29635 492
rect 29635 -884 29669 492
rect 29669 -884 29678 492
rect 29824 -884 29833 492
rect 29833 -884 29867 492
rect 29867 -884 29876 492
rect 30022 -884 30031 492
rect 30031 -884 30065 492
rect 30065 -884 30074 492
rect 30220 -884 30229 492
rect 30229 -884 30263 492
rect 30263 -884 30272 492
rect 30418 -884 30427 492
rect 30427 -884 30461 492
rect 30461 -884 30470 492
rect 30616 -884 30625 492
rect 30625 -884 30659 492
rect 30659 -884 30668 492
rect 30814 -884 30823 492
rect 30823 -884 30857 492
rect 30857 -884 30866 492
rect 31012 -884 31021 492
rect 31021 -884 31055 492
rect 31055 -884 31064 492
rect 31210 -884 31219 492
rect 31219 -884 31253 492
rect 31253 -884 31262 492
rect 31408 -884 31417 492
rect 31417 -884 31451 492
rect 31451 -884 31460 492
rect 31606 492 31658 493
rect 31606 -883 31615 492
rect 31615 -883 31649 492
rect 31649 -883 31658 492
rect 23062 -1081 23196 -947
rect 23062 -1285 23196 -1151
rect 23290 -2520 23299 -1144
rect 23299 -2520 23333 -1144
rect 23333 -2520 23342 -1144
rect 23488 -2520 23497 -1144
rect 23497 -2520 23531 -1144
rect 23531 -2520 23540 -1144
rect 23686 -2520 23695 -1144
rect 23695 -2520 23729 -1144
rect 23729 -2520 23738 -1144
rect 23884 -2520 23893 -1144
rect 23893 -2520 23927 -1144
rect 23927 -2520 23936 -1144
rect 24082 -2520 24091 -1144
rect 24091 -2520 24125 -1144
rect 24125 -2520 24134 -1144
rect 24280 -2520 24289 -1144
rect 24289 -2520 24323 -1144
rect 24323 -2520 24332 -1144
rect 24478 -2520 24487 -1144
rect 24487 -2520 24521 -1144
rect 24521 -2520 24530 -1144
rect 24676 -2520 24685 -1144
rect 24685 -2520 24719 -1144
rect 24719 -2520 24728 -1144
rect 24874 -2520 24883 -1144
rect 24883 -2520 24917 -1144
rect 24917 -2520 24926 -1144
rect 25072 -2520 25081 -1144
rect 25081 -2520 25115 -1144
rect 25115 -2520 25124 -1144
rect 25270 -2520 25279 -1144
rect 25279 -2520 25313 -1144
rect 25313 -2520 25322 -1144
rect 25468 -2520 25477 -1144
rect 25477 -2520 25511 -1144
rect 25511 -2520 25520 -1144
rect 25666 -2520 25675 -1144
rect 25675 -2520 25709 -1144
rect 25709 -2520 25718 -1144
rect 25864 -2520 25873 -1144
rect 25873 -2520 25907 -1144
rect 25907 -2520 25916 -1144
rect 26062 -2520 26071 -1144
rect 26071 -2520 26105 -1144
rect 26105 -2520 26114 -1144
rect 26260 -2520 26269 -1144
rect 26269 -2520 26303 -1144
rect 26303 -2520 26312 -1144
rect 26458 -2520 26467 -1144
rect 26467 -2520 26501 -1144
rect 26501 -2520 26510 -1144
rect 26656 -2520 26665 -1144
rect 26665 -2520 26699 -1144
rect 26699 -2520 26708 -1144
rect 26854 -2520 26863 -1144
rect 26863 -2520 26897 -1144
rect 26897 -2520 26906 -1144
rect 27052 -2520 27061 -1144
rect 27061 -2520 27095 -1144
rect 27095 -2520 27104 -1144
rect 27250 -2520 27259 -1144
rect 27259 -2520 27293 -1144
rect 27293 -2520 27302 -1144
rect 27448 -2520 27457 -1144
rect 27457 -2520 27491 -1144
rect 27491 -2520 27500 -1144
rect 27646 -2520 27655 -1144
rect 27655 -2520 27689 -1144
rect 27689 -2520 27698 -1144
rect 27844 -2520 27853 -1144
rect 27853 -2520 27887 -1144
rect 27887 -2520 27896 -1144
rect 28042 -2520 28051 -1144
rect 28051 -2520 28085 -1144
rect 28085 -2520 28094 -1144
rect 28240 -2520 28249 -1144
rect 28249 -2520 28283 -1144
rect 28283 -2520 28292 -1144
rect 28438 -2520 28447 -1144
rect 28447 -2520 28481 -1144
rect 28481 -2520 28490 -1144
rect 28636 -2520 28645 -1144
rect 28645 -2520 28679 -1144
rect 28679 -2520 28688 -1144
rect 28834 -2520 28843 -1144
rect 28843 -2520 28877 -1144
rect 28877 -2520 28886 -1144
rect 29032 -2520 29041 -1144
rect 29041 -2520 29075 -1144
rect 29075 -2520 29084 -1144
rect 29230 -2520 29239 -1144
rect 29239 -2520 29273 -1144
rect 29273 -2520 29282 -1144
rect 29428 -2520 29437 -1144
rect 29437 -2520 29471 -1144
rect 29471 -2520 29480 -1144
rect 29626 -2520 29635 -1144
rect 29635 -2520 29669 -1144
rect 29669 -2520 29678 -1144
rect 29824 -2520 29833 -1144
rect 29833 -2520 29867 -1144
rect 29867 -2520 29876 -1144
rect 30022 -2520 30031 -1144
rect 30031 -2520 30065 -1144
rect 30065 -2520 30074 -1144
rect 30220 -2520 30229 -1144
rect 30229 -2520 30263 -1144
rect 30263 -2520 30272 -1144
rect 30418 -2520 30427 -1144
rect 30427 -2520 30461 -1144
rect 30461 -2520 30470 -1144
rect 30616 -2520 30625 -1144
rect 30625 -2520 30659 -1144
rect 30659 -2520 30668 -1144
rect 30814 -2520 30823 -1144
rect 30823 -2520 30857 -1144
rect 30857 -2520 30866 -1144
rect 31012 -2520 31021 -1144
rect 31021 -2520 31055 -1144
rect 31055 -2520 31064 -1144
rect 31210 -2520 31219 -1144
rect 31219 -2520 31253 -1144
rect 31253 -2520 31262 -1144
rect 31408 -2520 31417 -1144
rect 31417 -2520 31451 -1144
rect 31451 -2520 31460 -1144
rect 31606 -1144 31658 -1143
rect 31606 -2519 31615 -1144
rect 31615 -2519 31649 -1144
rect 31649 -2519 31658 -1144
rect 23290 -4721 23299 -3345
rect 23299 -4721 23333 -3345
rect 23333 -4721 23342 -3345
rect 23488 -4721 23497 -3345
rect 23497 -4721 23531 -3345
rect 23531 -4721 23540 -3345
rect 23686 -4721 23695 -3345
rect 23695 -4721 23729 -3345
rect 23729 -4721 23738 -3345
rect 23884 -4721 23893 -3345
rect 23893 -4721 23927 -3345
rect 23927 -4721 23936 -3345
rect 24082 -4721 24091 -3345
rect 24091 -4721 24125 -3345
rect 24125 -4721 24134 -3345
rect 24280 -4721 24289 -3345
rect 24289 -4721 24323 -3345
rect 24323 -4721 24332 -3345
rect 24478 -4721 24487 -3345
rect 24487 -4721 24521 -3345
rect 24521 -4721 24530 -3345
rect 24676 -4721 24685 -3345
rect 24685 -4721 24719 -3345
rect 24719 -4721 24728 -3345
rect 24874 -4721 24883 -3345
rect 24883 -4721 24917 -3345
rect 24917 -4721 24926 -3345
rect 25072 -4721 25081 -3345
rect 25081 -4721 25115 -3345
rect 25115 -4721 25124 -3345
rect 25270 -4721 25279 -3345
rect 25279 -4721 25313 -3345
rect 25313 -4721 25322 -3345
rect 25468 -4721 25477 -3345
rect 25477 -4721 25511 -3345
rect 25511 -4721 25520 -3345
rect 25666 -4721 25675 -3345
rect 25675 -4721 25709 -3345
rect 25709 -4721 25718 -3345
rect 25864 -4721 25873 -3345
rect 25873 -4721 25907 -3345
rect 25907 -4721 25916 -3345
rect 26062 -4721 26071 -3345
rect 26071 -4721 26105 -3345
rect 26105 -4721 26114 -3345
rect 26260 -4721 26269 -3345
rect 26269 -4721 26303 -3345
rect 26303 -4721 26312 -3345
rect 26458 -4721 26467 -3345
rect 26467 -4721 26501 -3345
rect 26501 -4721 26510 -3345
rect 26656 -4721 26665 -3345
rect 26665 -4721 26699 -3345
rect 26699 -4721 26708 -3345
rect 26854 -4721 26863 -3345
rect 26863 -4721 26897 -3345
rect 26897 -4721 26906 -3345
rect 27052 -4721 27061 -3345
rect 27061 -4721 27095 -3345
rect 27095 -4721 27104 -3345
rect 27250 -4721 27259 -3345
rect 27259 -4721 27293 -3345
rect 27293 -4721 27302 -3345
rect 27448 -4721 27457 -3345
rect 27457 -4721 27491 -3345
rect 27491 -4721 27500 -3345
rect 27646 -4721 27655 -3345
rect 27655 -4721 27689 -3345
rect 27689 -4721 27698 -3345
rect 27844 -4721 27853 -3345
rect 27853 -4721 27887 -3345
rect 27887 -4721 27896 -3345
rect 28042 -4721 28051 -3345
rect 28051 -4721 28085 -3345
rect 28085 -4721 28094 -3345
rect 28240 -4721 28249 -3345
rect 28249 -4721 28283 -3345
rect 28283 -4721 28292 -3345
rect 28438 -4721 28447 -3345
rect 28447 -4721 28481 -3345
rect 28481 -4721 28490 -3345
rect 28636 -4721 28645 -3345
rect 28645 -4721 28679 -3345
rect 28679 -4721 28688 -3345
rect 28834 -4721 28843 -3345
rect 28843 -4721 28877 -3345
rect 28877 -4721 28886 -3345
rect 29032 -4721 29041 -3345
rect 29041 -4721 29075 -3345
rect 29075 -4721 29084 -3345
rect 29230 -4721 29239 -3345
rect 29239 -4721 29273 -3345
rect 29273 -4721 29282 -3345
rect 29428 -4721 29437 -3345
rect 29437 -4721 29471 -3345
rect 29471 -4721 29480 -3345
rect 29626 -4721 29635 -3345
rect 29635 -4721 29669 -3345
rect 29669 -4721 29678 -3345
rect 29824 -4721 29833 -3345
rect 29833 -4721 29867 -3345
rect 29867 -4721 29876 -3345
rect 30022 -4721 30031 -3345
rect 30031 -4721 30065 -3345
rect 30065 -4721 30074 -3345
rect 30220 -4721 30229 -3345
rect 30229 -4721 30263 -3345
rect 30263 -4721 30272 -3345
rect 30418 -4721 30427 -3345
rect 30427 -4721 30461 -3345
rect 30461 -4721 30470 -3345
rect 30616 -4721 30625 -3345
rect 30625 -4721 30659 -3345
rect 30659 -4721 30668 -3345
rect 30814 -4721 30823 -3345
rect 30823 -4721 30857 -3345
rect 30857 -4721 30866 -3345
rect 31012 -4721 31021 -3345
rect 31021 -4721 31055 -3345
rect 31055 -4721 31064 -3345
rect 31210 -4721 31219 -3345
rect 31219 -4721 31253 -3345
rect 31253 -4721 31262 -3345
rect 31408 -4721 31417 -3345
rect 31417 -4721 31451 -3345
rect 31451 -4721 31460 -3345
rect 31606 -3345 31658 -3344
rect 31606 -4720 31615 -3345
rect 31615 -4720 31649 -3345
rect 31649 -4720 31658 -3345
<< metal2 >>
rect -399 2128 -347 2134
rect -399 492 -347 752
rect -627 -743 -493 -733
rect -627 -887 -493 -877
rect -627 -947 -493 -937
rect -627 -1091 -493 -1081
rect -627 -1151 -493 -1141
rect -627 -1295 -493 -1285
rect -399 -1144 -347 -884
rect -399 -3345 -347 -2520
rect -399 -4731 -347 -4721
rect -201 2128 -149 2138
rect -201 492 -149 752
rect -201 -1144 -149 -884
rect -201 -3345 -149 -2520
rect -201 -4783 -149 -4721
rect -3 2128 49 2134
rect -3 492 49 752
rect -3 -1144 49 -884
rect -3 -3345 49 -2520
rect -3 -4731 49 -4721
rect 195 2128 247 2138
rect 195 492 247 752
rect 195 -1144 247 -884
rect 195 -3345 247 -2520
rect 195 -4783 247 -4721
rect 393 2128 445 2134
rect 393 492 445 752
rect 393 -1144 445 -884
rect 393 -3345 445 -2520
rect 393 -4731 445 -4721
rect 591 2128 643 2138
rect 591 492 643 752
rect 591 -1144 643 -884
rect 591 -3345 643 -2520
rect 591 -4783 643 -4721
rect 789 2128 841 2134
rect 789 492 841 752
rect 789 -1144 841 -884
rect 789 -3345 841 -2520
rect 789 -4731 841 -4721
rect 987 2128 1039 2138
rect 987 492 1039 752
rect 987 -1144 1039 -884
rect 987 -3345 1039 -2520
rect 987 -4783 1039 -4721
rect 1185 2128 1237 2134
rect 1185 492 1237 752
rect 1185 -1144 1237 -884
rect 1185 -3345 1237 -2520
rect 1185 -4731 1237 -4721
rect 1383 2128 1435 2138
rect 1383 492 1435 752
rect 1383 -1144 1435 -884
rect 1383 -3345 1435 -2520
rect 1383 -4783 1435 -4721
rect 1581 2128 1633 2134
rect 1581 492 1633 752
rect 1581 -1144 1633 -884
rect 1581 -3345 1633 -2520
rect 1581 -4731 1633 -4721
rect 1779 2128 1831 2138
rect 1779 492 1831 752
rect 1779 -1144 1831 -884
rect 1779 -3345 1831 -2520
rect 1779 -4783 1831 -4721
rect 1977 2128 2029 2134
rect 1977 492 2029 752
rect 1977 -1144 2029 -884
rect 1977 -3345 2029 -2520
rect 1977 -4731 2029 -4721
rect 2175 2128 2227 2138
rect 2175 492 2227 752
rect 2175 -1144 2227 -884
rect 2175 -3345 2227 -2520
rect 2175 -4783 2227 -4721
rect 2373 2128 2425 2134
rect 2373 492 2425 752
rect 2373 -1144 2425 -884
rect 2373 -3345 2425 -2520
rect 2373 -4731 2425 -4721
rect 2571 2128 2623 2138
rect 2571 492 2623 752
rect 2571 -1144 2623 -884
rect 2571 -3345 2623 -2520
rect 2571 -4783 2623 -4721
rect 2769 2128 2821 2134
rect 2769 492 2821 752
rect 2769 -1144 2821 -884
rect 2769 -3345 2821 -2520
rect 2769 -4731 2821 -4721
rect 2967 2128 3019 2138
rect 2967 492 3019 752
rect 2967 -1144 3019 -884
rect 2967 -3345 3019 -2520
rect 2967 -4783 3019 -4721
rect 3165 2128 3217 2134
rect 3165 492 3217 752
rect 3165 -1144 3217 -884
rect 3165 -3345 3217 -2520
rect 3165 -4731 3217 -4721
rect 3363 2128 3415 2138
rect 3363 492 3415 752
rect 3363 -1144 3415 -884
rect 3363 -3345 3415 -2520
rect 3363 -4783 3415 -4721
rect 3561 2128 3613 2134
rect 3561 492 3613 752
rect 3561 -1144 3613 -884
rect 3561 -3345 3613 -2520
rect 3561 -4731 3613 -4721
rect 3759 2128 3811 2138
rect 3759 492 3811 752
rect 3759 -1144 3811 -884
rect 3759 -3345 3811 -2520
rect 3759 -4783 3811 -4721
rect 3957 2128 4009 2134
rect 3957 492 4009 752
rect 3957 -1144 4009 -884
rect 3957 -3345 4009 -2520
rect 3957 -4731 4009 -4721
rect 4155 2128 4207 2138
rect 4155 492 4207 752
rect 4155 -1144 4207 -884
rect 4155 -3345 4207 -2520
rect 4155 -4783 4207 -4721
rect 4353 2128 4405 2134
rect 4353 492 4405 752
rect 4353 -1144 4405 -884
rect 4353 -3345 4405 -2520
rect 4353 -4731 4405 -4721
rect 4551 2128 4603 2138
rect 4551 492 4603 752
rect 4551 -1144 4603 -884
rect 4551 -3345 4603 -2520
rect 4551 -4783 4603 -4721
rect 4749 2128 4801 2134
rect 4749 492 4801 752
rect 4749 -1144 4801 -884
rect 4749 -3345 4801 -2520
rect 4749 -4731 4801 -4721
rect 4947 2128 4999 2138
rect 4947 492 4999 752
rect 4947 -1144 4999 -884
rect 4947 -3345 4999 -2520
rect 4947 -4783 4999 -4721
rect 5145 2128 5197 2134
rect 5145 492 5197 752
rect 5145 -1144 5197 -884
rect 5145 -3345 5197 -2520
rect 5145 -4731 5197 -4721
rect 5343 2128 5395 2138
rect 5343 492 5395 752
rect 5343 -1144 5395 -884
rect 5343 -3345 5395 -2520
rect 5343 -4783 5395 -4721
rect 5541 2128 5593 2134
rect 5541 492 5593 752
rect 5541 -1144 5593 -884
rect 5541 -3345 5593 -2520
rect 5541 -4731 5593 -4721
rect 5739 2128 5791 2138
rect 5739 492 5791 752
rect 5739 -1144 5791 -884
rect 5739 -3345 5791 -2520
rect 5739 -4783 5791 -4721
rect 5937 2128 5989 2134
rect 5937 492 5989 752
rect 5937 -1144 5989 -884
rect 5937 -3345 5989 -2520
rect 5937 -4731 5989 -4721
rect 6135 2128 6187 2138
rect 6135 492 6187 752
rect 6135 -1144 6187 -884
rect 6135 -3345 6187 -2520
rect 6135 -4783 6187 -4721
rect 6333 2128 6385 2134
rect 6333 492 6385 752
rect 6333 -1144 6385 -884
rect 6333 -3345 6385 -2520
rect 6333 -4731 6385 -4721
rect 6531 2128 6583 2138
rect 6531 492 6583 752
rect 6531 -1144 6583 -884
rect 6531 -3345 6583 -2520
rect 6531 -4783 6583 -4721
rect 6729 2128 6781 2134
rect 6729 492 6781 752
rect 6729 -1144 6781 -884
rect 6729 -3345 6781 -2520
rect 6729 -4731 6781 -4721
rect 6927 2128 6979 2138
rect 6927 492 6979 752
rect 6927 -1144 6979 -884
rect 6927 -3345 6979 -2520
rect 6927 -4783 6979 -4721
rect 7125 2128 7177 2134
rect 7125 492 7177 752
rect 7125 -1144 7177 -884
rect 7125 -3345 7177 -2520
rect 7125 -4731 7177 -4721
rect 7323 2128 7375 2138
rect 7323 492 7375 752
rect 7323 -1144 7375 -884
rect 7323 -3345 7375 -2520
rect 7323 -4783 7375 -4721
rect 7521 2128 7573 2134
rect 7521 492 7573 752
rect 7521 -1144 7573 -884
rect 7521 -3345 7573 -2520
rect 7521 -4731 7573 -4721
rect 7719 2128 7771 2138
rect 7719 492 7771 752
rect 7719 -1144 7771 -884
rect 7719 -3345 7771 -2520
rect 7719 -4783 7771 -4721
rect 7917 2129 7969 2135
rect 7917 493 7969 753
rect 11440 2128 11492 2134
rect 11440 492 11492 752
rect 7917 -1143 7969 -883
rect 8063 -743 8197 -733
rect 8063 -887 8197 -877
rect 11212 -743 11346 -733
rect 11212 -887 11346 -877
rect 8063 -947 8197 -937
rect 8063 -1091 8197 -1081
rect 11212 -947 11346 -937
rect 11212 -1091 11346 -1081
rect 8063 -1151 8197 -1141
rect 8063 -1295 8197 -1285
rect 11212 -1151 11346 -1141
rect 11212 -1295 11346 -1285
rect 11440 -1144 11492 -884
rect 7917 -3344 7969 -2519
rect 7917 -4730 7969 -4720
rect 11440 -3345 11492 -2520
rect 11440 -4731 11492 -4721
rect 11638 2128 11690 2138
rect 11638 492 11690 752
rect 11638 -1144 11690 -884
rect 11638 -3345 11690 -2520
rect 11638 -4783 11690 -4721
rect 11836 2128 11888 2134
rect 11836 492 11888 752
rect 11836 -1144 11888 -884
rect 11836 -3345 11888 -2520
rect 11836 -4731 11888 -4721
rect 12034 2128 12086 2138
rect 12034 492 12086 752
rect 12034 -1144 12086 -884
rect 12034 -3345 12086 -2520
rect 12034 -4783 12086 -4721
rect 12232 2128 12284 2134
rect 12232 492 12284 752
rect 12232 -1144 12284 -884
rect 12232 -3345 12284 -2520
rect 12232 -4731 12284 -4721
rect 12430 2128 12482 2138
rect 12430 492 12482 752
rect 12430 -1144 12482 -884
rect 12430 -3345 12482 -2520
rect 12430 -4783 12482 -4721
rect 12628 2128 12680 2134
rect 12628 492 12680 752
rect 12628 -1144 12680 -884
rect 12628 -3345 12680 -2520
rect 12628 -4731 12680 -4721
rect 12826 2128 12878 2138
rect 12826 492 12878 752
rect 12826 -1144 12878 -884
rect 12826 -3345 12878 -2520
rect 12826 -4783 12878 -4721
rect 13024 2128 13076 2134
rect 13024 492 13076 752
rect 13024 -1144 13076 -884
rect 13024 -3345 13076 -2520
rect 13024 -4731 13076 -4721
rect 13222 2128 13274 2138
rect 13222 492 13274 752
rect 13222 -1144 13274 -884
rect 13222 -3345 13274 -2520
rect 13222 -4783 13274 -4721
rect 13420 2128 13472 2134
rect 13420 492 13472 752
rect 13420 -1144 13472 -884
rect 13420 -3345 13472 -2520
rect 13420 -4731 13472 -4721
rect 13618 2128 13670 2138
rect 13618 492 13670 752
rect 13618 -1144 13670 -884
rect 13618 -3345 13670 -2520
rect 13618 -4783 13670 -4721
rect 13816 2128 13868 2134
rect 13816 492 13868 752
rect 13816 -1144 13868 -884
rect 13816 -3345 13868 -2520
rect 13816 -4731 13868 -4721
rect 14014 2128 14066 2138
rect 14014 492 14066 752
rect 14014 -1144 14066 -884
rect 14014 -3345 14066 -2520
rect 14014 -4783 14066 -4721
rect 14212 2128 14264 2134
rect 14212 492 14264 752
rect 14212 -1144 14264 -884
rect 14212 -3345 14264 -2520
rect 14212 -4731 14264 -4721
rect 14410 2128 14462 2138
rect 14410 492 14462 752
rect 14410 -1144 14462 -884
rect 14410 -3345 14462 -2520
rect 14410 -4783 14462 -4721
rect 14608 2128 14660 2134
rect 14608 492 14660 752
rect 14608 -1144 14660 -884
rect 14608 -3345 14660 -2520
rect 14608 -4731 14660 -4721
rect 14806 2128 14858 2138
rect 14806 492 14858 752
rect 14806 -1144 14858 -884
rect 14806 -3345 14858 -2520
rect 14806 -4783 14858 -4721
rect 15004 2128 15056 2134
rect 15004 492 15056 752
rect 15004 -1144 15056 -884
rect 15004 -3345 15056 -2520
rect 15004 -4731 15056 -4721
rect 15202 2128 15254 2138
rect 15202 492 15254 752
rect 15202 -1144 15254 -884
rect 15202 -3345 15254 -2520
rect 15202 -4783 15254 -4721
rect 15400 2128 15452 2134
rect 15400 492 15452 752
rect 15400 -1144 15452 -884
rect 15400 -3345 15452 -2520
rect 15400 -4731 15452 -4721
rect 15598 2128 15650 2138
rect 15598 492 15650 752
rect 15598 -1144 15650 -884
rect 15598 -3345 15650 -2520
rect 15598 -4783 15650 -4721
rect 15796 2128 15848 2134
rect 15796 492 15848 752
rect 15796 -1144 15848 -884
rect 15796 -3345 15848 -2520
rect 15796 -4731 15848 -4721
rect 15994 2128 16046 2138
rect 15994 492 16046 752
rect 15994 -1144 16046 -884
rect 15994 -3345 16046 -2520
rect 15994 -4783 16046 -4721
rect 16192 2128 16244 2134
rect 16192 492 16244 752
rect 16192 -1144 16244 -884
rect 16192 -3345 16244 -2520
rect 16192 -4731 16244 -4721
rect 16390 2128 16442 2138
rect 16390 492 16442 752
rect 16390 -1144 16442 -884
rect 16390 -3345 16442 -2520
rect 16390 -4783 16442 -4721
rect 16588 2128 16640 2134
rect 16588 492 16640 752
rect 16588 -1144 16640 -884
rect 16588 -3345 16640 -2520
rect 16588 -4731 16640 -4721
rect 16786 2128 16838 2138
rect 16786 492 16838 752
rect 16786 -1144 16838 -884
rect 16786 -3345 16838 -2520
rect 16786 -4783 16838 -4721
rect 16984 2128 17036 2134
rect 16984 492 17036 752
rect 16984 -1144 17036 -884
rect 16984 -3345 17036 -2520
rect 16984 -4731 17036 -4721
rect 17182 2128 17234 2138
rect 17182 492 17234 752
rect 17182 -1144 17234 -884
rect 17182 -3345 17234 -2520
rect 17182 -4783 17234 -4721
rect 17380 2128 17432 2134
rect 17380 492 17432 752
rect 17380 -1144 17432 -884
rect 17380 -3345 17432 -2520
rect 17380 -4731 17432 -4721
rect 17578 2128 17630 2138
rect 17578 492 17630 752
rect 17578 -1144 17630 -884
rect 17578 -3345 17630 -2520
rect 17578 -4783 17630 -4721
rect 17776 2128 17828 2134
rect 17776 492 17828 752
rect 17776 -1144 17828 -884
rect 17776 -3345 17828 -2520
rect 17776 -4731 17828 -4721
rect 17974 2128 18026 2138
rect 17974 492 18026 752
rect 17974 -1144 18026 -884
rect 17974 -3345 18026 -2520
rect 17974 -4783 18026 -4721
rect 18172 2128 18224 2134
rect 18172 492 18224 752
rect 18172 -1144 18224 -884
rect 18172 -3345 18224 -2520
rect 18172 -4731 18224 -4721
rect 18370 2128 18422 2138
rect 18370 492 18422 752
rect 18370 -1144 18422 -884
rect 18370 -3345 18422 -2520
rect 18370 -4783 18422 -4721
rect 18568 2128 18620 2134
rect 18568 492 18620 752
rect 18568 -1144 18620 -884
rect 18568 -3345 18620 -2520
rect 18568 -4731 18620 -4721
rect 18766 2128 18818 2138
rect 18766 492 18818 752
rect 18766 -1144 18818 -884
rect 18766 -3345 18818 -2520
rect 18766 -4783 18818 -4721
rect 18964 2128 19016 2134
rect 18964 492 19016 752
rect 18964 -1144 19016 -884
rect 18964 -3345 19016 -2520
rect 18964 -4731 19016 -4721
rect 19162 2128 19214 2138
rect 19162 492 19214 752
rect 19162 -1144 19214 -884
rect 19162 -3345 19214 -2520
rect 19162 -4783 19214 -4721
rect 19360 2128 19412 2134
rect 19360 492 19412 752
rect 19360 -1144 19412 -884
rect 19360 -3345 19412 -2520
rect 19360 -4731 19412 -4721
rect 19558 2128 19610 2138
rect 19558 492 19610 752
rect 19558 -1144 19610 -884
rect 19558 -3345 19610 -2520
rect 19558 -4783 19610 -4721
rect 19756 2129 19808 2135
rect 19756 493 19808 753
rect 23290 2128 23342 2134
rect 23290 492 23342 752
rect 19756 -1143 19808 -883
rect 19902 -743 20036 -733
rect 19902 -887 20036 -877
rect 23062 -743 23196 -733
rect 23062 -887 23196 -877
rect 19902 -947 20036 -937
rect 19902 -1091 20036 -1081
rect 23062 -947 23196 -937
rect 23062 -1091 23196 -1081
rect 19902 -1151 20036 -1141
rect 19902 -1295 20036 -1285
rect 23062 -1151 23196 -1141
rect 23062 -1295 23196 -1285
rect 23290 -1144 23342 -884
rect 19756 -3344 19808 -2519
rect 19756 -4730 19808 -4720
rect 23290 -3345 23342 -2520
rect 23290 -4731 23342 -4721
rect 23488 2128 23540 2138
rect 23488 492 23540 752
rect 23488 -1144 23540 -884
rect 23488 -3345 23540 -2520
rect 23488 -4783 23540 -4721
rect 23686 2128 23738 2134
rect 23686 492 23738 752
rect 23686 -1144 23738 -884
rect 23686 -3345 23738 -2520
rect 23686 -4731 23738 -4721
rect 23884 2128 23936 2138
rect 23884 492 23936 752
rect 23884 -1144 23936 -884
rect 23884 -3345 23936 -2520
rect 23884 -4783 23936 -4721
rect 24082 2128 24134 2134
rect 24082 492 24134 752
rect 24082 -1144 24134 -884
rect 24082 -3345 24134 -2520
rect 24082 -4731 24134 -4721
rect 24280 2128 24332 2138
rect 24280 492 24332 752
rect 24280 -1144 24332 -884
rect 24280 -3345 24332 -2520
rect 24280 -4783 24332 -4721
rect 24478 2128 24530 2134
rect 24478 492 24530 752
rect 24478 -1144 24530 -884
rect 24478 -3345 24530 -2520
rect 24478 -4731 24530 -4721
rect 24676 2128 24728 2138
rect 24676 492 24728 752
rect 24676 -1144 24728 -884
rect 24676 -3345 24728 -2520
rect 24676 -4783 24728 -4721
rect 24874 2128 24926 2134
rect 24874 492 24926 752
rect 24874 -1144 24926 -884
rect 24874 -3345 24926 -2520
rect 24874 -4731 24926 -4721
rect 25072 2128 25124 2138
rect 25072 492 25124 752
rect 25072 -1144 25124 -884
rect 25072 -3345 25124 -2520
rect 25072 -4783 25124 -4721
rect 25270 2128 25322 2134
rect 25270 492 25322 752
rect 25270 -1144 25322 -884
rect 25270 -3345 25322 -2520
rect 25270 -4731 25322 -4721
rect 25468 2128 25520 2138
rect 25468 492 25520 752
rect 25468 -1144 25520 -884
rect 25468 -3345 25520 -2520
rect 25468 -4783 25520 -4721
rect 25666 2128 25718 2134
rect 25666 492 25718 752
rect 25666 -1144 25718 -884
rect 25666 -3345 25718 -2520
rect 25666 -4731 25718 -4721
rect 25864 2128 25916 2138
rect 25864 492 25916 752
rect 25864 -1144 25916 -884
rect 25864 -3345 25916 -2520
rect 25864 -4783 25916 -4721
rect 26062 2128 26114 2134
rect 26062 492 26114 752
rect 26062 -1144 26114 -884
rect 26062 -3345 26114 -2520
rect 26062 -4731 26114 -4721
rect 26260 2128 26312 2138
rect 26260 492 26312 752
rect 26260 -1144 26312 -884
rect 26260 -3345 26312 -2520
rect 26260 -4783 26312 -4721
rect 26458 2128 26510 2134
rect 26458 492 26510 752
rect 26458 -1144 26510 -884
rect 26458 -3345 26510 -2520
rect 26458 -4731 26510 -4721
rect 26656 2128 26708 2138
rect 26656 492 26708 752
rect 26656 -1144 26708 -884
rect 26656 -3345 26708 -2520
rect 26656 -4783 26708 -4721
rect 26854 2128 26906 2134
rect 26854 492 26906 752
rect 26854 -1144 26906 -884
rect 26854 -3345 26906 -2520
rect 26854 -4731 26906 -4721
rect 27052 2128 27104 2138
rect 27052 492 27104 752
rect 27052 -1144 27104 -884
rect 27052 -3345 27104 -2520
rect 27052 -4783 27104 -4721
rect 27250 2128 27302 2134
rect 27250 492 27302 752
rect 27250 -1144 27302 -884
rect 27250 -3345 27302 -2520
rect 27250 -4731 27302 -4721
rect 27448 2128 27500 2138
rect 27448 492 27500 752
rect 27448 -1144 27500 -884
rect 27448 -3345 27500 -2520
rect 27448 -4783 27500 -4721
rect 27646 2128 27698 2134
rect 27646 492 27698 752
rect 27646 -1144 27698 -884
rect 27646 -3345 27698 -2520
rect 27646 -4731 27698 -4721
rect 27844 2128 27896 2138
rect 27844 492 27896 752
rect 27844 -1144 27896 -884
rect 27844 -3345 27896 -2520
rect 27844 -4783 27896 -4721
rect 28042 2128 28094 2134
rect 28042 492 28094 752
rect 28042 -1144 28094 -884
rect 28042 -3345 28094 -2520
rect 28042 -4731 28094 -4721
rect 28240 2128 28292 2138
rect 28240 492 28292 752
rect 28240 -1144 28292 -884
rect 28240 -3345 28292 -2520
rect 28240 -4783 28292 -4721
rect 28438 2128 28490 2134
rect 28438 492 28490 752
rect 28438 -1144 28490 -884
rect 28438 -3345 28490 -2520
rect 28438 -4731 28490 -4721
rect 28636 2128 28688 2138
rect 28636 492 28688 752
rect 28636 -1144 28688 -884
rect 28636 -3345 28688 -2520
rect 28636 -4783 28688 -4721
rect 28834 2128 28886 2134
rect 28834 492 28886 752
rect 28834 -1144 28886 -884
rect 28834 -3345 28886 -2520
rect 28834 -4731 28886 -4721
rect 29032 2128 29084 2138
rect 29032 492 29084 752
rect 29032 -1144 29084 -884
rect 29032 -3345 29084 -2520
rect 29032 -4783 29084 -4721
rect 29230 2128 29282 2134
rect 29230 492 29282 752
rect 29230 -1144 29282 -884
rect 29230 -3345 29282 -2520
rect 29230 -4731 29282 -4721
rect 29428 2128 29480 2138
rect 29428 492 29480 752
rect 29428 -1144 29480 -884
rect 29428 -3345 29480 -2520
rect 29428 -4783 29480 -4721
rect 29626 2128 29678 2134
rect 29626 492 29678 752
rect 29626 -1144 29678 -884
rect 29626 -3345 29678 -2520
rect 29626 -4731 29678 -4721
rect 29824 2128 29876 2138
rect 29824 492 29876 752
rect 29824 -1144 29876 -884
rect 29824 -3345 29876 -2520
rect 29824 -4783 29876 -4721
rect 30022 2128 30074 2134
rect 30022 492 30074 752
rect 30022 -1144 30074 -884
rect 30022 -3345 30074 -2520
rect 30022 -4731 30074 -4721
rect 30220 2128 30272 2138
rect 30220 492 30272 752
rect 30220 -1144 30272 -884
rect 30220 -3345 30272 -2520
rect 30220 -4783 30272 -4721
rect 30418 2128 30470 2134
rect 30418 492 30470 752
rect 30418 -1144 30470 -884
rect 30418 -3345 30470 -2520
rect 30418 -4731 30470 -4721
rect 30616 2128 30668 2138
rect 30616 492 30668 752
rect 30616 -1144 30668 -884
rect 30616 -3345 30668 -2520
rect 30616 -4783 30668 -4721
rect 30814 2128 30866 2134
rect 30814 492 30866 752
rect 30814 -1144 30866 -884
rect 30814 -3345 30866 -2520
rect 30814 -4731 30866 -4721
rect 31012 2128 31064 2138
rect 31012 492 31064 752
rect 31012 -1144 31064 -884
rect 31012 -3345 31064 -2520
rect 31012 -4783 31064 -4721
rect 31210 2128 31262 2134
rect 31210 492 31262 752
rect 31210 -1144 31262 -884
rect 31210 -3345 31262 -2520
rect 31210 -4731 31262 -4721
rect 31408 2128 31460 2138
rect 31408 492 31460 752
rect 31408 -1144 31460 -884
rect 31408 -3345 31460 -2520
rect 31408 -4783 31460 -4721
rect 31606 2129 31658 2135
rect 31606 493 31658 753
rect 31606 -1143 31658 -883
rect 31606 -3344 31658 -2519
rect 31606 -4730 31658 -4720
rect -225 -4805 -129 -4783
rect -225 -4861 -203 -4805
rect -147 -4861 -129 -4805
rect -225 -4879 -129 -4861
rect 171 -4805 267 -4783
rect 171 -4861 193 -4805
rect 249 -4861 267 -4805
rect 171 -4879 267 -4861
rect 567 -4805 663 -4783
rect 567 -4861 589 -4805
rect 645 -4861 663 -4805
rect 567 -4879 663 -4861
rect 963 -4805 1059 -4783
rect 963 -4861 985 -4805
rect 1041 -4861 1059 -4805
rect 963 -4879 1059 -4861
rect 1359 -4805 1455 -4783
rect 1359 -4861 1381 -4805
rect 1437 -4861 1455 -4805
rect 1359 -4879 1455 -4861
rect 1755 -4805 1851 -4783
rect 1755 -4861 1777 -4805
rect 1833 -4861 1851 -4805
rect 1755 -4879 1851 -4861
rect 2151 -4805 2247 -4783
rect 2151 -4861 2173 -4805
rect 2229 -4861 2247 -4805
rect 2151 -4879 2247 -4861
rect 2547 -4805 2643 -4783
rect 2547 -4861 2569 -4805
rect 2625 -4861 2643 -4805
rect 2547 -4879 2643 -4861
rect 2943 -4805 3039 -4783
rect 2943 -4861 2965 -4805
rect 3021 -4861 3039 -4805
rect 2943 -4879 3039 -4861
rect 3339 -4805 3435 -4783
rect 3339 -4861 3361 -4805
rect 3417 -4861 3435 -4805
rect 3339 -4879 3435 -4861
rect 3735 -4805 3831 -4783
rect 3735 -4861 3757 -4805
rect 3813 -4861 3831 -4805
rect 3735 -4879 3831 -4861
rect 4131 -4805 4227 -4783
rect 4131 -4861 4153 -4805
rect 4209 -4861 4227 -4805
rect 4131 -4879 4227 -4861
rect 4527 -4805 4623 -4783
rect 4527 -4861 4549 -4805
rect 4605 -4861 4623 -4805
rect 4527 -4879 4623 -4861
rect 4923 -4805 5019 -4783
rect 4923 -4861 4945 -4805
rect 5001 -4861 5019 -4805
rect 4923 -4879 5019 -4861
rect 5319 -4805 5415 -4783
rect 5319 -4861 5341 -4805
rect 5397 -4861 5415 -4805
rect 5319 -4879 5415 -4861
rect 5715 -4805 5811 -4783
rect 5715 -4861 5737 -4805
rect 5793 -4861 5811 -4805
rect 5715 -4879 5811 -4861
rect 6111 -4805 6207 -4783
rect 6111 -4861 6133 -4805
rect 6189 -4861 6207 -4805
rect 6111 -4879 6207 -4861
rect 6507 -4805 6603 -4783
rect 6507 -4861 6529 -4805
rect 6585 -4861 6603 -4805
rect 6507 -4879 6603 -4861
rect 6903 -4805 6999 -4783
rect 6903 -4861 6925 -4805
rect 6981 -4861 6999 -4805
rect 6903 -4879 6999 -4861
rect 7299 -4805 7395 -4783
rect 7299 -4861 7321 -4805
rect 7377 -4861 7395 -4805
rect 7299 -4879 7395 -4861
rect 7695 -4805 7791 -4783
rect 7695 -4861 7717 -4805
rect 7773 -4861 7791 -4805
rect 7695 -4879 7791 -4861
rect 11614 -4805 11710 -4783
rect 11614 -4861 11636 -4805
rect 11692 -4861 11710 -4805
rect 11614 -4879 11710 -4861
rect 12010 -4805 12106 -4783
rect 12010 -4861 12032 -4805
rect 12088 -4861 12106 -4805
rect 12010 -4879 12106 -4861
rect 12406 -4805 12502 -4783
rect 12406 -4861 12428 -4805
rect 12484 -4861 12502 -4805
rect 12406 -4879 12502 -4861
rect 12802 -4805 12898 -4783
rect 12802 -4861 12824 -4805
rect 12880 -4861 12898 -4805
rect 12802 -4879 12898 -4861
rect 13198 -4805 13294 -4783
rect 13198 -4861 13220 -4805
rect 13276 -4861 13294 -4805
rect 13198 -4879 13294 -4861
rect 13594 -4805 13690 -4783
rect 13594 -4861 13616 -4805
rect 13672 -4861 13690 -4805
rect 13594 -4879 13690 -4861
rect 13990 -4805 14086 -4783
rect 13990 -4861 14012 -4805
rect 14068 -4861 14086 -4805
rect 13990 -4879 14086 -4861
rect 14386 -4805 14482 -4783
rect 14386 -4861 14408 -4805
rect 14464 -4861 14482 -4805
rect 14386 -4879 14482 -4861
rect 14782 -4805 14878 -4783
rect 14782 -4861 14804 -4805
rect 14860 -4861 14878 -4805
rect 14782 -4879 14878 -4861
rect 15178 -4805 15274 -4783
rect 15178 -4861 15200 -4805
rect 15256 -4861 15274 -4805
rect 15178 -4879 15274 -4861
rect 15574 -4805 15670 -4783
rect 15574 -4861 15596 -4805
rect 15652 -4861 15670 -4805
rect 15574 -4879 15670 -4861
rect 15970 -4805 16066 -4783
rect 15970 -4861 15992 -4805
rect 16048 -4861 16066 -4805
rect 15970 -4879 16066 -4861
rect 16366 -4805 16462 -4783
rect 16366 -4861 16388 -4805
rect 16444 -4861 16462 -4805
rect 16366 -4879 16462 -4861
rect 16762 -4805 16858 -4783
rect 16762 -4861 16784 -4805
rect 16840 -4861 16858 -4805
rect 16762 -4879 16858 -4861
rect 17158 -4805 17254 -4783
rect 17158 -4861 17180 -4805
rect 17236 -4861 17254 -4805
rect 17158 -4879 17254 -4861
rect 17554 -4805 17650 -4783
rect 17554 -4861 17576 -4805
rect 17632 -4861 17650 -4805
rect 17554 -4879 17650 -4861
rect 17950 -4805 18046 -4783
rect 17950 -4861 17972 -4805
rect 18028 -4861 18046 -4805
rect 17950 -4879 18046 -4861
rect 18346 -4805 18442 -4783
rect 18346 -4861 18368 -4805
rect 18424 -4861 18442 -4805
rect 18346 -4879 18442 -4861
rect 18742 -4805 18838 -4783
rect 18742 -4861 18764 -4805
rect 18820 -4861 18838 -4805
rect 18742 -4879 18838 -4861
rect 19138 -4805 19234 -4783
rect 19138 -4861 19160 -4805
rect 19216 -4861 19234 -4805
rect 19138 -4879 19234 -4861
rect 19534 -4805 19630 -4783
rect 19534 -4861 19556 -4805
rect 19612 -4861 19630 -4805
rect 19534 -4879 19630 -4861
rect 23464 -4805 23560 -4783
rect 23464 -4861 23486 -4805
rect 23542 -4861 23560 -4805
rect 23464 -4879 23560 -4861
rect 23860 -4805 23956 -4783
rect 23860 -4861 23882 -4805
rect 23938 -4861 23956 -4805
rect 23860 -4879 23956 -4861
rect 24256 -4805 24352 -4783
rect 24256 -4861 24278 -4805
rect 24334 -4861 24352 -4805
rect 24256 -4879 24352 -4861
rect 24652 -4805 24748 -4783
rect 24652 -4861 24674 -4805
rect 24730 -4861 24748 -4805
rect 24652 -4879 24748 -4861
rect 25048 -4805 25144 -4783
rect 25048 -4861 25070 -4805
rect 25126 -4861 25144 -4805
rect 25048 -4879 25144 -4861
rect 25444 -4805 25540 -4783
rect 25444 -4861 25466 -4805
rect 25522 -4861 25540 -4805
rect 25444 -4879 25540 -4861
rect 25840 -4805 25936 -4783
rect 25840 -4861 25862 -4805
rect 25918 -4861 25936 -4805
rect 25840 -4879 25936 -4861
rect 26236 -4805 26332 -4783
rect 26236 -4861 26258 -4805
rect 26314 -4861 26332 -4805
rect 26236 -4879 26332 -4861
rect 26632 -4805 26728 -4783
rect 26632 -4861 26654 -4805
rect 26710 -4861 26728 -4805
rect 26632 -4879 26728 -4861
rect 27028 -4805 27124 -4783
rect 27028 -4861 27050 -4805
rect 27106 -4861 27124 -4805
rect 27028 -4879 27124 -4861
rect 27424 -4805 27520 -4783
rect 27424 -4861 27446 -4805
rect 27502 -4861 27520 -4805
rect 27424 -4879 27520 -4861
rect 27820 -4805 27916 -4783
rect 27820 -4861 27842 -4805
rect 27898 -4861 27916 -4805
rect 27820 -4879 27916 -4861
rect 28216 -4805 28312 -4783
rect 28216 -4861 28238 -4805
rect 28294 -4861 28312 -4805
rect 28216 -4879 28312 -4861
rect 28612 -4805 28708 -4783
rect 28612 -4861 28634 -4805
rect 28690 -4861 28708 -4805
rect 28612 -4879 28708 -4861
rect 29008 -4805 29104 -4783
rect 29008 -4861 29030 -4805
rect 29086 -4861 29104 -4805
rect 29008 -4879 29104 -4861
rect 29404 -4805 29500 -4783
rect 29404 -4861 29426 -4805
rect 29482 -4861 29500 -4805
rect 29404 -4879 29500 -4861
rect 29800 -4805 29896 -4783
rect 29800 -4861 29822 -4805
rect 29878 -4861 29896 -4805
rect 29800 -4879 29896 -4861
rect 30196 -4805 30292 -4783
rect 30196 -4861 30218 -4805
rect 30274 -4861 30292 -4805
rect 30196 -4879 30292 -4861
rect 30592 -4805 30688 -4783
rect 30592 -4861 30614 -4805
rect 30670 -4861 30688 -4805
rect 30592 -4879 30688 -4861
rect 30988 -4805 31084 -4783
rect 30988 -4861 31010 -4805
rect 31066 -4861 31084 -4805
rect 30988 -4879 31084 -4861
rect 31384 -4805 31480 -4783
rect 31384 -4861 31406 -4805
rect 31462 -4861 31480 -4805
rect 31384 -4879 31480 -4861
<< via2 >>
rect -627 -877 -493 -743
rect -627 -1081 -493 -947
rect -627 -1285 -493 -1151
rect 8063 -877 8197 -743
rect 11212 -877 11346 -743
rect 8063 -1081 8197 -947
rect 11212 -1081 11346 -947
rect 8063 -1285 8197 -1151
rect 11212 -1285 11346 -1151
rect 19902 -877 20036 -743
rect 23062 -877 23196 -743
rect 19902 -1081 20036 -947
rect 23062 -1081 23196 -947
rect 19902 -1285 20036 -1151
rect 23062 -1285 23196 -1151
rect -203 -4861 -147 -4805
rect 193 -4861 249 -4805
rect 589 -4861 645 -4805
rect 985 -4861 1041 -4805
rect 1381 -4861 1437 -4805
rect 1777 -4861 1833 -4805
rect 2173 -4861 2229 -4805
rect 2569 -4861 2625 -4805
rect 2965 -4861 3021 -4805
rect 3361 -4861 3417 -4805
rect 3757 -4861 3813 -4805
rect 4153 -4861 4209 -4805
rect 4549 -4861 4605 -4805
rect 4945 -4861 5001 -4805
rect 5341 -4861 5397 -4805
rect 5737 -4861 5793 -4805
rect 6133 -4861 6189 -4805
rect 6529 -4861 6585 -4805
rect 6925 -4861 6981 -4805
rect 7321 -4861 7377 -4805
rect 7717 -4861 7773 -4805
rect 11636 -4861 11692 -4805
rect 12032 -4861 12088 -4805
rect 12428 -4861 12484 -4805
rect 12824 -4861 12880 -4805
rect 13220 -4861 13276 -4805
rect 13616 -4861 13672 -4805
rect 14012 -4861 14068 -4805
rect 14408 -4861 14464 -4805
rect 14804 -4861 14860 -4805
rect 15200 -4861 15256 -4805
rect 15596 -4861 15652 -4805
rect 15992 -4861 16048 -4805
rect 16388 -4861 16444 -4805
rect 16784 -4861 16840 -4805
rect 17180 -4861 17236 -4805
rect 17576 -4861 17632 -4805
rect 17972 -4861 18028 -4805
rect 18368 -4861 18424 -4805
rect 18764 -4861 18820 -4805
rect 19160 -4861 19216 -4805
rect 19556 -4861 19612 -4805
rect 23486 -4861 23542 -4805
rect 23882 -4861 23938 -4805
rect 24278 -4861 24334 -4805
rect 24674 -4861 24730 -4805
rect 25070 -4861 25126 -4805
rect 25466 -4861 25522 -4805
rect 25862 -4861 25918 -4805
rect 26258 -4861 26314 -4805
rect 26654 -4861 26710 -4805
rect 27050 -4861 27106 -4805
rect 27446 -4861 27502 -4805
rect 27842 -4861 27898 -4805
rect 28238 -4861 28294 -4805
rect 28634 -4861 28690 -4805
rect 29030 -4861 29086 -4805
rect 29426 -4861 29482 -4805
rect 29822 -4861 29878 -4805
rect 30218 -4861 30274 -4805
rect 30614 -4861 30670 -4805
rect 31010 -4861 31066 -4805
rect 31406 -4861 31462 -4805
<< metal3 >>
rect -637 -743 -483 -738
rect -637 -877 -627 -743
rect -493 -877 -483 -743
rect -637 -882 -483 -877
rect 8053 -743 11356 -738
rect 8053 -877 8063 -743
rect 8197 -877 11212 -743
rect 11346 -877 11356 -743
rect -637 -947 -483 -942
rect -637 -1081 -627 -947
rect -493 -1081 -483 -947
rect -637 -1086 -483 -1081
rect 8053 -947 11356 -877
rect 19892 -743 23206 -738
rect 19892 -877 19902 -743
rect 20036 -877 23062 -743
rect 23196 -877 23206 -743
rect 19892 -882 23206 -877
rect 20036 -942 23062 -882
rect 8053 -1081 8063 -947
rect 8197 -1081 11212 -947
rect 11346 -1081 11356 -947
rect -637 -1151 -483 -1146
rect -637 -1285 -627 -1151
rect -493 -1285 -483 -1151
rect -637 -1290 -483 -1285
rect 8053 -1151 11356 -1081
rect 19892 -947 23206 -942
rect 19892 -1081 19902 -947
rect 20036 -1081 23062 -947
rect 23196 -1081 23206 -947
rect 19892 -1086 23206 -1081
rect 20036 -1146 23062 -1086
rect 8053 -1285 8063 -1151
rect 8197 -1285 11212 -1151
rect 11346 -1285 11356 -1151
rect 8053 -1290 11356 -1285
rect 19892 -1151 23206 -1146
rect 19892 -1285 19902 -1151
rect 20036 -1285 23062 -1151
rect 23196 -1285 23206 -1151
rect 19892 -1290 23206 -1285
rect -225 -4805 7791 -4783
rect -225 -4861 -203 -4805
rect -147 -4861 193 -4805
rect 249 -4861 589 -4805
rect 645 -4861 985 -4805
rect 1041 -4861 1381 -4805
rect 1437 -4861 1777 -4805
rect 1833 -4861 2173 -4805
rect 2229 -4861 2569 -4805
rect 2625 -4861 2965 -4805
rect 3021 -4861 3361 -4805
rect 3417 -4861 3757 -4805
rect 3813 -4861 4153 -4805
rect 4209 -4861 4549 -4805
rect 4605 -4861 4945 -4805
rect 5001 -4861 5341 -4805
rect 5397 -4861 5737 -4805
rect 5793 -4861 6133 -4805
rect 6189 -4861 6529 -4805
rect 6585 -4861 6925 -4805
rect 6981 -4861 7321 -4805
rect 7377 -4861 7717 -4805
rect 7773 -4861 7791 -4805
rect -225 -4879 7791 -4861
rect 11614 -4805 19630 -4783
rect 11614 -4861 11636 -4805
rect 11692 -4861 12032 -4805
rect 12088 -4861 12428 -4805
rect 12484 -4861 12824 -4805
rect 12880 -4861 13220 -4805
rect 13276 -4861 13616 -4805
rect 13672 -4861 14012 -4805
rect 14068 -4861 14408 -4805
rect 14464 -4861 14804 -4805
rect 14860 -4861 15200 -4805
rect 15256 -4861 15596 -4805
rect 15652 -4861 15992 -4805
rect 16048 -4861 16388 -4805
rect 16444 -4861 16784 -4805
rect 16840 -4861 17180 -4805
rect 17236 -4861 17576 -4805
rect 17632 -4861 17972 -4805
rect 18028 -4861 18368 -4805
rect 18424 -4861 18764 -4805
rect 18820 -4861 19160 -4805
rect 19216 -4861 19556 -4805
rect 19612 -4861 19630 -4805
rect 11614 -4879 19630 -4861
rect 23464 -4805 31480 -4783
rect 23464 -4861 23486 -4805
rect 23542 -4861 23882 -4805
rect 23938 -4861 24278 -4805
rect 24334 -4861 24674 -4805
rect 24730 -4861 25070 -4805
rect 25126 -4861 25466 -4805
rect 25522 -4861 25862 -4805
rect 25918 -4861 26258 -4805
rect 26314 -4861 26654 -4805
rect 26710 -4861 27050 -4805
rect 27106 -4861 27446 -4805
rect 27502 -4861 27842 -4805
rect 27898 -4861 28238 -4805
rect 28294 -4861 28634 -4805
rect 28690 -4861 29030 -4805
rect 29086 -4861 29426 -4805
rect 29482 -4861 29822 -4805
rect 29878 -4861 30218 -4805
rect 30274 -4861 30614 -4805
rect 30670 -4861 31010 -4805
rect 31066 -4861 31406 -4805
rect 31462 -4861 31480 -4805
rect 23464 -4879 31480 -4861
use sky130_fd_pr__pfet_01v8_ZYZ5C6  sky130_fd_pr__pfet_01v8_ZYZ5C6_0
timestamp 1615920820
transform 1 0 3785 0 1 1404
box -4223 -764 4223 798
use sky130_fd_pr__pfet_01v8_9JQ4XZ  sky130_fd_pr__pfet_01v8_9JQ4XZ_0
timestamp 1615920820
transform 1 0 3785 0 1 -1014
box -4223 -1618 4223 1618
use sky130_fd_pr__pfet_01v8_ZYZ5C6  sky130_fd_pr__pfet_01v8_ZYZ5C6_1
timestamp 1615920820
transform -1 0 3785 0 -1 -3997
box -4223 -764 4223 798
<< end >>
