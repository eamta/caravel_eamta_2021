magic
tech sky130A
magscale 1 2
timestamp 1615566114
<< nmos >>
rect -15 -96 15 84
<< ndiff >>
rect -73 72 -15 84
rect -73 -48 -61 72
rect -27 -48 -15 72
rect -73 -96 -15 -48
rect 15 72 73 84
rect 15 -48 27 72
rect 61 -48 73 72
rect 15 -96 73 -48
<< ndiffc >>
rect -61 -48 -27 72
rect 27 -48 61 72
<< poly >>
rect -15 84 15 110
rect -15 -122 15 -96
<< locali >>
rect -61 72 -27 88
rect -61 -100 -27 -48
rect 27 72 61 88
rect 27 -100 61 -48
<< viali >>
rect -61 -48 -27 72
rect 27 -48 61 72
<< metal1 >>
rect -67 72 -21 84
rect -67 -48 -61 72
rect -27 -48 -21 72
rect -67 -60 -21 -48
rect 21 72 67 84
rect 21 -48 27 72
rect 61 -48 67 72
rect 21 -60 67 -48
rect -67 -116 67 -88
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.9 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
