magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 3680 2021 3715 2055
rect 3681 2002 3715 2021
rect 4067 2002 4120 2003
rect 3511 1953 3569 1959
rect 3511 1919 3523 1953
rect 3511 1913 3569 1919
rect 1888 1797 1923 1831
rect 418 1763 453 1781
rect 382 1748 453 1763
rect 733 1748 768 1782
rect 1889 1778 1923 1797
rect 195 1625 253 1631
rect 195 1591 207 1625
rect 195 1585 253 1591
rect 382 1510 452 1748
rect 734 1729 768 1748
rect 1908 1735 1923 1778
rect 753 1686 768 1729
rect 564 1680 622 1686
rect 564 1646 576 1680
rect 564 1640 622 1646
rect 0 1472 452 1510
rect 532 1472 566 1506
rect 620 1472 654 1506
rect 734 1472 768 1686
rect 787 1695 822 1729
rect 787 1472 821 1695
rect 933 1627 991 1633
rect 933 1593 945 1627
rect 1103 1604 1137 1633
rect 933 1587 991 1593
rect 1103 1568 1173 1604
rect 1103 1534 1191 1568
rect 1471 1534 1506 1568
rect 1103 1510 1190 1534
rect 1472 1515 1506 1534
rect 1537 1551 1542 1604
rect 1573 1551 1607 1735
rect 1719 1729 1777 1735
rect 1719 1695 1731 1729
rect 1719 1689 1777 1695
rect 1889 1569 1923 1735
rect 1942 1744 1977 1778
rect 2257 1744 2292 1778
rect 1889 1551 1929 1569
rect 1537 1536 1929 1551
rect 1537 1515 1928 1536
rect 1491 1510 1506 1515
rect 1525 1510 1928 1515
rect 901 1472 935 1506
rect 989 1472 1023 1506
rect 1103 1472 1928 1510
rect 1942 1472 1976 1744
rect 2258 1725 2292 1744
rect 2277 1697 2292 1725
rect 2311 1697 2346 1725
rect 2407 1697 2565 1725
rect 2359 1691 2565 1697
rect 2626 1691 2661 1725
rect 2088 1676 2146 1682
rect 2088 1642 2100 1676
rect 2258 1663 2292 1682
rect 2359 1663 2517 1691
rect 2088 1636 2146 1642
rect 2056 1570 2090 1599
rect 1990 1536 2010 1570
rect 2044 1536 2190 1570
rect 2224 1536 2244 1570
rect 2044 1502 2133 1515
rect 2176 1506 2178 1536
rect 2185 1506 2190 1536
rect 2018 1472 2133 1502
rect 2144 1472 2206 1506
rect -1334 1421 -1299 1455
rect -1333 1402 -1299 1421
rect 0 1438 2206 1472
rect 2210 1472 2244 1536
rect 2210 1438 2212 1472
rect 2224 1438 2248 1472
rect -947 1402 -894 1403
rect -1503 1353 -1445 1359
rect -1503 1319 -1491 1353
rect -1503 1313 -1445 1319
rect -1685 1214 -1387 1267
rect -1314 1214 -1299 1402
rect -1280 1368 -1245 1402
rect -965 1368 -894 1402
rect -1280 1214 -1246 1368
rect -964 1367 -894 1368
rect -947 1333 -876 1367
rect -596 1333 -561 1367
rect -1134 1300 -1076 1306
rect -1134 1266 -1122 1300
rect -1134 1260 -1076 1266
rect -1685 1161 -1018 1214
rect -947 1161 -877 1333
rect -595 1314 -561 1333
rect 0 1366 452 1438
rect 520 1419 560 1438
rect 598 1419 666 1438
rect 536 1400 650 1406
rect 576 1384 620 1390
rect 545 1372 657 1384
rect 464 1366 480 1372
rect 545 1369 660 1372
rect 0 1356 490 1366
rect 0 1346 496 1356
rect 0 1340 452 1346
rect 0 1332 444 1340
rect -576 1271 -561 1314
rect -765 1265 -707 1271
rect -765 1231 -753 1265
rect -765 1225 -707 1231
rect -1685 1125 -877 1161
rect -1685 1106 -685 1125
rect -1685 1091 -675 1106
rect -1685 1029 -877 1091
rect -809 1057 -796 1070
rect -1685 1023 -831 1029
rect -1685 989 -877 1023
rect -831 989 -827 1023
rect -809 1004 -793 1057
rect -797 1000 -793 1004
rect -719 1000 -675 1091
rect -595 1072 -561 1271
rect -542 1280 -507 1314
rect -227 1280 -192 1314
rect 0 1297 435 1332
rect -542 1072 -508 1280
rect -226 1261 -192 1280
rect -396 1212 -338 1218
rect -396 1178 -384 1212
rect -396 1172 -338 1178
rect -666 1004 -641 1072
rect -595 1038 -316 1072
rect -1685 983 -831 989
rect -1685 964 -877 983
rect -1685 917 -853 964
rect -719 963 -685 1000
rect -765 957 -685 963
rect -1685 891 -877 917
rect -803 906 -799 946
rect -769 938 -740 957
rect -719 938 -685 957
rect -769 923 -685 938
rect -765 917 -685 923
rect -719 910 -685 917
rect -1654 872 -1625 891
rect -1571 880 -1537 891
rect -1457 872 -1423 891
rect -1404 872 -1370 891
rect -1316 872 -877 891
rect -833 872 -799 906
rect -793 889 -679 910
rect -719 872 -685 889
rect -666 872 -632 1004
rect -595 872 -561 1038
rect -542 976 -508 1038
rect -350 1037 -316 1038
rect -207 1037 -192 1261
rect -173 1227 -138 1261
rect 13 1253 435 1297
rect 446 1270 452 1340
rect 470 1340 496 1346
rect 470 1322 490 1340
rect 560 1338 660 1369
rect 665 1356 686 1384
rect 734 1366 768 1438
rect 787 1384 821 1438
rect 926 1410 935 1438
rect 872 1390 901 1396
rect 918 1390 947 1410
rect 872 1384 947 1390
rect 702 1356 768 1366
rect 696 1346 768 1356
rect 696 1340 733 1346
rect 560 1332 622 1338
rect 560 1322 598 1332
rect 640 1306 660 1338
rect 712 1322 733 1340
rect 734 1340 768 1346
rect 734 1332 746 1340
rect 747 1332 768 1340
rect 734 1322 768 1332
rect 734 1270 746 1322
rect 446 1259 491 1270
rect 36 1227 177 1253
rect 418 1236 422 1253
rect 446 1247 480 1259
rect 435 1236 491 1247
rect 540 1236 686 1270
rect 701 1259 746 1270
rect 712 1247 746 1259
rect 747 1247 768 1322
rect 701 1236 768 1247
rect 772 1236 822 1384
rect 872 1378 935 1384
rect 872 1372 901 1378
rect 926 1362 935 1378
rect 960 1367 969 1438
rect 1010 1390 1035 1438
rect 989 1384 1035 1390
rect 1103 1384 1928 1438
rect 1942 1415 1976 1438
rect 2044 1434 2120 1438
rect 2044 1415 2102 1434
rect 2130 1415 2190 1438
rect 1942 1402 2164 1415
rect 2176 1411 2178 1415
rect 2172 1402 2174 1410
rect 1942 1400 2174 1402
rect 989 1378 1023 1384
rect 949 1366 977 1367
rect 1064 1366 1089 1384
rect 895 1306 906 1353
rect 948 1325 1006 1366
rect 933 1319 1006 1325
rect 929 1285 1006 1319
rect 933 1279 995 1285
rect 948 1269 995 1279
rect -173 1037 -139 1227
rect -27 1163 31 1165
rect 48 1163 69 1193
rect 143 1163 177 1227
rect 364 1225 422 1236
rect 285 1204 422 1225
rect 540 1204 598 1236
rect 628 1204 686 1236
rect 772 1217 821 1236
rect 1103 1232 1940 1384
rect 1942 1366 1976 1400
rect 2008 1387 2010 1391
rect 2022 1387 2042 1391
rect 2066 1387 2130 1400
rect 2172 1387 2174 1400
rect 1996 1366 2049 1387
rect 2066 1384 2142 1387
rect 2066 1372 2181 1384
rect 1942 1356 2049 1366
rect 2050 1368 2181 1372
rect 2050 1356 2072 1368
rect 1942 1346 2072 1356
rect 1942 1322 1987 1346
rect 1996 1322 2072 1346
rect 2084 1356 2181 1368
rect 2084 1334 2150 1356
rect 1942 1266 1976 1322
rect 1996 1266 2002 1322
rect 2008 1300 2042 1322
rect 2050 1306 2072 1322
rect 2096 1322 2160 1334
rect 2096 1318 2150 1322
rect 2004 1266 2042 1300
rect 2096 1266 2130 1318
rect 2210 1306 2248 1438
rect 2210 1266 2244 1306
rect 2258 1266 2297 1663
rect 1942 1232 2260 1266
rect 1103 1217 1928 1232
rect 772 1212 1006 1217
rect 1064 1212 1928 1217
rect 772 1198 1928 1212
rect 1996 1222 2002 1232
rect 1996 1207 2017 1222
rect 2096 1219 2114 1232
rect 364 1188 366 1194
rect 322 1178 334 1188
rect 364 1178 376 1188
rect 772 1183 1911 1198
rect 316 1174 344 1178
rect 354 1174 382 1178
rect 316 1163 382 1174
rect 418 1171 491 1182
rect 540 1179 686 1182
rect 523 1178 553 1179
rect 418 1163 480 1171
rect -27 1159 480 1163
rect 522 1159 554 1178
rect 587 1171 639 1179
rect 701 1178 768 1182
rect 772 1178 822 1183
rect 1120 1178 1911 1183
rect 701 1171 1911 1178
rect 2054 1176 2084 1207
rect 598 1159 628 1171
rect 712 1159 746 1171
rect -27 1125 -15 1159
rect 2 1154 491 1159
rect 522 1154 565 1159
rect 2 1148 565 1154
rect 587 1148 639 1159
rect 701 1148 746 1159
rect 2 1136 452 1148
rect 522 1144 533 1148
rect 543 1144 564 1148
rect 553 1138 564 1144
rect 523 1136 564 1138
rect 2 1127 582 1136
rect 13 1125 582 1127
rect -27 1119 582 1125
rect 13 1100 582 1119
rect 628 1110 630 1116
rect 586 1100 598 1110
rect 628 1100 640 1110
rect 13 1084 646 1100
rect 734 1086 746 1148
rect 747 1144 1911 1171
rect 747 1086 768 1144
rect 13 1066 640 1084
rect 13 1060 610 1066
rect 626 1060 640 1066
rect 13 1056 640 1060
rect 13 1050 630 1056
rect 13 1040 626 1050
rect 13 1037 595 1040
rect -350 1018 595 1037
rect 608 1030 626 1040
rect -440 1004 -427 1017
rect -542 970 -462 976
rect -542 938 -508 970
rect -462 938 -458 970
rect -440 951 -424 1004
rect -428 947 -424 951
rect -350 986 582 1018
rect -350 976 250 986
rect 338 982 354 986
rect 365 982 582 986
rect -350 975 264 976
rect -350 948 319 975
rect 338 964 582 982
rect 342 958 582 964
rect 365 948 582 958
rect -542 936 -458 938
rect -350 942 297 948
rect 304 942 582 948
rect -350 941 582 942
rect -542 930 -462 936
rect -542 911 -508 930
rect -350 926 297 941
rect 304 931 582 941
rect 608 984 643 999
rect 608 931 628 984
rect 734 931 768 1086
rect 772 1129 822 1144
rect 1120 1129 1911 1144
rect 772 1110 1911 1129
rect 2036 1166 2084 1176
rect 2086 1166 2133 1207
rect 2036 1126 2133 1166
rect 2036 1120 2098 1126
rect 772 1095 1006 1110
rect 1120 1100 1911 1110
rect 1917 1100 1928 1111
rect 2036 1110 2084 1120
rect 772 1055 822 1095
rect 1120 1094 1928 1100
rect 772 1024 909 1055
rect 979 1043 1006 1074
rect 948 1033 1006 1043
rect 933 1024 1006 1033
rect 787 1018 821 1024
rect 860 1018 862 1024
rect 787 1008 830 1018
rect 860 1008 872 1018
rect 787 992 878 1008
rect 933 993 945 1024
rect 948 993 995 1024
rect 1122 1022 1137 1094
rect 1388 1076 1398 1094
rect 1408 1090 1436 1094
rect 1410 1084 1436 1090
rect 1410 1076 1430 1084
rect 1388 1066 1430 1076
rect 1404 1056 1430 1066
rect 1489 1058 1928 1094
rect 2210 1058 2260 1232
rect 1404 1050 1420 1056
rect 1489 1047 2013 1058
rect 1489 1042 2002 1047
rect 2026 1042 2260 1058
rect 1489 1041 2260 1042
rect 1894 1024 2260 1041
rect 2263 1097 2297 1266
rect 2311 1348 2345 1663
rect 2437 1611 2453 1623
rect 2437 1601 2457 1611
rect 2437 1595 2453 1601
rect 2421 1580 2423 1589
rect 2431 1580 2455 1595
rect 2469 1589 2493 1623
rect 2593 1601 2613 1691
rect 2405 1561 2471 1580
rect 2409 1555 2467 1561
rect 2425 1542 2459 1546
rect 2471 1542 2495 1545
rect 2513 1542 2533 1546
rect 2413 1530 2471 1542
rect 2507 1530 2533 1542
rect 2413 1527 2468 1530
rect 2377 1514 2379 1518
rect 2391 1514 2411 1518
rect 2365 1510 2417 1514
rect 2419 1510 2459 1527
rect 2365 1472 2411 1510
rect 2425 1472 2459 1510
rect 2465 1514 2499 1518
rect 2465 1510 2505 1514
rect 2507 1510 2537 1530
rect 2465 1472 2499 1510
rect 2513 1506 2537 1510
rect 2545 1506 2547 1546
rect 2513 1472 2547 1506
rect 2554 1472 2559 1542
rect 2579 1472 2613 1601
rect 2627 1644 2661 1691
rect 2680 1644 2715 1672
rect 2776 1644 2934 1672
rect 3511 1663 3569 1669
rect 2627 1610 2667 1644
rect 2728 1638 2934 1644
rect 2995 1638 3030 1655
rect 2728 1610 2886 1638
rect 2627 1472 2666 1610
rect 2680 1483 2714 1610
rect 2806 1558 2822 1570
rect 2806 1548 2826 1558
rect 2806 1542 2822 1548
rect 2790 1527 2792 1536
rect 2800 1527 2824 1542
rect 2838 1538 2862 1570
rect 2962 1548 2982 1638
rect 2836 1530 2884 1538
rect 2774 1510 2840 1527
rect 2774 1508 2912 1510
rect 2836 1506 2912 1508
rect 2794 1489 2828 1506
rect 2836 1502 2916 1506
rect 2840 1489 2864 1492
rect 2782 1483 2840 1489
rect 2882 1483 2916 1502
rect 2680 1472 2916 1483
rect 2923 1472 2928 1489
rect 2948 1472 2982 1548
rect 2996 1637 3030 1638
rect 2996 1601 3066 1637
rect 3511 1629 3523 1663
rect 3511 1623 3569 1629
rect 2996 1567 3084 1601
rect 2996 1510 3083 1567
rect 3461 1548 3619 1561
rect 3700 1548 3715 2002
rect 3734 1968 3769 2002
rect 4049 1968 4120 2002
rect 3734 1548 3768 1968
rect 4050 1967 4120 1968
rect 4067 1933 4138 1967
rect 4418 1933 4453 1967
rect 3880 1900 3938 1906
rect 3880 1866 3892 1900
rect 3880 1860 3938 1866
rect 3880 1610 3938 1616
rect 3880 1576 3892 1610
rect 3880 1570 3938 1576
rect 3461 1527 3672 1548
rect 3384 1510 3399 1527
rect 3418 1526 3453 1527
rect 3514 1526 3672 1527
rect 4067 1531 4137 1933
rect 4419 1914 4453 1933
rect 4249 1865 4307 1871
rect 4249 1831 4261 1865
rect 4249 1825 4307 1831
rect 4249 1557 4307 1563
rect 3418 1514 3734 1526
rect 3418 1510 3452 1514
rect 2996 1508 3964 1510
rect 2996 1495 3988 1508
rect 2996 1472 4041 1495
rect 2352 1461 4041 1472
rect 4067 1478 4173 1531
rect 4249 1523 4261 1557
rect 4249 1517 4307 1523
rect 4438 1478 4453 1914
rect 4472 1880 4507 1914
rect 4787 1880 4822 1914
rect 4472 1478 4506 1880
rect 4788 1861 4822 1880
rect 4618 1812 4676 1818
rect 4618 1778 4630 1812
rect 4618 1772 4676 1778
rect 4618 1504 4676 1510
rect 2352 1438 3964 1461
rect 2365 1400 2411 1438
rect 2425 1400 2459 1438
rect 2365 1374 2417 1400
rect 2419 1374 2459 1400
rect 2465 1402 2499 1438
rect 2513 1402 2537 1438
rect 2545 1402 2547 1438
rect 2554 1402 2559 1438
rect 2365 1362 2445 1374
rect 2365 1348 2420 1362
rect 2425 1358 2445 1362
rect 2432 1349 2445 1358
rect 2465 1362 2559 1402
rect 2465 1349 2511 1362
rect 2513 1358 2547 1362
rect 2432 1348 2511 1349
rect 2311 1320 2351 1348
rect 2377 1334 2417 1348
rect 2377 1320 2411 1334
rect 2311 1286 2411 1320
rect 2311 1213 2351 1286
rect 2377 1247 2411 1286
rect 2373 1213 2411 1247
rect 2423 1315 2511 1348
rect 2532 1336 2565 1348
rect 2532 1315 2578 1336
rect 2423 1281 2578 1315
rect 2423 1265 2511 1281
rect 2423 1213 2453 1265
rect 2496 1250 2511 1265
rect 2532 1265 2534 1281
rect 2544 1265 2578 1281
rect 2465 1213 2499 1247
rect 2532 1236 2578 1265
rect 2532 1213 2565 1236
rect 2579 1213 2613 1438
rect 2627 1213 2666 1438
rect 2311 1179 2511 1213
rect 2532 1179 2666 1213
rect 2332 1168 2351 1179
rect 2390 1169 2411 1179
rect 2423 1169 2453 1179
rect 2377 1168 2411 1169
rect 2420 1168 2453 1169
rect 2532 1168 2565 1179
rect 2377 1166 2423 1168
rect 2375 1154 2423 1166
rect 2423 1131 2453 1154
rect 2421 1113 2455 1131
rect 2579 1116 2613 1179
rect 2409 1107 2467 1113
rect 2409 1097 2421 1107
rect 2579 1097 2630 1116
rect 2263 1063 2314 1097
rect 2379 1086 2482 1097
rect 2549 1086 2630 1097
rect 2390 1074 2471 1086
rect 2560 1082 2630 1086
rect 2379 1063 2482 1074
rect 2560 1066 2613 1082
rect 1103 1004 1137 1022
rect 2202 1016 2204 1022
rect 2160 1008 2172 1016
rect 2202 1008 2214 1016
rect 787 931 821 992
rect 828 984 872 992
rect 933 987 991 993
rect 1103 986 1542 1004
rect 828 974 1057 984
rect 1103 974 1540 986
rect 1860 974 2220 1008
rect 2263 1005 2297 1063
rect 860 964 874 974
rect 1103 968 1173 974
rect 2202 970 2214 974
rect 2263 971 2298 1005
rect 2379 994 2482 1005
rect 2390 990 2471 994
rect 2390 982 2512 990
rect 2379 976 2523 982
rect 2590 976 2613 1066
rect 2632 1044 2666 1179
rect 2680 1214 2714 1438
rect 2734 1400 2780 1438
rect 2794 1400 2828 1438
rect 2734 1367 2786 1400
rect 2788 1367 2828 1400
rect 2834 1404 2868 1438
rect 2834 1400 2870 1404
rect 2882 1400 2906 1438
rect 2914 1404 2916 1438
rect 2834 1367 2874 1400
rect 2876 1367 2906 1400
rect 2923 1389 2928 1438
rect 2917 1370 2928 1389
rect 2734 1354 2906 1367
rect 2914 1354 2928 1370
rect 2734 1348 2928 1354
rect 2746 1336 2920 1348
rect 2720 1321 2920 1336
rect 2720 1309 2902 1321
rect 2914 1309 2920 1321
rect 2720 1281 2792 1309
rect 2794 1305 2920 1309
rect 2720 1236 2780 1281
rect 2786 1268 2792 1281
rect 2802 1281 2920 1305
rect 2802 1278 2870 1281
rect 2872 1278 2920 1281
rect 2802 1270 2920 1278
rect 2948 1339 2982 1438
rect 2996 1399 3964 1438
rect 2996 1383 3991 1399
rect 4067 1385 4542 1478
rect 4618 1470 4630 1504
rect 4618 1464 4676 1470
rect 4807 1407 4822 1861
rect 4841 1827 4876 1861
rect 4841 1407 4875 1827
rect 4987 1759 5045 1765
rect 4987 1725 4999 1759
rect 5157 1736 5191 1754
rect 4987 1719 5045 1725
rect 5157 1700 5227 1736
rect 5174 1666 5245 1700
rect 4987 1451 5045 1457
rect 4987 1417 4999 1451
rect 4987 1411 5045 1417
rect 4621 1402 4779 1407
rect 2996 1359 3975 1383
rect 2996 1353 3991 1359
rect 2996 1339 3964 1353
rect 2804 1262 2919 1270
rect 2680 1168 2734 1214
rect 2746 1194 2780 1236
rect 2742 1168 2780 1194
rect 2680 1160 2714 1168
rect 2734 1160 2780 1168
rect 2822 1228 2919 1262
rect 2822 1214 2888 1228
rect 2822 1212 2932 1214
rect 2822 1194 2836 1212
rect 2822 1160 2868 1194
rect 2880 1168 2932 1212
rect 2948 1197 3964 1339
rect 4122 1288 4137 1385
rect 4156 1288 4190 1385
rect 4302 1340 4360 1346
rect 4436 1345 4542 1385
rect 4568 1373 4779 1402
rect 4840 1373 4875 1407
rect 4568 1368 4731 1373
rect 4573 1345 4731 1368
rect 4302 1306 4314 1340
rect 4436 1332 4559 1345
rect 4302 1300 4360 1306
rect 4441 1288 4559 1332
rect 4072 1197 4559 1288
rect 4651 1293 4667 1305
rect 4651 1283 4671 1293
rect 4651 1277 4667 1283
rect 4635 1262 4637 1271
rect 4645 1262 4669 1277
rect 4683 1271 4707 1305
rect 4807 1278 4827 1373
rect 4619 1243 4685 1262
rect 4623 1237 4681 1243
rect 4639 1224 4673 1228
rect 4685 1224 4709 1227
rect 4727 1224 4747 1228
rect 4627 1212 4685 1224
rect 4721 1212 4747 1224
rect 4627 1209 4682 1212
rect 2948 1163 4035 1197
rect 4069 1163 4559 1197
rect 4591 1196 4593 1200
rect 4605 1196 4625 1200
rect 2948 1160 3964 1163
rect 2680 1143 3964 1160
rect 2680 1126 2720 1143
rect 2734 1141 3964 1143
rect 2734 1132 3351 1141
rect 2734 1129 3083 1132
rect 3111 1129 3149 1132
rect 3203 1129 3240 1132
rect 2734 1126 3069 1129
rect 2822 1116 2836 1126
rect 2948 1116 3069 1126
rect 2822 1101 2851 1116
rect 2912 1092 3066 1116
rect 3078 1107 3083 1129
rect 3103 1114 3161 1129
rect 3191 1116 3249 1129
rect 3103 1107 3149 1114
rect 3156 1107 3161 1114
rect 3172 1107 3249 1116
rect 3264 1107 3271 1132
rect 3283 1107 3298 1132
rect 3317 1107 3351 1132
rect 3365 1107 3404 1141
rect 2912 1082 2928 1092
rect 2948 1090 3066 1092
rect 3103 1096 3263 1107
rect 2774 1060 2778 1070
rect 2790 1060 2824 1078
rect 2948 1066 3035 1090
rect 3049 1084 3050 1090
rect 3103 1084 3252 1096
rect 3049 1082 3061 1084
rect 3049 1078 3069 1082
rect 3103 1078 3263 1084
rect 3049 1073 3264 1078
rect 3317 1073 3337 1107
rect 3156 1066 3161 1073
rect 3191 1066 3249 1073
rect 2774 1054 2836 1060
rect 2774 1044 2790 1054
rect 2948 1044 2962 1066
rect 2632 1033 2758 1044
rect 2763 1033 2851 1044
rect 2921 1033 2962 1044
rect 2632 1021 2666 1033
rect 2670 1021 2758 1033
rect 2774 1021 2840 1033
rect 2932 1021 2962 1033
rect 2632 1014 2758 1021
rect 2632 976 2647 1014
rect 2659 1010 2758 1014
rect 2763 1010 2851 1021
rect 2921 1010 2962 1021
rect 2659 983 2666 1010
rect 2774 1004 2778 1010
rect 2948 976 2962 1010
rect 2379 971 2579 976
rect 860 958 862 964
rect 867 962 874 964
rect 901 946 935 950
rect 895 940 947 946
rect 989 940 1023 950
rect 1120 940 1506 968
rect 1894 951 2244 970
rect 1858 940 2244 951
rect 895 934 902 940
rect 903 931 947 940
rect 304 930 827 931
rect 334 926 827 930
rect -350 914 827 926
rect -542 910 -484 911
rect -350 910 231 914
rect 239 910 250 914
rect 251 910 291 914
rect 298 910 356 914
rect 365 910 827 914
rect -548 906 -434 910
rect -350 906 827 910
rect 918 906 947 931
rect 1120 934 1201 940
rect 1225 934 1281 940
rect 1377 934 1429 940
rect 1120 910 1190 934
rect 1256 910 1270 924
rect 1388 910 1406 924
rect 1502 910 1506 940
rect 1526 915 1546 940
rect 1858 915 1911 940
rect 1957 936 2013 940
rect 2084 936 2129 940
rect 2161 936 2213 940
rect 1525 910 1911 915
rect 1120 906 1911 910
rect -552 902 -430 906
rect -384 904 827 906
rect -552 872 -484 902
rect -464 872 -430 902
rect -400 872 -396 904
rect -384 872 -371 904
rect -350 878 827 904
rect 901 878 947 906
rect 989 878 1023 906
rect 1103 878 1911 906
rect 1994 884 2002 926
rect 2084 906 2094 936
rect 2108 916 2128 936
rect 2104 906 2128 916
rect 2114 902 2128 906
rect 2018 896 2128 902
rect 2018 884 2120 896
rect 2210 884 2213 936
rect -350 874 1911 878
rect 1928 874 2213 884
rect -350 872 2213 874
rect -1654 870 -418 872
rect -411 870 2213 872
rect -1654 868 2213 870
rect -1654 864 -1583 868
rect -1627 859 -1583 864
rect -1575 861 2213 868
rect 2229 884 2244 940
rect 2263 888 2297 971
rect 2371 927 2378 971
rect 2405 961 2421 971
rect 2464 961 2579 971
rect 2409 955 2579 961
rect 2464 952 2579 955
rect 2444 940 2579 952
rect 2423 914 2453 924
rect 2464 914 2579 940
rect 2375 902 2423 914
rect 2453 909 2579 914
rect 2464 908 2579 909
rect 2590 974 2647 976
rect 2590 948 2632 974
rect 2590 908 2647 948
rect 2666 908 2962 976
rect 2965 1044 3035 1066
rect 3222 1054 3249 1066
rect 3207 1044 3249 1054
rect 3264 1044 3271 1073
rect 2965 1039 3115 1044
rect 3149 1039 3203 1044
rect 3207 1039 3264 1044
rect 2965 946 3035 1039
rect 3222 1035 3251 1039
rect 3109 1010 3251 1035
rect 3147 1001 3205 1007
rect 3143 976 3209 1001
rect 3147 967 3159 976
rect 3147 961 3205 967
rect 3052 946 3054 961
rect 3222 951 3251 1010
rect 2965 940 3054 946
rect 2965 908 3035 940
rect 2465 906 2499 908
rect 2377 899 2423 902
rect 2263 884 2365 888
rect -1575 859 2210 861
rect -1627 849 2210 859
rect -1627 838 2213 849
rect -1620 830 -1591 838
rect -1624 804 -1565 821
rect -1624 783 -1574 804
rect -1566 787 -1565 804
rect -1632 771 -1574 783
rect -1532 771 -1531 787
rect -1632 768 -1631 771
rect -1620 749 -1586 771
rect -1457 719 -1423 838
rect -1632 685 -1486 719
rect -1454 685 -1423 719
rect -1420 666 -1370 838
rect -1302 815 -1232 837
rect -1290 811 -1264 815
rect -1216 809 -1214 838
rect -1196 815 -1156 837
rect -1324 777 -1298 787
rect -1220 783 -1178 802
rect -1174 783 -1154 809
rect -1293 768 -1286 783
rect -1246 734 -1239 768
rect -1232 734 -1173 783
rect -1232 718 -1196 734
rect -1232 703 -1217 718
rect -1122 700 -1098 787
rect -1132 666 -1098 700
rect -1088 666 -1054 838
rect -1420 651 -1286 666
rect -1404 632 -1286 651
rect -1232 632 -1086 666
rect -1069 632 -1054 666
rect -1035 748 -1001 838
rect -911 821 -632 838
rect -586 821 -561 838
rect -933 762 -875 802
rect -868 762 -787 802
rect -833 758 -799 762
rect -1035 632 -1000 748
rect -890 733 -868 748
rect -875 731 -868 733
rect -893 721 -868 731
rect -814 736 -796 748
rect -814 724 -768 736
rect -893 715 -831 721
rect -893 681 -868 715
rect -836 681 -827 715
rect -814 681 -793 724
rect -893 675 -831 681
rect -893 665 -868 675
rect -883 650 -868 665
rect -814 650 -812 681
rect -802 647 -793 681
rect -719 670 -680 821
rect -1220 599 -1186 632
rect -1035 598 -1020 632
rect -1014 613 -1001 632
rect -719 613 -685 670
rect -1014 579 -868 613
rect -814 579 -685 613
rect -666 614 -632 821
rect -552 802 -508 838
rect -480 802 -430 836
rect -350 816 2054 838
rect 2062 816 2072 825
rect 2084 816 2213 838
rect 2229 820 2365 884
rect 2390 824 2420 899
rect 2377 820 2420 824
rect 2465 820 2499 824
rect 2229 816 2328 820
rect -350 802 1928 816
rect -564 784 1928 802
rect 1930 804 2008 816
rect 2026 815 2084 816
rect 2014 804 2164 815
rect 1930 800 2164 804
rect 1930 788 2008 800
rect 1940 787 2012 788
rect 2026 787 2040 800
rect 2054 787 2084 800
rect 2096 787 2106 791
rect 1940 784 2142 787
rect 2210 784 2248 816
rect 2260 784 2328 816
rect 2332 790 2351 820
rect 2365 806 2499 820
rect 2532 806 2565 908
rect 2365 790 2500 806
rect -564 768 1940 784
rect -564 767 -526 768
rect -626 636 -598 736
rect -591 720 -580 748
rect -564 734 -510 767
rect -564 709 -506 734
rect -464 721 -430 754
rect -429 748 -418 768
rect -350 748 1940 768
rect -418 743 -414 748
rect -384 743 1940 748
rect -350 736 1940 743
rect -372 734 1940 736
rect -350 726 1940 734
rect 1968 726 2260 784
rect 2263 756 2282 784
rect 2332 756 2500 790
rect -556 684 -506 709
rect -472 696 -427 709
rect -544 670 -510 684
rect -472 670 -426 696
rect -350 672 1928 726
rect 1968 722 2072 726
rect 1940 672 1968 698
rect 1996 672 2002 722
rect 2008 672 2042 722
rect 2062 706 2072 722
rect 2096 722 2160 726
rect 2096 672 2130 722
rect 2210 672 2260 726
rect -472 668 -427 670
rect -520 662 -427 668
rect -524 636 -427 662
rect -520 628 -508 636
rect -472 628 -427 636
rect -350 647 1940 672
rect 1957 661 2260 672
rect 1968 649 2260 661
rect 1957 647 2260 649
rect -350 638 2260 647
rect -350 629 1940 638
rect 1996 629 2026 638
rect 2096 629 2114 638
rect 2210 629 2260 638
rect 2263 726 2282 754
rect 2332 731 2351 756
rect 2365 731 2478 756
rect 2332 730 2478 731
rect 2263 629 2297 726
rect 2390 706 2420 730
rect 2377 704 2420 706
rect 2326 672 2365 698
rect 2377 672 2411 704
rect 2432 672 2445 730
rect 2532 729 2578 806
rect 2579 729 2613 908
rect 2632 729 2666 908
rect 2738 902 2836 908
rect 2738 861 2834 902
rect 2874 861 2875 908
rect 2948 899 3035 908
rect 3283 899 3298 1073
rect 3317 899 3332 1073
rect 2948 865 3108 899
rect 3211 888 3263 899
rect 3222 876 3252 888
rect 3211 874 3263 876
rect 3336 874 3351 1073
rect 3110 865 3351 874
rect 3370 906 3404 1107
rect 3418 1054 3452 1141
rect 3482 1131 3486 1141
rect 3538 1139 3562 1141
rect 3576 1139 3600 1141
rect 3533 1106 3626 1139
rect 3640 1106 3668 1141
rect 3533 1098 3578 1106
rect 3533 1097 3560 1098
rect 3591 1097 3640 1098
rect 3575 1088 3641 1097
rect 3700 1088 3720 1141
rect 3480 1076 3518 1088
rect 3572 1081 3640 1088
rect 3572 1076 3602 1081
rect 3472 1064 3518 1076
rect 3472 1054 3486 1064
rect 3560 1061 3618 1076
rect 3572 1054 3618 1061
rect 3625 1054 3640 1081
rect 3686 1054 3720 1088
rect 3734 1054 3773 1141
rect 3418 1043 3681 1054
rect 3418 1031 3670 1043
rect 3418 1020 3618 1031
rect 3629 1020 3681 1031
rect 3686 1020 3706 1054
rect 3739 1048 3773 1054
rect 3720 1020 3773 1048
rect 3472 1011 3558 1020
rect 3705 1014 3720 1020
rect 3739 1014 3773 1020
rect 3470 986 3558 1011
rect 3720 986 3773 1014
rect 3486 961 3530 986
rect 3536 948 3546 979
rect 3528 944 3558 948
rect 3512 914 3578 944
rect 3482 906 3516 910
rect 3370 865 3405 906
rect 3482 894 3528 906
rect 3582 894 3593 906
rect 3594 894 3612 910
rect 3482 880 3612 894
rect 3686 906 3720 960
rect 2734 839 2766 861
rect 2822 846 2851 861
rect 2822 839 2836 846
rect 2874 839 2880 861
rect 2734 792 2880 839
rect 2948 829 3018 865
rect 3370 846 3404 865
rect 3686 846 3728 906
rect 3370 831 3528 846
rect 2734 790 2792 792
rect 2720 756 2792 790
rect 2802 756 2880 792
rect 2886 756 2902 790
rect 2734 729 2780 756
rect 2786 740 2792 756
rect 2822 740 2852 756
rect 2532 728 2780 729
rect 2874 729 2880 756
rect 2914 740 2920 806
rect 2948 757 2982 829
rect 3018 757 3086 829
rect 3382 812 3528 831
rect 3582 812 3728 846
rect 3705 759 3728 812
rect 3739 793 3773 986
rect 3787 1014 3821 1141
rect 3840 1111 3870 1141
rect 4021 1137 4023 1163
rect 4030 1141 4035 1163
rect 4055 1141 4559 1163
rect 3895 1111 3916 1137
rect 3881 1103 3916 1111
rect 4055 1103 4057 1141
rect 3881 1095 3969 1103
rect 3881 1061 3931 1095
rect 3945 1069 3969 1095
rect 3881 1045 3916 1061
rect 3849 1023 3887 1035
rect 3899 1023 3916 1045
rect 4069 1035 4559 1141
rect 3841 1014 3893 1023
rect 3787 1001 3893 1014
rect 3907 1010 3916 1023
rect 3904 1001 3921 1010
rect 3941 1001 3975 1035
rect 3787 967 3987 1001
rect 4055 967 4559 1035
rect 3793 964 3893 967
rect 3819 948 3893 964
rect 3904 964 3975 967
rect 3904 952 3921 964
rect 3841 933 3893 948
rect 3907 933 3916 952
rect 3840 929 3878 933
rect 3840 911 3870 929
rect 3899 911 3916 933
rect 3941 945 3975 964
rect 3941 929 3950 945
rect 3881 901 3916 911
rect 3881 895 3943 901
rect 4072 895 4559 967
rect 4579 1016 4631 1196
rect 4633 1044 4673 1209
rect 4639 1040 4673 1044
rect 4679 1196 4713 1200
rect 4679 1044 4719 1196
rect 4721 1056 4751 1212
rect 4721 1044 4747 1056
rect 4679 1031 4725 1044
rect 4727 1040 4747 1044
rect 4759 1040 4761 1228
rect 4768 1044 4773 1224
rect 4793 1044 4827 1278
rect 4579 1006 4625 1016
rect 4579 895 4613 1006
rect 4649 997 4725 1031
rect 4793 1006 4795 1044
rect 4667 963 4747 997
rect 4667 947 4725 963
rect 4710 932 4725 947
rect 4807 929 4827 1044
rect 4679 895 4713 929
rect 4793 895 4827 929
rect 4841 1349 4875 1373
rect 5174 1390 5244 1666
rect 5356 1598 5414 1604
rect 5356 1564 5368 1598
rect 5356 1558 5414 1564
rect 5356 1398 5414 1404
rect 4894 1349 4929 1354
rect 4990 1349 5148 1354
rect 4841 1292 4881 1349
rect 4937 1320 5148 1349
rect 4937 1315 5100 1320
rect 4942 1292 5100 1315
rect 4841 895 4880 1292
rect 3881 861 3912 895
rect 4072 878 4565 895
rect 3881 855 3943 861
rect 3881 845 3912 855
rect 3794 816 3807 820
rect 3782 793 3827 816
rect 3739 759 3928 793
rect 4072 759 4142 878
rect 4254 842 4312 848
rect 4254 808 4266 842
rect 4254 802 4312 808
rect 2948 739 3108 757
rect 2948 729 3020 739
rect 2874 728 3020 729
rect 3050 728 3108 739
rect 3164 730 3310 757
rect 3382 738 3394 757
rect 2465 672 2499 706
rect 2545 698 2578 728
rect 2579 698 2613 728
rect 2632 698 2666 728
rect 2764 718 2780 728
rect 2511 672 2734 698
rect 2746 672 2780 706
rect 2834 672 2868 706
rect 2948 703 3018 728
rect 3382 726 3405 738
rect 3705 725 3716 759
rect 3882 722 3916 759
rect 4072 723 4125 759
rect 4443 706 4458 878
rect 4477 779 4511 878
rect 4525 861 4565 878
rect 4579 861 4725 895
rect 4793 861 4813 895
rect 4635 795 4669 813
rect 4623 789 4681 795
rect 4623 779 4635 789
rect 4477 745 4512 779
rect 4608 768 4696 779
rect 4619 756 4685 768
rect 4608 745 4696 756
rect 2948 702 2962 703
rect 2965 702 3061 703
rect 2948 698 3036 702
rect 2880 672 3036 698
rect 3050 692 3061 702
rect 3097 693 3263 703
rect 3097 672 3255 693
rect 2352 639 2511 672
rect 2579 639 2613 672
rect 2632 639 2666 672
rect 2712 639 2880 672
rect 2948 639 3268 672
rect 3316 669 3351 703
rect 4477 687 4511 745
rect 2352 638 3268 639
rect 3283 638 3284 669
rect 3317 638 3351 669
rect 3439 651 3899 672
rect 4477 653 4512 687
rect 4608 676 4696 687
rect 4619 664 4685 676
rect 4608 653 4696 664
rect -520 622 -458 628
rect -472 614 -458 622
rect -350 614 2303 629
rect -666 568 -580 614
rect -472 568 -414 614
rect -384 576 2303 614
rect 2365 576 2423 594
rect 2453 576 2511 594
rect 2598 576 2613 638
rect 2632 576 2666 638
rect -384 568 2672 576
rect -666 537 -638 568
rect -350 560 2672 568
rect -632 543 -580 560
rect -555 549 -499 560
rect -472 554 -350 560
rect -472 550 -346 554
rect -333 550 2672 560
rect -544 537 -510 549
rect -472 543 2672 550
rect -666 526 -627 537
rect -555 526 -499 537
rect -468 532 2672 543
rect -468 526 -280 532
rect -333 516 -280 526
rect -736 482 -732 516
rect -434 492 -280 516
rect -201 496 -83 507
rect -333 490 -280 492
rect -297 484 -296 490
rect -190 484 -94 496
rect 0 494 2672 532
rect -297 478 -285 484
rect -201 478 -83 484
rect -297 473 -82 478
rect -626 410 -624 444
rect -331 439 -82 444
rect 0 437 1213 494
rect 1281 444 1285 494
rect 1312 459 1339 494
rect 1388 466 1427 494
rect 1297 444 1339 459
rect 1293 440 1327 442
rect 1381 440 1415 442
rect 1489 441 2672 494
rect 36 386 1213 437
rect 1259 406 1449 408
rect -852 340 -848 374
rect -294 346 -292 374
rect -326 340 -292 346
rect 216 342 226 376
rect 240 342 260 376
rect 441 374 527 386
rect 598 378 628 386
rect 712 378 746 386
rect 587 374 639 378
rect 701 374 757 378
rect 776 374 791 386
rect 441 367 791 374
rect 810 382 844 386
rect 852 384 872 386
rect 850 382 872 384
rect 918 382 1052 386
rect 1126 382 1213 386
rect 810 374 1213 382
rect 810 348 844 374
rect 860 364 872 374
rect 860 358 862 364
rect 1126 348 1213 374
rect 1325 397 1383 403
rect 1325 363 1337 397
rect 1325 357 1383 363
rect 810 340 1213 348
rect 1388 347 1418 386
rect 1502 378 1529 441
rect 1495 340 1529 378
rect 1548 378 1563 441
rect 1650 402 1665 441
rect 1648 391 1665 402
rect 1738 406 1766 441
rect 1738 391 1781 406
rect 430 337 871 340
rect 907 337 959 340
rect 1111 337 1213 340
rect 430 333 860 337
rect 446 306 456 333
rect 470 306 490 333
rect 810 325 860 333
rect 918 325 948 337
rect 810 314 871 325
rect 907 314 959 325
rect 1120 319 1213 337
rect 999 314 1213 319
rect 1120 306 1132 314
rect 1142 310 1204 314
rect 1142 306 1213 310
rect 1486 306 1495 329
rect 1502 306 1546 340
rect 1548 306 1574 378
rect 1648 360 1650 391
rect 1864 386 2672 441
rect 2778 454 2836 460
rect 2778 420 2790 454
rect 2778 414 2836 420
rect 1656 374 1790 378
rect 1690 344 1692 360
rect 1690 340 1756 344
rect 1143 295 1213 306
rect 1064 282 1080 288
rect 1143 284 1308 295
rect 1377 284 1429 295
rect 1452 284 1495 295
rect 1502 284 1529 306
rect 1046 272 1090 282
rect 1046 262 1096 272
rect 1070 256 1096 262
rect 1070 254 1090 256
rect 1046 238 1090 254
rect -582 192 -580 230
rect 1064 228 1090 238
rect 1064 222 1080 228
rect 1143 225 1544 284
rect -544 156 -542 192
rect 178 188 182 216
rect 216 164 226 188
rect 240 164 260 188
rect 216 154 260 164
rect 276 154 288 216
rect 408 188 422 216
rect 674 188 686 216
rect 446 164 460 188
rect 470 164 490 188
rect 446 154 490 164
rect 712 164 724 188
rect 736 164 756 188
rect 712 154 756 164
rect 772 154 784 216
rect 1198 188 1210 216
rect 1464 188 1476 216
rect 1512 204 1544 225
rect 1548 238 1563 306
rect 1690 294 1692 340
rect 1864 242 1951 386
rect 1997 305 2002 386
rect 2025 333 2030 386
rect 2107 359 2114 386
rect 2118 359 2156 378
rect 2170 374 2220 386
rect 2100 345 2156 359
rect 2084 333 2156 345
rect 2157 333 2165 374
rect 2202 364 2214 374
rect 2202 358 2204 364
rect 2227 335 2672 386
rect 2025 329 2071 333
rect 2084 329 2165 333
rect 2084 325 2087 329
rect 2108 325 2128 329
rect 2025 306 2134 325
rect 1997 301 2187 305
rect 2059 272 2125 291
rect 2252 270 2267 335
rect 1609 238 1661 242
rect 1721 238 1777 242
rect 1841 238 1951 242
rect 1548 208 1951 238
rect 1562 204 1574 208
rect 1694 204 1776 208
rect 1794 204 1804 208
rect 1512 188 1608 204
rect 1236 164 1248 188
rect 1260 164 1280 188
rect 1236 154 1280 164
rect 1502 174 1608 188
rect 1662 174 1840 204
rect 1881 189 1951 208
rect 1968 189 1985 204
rect 2026 189 2040 216
rect 2233 189 2267 270
rect 1881 188 2267 189
rect 1502 172 1546 174
rect 1502 164 1514 172
rect 1526 164 1546 172
rect 1502 154 1546 164
rect 1562 154 1574 174
rect 1708 172 1776 174
rect 1732 164 1746 172
rect 1756 164 1776 172
rect 1732 154 1776 164
rect 1794 154 1804 174
rect 1881 172 1940 188
rect 1957 178 2267 188
rect 1917 155 1940 172
rect 1968 155 2267 178
rect 2286 155 2320 335
rect 2596 282 2672 335
rect 2965 318 3035 638
rect 3317 607 3318 638
rect 3159 600 3193 601
rect 3147 401 3205 407
rect 3147 367 3159 401
rect 3147 361 3205 367
rect 2965 282 3018 318
rect 3336 265 3351 638
rect 3370 616 3405 650
rect 3439 638 3923 651
rect 3466 616 3624 638
rect 3685 616 3720 638
rect 4108 633 4143 651
rect 3370 265 3404 616
rect 3686 597 3720 616
rect 4072 618 4143 633
rect 2432 238 2490 244
rect 2432 204 2444 238
rect 3370 231 3385 265
rect 3705 212 3720 597
rect 3739 563 3774 597
rect 3739 212 3773 563
rect 3885 495 3943 501
rect 3885 461 3897 495
rect 3885 455 3943 461
rect 3885 295 3943 301
rect 3885 261 3897 295
rect 3885 255 3943 261
rect 2432 198 2490 204
rect 3739 178 3754 212
rect 4072 159 4142 618
rect 4254 550 4312 556
rect 4254 516 4266 550
rect 4254 510 4312 516
rect 4254 242 4312 248
rect 4254 208 4266 242
rect 4254 202 4312 208
rect 1968 154 2012 155
rect 2026 154 2040 155
rect 234 144 260 154
rect 464 144 490 154
rect 730 144 756 154
rect 1254 144 1280 154
rect 1520 144 1546 154
rect 1750 144 1776 154
rect 1986 144 2012 154
rect 234 138 250 144
rect 464 138 480 144
rect 730 138 746 144
rect 1254 138 1270 144
rect 1520 138 1536 144
rect 1750 138 1766 144
rect 1986 138 2002 144
rect 2286 126 2314 155
rect -1696 102 -1632 126
rect 2286 121 2301 126
rect 4072 123 4125 159
rect 4443 106 4458 652
rect 4477 106 4511 653
rect 4623 643 4635 653
rect 4623 637 4681 643
rect 4623 189 4681 195
rect 4623 155 4635 189
rect 4623 149 4681 155
rect -1668 74 -1632 98
rect 4477 72 4492 106
rect 4812 53 4827 861
rect 4846 726 4880 895
rect 4894 842 4928 1292
rect 5020 1240 5036 1252
rect 5020 1230 5040 1240
rect 5020 1224 5036 1230
rect 5004 1209 5006 1218
rect 5014 1209 5038 1224
rect 5052 1218 5076 1252
rect 5174 1226 5280 1390
rect 5356 1364 5368 1398
rect 5356 1358 5414 1364
rect 5176 1225 5196 1226
rect 4988 1190 5054 1209
rect 4992 1184 5050 1190
rect 5008 1171 5042 1175
rect 5054 1171 5078 1174
rect 5096 1171 5116 1175
rect 4996 1159 5054 1171
rect 5090 1159 5116 1171
rect 4996 1156 5051 1159
rect 4960 1143 4962 1147
rect 4974 1143 4994 1147
rect 4948 963 5000 1143
rect 5002 991 5042 1156
rect 5008 987 5042 991
rect 5048 1143 5082 1147
rect 5048 991 5088 1143
rect 5090 1003 5120 1159
rect 5090 991 5116 1003
rect 5048 978 5094 991
rect 5096 987 5116 991
rect 5128 987 5130 1175
rect 5137 991 5142 1171
rect 5162 1021 5196 1225
rect 5210 1193 5280 1226
rect 5210 1159 5298 1193
rect 5578 1159 5613 1193
rect 5210 1021 5297 1159
rect 5579 1140 5613 1159
rect 5409 1091 5467 1097
rect 5409 1057 5421 1091
rect 5409 1051 5467 1057
rect 5598 1039 5613 1140
rect 5162 991 5297 1021
rect 4948 953 4994 963
rect 4948 842 4982 953
rect 5018 944 5094 978
rect 5162 953 5164 991
rect 5176 985 5297 991
rect 5377 985 5411 1023
rect 5176 951 5280 985
rect 5311 951 5331 985
rect 5365 951 5511 985
rect 5545 951 5565 985
rect 5036 910 5116 944
rect 5036 894 5094 910
rect 5079 879 5094 894
rect 5176 876 5297 951
rect 5377 925 5411 951
rect 5497 925 5499 951
rect 5506 929 5511 951
rect 5531 929 5565 951
rect 5531 891 5533 929
rect 5389 883 5405 891
rect 5048 842 5082 876
rect 4894 808 4934 842
rect 4948 808 5094 842
rect 5162 808 5297 876
rect 5383 849 5407 883
rect 5421 857 5445 891
rect 5545 823 5565 929
rect 5325 811 5363 823
rect 5179 789 5297 808
rect 5317 799 5363 811
rect 5317 789 5351 799
rect 5417 789 5451 823
rect 5531 789 5565 823
rect 5579 932 5613 1039
rect 5632 1106 5667 1140
rect 5632 932 5666 1106
rect 5778 1038 5836 1044
rect 5778 1004 5790 1038
rect 5778 998 5836 1004
rect 5746 932 5780 970
rect 5917 932 6018 1023
rect 5579 898 5619 932
rect 5632 898 5647 932
rect 5680 898 5700 932
rect 5734 898 5880 932
rect 5914 898 6018 932
rect 5579 789 5618 898
rect 5179 772 5303 789
rect 5004 742 5038 760
rect 4992 736 5050 742
rect 4992 726 5004 736
rect 4846 692 4881 726
rect 4977 715 5065 726
rect 4988 703 5054 715
rect 4977 692 5065 703
rect 4846 634 4880 692
rect 4846 600 4881 634
rect 4977 623 5065 634
rect 4988 611 5054 623
rect 4977 600 5065 611
rect 4846 53 4880 600
rect 4992 590 5004 600
rect 4992 584 5050 590
rect 5179 581 5249 772
rect 5263 755 5303 772
rect 5317 755 5463 789
rect 5531 755 5551 789
rect 5361 683 5419 689
rect 5361 649 5373 683
rect 5361 643 5419 649
rect 5179 547 5250 581
rect 5550 547 5565 755
rect 5584 547 5618 789
rect 5632 736 5666 898
rect 5746 872 5780 898
rect 5866 872 5868 898
rect 5875 876 5880 898
rect 5900 876 6018 898
rect 5900 838 5902 876
rect 5758 830 5774 838
rect 5752 796 5776 830
rect 5790 804 5814 838
rect 5914 770 6018 876
rect 6099 885 6157 891
rect 6099 851 6111 885
rect 6269 862 6303 880
rect 6099 845 6157 851
rect 6269 826 6339 862
rect 5694 758 5732 770
rect 5686 746 5732 758
rect 5686 736 5720 746
rect 5786 736 5820 770
rect 5632 702 5672 736
rect 5686 702 5832 736
rect 5900 702 6018 770
rect 5917 666 6018 702
rect 6286 792 6357 826
rect 6637 792 6672 826
rect 7060 809 7095 827
rect 5730 630 5788 636
rect 5730 596 5742 630
rect 5730 590 5788 596
rect 5179 511 5232 547
rect 5584 513 5599 547
rect 5917 494 5987 666
rect 6099 577 6157 583
rect 6099 543 6111 577
rect 6099 537 6157 543
rect 5917 458 5970 494
rect 5162 421 5196 439
rect 6286 422 6356 792
rect 6638 773 6672 792
rect 7024 794 7095 809
rect 7375 794 7410 828
rect 6468 724 6526 730
rect 6468 690 6480 724
rect 6468 684 6526 690
rect 6468 524 6526 530
rect 6468 490 6480 524
rect 6468 484 6526 490
rect 5162 385 5232 421
rect 6286 388 6357 422
rect 6657 388 6672 773
rect 6691 739 6726 773
rect 6691 388 6725 739
rect 6837 671 6895 677
rect 6837 637 6849 671
rect 6837 631 6895 637
rect 6837 471 6895 477
rect 6837 437 6849 471
rect 6837 431 6895 437
rect 5179 351 5250 385
rect 5530 351 5565 385
rect 5953 368 5988 386
rect 4992 136 5050 142
rect 4992 102 5004 136
rect 4992 96 5050 102
rect 4846 19 4861 53
rect 5179 0 5249 351
rect 5531 332 5565 351
rect 5917 353 5988 368
rect 5361 283 5419 289
rect 5361 249 5373 283
rect 5361 243 5419 249
rect 5361 83 5419 89
rect 5361 49 5373 83
rect 5361 43 5419 49
rect 5179 -36 5232 0
rect 5550 -53 5565 332
rect 5584 298 5619 332
rect 5584 -53 5618 298
rect 5730 230 5788 236
rect 5730 196 5742 230
rect 5730 190 5788 196
rect 5730 30 5788 36
rect 5730 -4 5742 30
rect 5730 -10 5788 -4
rect 5584 -87 5599 -53
rect 5917 -106 5987 353
rect 6286 352 6339 388
rect 6691 354 6706 388
rect 7024 335 7094 794
rect 7376 775 7410 794
rect 7206 726 7264 732
rect 7206 692 7218 726
rect 7206 686 7264 692
rect 7206 418 7264 424
rect 7206 384 7218 418
rect 7206 378 7264 384
rect 7024 299 7077 335
rect 6099 285 6157 291
rect 6099 251 6111 285
rect 7395 282 7410 775
rect 7429 741 7464 775
rect 6269 262 6303 280
rect 7429 263 7463 741
rect 7575 673 7633 679
rect 7575 639 7587 673
rect 7745 650 7779 668
rect 7575 633 7633 639
rect 7745 614 7815 650
rect 7762 580 7833 614
rect 7575 365 7633 371
rect 7575 331 7587 365
rect 7575 325 7633 331
rect 6099 245 6157 251
rect 6269 226 6339 262
rect 7429 229 7464 263
rect 6286 192 6357 226
rect 6637 192 6672 226
rect 7060 209 7095 227
rect 6099 -23 6157 -17
rect 6099 -57 6111 -23
rect 6099 -63 6157 -57
rect 5917 -142 5970 -106
rect 6286 -159 6356 192
rect 6638 173 6672 192
rect 7024 194 7095 209
rect 7375 194 7410 228
rect 6468 124 6526 130
rect 6468 90 6480 124
rect 6468 84 6526 90
rect 6468 -76 6526 -70
rect 6468 -110 6480 -76
rect 6468 -116 6526 -110
rect 6286 -195 6339 -159
rect 6657 -212 6672 173
rect 6691 139 6726 173
rect 6691 -212 6725 139
rect 6837 71 6895 77
rect 6837 37 6849 71
rect 6837 31 6895 37
rect 6837 -129 6895 -123
rect 6837 -163 6849 -129
rect 6837 -169 6895 -163
rect 6691 -246 6706 -212
rect 7024 -265 7094 194
rect 7376 175 7410 194
rect 7762 210 7832 580
rect 7944 512 8002 518
rect 7944 478 7956 512
rect 7944 472 8002 478
rect 7944 312 8002 318
rect 7944 278 7956 312
rect 7944 272 8002 278
rect 7762 176 7833 210
rect 7206 126 7264 132
rect 7206 92 7218 126
rect 7206 86 7264 92
rect 7206 -182 7264 -176
rect 7206 -216 7218 -182
rect 7206 -222 7264 -216
rect 7024 -301 7077 -265
rect 7395 -318 7410 175
rect 7429 141 7464 175
rect 7429 -318 7463 141
rect 7762 140 7815 176
rect 7575 73 7633 79
rect 7575 39 7587 73
rect 7745 50 7779 68
rect 7575 33 7633 39
rect 7745 14 7815 50
rect 7762 -20 7833 14
rect 7575 -235 7633 -229
rect 7575 -269 7587 -235
rect 7575 -275 7633 -269
rect 7429 -352 7444 -318
rect 7762 -371 7832 -20
rect 7944 -88 8002 -82
rect 7944 -122 7956 -88
rect 7944 -128 8002 -122
rect 7944 -288 8002 -282
rect 7944 -322 7956 -288
rect 7944 -328 8002 -322
rect 7762 -407 7815 -371
<< metal1 >>
rect -1668 877 2296 910
rect -29 574 2003 607
rect -429 573 12 574
rect -1529 541 12 573
rect -1529 381 -1494 541
rect -434 517 -368 541
rect 1967 540 2003 574
rect -434 513 -383 517
rect -1282 493 -1212 499
rect -1282 481 -1276 493
rect -1409 447 -1276 481
rect -1282 435 -1276 447
rect -1218 481 -1212 493
rect -418 488 -383 513
rect 120 512 190 518
rect -1218 447 -518 481
rect 120 454 126 512
rect 184 454 190 512
rect 120 448 190 454
rect -1218 435 -1212 447
rect -1282 429 -1212 435
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect -552 373 -518 447
rect -552 339 -296 373
rect -49 342 223 373
rect 810 367 880 373
rect -49 266 -18 342
rect 810 309 816 367
rect 874 309 880 367
rect 810 303 880 309
rect 1967 305 2002 540
rect 2226 318 2296 324
rect 2226 305 2232 318
rect -542 235 -18 266
rect 1967 271 2232 305
rect -542 184 -511 235
rect 0 33 200 200
rect 1967 185 2002 271
rect 2226 260 2232 271
rect 2290 260 2296 318
rect 2226 254 2296 260
rect -1668 0 2296 33
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
<< via1 >>
rect -1276 435 -1218 493
rect 126 454 184 512
rect -1110 352 -1052 410
rect 816 309 874 367
rect 2232 260 2290 318
<< metal2 >>
rect 120 512 190 910
rect -1282 493 -1212 498
rect -1282 435 -1276 493
rect -1218 435 -1212 493
rect -1282 429 -1212 435
rect 120 454 126 512
rect 184 454 190 512
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect 120 0 190 454
rect 810 367 880 910
rect 810 309 816 367
rect 874 309 880 367
rect 810 0 880 309
rect 2226 318 2296 324
rect 2226 260 2232 318
rect 2290 260 2296 318
rect 2226 254 2296 260
use and_scan  and_scan_0
timestamp 1624053917
transform 1 0 -1632 0 1 344
box -53 -2800 2214 1147
use and_scan  XAND1
timestamp 1624053917
transform 1 0 3382 0 1 944
box -53 -2800 2214 1147
use xor_scan  xor_scan_0
timestamp 1624053917
transform 1 0 -1756 0 1 102
box -53 -2800 4428 1165
use xor_scan  XXOR1
timestamp 1624053917
transform 1 0 1590 0 1 702
box -53 -2800 4428 1165
use dffc_scan  dffc_scan_0
timestamp 1624053917
transform 1 0 66 0 1 106
box -66 -3600 8118 1112
use dffc_scan  xDFFC1
timestamp 1624053917
transform 1 0 66 0 1 706
box -66 -3600 8118 1112
<< labels >>
rlabel metal2 845 910 845 910 1 CLR
rlabel metal2 2296 288 2296 288 3 Dn
rlabel metal2 157 910 157 910 1 CLK
rlabel metal2 -1246 498 -1246 498 1 CE
rlabel metal2 -1081 346 -1081 346 5 Sout
rlabel metal1 260 910 260 910 1 VDD
rlabel metal1 226 0 226 0 5 VSS
rlabel metal1 15 16 15 16 5 VSS
rlabel space 15 852 15 852 5 VDD
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Dn
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 CE
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLR
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLK
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Sout
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 {}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 VDD
port 9 nsew
<< end >>
