magic
tech sky130A
magscale 1 2
timestamp 1616195620
<< nwell >>
rect -354 820 647 821
rect -355 384 647 820
rect -355 381 -354 384
rect -342 381 647 384
<< psubdiff >>
rect -269 -117 -245 -83
rect 555 -117 579 -83
<< nsubdiff >>
rect -273 751 43 785
rect 353 751 576 785
<< psubdiffcont >>
rect -245 -117 555 -83
<< nsubdiffcont >>
rect 43 751 353 785
<< poly >>
rect 43 691 352 721
rect -260 428 -230 649
rect -60 428 -30 649
rect -260 398 -30 428
rect -260 384 -230 398
rect -295 368 -230 384
rect -295 334 -285 368
rect -251 334 -230 368
rect -295 318 -230 334
rect -260 -39 -230 318
rect -66 318 -12 333
rect 43 318 73 691
rect 146 363 176 649
rect 234 375 264 649
rect 322 417 352 691
rect 522 375 552 649
rect -66 317 73 318
rect -66 283 -56 317
rect -22 288 73 317
rect 138 347 192 363
rect 138 313 148 347
rect 182 313 192 347
rect 234 345 552 375
rect 138 297 192 313
rect -22 283 -12 288
rect -66 267 -12 283
rect -54 23 -24 267
rect 146 5 176 297
rect 522 276 552 345
rect 522 260 624 276
rect 234 -39 264 237
rect 322 5 352 237
rect 522 226 580 260
rect 614 226 624 260
rect 522 210 624 226
rect 522 5 552 210
rect 322 -25 552 5
rect -260 -69 264 -39
<< polycont >>
rect -285 334 -251 368
rect -56 283 -22 317
rect 148 313 182 347
rect 580 226 614 260
<< locali >>
rect -295 368 -241 384
rect -295 334 -285 368
rect -251 334 -241 368
rect -295 318 -241 334
rect 138 347 192 363
rect -66 317 -12 333
rect -66 283 -56 317
rect -22 283 -12 317
rect 138 313 148 347
rect 182 313 192 347
rect 138 297 192 313
rect -66 267 -12 283
rect 570 260 624 276
rect 570 226 580 260
rect 614 226 624 260
rect 570 210 624 226
<< viali >>
rect -273 751 43 785
rect 43 751 353 785
rect 353 751 576 785
rect -285 334 -251 368
rect -56 283 -22 317
rect 148 313 182 347
rect 580 226 614 260
rect -270 -117 -245 -83
rect -245 -117 555 -83
rect 555 -117 580 -83
rect -270 -118 580 -117
<< metal1 >>
rect -354 785 647 821
rect -354 751 -273 785
rect 576 751 647 785
rect -354 745 647 751
rect -301 638 -270 745
rect -309 559 -270 638
rect -109 624 -69 745
rect -109 611 -68 624
rect -309 452 -271 559
rect -220 452 -180 611
rect -108 459 -68 611
rect -21 587 19 617
rect 99 587 139 619
rect -21 483 139 587
rect -21 475 24 483
rect 95 475 139 483
rect 187 481 227 621
rect 362 617 402 745
rect -21 452 19 475
rect 99 454 139 475
rect 184 456 227 481
rect 361 608 402 617
rect -223 446 -180 452
rect -223 445 -195 446
rect -223 443 -189 445
rect 184 443 224 456
rect 361 452 401 608
rect 471 485 511 622
rect 567 616 598 745
rect 471 457 512 485
rect -342 368 -241 384
rect -342 334 -285 368
rect -251 334 -241 368
rect -342 318 -241 334
rect -212 316 -184 443
rect 182 433 224 443
rect 472 437 512 457
rect 564 451 604 616
rect 182 415 210 433
rect 56 387 210 415
rect 56 355 84 387
rect -66 317 -12 333
rect -66 316 -56 317
rect -212 287 -56 316
rect -310 46 -274 135
rect -212 133 -184 287
rect -66 283 -56 287
rect -22 283 -12 317
rect 31 303 41 355
rect 93 303 103 355
rect 138 347 192 359
rect 138 313 148 347
rect 182 327 192 347
rect 476 327 507 437
rect 182 313 507 327
rect -66 267 -12 283
rect 56 269 84 303
rect 138 299 507 313
rect 138 297 192 299
rect 56 239 210 269
rect -217 132 -186 133
rect -310 -76 -279 46
rect -222 45 -186 132
rect -107 77 -61 227
rect 182 217 210 239
rect 182 211 231 217
rect -103 -76 -63 77
rect -6 -7 24 157
rect 89 27 137 202
rect 183 42 231 211
rect 101 -7 131 27
rect 270 25 318 200
rect 358 32 406 207
rect 476 154 507 299
rect 570 260 625 276
rect 570 226 580 260
rect 614 226 625 260
rect 570 210 625 226
rect 473 33 513 154
rect 278 -7 308 25
rect -6 -35 308 -7
rect 362 -76 402 32
rect 561 30 601 113
rect 565 -76 596 30
rect -355 -83 647 -76
rect -355 -118 -270 -83
rect 580 -118 647 -83
rect -355 -124 647 -118
<< via1 >>
rect 41 303 93 355
<< metal2 >>
rect 31 355 103 365
rect 31 303 41 355
rect 93 303 103 355
rect 31 293 103 303
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615298455
transform 1 0 -245 0 1 88
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_0
timestamp 1614978561
transform 1 0 -39 0 1 139
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_1
timestamp 1614978561
transform 1 0 161 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_2
timestamp 1614978561
transform 1 0 249 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_3
timestamp 1614978561
transform 1 0 337 0 1 121
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_1
timestamp 1615298455
transform 1 0 537 0 1 76
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_0
timestamp 1614978561
transform 1 0 -45 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_4
timestamp 1614978561
transform 1 0 -245 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_1
timestamp 1614978561
transform 1 0 161 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_2
timestamp 1614978561
transform 1 0 249 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_3
timestamp 1614978561
transform 1 0 337 0 1 533
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_5
timestamp 1614978561
transform 1 0 537 0 1 533
box -109 -152 109 152
<< labels >>
rlabel metal1 -354 -124 646 -76 1 vss
rlabel nwell -354 745 646 821 1 vdd
rlabel metal2 31 293 103 365 1 out
rlabel metal1 570 210 625 276 1 in1
rlabel metal1 -342 318 -241 384 1 in2
<< end >>
