magic
tech sky130A
magscale 1 2
timestamp 1616600406
<< error_p >>
rect -2920 345 -2862 351
rect -2802 345 -2744 351
rect -2684 345 -2626 351
rect -2566 345 -2508 351
rect -2448 345 -2390 351
rect -2330 345 -2272 351
rect -2212 345 -2154 351
rect -2094 345 -2036 351
rect -1976 345 -1918 351
rect -1858 345 -1800 351
rect -1740 345 -1682 351
rect -1622 345 -1564 351
rect -1504 345 -1446 351
rect -1386 345 -1328 351
rect -1268 345 -1210 351
rect -1150 345 -1092 351
rect -1032 345 -974 351
rect -914 345 -856 351
rect -796 345 -738 351
rect -678 345 -620 351
rect -560 345 -502 351
rect -442 345 -384 351
rect -324 345 -266 351
rect -206 345 -148 351
rect -88 345 -30 351
rect 30 345 88 351
rect 148 345 206 351
rect 266 345 324 351
rect 384 345 442 351
rect 502 345 560 351
rect 620 345 678 351
rect 738 345 796 351
rect 856 345 914 351
rect 974 345 1032 351
rect 1092 345 1150 351
rect 1210 345 1268 351
rect 1328 345 1386 351
rect 1446 345 1504 351
rect 1564 345 1622 351
rect 1682 345 1740 351
rect 1800 345 1858 351
rect 1918 345 1976 351
rect 2036 345 2094 351
rect 2154 345 2212 351
rect 2272 345 2330 351
rect 2390 345 2448 351
rect 2508 345 2566 351
rect 2626 345 2684 351
rect 2744 345 2802 351
rect 2862 345 2920 351
rect -2920 311 -2908 345
rect -2802 311 -2790 345
rect -2684 311 -2672 345
rect -2566 311 -2554 345
rect -2448 311 -2436 345
rect -2330 311 -2318 345
rect -2212 311 -2200 345
rect -2094 311 -2082 345
rect -1976 311 -1964 345
rect -1858 311 -1846 345
rect -1740 311 -1728 345
rect -1622 311 -1610 345
rect -1504 311 -1492 345
rect -1386 311 -1374 345
rect -1268 311 -1256 345
rect -1150 311 -1138 345
rect -1032 311 -1020 345
rect -914 311 -902 345
rect -796 311 -784 345
rect -678 311 -666 345
rect -560 311 -548 345
rect -442 311 -430 345
rect -324 311 -312 345
rect -206 311 -194 345
rect -88 311 -76 345
rect 30 311 42 345
rect 148 311 160 345
rect 266 311 278 345
rect 384 311 396 345
rect 502 311 514 345
rect 620 311 632 345
rect 738 311 750 345
rect 856 311 868 345
rect 974 311 986 345
rect 1092 311 1104 345
rect 1210 311 1222 345
rect 1328 311 1340 345
rect 1446 311 1458 345
rect 1564 311 1576 345
rect 1682 311 1694 345
rect 1800 311 1812 345
rect 1918 311 1930 345
rect 2036 311 2048 345
rect 2154 311 2166 345
rect 2272 311 2284 345
rect 2390 311 2402 345
rect 2508 311 2520 345
rect 2626 311 2638 345
rect 2744 311 2756 345
rect 2862 311 2874 345
rect -2920 305 -2862 311
rect -2802 305 -2744 311
rect -2684 305 -2626 311
rect -2566 305 -2508 311
rect -2448 305 -2390 311
rect -2330 305 -2272 311
rect -2212 305 -2154 311
rect -2094 305 -2036 311
rect -1976 305 -1918 311
rect -1858 305 -1800 311
rect -1740 305 -1682 311
rect -1622 305 -1564 311
rect -1504 305 -1446 311
rect -1386 305 -1328 311
rect -1268 305 -1210 311
rect -1150 305 -1092 311
rect -1032 305 -974 311
rect -914 305 -856 311
rect -796 305 -738 311
rect -678 305 -620 311
rect -560 305 -502 311
rect -442 305 -384 311
rect -324 305 -266 311
rect -206 305 -148 311
rect -88 305 -30 311
rect 30 305 88 311
rect 148 305 206 311
rect 266 305 324 311
rect 384 305 442 311
rect 502 305 560 311
rect 620 305 678 311
rect 738 305 796 311
rect 856 305 914 311
rect 974 305 1032 311
rect 1092 305 1150 311
rect 1210 305 1268 311
rect 1328 305 1386 311
rect 1446 305 1504 311
rect 1564 305 1622 311
rect 1682 305 1740 311
rect 1800 305 1858 311
rect 1918 305 1976 311
rect 2036 305 2094 311
rect 2154 305 2212 311
rect 2272 305 2330 311
rect 2390 305 2448 311
rect 2508 305 2566 311
rect 2626 305 2684 311
rect 2744 305 2802 311
rect 2862 305 2920 311
<< nwell >>
rect -3117 -484 3117 484
<< pmos >>
rect -2921 -336 -2861 264
rect -2803 -336 -2743 264
rect -2685 -336 -2625 264
rect -2567 -336 -2507 264
rect -2449 -336 -2389 264
rect -2331 -336 -2271 264
rect -2213 -336 -2153 264
rect -2095 -336 -2035 264
rect -1977 -336 -1917 264
rect -1859 -336 -1799 264
rect -1741 -336 -1681 264
rect -1623 -336 -1563 264
rect -1505 -336 -1445 264
rect -1387 -336 -1327 264
rect -1269 -336 -1209 264
rect -1151 -336 -1091 264
rect -1033 -336 -973 264
rect -915 -336 -855 264
rect -797 -336 -737 264
rect -679 -336 -619 264
rect -561 -336 -501 264
rect -443 -336 -383 264
rect -325 -336 -265 264
rect -207 -336 -147 264
rect -89 -336 -29 264
rect 29 -336 89 264
rect 147 -336 207 264
rect 265 -336 325 264
rect 383 -336 443 264
rect 501 -336 561 264
rect 619 -336 679 264
rect 737 -336 797 264
rect 855 -336 915 264
rect 973 -336 1033 264
rect 1091 -336 1151 264
rect 1209 -336 1269 264
rect 1327 -336 1387 264
rect 1445 -336 1505 264
rect 1563 -336 1623 264
rect 1681 -336 1741 264
rect 1799 -336 1859 264
rect 1917 -336 1977 264
rect 2035 -336 2095 264
rect 2153 -336 2213 264
rect 2271 -336 2331 264
rect 2389 -336 2449 264
rect 2507 -336 2567 264
rect 2625 -336 2685 264
rect 2743 -336 2803 264
rect 2861 -336 2921 264
<< pdiff >>
rect -2979 252 -2921 264
rect -2979 -324 -2967 252
rect -2933 -324 -2921 252
rect -2979 -336 -2921 -324
rect -2861 252 -2803 264
rect -2861 -324 -2849 252
rect -2815 -324 -2803 252
rect -2861 -336 -2803 -324
rect -2743 252 -2685 264
rect -2743 -324 -2731 252
rect -2697 -324 -2685 252
rect -2743 -336 -2685 -324
rect -2625 252 -2567 264
rect -2625 -324 -2613 252
rect -2579 -324 -2567 252
rect -2625 -336 -2567 -324
rect -2507 252 -2449 264
rect -2507 -324 -2495 252
rect -2461 -324 -2449 252
rect -2507 -336 -2449 -324
rect -2389 252 -2331 264
rect -2389 -324 -2377 252
rect -2343 -324 -2331 252
rect -2389 -336 -2331 -324
rect -2271 252 -2213 264
rect -2271 -324 -2259 252
rect -2225 -324 -2213 252
rect -2271 -336 -2213 -324
rect -2153 252 -2095 264
rect -2153 -324 -2141 252
rect -2107 -324 -2095 252
rect -2153 -336 -2095 -324
rect -2035 252 -1977 264
rect -2035 -324 -2023 252
rect -1989 -324 -1977 252
rect -2035 -336 -1977 -324
rect -1917 252 -1859 264
rect -1917 -324 -1905 252
rect -1871 -324 -1859 252
rect -1917 -336 -1859 -324
rect -1799 252 -1741 264
rect -1799 -324 -1787 252
rect -1753 -324 -1741 252
rect -1799 -336 -1741 -324
rect -1681 252 -1623 264
rect -1681 -324 -1669 252
rect -1635 -324 -1623 252
rect -1681 -336 -1623 -324
rect -1563 252 -1505 264
rect -1563 -324 -1551 252
rect -1517 -324 -1505 252
rect -1563 -336 -1505 -324
rect -1445 252 -1387 264
rect -1445 -324 -1433 252
rect -1399 -324 -1387 252
rect -1445 -336 -1387 -324
rect -1327 252 -1269 264
rect -1327 -324 -1315 252
rect -1281 -324 -1269 252
rect -1327 -336 -1269 -324
rect -1209 252 -1151 264
rect -1209 -324 -1197 252
rect -1163 -324 -1151 252
rect -1209 -336 -1151 -324
rect -1091 252 -1033 264
rect -1091 -324 -1079 252
rect -1045 -324 -1033 252
rect -1091 -336 -1033 -324
rect -973 252 -915 264
rect -973 -324 -961 252
rect -927 -324 -915 252
rect -973 -336 -915 -324
rect -855 252 -797 264
rect -855 -324 -843 252
rect -809 -324 -797 252
rect -855 -336 -797 -324
rect -737 252 -679 264
rect -737 -324 -725 252
rect -691 -324 -679 252
rect -737 -336 -679 -324
rect -619 252 -561 264
rect -619 -324 -607 252
rect -573 -324 -561 252
rect -619 -336 -561 -324
rect -501 252 -443 264
rect -501 -324 -489 252
rect -455 -324 -443 252
rect -501 -336 -443 -324
rect -383 252 -325 264
rect -383 -324 -371 252
rect -337 -324 -325 252
rect -383 -336 -325 -324
rect -265 252 -207 264
rect -265 -324 -253 252
rect -219 -324 -207 252
rect -265 -336 -207 -324
rect -147 252 -89 264
rect -147 -324 -135 252
rect -101 -324 -89 252
rect -147 -336 -89 -324
rect -29 252 29 264
rect -29 -324 -17 252
rect 17 -324 29 252
rect -29 -336 29 -324
rect 89 252 147 264
rect 89 -324 101 252
rect 135 -324 147 252
rect 89 -336 147 -324
rect 207 252 265 264
rect 207 -324 219 252
rect 253 -324 265 252
rect 207 -336 265 -324
rect 325 252 383 264
rect 325 -324 337 252
rect 371 -324 383 252
rect 325 -336 383 -324
rect 443 252 501 264
rect 443 -324 455 252
rect 489 -324 501 252
rect 443 -336 501 -324
rect 561 252 619 264
rect 561 -324 573 252
rect 607 -324 619 252
rect 561 -336 619 -324
rect 679 252 737 264
rect 679 -324 691 252
rect 725 -324 737 252
rect 679 -336 737 -324
rect 797 252 855 264
rect 797 -324 809 252
rect 843 -324 855 252
rect 797 -336 855 -324
rect 915 252 973 264
rect 915 -324 927 252
rect 961 -324 973 252
rect 915 -336 973 -324
rect 1033 252 1091 264
rect 1033 -324 1045 252
rect 1079 -324 1091 252
rect 1033 -336 1091 -324
rect 1151 252 1209 264
rect 1151 -324 1163 252
rect 1197 -324 1209 252
rect 1151 -336 1209 -324
rect 1269 252 1327 264
rect 1269 -324 1281 252
rect 1315 -324 1327 252
rect 1269 -336 1327 -324
rect 1387 252 1445 264
rect 1387 -324 1399 252
rect 1433 -324 1445 252
rect 1387 -336 1445 -324
rect 1505 252 1563 264
rect 1505 -324 1517 252
rect 1551 -324 1563 252
rect 1505 -336 1563 -324
rect 1623 252 1681 264
rect 1623 -324 1635 252
rect 1669 -324 1681 252
rect 1623 -336 1681 -324
rect 1741 252 1799 264
rect 1741 -324 1753 252
rect 1787 -324 1799 252
rect 1741 -336 1799 -324
rect 1859 252 1917 264
rect 1859 -324 1871 252
rect 1905 -324 1917 252
rect 1859 -336 1917 -324
rect 1977 252 2035 264
rect 1977 -324 1989 252
rect 2023 -324 2035 252
rect 1977 -336 2035 -324
rect 2095 252 2153 264
rect 2095 -324 2107 252
rect 2141 -324 2153 252
rect 2095 -336 2153 -324
rect 2213 252 2271 264
rect 2213 -324 2225 252
rect 2259 -324 2271 252
rect 2213 -336 2271 -324
rect 2331 252 2389 264
rect 2331 -324 2343 252
rect 2377 -324 2389 252
rect 2331 -336 2389 -324
rect 2449 252 2507 264
rect 2449 -324 2461 252
rect 2495 -324 2507 252
rect 2449 -336 2507 -324
rect 2567 252 2625 264
rect 2567 -324 2579 252
rect 2613 -324 2625 252
rect 2567 -336 2625 -324
rect 2685 252 2743 264
rect 2685 -324 2697 252
rect 2731 -324 2743 252
rect 2685 -336 2743 -324
rect 2803 252 2861 264
rect 2803 -324 2815 252
rect 2849 -324 2861 252
rect 2803 -336 2861 -324
rect 2921 252 2979 264
rect 2921 -324 2933 252
rect 2967 -324 2979 252
rect 2921 -336 2979 -324
<< pdiffc >>
rect -2967 -324 -2933 252
rect -2849 -324 -2815 252
rect -2731 -324 -2697 252
rect -2613 -324 -2579 252
rect -2495 -324 -2461 252
rect -2377 -324 -2343 252
rect -2259 -324 -2225 252
rect -2141 -324 -2107 252
rect -2023 -324 -1989 252
rect -1905 -324 -1871 252
rect -1787 -324 -1753 252
rect -1669 -324 -1635 252
rect -1551 -324 -1517 252
rect -1433 -324 -1399 252
rect -1315 -324 -1281 252
rect -1197 -324 -1163 252
rect -1079 -324 -1045 252
rect -961 -324 -927 252
rect -843 -324 -809 252
rect -725 -324 -691 252
rect -607 -324 -573 252
rect -489 -324 -455 252
rect -371 -324 -337 252
rect -253 -324 -219 252
rect -135 -324 -101 252
rect -17 -324 17 252
rect 101 -324 135 252
rect 219 -324 253 252
rect 337 -324 371 252
rect 455 -324 489 252
rect 573 -324 607 252
rect 691 -324 725 252
rect 809 -324 843 252
rect 927 -324 961 252
rect 1045 -324 1079 252
rect 1163 -324 1197 252
rect 1281 -324 1315 252
rect 1399 -324 1433 252
rect 1517 -324 1551 252
rect 1635 -324 1669 252
rect 1753 -324 1787 252
rect 1871 -324 1905 252
rect 1989 -324 2023 252
rect 2107 -324 2141 252
rect 2225 -324 2259 252
rect 2343 -324 2377 252
rect 2461 -324 2495 252
rect 2579 -324 2613 252
rect 2697 -324 2731 252
rect 2815 -324 2849 252
rect 2933 -324 2967 252
<< nsubdiff >>
rect -3081 414 -2985 448
rect 2985 414 3081 448
rect -3081 351 -3047 414
rect 3047 351 3081 414
rect -3081 -414 -3047 -351
rect 3047 -414 3081 -351
rect -3081 -448 -2985 -414
rect 2985 -448 3081 -414
<< nsubdiffcont >>
rect -2985 414 2985 448
rect -3081 -351 -3047 351
rect 3047 -351 3081 351
rect -2985 -448 2985 -414
<< poly >>
rect -2924 345 -2858 361
rect -2924 311 -2908 345
rect -2874 311 -2858 345
rect -2924 295 -2858 311
rect -2806 345 -2740 361
rect -2806 311 -2790 345
rect -2756 311 -2740 345
rect -2806 295 -2740 311
rect -2688 345 -2622 361
rect -2688 311 -2672 345
rect -2638 311 -2622 345
rect -2688 295 -2622 311
rect -2570 345 -2504 361
rect -2570 311 -2554 345
rect -2520 311 -2504 345
rect -2570 295 -2504 311
rect -2452 345 -2386 361
rect -2452 311 -2436 345
rect -2402 311 -2386 345
rect -2452 295 -2386 311
rect -2334 345 -2268 361
rect -2334 311 -2318 345
rect -2284 311 -2268 345
rect -2334 295 -2268 311
rect -2216 345 -2150 361
rect -2216 311 -2200 345
rect -2166 311 -2150 345
rect -2216 295 -2150 311
rect -2098 345 -2032 361
rect -2098 311 -2082 345
rect -2048 311 -2032 345
rect -2098 295 -2032 311
rect -1980 345 -1914 361
rect -1980 311 -1964 345
rect -1930 311 -1914 345
rect -1980 295 -1914 311
rect -1862 345 -1796 361
rect -1862 311 -1846 345
rect -1812 311 -1796 345
rect -1862 295 -1796 311
rect -1744 345 -1678 361
rect -1744 311 -1728 345
rect -1694 311 -1678 345
rect -1744 295 -1678 311
rect -1626 345 -1560 361
rect -1626 311 -1610 345
rect -1576 311 -1560 345
rect -1626 295 -1560 311
rect -1508 345 -1442 361
rect -1508 311 -1492 345
rect -1458 311 -1442 345
rect -1508 295 -1442 311
rect -1390 345 -1324 361
rect -1390 311 -1374 345
rect -1340 311 -1324 345
rect -1390 295 -1324 311
rect -1272 345 -1206 361
rect -1272 311 -1256 345
rect -1222 311 -1206 345
rect -1272 295 -1206 311
rect -1154 345 -1088 361
rect -1154 311 -1138 345
rect -1104 311 -1088 345
rect -1154 295 -1088 311
rect -1036 345 -970 361
rect -1036 311 -1020 345
rect -986 311 -970 345
rect -1036 295 -970 311
rect -918 345 -852 361
rect -918 311 -902 345
rect -868 311 -852 345
rect -918 295 -852 311
rect -800 345 -734 361
rect -800 311 -784 345
rect -750 311 -734 345
rect -800 295 -734 311
rect -682 345 -616 361
rect -682 311 -666 345
rect -632 311 -616 345
rect -682 295 -616 311
rect -564 345 -498 361
rect -564 311 -548 345
rect -514 311 -498 345
rect -564 295 -498 311
rect -446 345 -380 361
rect -446 311 -430 345
rect -396 311 -380 345
rect -446 295 -380 311
rect -328 345 -262 361
rect -328 311 -312 345
rect -278 311 -262 345
rect -328 295 -262 311
rect -210 345 -144 361
rect -210 311 -194 345
rect -160 311 -144 345
rect -210 295 -144 311
rect -92 345 -26 361
rect -92 311 -76 345
rect -42 311 -26 345
rect -92 295 -26 311
rect 26 345 92 361
rect 26 311 42 345
rect 76 311 92 345
rect 26 295 92 311
rect 144 345 210 361
rect 144 311 160 345
rect 194 311 210 345
rect 144 295 210 311
rect 262 345 328 361
rect 262 311 278 345
rect 312 311 328 345
rect 262 295 328 311
rect 380 345 446 361
rect 380 311 396 345
rect 430 311 446 345
rect 380 295 446 311
rect 498 345 564 361
rect 498 311 514 345
rect 548 311 564 345
rect 498 295 564 311
rect 616 345 682 361
rect 616 311 632 345
rect 666 311 682 345
rect 616 295 682 311
rect 734 345 800 361
rect 734 311 750 345
rect 784 311 800 345
rect 734 295 800 311
rect 852 345 918 361
rect 852 311 868 345
rect 902 311 918 345
rect 852 295 918 311
rect 970 345 1036 361
rect 970 311 986 345
rect 1020 311 1036 345
rect 970 295 1036 311
rect 1088 345 1154 361
rect 1088 311 1104 345
rect 1138 311 1154 345
rect 1088 295 1154 311
rect 1206 345 1272 361
rect 1206 311 1222 345
rect 1256 311 1272 345
rect 1206 295 1272 311
rect 1324 345 1390 361
rect 1324 311 1340 345
rect 1374 311 1390 345
rect 1324 295 1390 311
rect 1442 345 1508 361
rect 1442 311 1458 345
rect 1492 311 1508 345
rect 1442 295 1508 311
rect 1560 345 1626 361
rect 1560 311 1576 345
rect 1610 311 1626 345
rect 1560 295 1626 311
rect 1678 345 1744 361
rect 1678 311 1694 345
rect 1728 311 1744 345
rect 1678 295 1744 311
rect 1796 345 1862 361
rect 1796 311 1812 345
rect 1846 311 1862 345
rect 1796 295 1862 311
rect 1914 345 1980 361
rect 1914 311 1930 345
rect 1964 311 1980 345
rect 1914 295 1980 311
rect 2032 345 2098 361
rect 2032 311 2048 345
rect 2082 311 2098 345
rect 2032 295 2098 311
rect 2150 345 2216 361
rect 2150 311 2166 345
rect 2200 311 2216 345
rect 2150 295 2216 311
rect 2268 345 2334 361
rect 2268 311 2284 345
rect 2318 311 2334 345
rect 2268 295 2334 311
rect 2386 345 2452 361
rect 2386 311 2402 345
rect 2436 311 2452 345
rect 2386 295 2452 311
rect 2504 345 2570 361
rect 2504 311 2520 345
rect 2554 311 2570 345
rect 2504 295 2570 311
rect 2622 345 2688 361
rect 2622 311 2638 345
rect 2672 311 2688 345
rect 2622 295 2688 311
rect 2740 345 2806 361
rect 2740 311 2756 345
rect 2790 311 2806 345
rect 2740 295 2806 311
rect 2858 345 2924 361
rect 2858 311 2874 345
rect 2908 311 2924 345
rect 2858 295 2924 311
rect -2921 264 -2861 295
rect -2803 264 -2743 295
rect -2685 264 -2625 295
rect -2567 264 -2507 295
rect -2449 264 -2389 295
rect -2331 264 -2271 295
rect -2213 264 -2153 295
rect -2095 264 -2035 295
rect -1977 264 -1917 295
rect -1859 264 -1799 295
rect -1741 264 -1681 295
rect -1623 264 -1563 295
rect -1505 264 -1445 295
rect -1387 264 -1327 295
rect -1269 264 -1209 295
rect -1151 264 -1091 295
rect -1033 264 -973 295
rect -915 264 -855 295
rect -797 264 -737 295
rect -679 264 -619 295
rect -561 264 -501 295
rect -443 264 -383 295
rect -325 264 -265 295
rect -207 264 -147 295
rect -89 264 -29 295
rect 29 264 89 295
rect 147 264 207 295
rect 265 264 325 295
rect 383 264 443 295
rect 501 264 561 295
rect 619 264 679 295
rect 737 264 797 295
rect 855 264 915 295
rect 973 264 1033 295
rect 1091 264 1151 295
rect 1209 264 1269 295
rect 1327 264 1387 295
rect 1445 264 1505 295
rect 1563 264 1623 295
rect 1681 264 1741 295
rect 1799 264 1859 295
rect 1917 264 1977 295
rect 2035 264 2095 295
rect 2153 264 2213 295
rect 2271 264 2331 295
rect 2389 264 2449 295
rect 2507 264 2567 295
rect 2625 264 2685 295
rect 2743 264 2803 295
rect 2861 264 2921 295
rect -2921 -362 -2861 -336
rect -2803 -362 -2743 -336
rect -2685 -362 -2625 -336
rect -2567 -362 -2507 -336
rect -2449 -362 -2389 -336
rect -2331 -362 -2271 -336
rect -2213 -362 -2153 -336
rect -2095 -362 -2035 -336
rect -1977 -362 -1917 -336
rect -1859 -362 -1799 -336
rect -1741 -362 -1681 -336
rect -1623 -362 -1563 -336
rect -1505 -362 -1445 -336
rect -1387 -362 -1327 -336
rect -1269 -362 -1209 -336
rect -1151 -362 -1091 -336
rect -1033 -362 -973 -336
rect -915 -362 -855 -336
rect -797 -362 -737 -336
rect -679 -362 -619 -336
rect -561 -362 -501 -336
rect -443 -362 -383 -336
rect -325 -362 -265 -336
rect -207 -362 -147 -336
rect -89 -362 -29 -336
rect 29 -362 89 -336
rect 147 -362 207 -336
rect 265 -362 325 -336
rect 383 -362 443 -336
rect 501 -362 561 -336
rect 619 -362 679 -336
rect 737 -362 797 -336
rect 855 -362 915 -336
rect 973 -362 1033 -336
rect 1091 -362 1151 -336
rect 1209 -362 1269 -336
rect 1327 -362 1387 -336
rect 1445 -362 1505 -336
rect 1563 -362 1623 -336
rect 1681 -362 1741 -336
rect 1799 -362 1859 -336
rect 1917 -362 1977 -336
rect 2035 -362 2095 -336
rect 2153 -362 2213 -336
rect 2271 -362 2331 -336
rect 2389 -362 2449 -336
rect 2507 -362 2567 -336
rect 2625 -362 2685 -336
rect 2743 -362 2803 -336
rect 2861 -362 2921 -336
<< polycont >>
rect -2908 311 -2874 345
rect -2790 311 -2756 345
rect -2672 311 -2638 345
rect -2554 311 -2520 345
rect -2436 311 -2402 345
rect -2318 311 -2284 345
rect -2200 311 -2166 345
rect -2082 311 -2048 345
rect -1964 311 -1930 345
rect -1846 311 -1812 345
rect -1728 311 -1694 345
rect -1610 311 -1576 345
rect -1492 311 -1458 345
rect -1374 311 -1340 345
rect -1256 311 -1222 345
rect -1138 311 -1104 345
rect -1020 311 -986 345
rect -902 311 -868 345
rect -784 311 -750 345
rect -666 311 -632 345
rect -548 311 -514 345
rect -430 311 -396 345
rect -312 311 -278 345
rect -194 311 -160 345
rect -76 311 -42 345
rect 42 311 76 345
rect 160 311 194 345
rect 278 311 312 345
rect 396 311 430 345
rect 514 311 548 345
rect 632 311 666 345
rect 750 311 784 345
rect 868 311 902 345
rect 986 311 1020 345
rect 1104 311 1138 345
rect 1222 311 1256 345
rect 1340 311 1374 345
rect 1458 311 1492 345
rect 1576 311 1610 345
rect 1694 311 1728 345
rect 1812 311 1846 345
rect 1930 311 1964 345
rect 2048 311 2082 345
rect 2166 311 2200 345
rect 2284 311 2318 345
rect 2402 311 2436 345
rect 2520 311 2554 345
rect 2638 311 2672 345
rect 2756 311 2790 345
rect 2874 311 2908 345
<< locali >>
rect -3081 414 -2985 448
rect 2985 414 3081 448
rect -3081 351 -3047 414
rect 3047 351 3081 414
rect -2924 311 -2908 345
rect -2874 311 -2858 345
rect -2806 311 -2790 345
rect -2756 311 -2740 345
rect -2688 311 -2672 345
rect -2638 311 -2622 345
rect -2570 311 -2554 345
rect -2520 311 -2504 345
rect -2452 311 -2436 345
rect -2402 311 -2386 345
rect -2334 311 -2318 345
rect -2284 311 -2268 345
rect -2216 311 -2200 345
rect -2166 311 -2150 345
rect -2098 311 -2082 345
rect -2048 311 -2032 345
rect -1980 311 -1964 345
rect -1930 311 -1914 345
rect -1862 311 -1846 345
rect -1812 311 -1796 345
rect -1744 311 -1728 345
rect -1694 311 -1678 345
rect -1626 311 -1610 345
rect -1576 311 -1560 345
rect -1508 311 -1492 345
rect -1458 311 -1442 345
rect -1390 311 -1374 345
rect -1340 311 -1324 345
rect -1272 311 -1256 345
rect -1222 311 -1206 345
rect -1154 311 -1138 345
rect -1104 311 -1088 345
rect -1036 311 -1020 345
rect -986 311 -970 345
rect -918 311 -902 345
rect -868 311 -852 345
rect -800 311 -784 345
rect -750 311 -734 345
rect -682 311 -666 345
rect -632 311 -616 345
rect -564 311 -548 345
rect -514 311 -498 345
rect -446 311 -430 345
rect -396 311 -380 345
rect -328 311 -312 345
rect -278 311 -262 345
rect -210 311 -194 345
rect -160 311 -144 345
rect -92 311 -76 345
rect -42 311 -26 345
rect 26 311 42 345
rect 76 311 92 345
rect 144 311 160 345
rect 194 311 210 345
rect 262 311 278 345
rect 312 311 328 345
rect 380 311 396 345
rect 430 311 446 345
rect 498 311 514 345
rect 548 311 564 345
rect 616 311 632 345
rect 666 311 682 345
rect 734 311 750 345
rect 784 311 800 345
rect 852 311 868 345
rect 902 311 918 345
rect 970 311 986 345
rect 1020 311 1036 345
rect 1088 311 1104 345
rect 1138 311 1154 345
rect 1206 311 1222 345
rect 1256 311 1272 345
rect 1324 311 1340 345
rect 1374 311 1390 345
rect 1442 311 1458 345
rect 1492 311 1508 345
rect 1560 311 1576 345
rect 1610 311 1626 345
rect 1678 311 1694 345
rect 1728 311 1744 345
rect 1796 311 1812 345
rect 1846 311 1862 345
rect 1914 311 1930 345
rect 1964 311 1980 345
rect 2032 311 2048 345
rect 2082 311 2098 345
rect 2150 311 2166 345
rect 2200 311 2216 345
rect 2268 311 2284 345
rect 2318 311 2334 345
rect 2386 311 2402 345
rect 2436 311 2452 345
rect 2504 311 2520 345
rect 2554 311 2570 345
rect 2622 311 2638 345
rect 2672 311 2688 345
rect 2740 311 2756 345
rect 2790 311 2806 345
rect 2858 311 2874 345
rect 2908 311 2924 345
rect -2967 252 -2933 268
rect -2967 -340 -2933 -324
rect -2849 252 -2815 268
rect -2849 -340 -2815 -324
rect -2731 252 -2697 268
rect -2731 -340 -2697 -324
rect -2613 252 -2579 268
rect -2613 -340 -2579 -324
rect -2495 252 -2461 268
rect -2495 -340 -2461 -324
rect -2377 252 -2343 268
rect -2377 -340 -2343 -324
rect -2259 252 -2225 268
rect -2259 -340 -2225 -324
rect -2141 252 -2107 268
rect -2141 -340 -2107 -324
rect -2023 252 -1989 268
rect -2023 -340 -1989 -324
rect -1905 252 -1871 268
rect -1905 -340 -1871 -324
rect -1787 252 -1753 268
rect -1787 -340 -1753 -324
rect -1669 252 -1635 268
rect -1669 -340 -1635 -324
rect -1551 252 -1517 268
rect -1551 -340 -1517 -324
rect -1433 252 -1399 268
rect -1433 -340 -1399 -324
rect -1315 252 -1281 268
rect -1315 -340 -1281 -324
rect -1197 252 -1163 268
rect -1197 -340 -1163 -324
rect -1079 252 -1045 268
rect -1079 -340 -1045 -324
rect -961 252 -927 268
rect -961 -340 -927 -324
rect -843 252 -809 268
rect -843 -340 -809 -324
rect -725 252 -691 268
rect -725 -340 -691 -324
rect -607 252 -573 268
rect -607 -340 -573 -324
rect -489 252 -455 268
rect -489 -340 -455 -324
rect -371 252 -337 268
rect -371 -340 -337 -324
rect -253 252 -219 268
rect -253 -340 -219 -324
rect -135 252 -101 268
rect -135 -340 -101 -324
rect -17 252 17 268
rect -17 -340 17 -324
rect 101 252 135 268
rect 101 -340 135 -324
rect 219 252 253 268
rect 219 -340 253 -324
rect 337 252 371 268
rect 337 -340 371 -324
rect 455 252 489 268
rect 455 -340 489 -324
rect 573 252 607 268
rect 573 -340 607 -324
rect 691 252 725 268
rect 691 -340 725 -324
rect 809 252 843 268
rect 809 -340 843 -324
rect 927 252 961 268
rect 927 -340 961 -324
rect 1045 252 1079 268
rect 1045 -340 1079 -324
rect 1163 252 1197 268
rect 1163 -340 1197 -324
rect 1281 252 1315 268
rect 1281 -340 1315 -324
rect 1399 252 1433 268
rect 1399 -340 1433 -324
rect 1517 252 1551 268
rect 1517 -340 1551 -324
rect 1635 252 1669 268
rect 1635 -340 1669 -324
rect 1753 252 1787 268
rect 1753 -340 1787 -324
rect 1871 252 1905 268
rect 1871 -340 1905 -324
rect 1989 252 2023 268
rect 1989 -340 2023 -324
rect 2107 252 2141 268
rect 2107 -340 2141 -324
rect 2225 252 2259 268
rect 2225 -340 2259 -324
rect 2343 252 2377 268
rect 2343 -340 2377 -324
rect 2461 252 2495 268
rect 2461 -340 2495 -324
rect 2579 252 2613 268
rect 2579 -340 2613 -324
rect 2697 252 2731 268
rect 2697 -340 2731 -324
rect 2815 252 2849 268
rect 2815 -340 2849 -324
rect 2933 252 2967 268
rect 2933 -340 2967 -324
rect -3081 -414 -3047 -351
rect 3047 -414 3081 -351
rect -3081 -448 -2985 -414
rect 2985 -448 3081 -414
<< viali >>
rect -2908 311 -2874 345
rect -2790 311 -2756 345
rect -2672 311 -2638 345
rect -2554 311 -2520 345
rect -2436 311 -2402 345
rect -2318 311 -2284 345
rect -2200 311 -2166 345
rect -2082 311 -2048 345
rect -1964 311 -1930 345
rect -1846 311 -1812 345
rect -1728 311 -1694 345
rect -1610 311 -1576 345
rect -1492 311 -1458 345
rect -1374 311 -1340 345
rect -1256 311 -1222 345
rect -1138 311 -1104 345
rect -1020 311 -986 345
rect -902 311 -868 345
rect -784 311 -750 345
rect -666 311 -632 345
rect -548 311 -514 345
rect -430 311 -396 345
rect -312 311 -278 345
rect -194 311 -160 345
rect -76 311 -42 345
rect 42 311 76 345
rect 160 311 194 345
rect 278 311 312 345
rect 396 311 430 345
rect 514 311 548 345
rect 632 311 666 345
rect 750 311 784 345
rect 868 311 902 345
rect 986 311 1020 345
rect 1104 311 1138 345
rect 1222 311 1256 345
rect 1340 311 1374 345
rect 1458 311 1492 345
rect 1576 311 1610 345
rect 1694 311 1728 345
rect 1812 311 1846 345
rect 1930 311 1964 345
rect 2048 311 2082 345
rect 2166 311 2200 345
rect 2284 311 2318 345
rect 2402 311 2436 345
rect 2520 311 2554 345
rect 2638 311 2672 345
rect 2756 311 2790 345
rect 2874 311 2908 345
rect -2967 -324 -2933 252
rect -2849 -324 -2815 252
rect -2731 -324 -2697 252
rect -2613 -324 -2579 252
rect -2495 -324 -2461 252
rect -2377 -324 -2343 252
rect -2259 -324 -2225 252
rect -2141 -324 -2107 252
rect -2023 -324 -1989 252
rect -1905 -324 -1871 252
rect -1787 -324 -1753 252
rect -1669 -324 -1635 252
rect -1551 -324 -1517 252
rect -1433 -324 -1399 252
rect -1315 -324 -1281 252
rect -1197 -324 -1163 252
rect -1079 -324 -1045 252
rect -961 -324 -927 252
rect -843 -324 -809 252
rect -725 -324 -691 252
rect -607 -324 -573 252
rect -489 -324 -455 252
rect -371 -324 -337 252
rect -253 -324 -219 252
rect -135 -324 -101 252
rect -17 -324 17 252
rect 101 -324 135 252
rect 219 -324 253 252
rect 337 -324 371 252
rect 455 -324 489 252
rect 573 -324 607 252
rect 691 -324 725 252
rect 809 -324 843 252
rect 927 -324 961 252
rect 1045 -324 1079 252
rect 1163 -324 1197 252
rect 1281 -324 1315 252
rect 1399 -324 1433 252
rect 1517 -324 1551 252
rect 1635 -324 1669 252
rect 1753 -324 1787 252
rect 1871 -324 1905 252
rect 1989 -324 2023 252
rect 2107 -324 2141 252
rect 2225 -324 2259 252
rect 2343 -324 2377 252
rect 2461 -324 2495 252
rect 2579 -324 2613 252
rect 2697 -324 2731 252
rect 2815 -324 2849 252
rect 2933 -324 2967 252
<< metal1 >>
rect -2920 345 -2862 351
rect -2920 311 -2908 345
rect -2874 311 -2862 345
rect -2920 305 -2862 311
rect -2802 345 -2744 351
rect -2802 311 -2790 345
rect -2756 311 -2744 345
rect -2802 305 -2744 311
rect -2684 345 -2626 351
rect -2684 311 -2672 345
rect -2638 311 -2626 345
rect -2684 305 -2626 311
rect -2566 345 -2508 351
rect -2566 311 -2554 345
rect -2520 311 -2508 345
rect -2566 305 -2508 311
rect -2448 345 -2390 351
rect -2448 311 -2436 345
rect -2402 311 -2390 345
rect -2448 305 -2390 311
rect -2330 345 -2272 351
rect -2330 311 -2318 345
rect -2284 311 -2272 345
rect -2330 305 -2272 311
rect -2212 345 -2154 351
rect -2212 311 -2200 345
rect -2166 311 -2154 345
rect -2212 305 -2154 311
rect -2094 345 -2036 351
rect -2094 311 -2082 345
rect -2048 311 -2036 345
rect -2094 305 -2036 311
rect -1976 345 -1918 351
rect -1976 311 -1964 345
rect -1930 311 -1918 345
rect -1976 305 -1918 311
rect -1858 345 -1800 351
rect -1858 311 -1846 345
rect -1812 311 -1800 345
rect -1858 305 -1800 311
rect -1740 345 -1682 351
rect -1740 311 -1728 345
rect -1694 311 -1682 345
rect -1740 305 -1682 311
rect -1622 345 -1564 351
rect -1622 311 -1610 345
rect -1576 311 -1564 345
rect -1622 305 -1564 311
rect -1504 345 -1446 351
rect -1504 311 -1492 345
rect -1458 311 -1446 345
rect -1504 305 -1446 311
rect -1386 345 -1328 351
rect -1386 311 -1374 345
rect -1340 311 -1328 345
rect -1386 305 -1328 311
rect -1268 345 -1210 351
rect -1268 311 -1256 345
rect -1222 311 -1210 345
rect -1268 305 -1210 311
rect -1150 345 -1092 351
rect -1150 311 -1138 345
rect -1104 311 -1092 345
rect -1150 305 -1092 311
rect -1032 345 -974 351
rect -1032 311 -1020 345
rect -986 311 -974 345
rect -1032 305 -974 311
rect -914 345 -856 351
rect -914 311 -902 345
rect -868 311 -856 345
rect -914 305 -856 311
rect -796 345 -738 351
rect -796 311 -784 345
rect -750 311 -738 345
rect -796 305 -738 311
rect -678 345 -620 351
rect -678 311 -666 345
rect -632 311 -620 345
rect -678 305 -620 311
rect -560 345 -502 351
rect -560 311 -548 345
rect -514 311 -502 345
rect -560 305 -502 311
rect -442 345 -384 351
rect -442 311 -430 345
rect -396 311 -384 345
rect -442 305 -384 311
rect -324 345 -266 351
rect -324 311 -312 345
rect -278 311 -266 345
rect -324 305 -266 311
rect -206 345 -148 351
rect -206 311 -194 345
rect -160 311 -148 345
rect -206 305 -148 311
rect -88 345 -30 351
rect -88 311 -76 345
rect -42 311 -30 345
rect -88 305 -30 311
rect 30 345 88 351
rect 30 311 42 345
rect 76 311 88 345
rect 30 305 88 311
rect 148 345 206 351
rect 148 311 160 345
rect 194 311 206 345
rect 148 305 206 311
rect 266 345 324 351
rect 266 311 278 345
rect 312 311 324 345
rect 266 305 324 311
rect 384 345 442 351
rect 384 311 396 345
rect 430 311 442 345
rect 384 305 442 311
rect 502 345 560 351
rect 502 311 514 345
rect 548 311 560 345
rect 502 305 560 311
rect 620 345 678 351
rect 620 311 632 345
rect 666 311 678 345
rect 620 305 678 311
rect 738 345 796 351
rect 738 311 750 345
rect 784 311 796 345
rect 738 305 796 311
rect 856 345 914 351
rect 856 311 868 345
rect 902 311 914 345
rect 856 305 914 311
rect 974 345 1032 351
rect 974 311 986 345
rect 1020 311 1032 345
rect 974 305 1032 311
rect 1092 345 1150 351
rect 1092 311 1104 345
rect 1138 311 1150 345
rect 1092 305 1150 311
rect 1210 345 1268 351
rect 1210 311 1222 345
rect 1256 311 1268 345
rect 1210 305 1268 311
rect 1328 345 1386 351
rect 1328 311 1340 345
rect 1374 311 1386 345
rect 1328 305 1386 311
rect 1446 345 1504 351
rect 1446 311 1458 345
rect 1492 311 1504 345
rect 1446 305 1504 311
rect 1564 345 1622 351
rect 1564 311 1576 345
rect 1610 311 1622 345
rect 1564 305 1622 311
rect 1682 345 1740 351
rect 1682 311 1694 345
rect 1728 311 1740 345
rect 1682 305 1740 311
rect 1800 345 1858 351
rect 1800 311 1812 345
rect 1846 311 1858 345
rect 1800 305 1858 311
rect 1918 345 1976 351
rect 1918 311 1930 345
rect 1964 311 1976 345
rect 1918 305 1976 311
rect 2036 345 2094 351
rect 2036 311 2048 345
rect 2082 311 2094 345
rect 2036 305 2094 311
rect 2154 345 2212 351
rect 2154 311 2166 345
rect 2200 311 2212 345
rect 2154 305 2212 311
rect 2272 345 2330 351
rect 2272 311 2284 345
rect 2318 311 2330 345
rect 2272 305 2330 311
rect 2390 345 2448 351
rect 2390 311 2402 345
rect 2436 311 2448 345
rect 2390 305 2448 311
rect 2508 345 2566 351
rect 2508 311 2520 345
rect 2554 311 2566 345
rect 2508 305 2566 311
rect 2626 345 2684 351
rect 2626 311 2638 345
rect 2672 311 2684 345
rect 2626 305 2684 311
rect 2744 345 2802 351
rect 2744 311 2756 345
rect 2790 311 2802 345
rect 2744 305 2802 311
rect 2862 345 2920 351
rect 2862 311 2874 345
rect 2908 311 2920 345
rect 2862 305 2920 311
rect -2973 252 -2927 264
rect -2973 -324 -2967 252
rect -2933 -324 -2927 252
rect -2973 -336 -2927 -324
rect -2855 252 -2809 264
rect -2855 -324 -2849 252
rect -2815 -324 -2809 252
rect -2855 -336 -2809 -324
rect -2737 252 -2691 264
rect -2737 -324 -2731 252
rect -2697 -324 -2691 252
rect -2737 -336 -2691 -324
rect -2619 252 -2573 264
rect -2619 -324 -2613 252
rect -2579 -324 -2573 252
rect -2619 -336 -2573 -324
rect -2501 252 -2455 264
rect -2501 -324 -2495 252
rect -2461 -324 -2455 252
rect -2501 -336 -2455 -324
rect -2383 252 -2337 264
rect -2383 -324 -2377 252
rect -2343 -324 -2337 252
rect -2383 -336 -2337 -324
rect -2265 252 -2219 264
rect -2265 -324 -2259 252
rect -2225 -324 -2219 252
rect -2265 -336 -2219 -324
rect -2147 252 -2101 264
rect -2147 -324 -2141 252
rect -2107 -324 -2101 252
rect -2147 -336 -2101 -324
rect -2029 252 -1983 264
rect -2029 -324 -2023 252
rect -1989 -324 -1983 252
rect -2029 -336 -1983 -324
rect -1911 252 -1865 264
rect -1911 -324 -1905 252
rect -1871 -324 -1865 252
rect -1911 -336 -1865 -324
rect -1793 252 -1747 264
rect -1793 -324 -1787 252
rect -1753 -324 -1747 252
rect -1793 -336 -1747 -324
rect -1675 252 -1629 264
rect -1675 -324 -1669 252
rect -1635 -324 -1629 252
rect -1675 -336 -1629 -324
rect -1557 252 -1511 264
rect -1557 -324 -1551 252
rect -1517 -324 -1511 252
rect -1557 -336 -1511 -324
rect -1439 252 -1393 264
rect -1439 -324 -1433 252
rect -1399 -324 -1393 252
rect -1439 -336 -1393 -324
rect -1321 252 -1275 264
rect -1321 -324 -1315 252
rect -1281 -324 -1275 252
rect -1321 -336 -1275 -324
rect -1203 252 -1157 264
rect -1203 -324 -1197 252
rect -1163 -324 -1157 252
rect -1203 -336 -1157 -324
rect -1085 252 -1039 264
rect -1085 -324 -1079 252
rect -1045 -324 -1039 252
rect -1085 -336 -1039 -324
rect -967 252 -921 264
rect -967 -324 -961 252
rect -927 -324 -921 252
rect -967 -336 -921 -324
rect -849 252 -803 264
rect -849 -324 -843 252
rect -809 -324 -803 252
rect -849 -336 -803 -324
rect -731 252 -685 264
rect -731 -324 -725 252
rect -691 -324 -685 252
rect -731 -336 -685 -324
rect -613 252 -567 264
rect -613 -324 -607 252
rect -573 -324 -567 252
rect -613 -336 -567 -324
rect -495 252 -449 264
rect -495 -324 -489 252
rect -455 -324 -449 252
rect -495 -336 -449 -324
rect -377 252 -331 264
rect -377 -324 -371 252
rect -337 -324 -331 252
rect -377 -336 -331 -324
rect -259 252 -213 264
rect -259 -324 -253 252
rect -219 -324 -213 252
rect -259 -336 -213 -324
rect -141 252 -95 264
rect -141 -324 -135 252
rect -101 -324 -95 252
rect -141 -336 -95 -324
rect -23 252 23 264
rect -23 -324 -17 252
rect 17 -324 23 252
rect -23 -336 23 -324
rect 95 252 141 264
rect 95 -324 101 252
rect 135 -324 141 252
rect 95 -336 141 -324
rect 213 252 259 264
rect 213 -324 219 252
rect 253 -324 259 252
rect 213 -336 259 -324
rect 331 252 377 264
rect 331 -324 337 252
rect 371 -324 377 252
rect 331 -336 377 -324
rect 449 252 495 264
rect 449 -324 455 252
rect 489 -324 495 252
rect 449 -336 495 -324
rect 567 252 613 264
rect 567 -324 573 252
rect 607 -324 613 252
rect 567 -336 613 -324
rect 685 252 731 264
rect 685 -324 691 252
rect 725 -324 731 252
rect 685 -336 731 -324
rect 803 252 849 264
rect 803 -324 809 252
rect 843 -324 849 252
rect 803 -336 849 -324
rect 921 252 967 264
rect 921 -324 927 252
rect 961 -324 967 252
rect 921 -336 967 -324
rect 1039 252 1085 264
rect 1039 -324 1045 252
rect 1079 -324 1085 252
rect 1039 -336 1085 -324
rect 1157 252 1203 264
rect 1157 -324 1163 252
rect 1197 -324 1203 252
rect 1157 -336 1203 -324
rect 1275 252 1321 264
rect 1275 -324 1281 252
rect 1315 -324 1321 252
rect 1275 -336 1321 -324
rect 1393 252 1439 264
rect 1393 -324 1399 252
rect 1433 -324 1439 252
rect 1393 -336 1439 -324
rect 1511 252 1557 264
rect 1511 -324 1517 252
rect 1551 -324 1557 252
rect 1511 -336 1557 -324
rect 1629 252 1675 264
rect 1629 -324 1635 252
rect 1669 -324 1675 252
rect 1629 -336 1675 -324
rect 1747 252 1793 264
rect 1747 -324 1753 252
rect 1787 -324 1793 252
rect 1747 -336 1793 -324
rect 1865 252 1911 264
rect 1865 -324 1871 252
rect 1905 -324 1911 252
rect 1865 -336 1911 -324
rect 1983 252 2029 264
rect 1983 -324 1989 252
rect 2023 -324 2029 252
rect 1983 -336 2029 -324
rect 2101 252 2147 264
rect 2101 -324 2107 252
rect 2141 -324 2147 252
rect 2101 -336 2147 -324
rect 2219 252 2265 264
rect 2219 -324 2225 252
rect 2259 -324 2265 252
rect 2219 -336 2265 -324
rect 2337 252 2383 264
rect 2337 -324 2343 252
rect 2377 -324 2383 252
rect 2337 -336 2383 -324
rect 2455 252 2501 264
rect 2455 -324 2461 252
rect 2495 -324 2501 252
rect 2455 -336 2501 -324
rect 2573 252 2619 264
rect 2573 -324 2579 252
rect 2613 -324 2619 252
rect 2573 -336 2619 -324
rect 2691 252 2737 264
rect 2691 -324 2697 252
rect 2731 -324 2737 252
rect 2691 -336 2737 -324
rect 2809 252 2855 264
rect 2809 -324 2815 252
rect 2849 -324 2855 252
rect 2809 -336 2855 -324
rect 2927 252 2973 264
rect 2927 -324 2933 252
rect 2967 -324 2973 252
rect 2927 -336 2973 -324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -431 3064 431
string parameters w 3 l 0.3 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
