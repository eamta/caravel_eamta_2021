magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect -10 906 17 924
rect 129 919 187 925
rect 129 908 141 919
rect 129 906 175 908
rect 316 906 386 1042
rect 498 974 556 980
rect 498 940 510 974
rect 668 951 702 969
rect 1090 951 1125 969
rect 498 934 556 940
rect 668 915 738 951
rect 1054 936 1125 951
rect 1405 936 1440 970
rect -28 870 386 906
rect 685 906 817 915
rect 466 870 500 904
rect 554 870 588 904
rect -28 836 622 870
rect -28 564 386 836
rect 585 798 600 813
rect 542 768 600 798
rect 454 713 512 746
rect 520 713 528 754
rect 542 746 570 768
rect 585 753 600 768
rect 668 798 679 809
rect 685 798 864 906
rect 668 768 864 798
rect 867 813 925 819
rect 867 779 892 813
rect 867 773 925 779
rect 668 757 679 768
rect 540 713 600 746
rect 466 709 500 713
rect 512 700 528 713
rect 554 709 588 713
rect 406 564 420 696
rect 432 692 440 696
rect 476 692 528 700
rect 582 692 616 696
rect 432 685 446 692
rect 432 680 440 685
rect 476 666 540 692
rect 544 675 616 692
rect 668 694 682 746
rect 685 694 864 768
rect 544 666 594 675
rect 494 632 594 666
rect 494 616 540 632
rect 548 626 556 632
rect 576 598 594 632
rect 668 564 864 694
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect -28 547 628 564
rect 352 530 628 547
rect 682 530 864 564
rect 494 508 528 530
rect 685 441 864 530
rect 1054 477 1124 936
rect 1406 917 1440 936
rect 1236 868 1294 874
rect 1236 834 1248 868
rect 1236 828 1294 834
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1054 388 1118 441
rect 1425 424 1440 917
rect 1459 883 1494 917
rect 1774 883 1809 917
rect 1459 424 1493 883
rect 1775 864 1809 883
rect 1605 815 1663 821
rect 1605 781 1617 815
rect 1605 775 1663 781
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1794 371 1809 864
rect 1828 830 1863 864
rect 2143 830 2178 864
rect 1828 371 1862 830
rect 2144 811 2178 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2163 318 2178 811
rect 2197 777 2232 811
rect 2512 777 2547 794
rect 2197 318 2231 777
rect 2513 776 2547 777
rect 2513 740 2583 776
rect 2343 709 2401 715
rect 2343 675 2355 709
rect 2530 706 2601 740
rect 2881 706 2916 740
rect 2343 669 2401 675
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2530 265 2600 706
rect 2882 687 2916 706
rect 2712 638 2770 644
rect 2712 604 2724 638
rect 2712 598 2770 604
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
rect 196 54 200 200
rect 224 82 228 228
rect 2901 212 2916 687
rect 2935 653 2970 687
rect 3250 653 3285 687
rect 2935 212 2969 653
rect 3251 634 3285 653
rect 3081 585 3139 591
rect 3081 551 3093 585
rect 3081 545 3139 551
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3270 159 3285 634
rect 3304 600 3339 634
rect 3619 600 3654 634
rect 3304 159 3338 600
rect 3620 581 3654 600
rect 4006 581 4059 582
rect 3450 532 3508 538
rect 3450 498 3462 532
rect 3450 492 3508 498
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 581
rect 3673 547 3708 581
rect 3988 547 4059 581
rect 3673 106 3707 547
rect 3989 546 4059 547
rect 4006 512 4077 546
rect 3819 479 3877 485
rect 3819 445 3831 479
rect 3819 439 3877 445
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4006 53 4076 512
rect 4188 444 4246 450
rect 4188 410 4200 444
rect 4188 404 4246 410
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4006 17 4059 53
<< nwell >>
rect -28 366 864 906
<< psubdiff >>
rect 54 -66 78 -32
rect 750 -66 774 -32
<< nsubdiff >>
rect 44 836 252 870
rect 598 836 764 870
<< psubdiffcont >>
rect 78 -66 750 -32
<< nsubdiffcont >>
rect 252 836 598 870
<< poly >>
rect 540 768 770 798
rect 540 692 570 768
rect 76 496 106 692
rect 76 466 306 496
rect 76 422 106 466
rect 364 424 394 514
rect -28 392 106 422
rect 76 308 106 392
rect 180 408 394 424
rect 180 374 196 408
rect 230 394 394 408
rect 452 432 482 514
rect 740 492 770 768
rect 646 462 770 492
rect 452 416 590 432
rect 452 402 540 416
rect 230 374 246 394
rect 180 358 246 374
rect 364 360 394 394
rect 524 382 540 402
rect 574 382 590 416
rect 524 366 590 382
rect 364 330 482 360
rect 76 278 306 308
rect -28 14 2 242
rect 76 86 106 278
rect 452 262 482 330
rect 540 262 570 366
rect 646 232 676 462
rect 718 338 784 354
rect 718 304 734 338
rect 768 304 784 338
rect 718 274 864 304
rect 646 202 770 232
rect 364 14 394 108
rect 740 14 770 202
rect -28 -16 770 14
<< polycont >>
rect 196 374 230 408
rect 540 382 574 416
rect 734 304 768 338
<< locali >>
rect 180 374 196 408
rect 230 374 246 408
rect 524 382 540 416
rect 574 382 590 416
rect 718 304 734 338
rect 768 304 784 338
<< viali >>
rect 16 836 252 870
rect 252 836 598 870
rect 598 836 814 870
rect 196 374 230 408
rect 540 382 574 416
rect 734 304 768 338
rect 42 -66 78 -32
rect 78 -66 750 -32
rect 750 -66 790 -32
<< metal1 >>
rect -28 870 864 878
rect -28 836 16 870
rect 814 836 864 870
rect -28 782 864 836
rect 30 524 64 782
rect 118 408 152 680
rect 230 524 264 782
rect 318 720 528 754
rect 318 680 352 720
rect 494 680 528 720
rect 180 408 246 424
rect 118 374 196 408
rect 230 374 246 408
rect 118 200 152 374
rect 180 358 246 374
rect 406 324 440 680
rect 582 524 616 782
rect 694 432 728 676
rect 782 520 816 782
rect 524 416 846 432
rect 524 382 540 416
rect 574 398 846 416
rect 574 382 590 398
rect 524 366 590 382
rect 718 338 784 354
rect 718 324 734 338
rect 406 304 734 324
rect 768 304 784 338
rect 406 290 784 304
rect 0 16 200 200
rect 230 16 264 234
rect 406 94 440 290
rect 718 288 784 290
rect 582 16 616 238
rect 812 202 846 398
rect 694 168 846 202
rect 694 64 728 168
rect 782 16 816 128
rect -28 -32 864 16
rect -28 -66 42 -32
rect 790 -66 864 -32
rect -28 -72 864 -66
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_01v8_J83WCX  sky130_fd_pr__nfet_01v8_J83WCX_0
timestamp 1615216760
transform 1 0 91 0 1 188
box -73 -102 73 40
use sky130_fd_pr__nfet_01v8_H7KMG3  sky130_fd_pr__nfet_01v8_H7KMG3_2
timestamp 1615216760
transform 1 0 467 0 1 203
box -73 -147 73 85
use sky130_fd_pr__nfet_01v8_H7KMG3  sky130_fd_pr__nfet_01v8_H7KMG3_1
timestamp 1615216760
transform 1 0 379 0 1 203
box -73 -147 73 85
use sky130_fd_pr__nfet_01v8_H7KMG3  sky130_fd_pr__nfet_01v8_H7KMG3_0
timestamp 1615216760
transform 1 0 291 0 1 203
box -73 -147 73 85
use sky130_fd_pr__nfet_01v8_H7KMG3  sky130_fd_pr__nfet_01v8_H7KMG3_3
timestamp 1615216760
transform 1 0 555 0 1 203
box -73 -147 73 85
use sky130_fd_pr__nfet_01v8_J83WCX  sky130_fd_pr__nfet_01v8_J83WCX_1
timestamp 1615216760
transform 1 0 755 0 1 126
box -73 -102 73 40
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 1634 0 1 644
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM7
timestamp 1624053917
transform 1 0 2372 0 1 538
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM6
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_L9ESED  XM10
timestamp 1624053917
transform 1 0 3110 0 1 423
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM9
timestamp 1624053917
transform 1 0 2741 0 1 476
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_XSLFBL  XM8
timestamp 1624053917
transform 1 0 4217 0 1 273
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_L9ESED  XM12
timestamp 1624053917
transform 1 0 3848 0 1 317
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM11
timestamp 1624053917
transform 1 0 3479 0 1 370
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_1
timestamp 1615394250
transform 1 0 291 0 1 602
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_0
timestamp 1615394250
transform 1 0 91 0 1 664
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_2
timestamp 1615394250
transform 1 0 379 0 1 602
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_3
timestamp 1615394250
transform 1 0 467 0 1 602
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_4
timestamp 1615394250
transform 1 0 555 0 1 602
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AY9XA  sky130_fd_pr__pfet_01v8_5AY9XA_5
timestamp 1615394250
transform 1 0 755 0 1 604
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM1
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM4
timestamp 1624053917
transform 1 0 1265 0 1 697
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM3
timestamp 1624053917
transform 1 0 896 0 1 696
box -211 -255 211 255
<< labels >>
rlabel poly -28 -16 2 242 1 in2
rlabel metal1 42 -66 790 -32 1 vss
rlabel poly 718 274 864 304 1 out
rlabel metal1 -22 834 8 868 1 vdd
rlabel poly -28 392 106 422 1 in1
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 in2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 in1
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
<< end >>
