magic
tech sky130A
magscale 1 2
timestamp 1616185029
<< error_p >>
rect -2920 -311 -2862 -305
rect -2802 -311 -2744 -305
rect -2684 -311 -2626 -305
rect -2566 -311 -2508 -305
rect -2448 -311 -2390 -305
rect -2330 -311 -2272 -305
rect -2212 -311 -2154 -305
rect -2094 -311 -2036 -305
rect -1976 -311 -1918 -305
rect -1858 -311 -1800 -305
rect -1740 -311 -1682 -305
rect -1622 -311 -1564 -305
rect -1504 -311 -1446 -305
rect -1386 -311 -1328 -305
rect -1268 -311 -1210 -305
rect -1150 -311 -1092 -305
rect -1032 -311 -974 -305
rect -914 -311 -856 -305
rect -796 -311 -738 -305
rect -678 -311 -620 -305
rect -560 -311 -502 -305
rect -442 -311 -384 -305
rect -324 -311 -266 -305
rect -206 -311 -148 -305
rect -88 -311 -30 -305
rect 30 -311 88 -305
rect 148 -311 206 -305
rect 266 -311 324 -305
rect 384 -311 442 -305
rect 502 -311 560 -305
rect 620 -311 678 -305
rect 738 -311 796 -305
rect 856 -311 914 -305
rect 974 -311 1032 -305
rect 1092 -311 1150 -305
rect 1210 -311 1268 -305
rect 1328 -311 1386 -305
rect 1446 -311 1504 -305
rect 1564 -311 1622 -305
rect 1682 -311 1740 -305
rect 1800 -311 1858 -305
rect 1918 -311 1976 -305
rect 2036 -311 2094 -305
rect 2154 -311 2212 -305
rect 2272 -311 2330 -305
rect 2390 -311 2448 -305
rect 2508 -311 2566 -305
rect 2626 -311 2684 -305
rect 2744 -311 2802 -305
rect 2862 -311 2920 -305
rect -2920 -345 -2908 -311
rect -2802 -345 -2790 -311
rect -2684 -345 -2672 -311
rect -2566 -345 -2554 -311
rect -2448 -345 -2436 -311
rect -2330 -345 -2318 -311
rect -2212 -345 -2200 -311
rect -2094 -345 -2082 -311
rect -1976 -345 -1964 -311
rect -1858 -345 -1846 -311
rect -1740 -345 -1728 -311
rect -1622 -345 -1610 -311
rect -1504 -345 -1492 -311
rect -1386 -345 -1374 -311
rect -1268 -345 -1256 -311
rect -1150 -345 -1138 -311
rect -1032 -345 -1020 -311
rect -914 -345 -902 -311
rect -796 -345 -784 -311
rect -678 -345 -666 -311
rect -560 -345 -548 -311
rect -442 -345 -430 -311
rect -324 -345 -312 -311
rect -206 -345 -194 -311
rect -88 -345 -76 -311
rect 30 -345 42 -311
rect 148 -345 160 -311
rect 266 -345 278 -311
rect 384 -345 396 -311
rect 502 -345 514 -311
rect 620 -345 632 -311
rect 738 -345 750 -311
rect 856 -345 868 -311
rect 974 -345 986 -311
rect 1092 -345 1104 -311
rect 1210 -345 1222 -311
rect 1328 -345 1340 -311
rect 1446 -345 1458 -311
rect 1564 -345 1576 -311
rect 1682 -345 1694 -311
rect 1800 -345 1812 -311
rect 1918 -345 1930 -311
rect 2036 -345 2048 -311
rect 2154 -345 2166 -311
rect 2272 -345 2284 -311
rect 2390 -345 2402 -311
rect 2508 -345 2520 -311
rect 2626 -345 2638 -311
rect 2744 -345 2756 -311
rect 2862 -345 2874 -311
rect -2920 -351 -2862 -345
rect -2802 -351 -2744 -345
rect -2684 -351 -2626 -345
rect -2566 -351 -2508 -345
rect -2448 -351 -2390 -345
rect -2330 -351 -2272 -345
rect -2212 -351 -2154 -345
rect -2094 -351 -2036 -345
rect -1976 -351 -1918 -345
rect -1858 -351 -1800 -345
rect -1740 -351 -1682 -345
rect -1622 -351 -1564 -345
rect -1504 -351 -1446 -345
rect -1386 -351 -1328 -345
rect -1268 -351 -1210 -345
rect -1150 -351 -1092 -345
rect -1032 -351 -974 -345
rect -914 -351 -856 -345
rect -796 -351 -738 -345
rect -678 -351 -620 -345
rect -560 -351 -502 -345
rect -442 -351 -384 -345
rect -324 -351 -266 -345
rect -206 -351 -148 -345
rect -88 -351 -30 -345
rect 30 -351 88 -345
rect 148 -351 206 -345
rect 266 -351 324 -345
rect 384 -351 442 -345
rect 502 -351 560 -345
rect 620 -351 678 -345
rect 738 -351 796 -345
rect 856 -351 914 -345
rect 974 -351 1032 -345
rect 1092 -351 1150 -345
rect 1210 -351 1268 -345
rect 1328 -351 1386 -345
rect 1446 -351 1504 -345
rect 1564 -351 1622 -345
rect 1682 -351 1740 -345
rect 1800 -351 1858 -345
rect 1918 -351 1976 -345
rect 2036 -351 2094 -345
rect 2154 -351 2212 -345
rect 2272 -351 2330 -345
rect 2390 -351 2448 -345
rect 2508 -351 2566 -345
rect 2626 -351 2684 -345
rect 2744 -351 2802 -345
rect 2862 -351 2920 -345
<< nwell >>
rect -3117 -484 3117 484
<< pmos >>
rect -2921 -264 -2861 336
rect -2803 -264 -2743 336
rect -2685 -264 -2625 336
rect -2567 -264 -2507 336
rect -2449 -264 -2389 336
rect -2331 -264 -2271 336
rect -2213 -264 -2153 336
rect -2095 -264 -2035 336
rect -1977 -264 -1917 336
rect -1859 -264 -1799 336
rect -1741 -264 -1681 336
rect -1623 -264 -1563 336
rect -1505 -264 -1445 336
rect -1387 -264 -1327 336
rect -1269 -264 -1209 336
rect -1151 -264 -1091 336
rect -1033 -264 -973 336
rect -915 -264 -855 336
rect -797 -264 -737 336
rect -679 -264 -619 336
rect -561 -264 -501 336
rect -443 -264 -383 336
rect -325 -264 -265 336
rect -207 -264 -147 336
rect -89 -264 -29 336
rect 29 -264 89 336
rect 147 -264 207 336
rect 265 -264 325 336
rect 383 -264 443 336
rect 501 -264 561 336
rect 619 -264 679 336
rect 737 -264 797 336
rect 855 -264 915 336
rect 973 -264 1033 336
rect 1091 -264 1151 336
rect 1209 -264 1269 336
rect 1327 -264 1387 336
rect 1445 -264 1505 336
rect 1563 -264 1623 336
rect 1681 -264 1741 336
rect 1799 -264 1859 336
rect 1917 -264 1977 336
rect 2035 -264 2095 336
rect 2153 -264 2213 336
rect 2271 -264 2331 336
rect 2389 -264 2449 336
rect 2507 -264 2567 336
rect 2625 -264 2685 336
rect 2743 -264 2803 336
rect 2861 -264 2921 336
<< pdiff >>
rect -2979 324 -2921 336
rect -2979 -252 -2967 324
rect -2933 -252 -2921 324
rect -2979 -264 -2921 -252
rect -2861 324 -2803 336
rect -2861 -252 -2849 324
rect -2815 -252 -2803 324
rect -2861 -264 -2803 -252
rect -2743 324 -2685 336
rect -2743 -252 -2731 324
rect -2697 -252 -2685 324
rect -2743 -264 -2685 -252
rect -2625 324 -2567 336
rect -2625 -252 -2613 324
rect -2579 -252 -2567 324
rect -2625 -264 -2567 -252
rect -2507 324 -2449 336
rect -2507 -252 -2495 324
rect -2461 -252 -2449 324
rect -2507 -264 -2449 -252
rect -2389 324 -2331 336
rect -2389 -252 -2377 324
rect -2343 -252 -2331 324
rect -2389 -264 -2331 -252
rect -2271 324 -2213 336
rect -2271 -252 -2259 324
rect -2225 -252 -2213 324
rect -2271 -264 -2213 -252
rect -2153 324 -2095 336
rect -2153 -252 -2141 324
rect -2107 -252 -2095 324
rect -2153 -264 -2095 -252
rect -2035 324 -1977 336
rect -2035 -252 -2023 324
rect -1989 -252 -1977 324
rect -2035 -264 -1977 -252
rect -1917 324 -1859 336
rect -1917 -252 -1905 324
rect -1871 -252 -1859 324
rect -1917 -264 -1859 -252
rect -1799 324 -1741 336
rect -1799 -252 -1787 324
rect -1753 -252 -1741 324
rect -1799 -264 -1741 -252
rect -1681 324 -1623 336
rect -1681 -252 -1669 324
rect -1635 -252 -1623 324
rect -1681 -264 -1623 -252
rect -1563 324 -1505 336
rect -1563 -252 -1551 324
rect -1517 -252 -1505 324
rect -1563 -264 -1505 -252
rect -1445 324 -1387 336
rect -1445 -252 -1433 324
rect -1399 -252 -1387 324
rect -1445 -264 -1387 -252
rect -1327 324 -1269 336
rect -1327 -252 -1315 324
rect -1281 -252 -1269 324
rect -1327 -264 -1269 -252
rect -1209 324 -1151 336
rect -1209 -252 -1197 324
rect -1163 -252 -1151 324
rect -1209 -264 -1151 -252
rect -1091 324 -1033 336
rect -1091 -252 -1079 324
rect -1045 -252 -1033 324
rect -1091 -264 -1033 -252
rect -973 324 -915 336
rect -973 -252 -961 324
rect -927 -252 -915 324
rect -973 -264 -915 -252
rect -855 324 -797 336
rect -855 -252 -843 324
rect -809 -252 -797 324
rect -855 -264 -797 -252
rect -737 324 -679 336
rect -737 -252 -725 324
rect -691 -252 -679 324
rect -737 -264 -679 -252
rect -619 324 -561 336
rect -619 -252 -607 324
rect -573 -252 -561 324
rect -619 -264 -561 -252
rect -501 324 -443 336
rect -501 -252 -489 324
rect -455 -252 -443 324
rect -501 -264 -443 -252
rect -383 324 -325 336
rect -383 -252 -371 324
rect -337 -252 -325 324
rect -383 -264 -325 -252
rect -265 324 -207 336
rect -265 -252 -253 324
rect -219 -252 -207 324
rect -265 -264 -207 -252
rect -147 324 -89 336
rect -147 -252 -135 324
rect -101 -252 -89 324
rect -147 -264 -89 -252
rect -29 324 29 336
rect -29 -252 -17 324
rect 17 -252 29 324
rect -29 -264 29 -252
rect 89 324 147 336
rect 89 -252 101 324
rect 135 -252 147 324
rect 89 -264 147 -252
rect 207 324 265 336
rect 207 -252 219 324
rect 253 -252 265 324
rect 207 -264 265 -252
rect 325 324 383 336
rect 325 -252 337 324
rect 371 -252 383 324
rect 325 -264 383 -252
rect 443 324 501 336
rect 443 -252 455 324
rect 489 -252 501 324
rect 443 -264 501 -252
rect 561 324 619 336
rect 561 -252 573 324
rect 607 -252 619 324
rect 561 -264 619 -252
rect 679 324 737 336
rect 679 -252 691 324
rect 725 -252 737 324
rect 679 -264 737 -252
rect 797 324 855 336
rect 797 -252 809 324
rect 843 -252 855 324
rect 797 -264 855 -252
rect 915 324 973 336
rect 915 -252 927 324
rect 961 -252 973 324
rect 915 -264 973 -252
rect 1033 324 1091 336
rect 1033 -252 1045 324
rect 1079 -252 1091 324
rect 1033 -264 1091 -252
rect 1151 324 1209 336
rect 1151 -252 1163 324
rect 1197 -252 1209 324
rect 1151 -264 1209 -252
rect 1269 324 1327 336
rect 1269 -252 1281 324
rect 1315 -252 1327 324
rect 1269 -264 1327 -252
rect 1387 324 1445 336
rect 1387 -252 1399 324
rect 1433 -252 1445 324
rect 1387 -264 1445 -252
rect 1505 324 1563 336
rect 1505 -252 1517 324
rect 1551 -252 1563 324
rect 1505 -264 1563 -252
rect 1623 324 1681 336
rect 1623 -252 1635 324
rect 1669 -252 1681 324
rect 1623 -264 1681 -252
rect 1741 324 1799 336
rect 1741 -252 1753 324
rect 1787 -252 1799 324
rect 1741 -264 1799 -252
rect 1859 324 1917 336
rect 1859 -252 1871 324
rect 1905 -252 1917 324
rect 1859 -264 1917 -252
rect 1977 324 2035 336
rect 1977 -252 1989 324
rect 2023 -252 2035 324
rect 1977 -264 2035 -252
rect 2095 324 2153 336
rect 2095 -252 2107 324
rect 2141 -252 2153 324
rect 2095 -264 2153 -252
rect 2213 324 2271 336
rect 2213 -252 2225 324
rect 2259 -252 2271 324
rect 2213 -264 2271 -252
rect 2331 324 2389 336
rect 2331 -252 2343 324
rect 2377 -252 2389 324
rect 2331 -264 2389 -252
rect 2449 324 2507 336
rect 2449 -252 2461 324
rect 2495 -252 2507 324
rect 2449 -264 2507 -252
rect 2567 324 2625 336
rect 2567 -252 2579 324
rect 2613 -252 2625 324
rect 2567 -264 2625 -252
rect 2685 324 2743 336
rect 2685 -252 2697 324
rect 2731 -252 2743 324
rect 2685 -264 2743 -252
rect 2803 324 2861 336
rect 2803 -252 2815 324
rect 2849 -252 2861 324
rect 2803 -264 2861 -252
rect 2921 324 2979 336
rect 2921 -252 2933 324
rect 2967 -252 2979 324
rect 2921 -264 2979 -252
<< pdiffc >>
rect -2967 -252 -2933 324
rect -2849 -252 -2815 324
rect -2731 -252 -2697 324
rect -2613 -252 -2579 324
rect -2495 -252 -2461 324
rect -2377 -252 -2343 324
rect -2259 -252 -2225 324
rect -2141 -252 -2107 324
rect -2023 -252 -1989 324
rect -1905 -252 -1871 324
rect -1787 -252 -1753 324
rect -1669 -252 -1635 324
rect -1551 -252 -1517 324
rect -1433 -252 -1399 324
rect -1315 -252 -1281 324
rect -1197 -252 -1163 324
rect -1079 -252 -1045 324
rect -961 -252 -927 324
rect -843 -252 -809 324
rect -725 -252 -691 324
rect -607 -252 -573 324
rect -489 -252 -455 324
rect -371 -252 -337 324
rect -253 -252 -219 324
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
rect 219 -252 253 324
rect 337 -252 371 324
rect 455 -252 489 324
rect 573 -252 607 324
rect 691 -252 725 324
rect 809 -252 843 324
rect 927 -252 961 324
rect 1045 -252 1079 324
rect 1163 -252 1197 324
rect 1281 -252 1315 324
rect 1399 -252 1433 324
rect 1517 -252 1551 324
rect 1635 -252 1669 324
rect 1753 -252 1787 324
rect 1871 -252 1905 324
rect 1989 -252 2023 324
rect 2107 -252 2141 324
rect 2225 -252 2259 324
rect 2343 -252 2377 324
rect 2461 -252 2495 324
rect 2579 -252 2613 324
rect 2697 -252 2731 324
rect 2815 -252 2849 324
rect 2933 -252 2967 324
<< nsubdiff >>
rect -3081 414 -2985 448
rect 2985 414 3081 448
rect -3081 351 -3047 414
rect 3047 351 3081 414
rect -3081 -414 -3047 -351
rect 3047 -414 3081 -351
rect -3081 -448 -2985 -414
rect 2985 -448 3081 -414
<< nsubdiffcont >>
rect -2985 414 2985 448
rect -3081 -351 -3047 351
rect 3047 -351 3081 351
rect -2985 -448 2985 -414
<< poly >>
rect -2921 336 -2861 362
rect -2803 336 -2743 362
rect -2685 336 -2625 362
rect -2567 336 -2507 362
rect -2449 336 -2389 362
rect -2331 336 -2271 362
rect -2213 336 -2153 362
rect -2095 336 -2035 362
rect -1977 336 -1917 362
rect -1859 336 -1799 362
rect -1741 336 -1681 362
rect -1623 336 -1563 362
rect -1505 336 -1445 362
rect -1387 336 -1327 362
rect -1269 336 -1209 362
rect -1151 336 -1091 362
rect -1033 336 -973 362
rect -915 336 -855 362
rect -797 336 -737 362
rect -679 336 -619 362
rect -561 336 -501 362
rect -443 336 -383 362
rect -325 336 -265 362
rect -207 336 -147 362
rect -89 336 -29 362
rect 29 336 89 362
rect 147 336 207 362
rect 265 336 325 362
rect 383 336 443 362
rect 501 336 561 362
rect 619 336 679 362
rect 737 336 797 362
rect 855 336 915 362
rect 973 336 1033 362
rect 1091 336 1151 362
rect 1209 336 1269 362
rect 1327 336 1387 362
rect 1445 336 1505 362
rect 1563 336 1623 362
rect 1681 336 1741 362
rect 1799 336 1859 362
rect 1917 336 1977 362
rect 2035 336 2095 362
rect 2153 336 2213 362
rect 2271 336 2331 362
rect 2389 336 2449 362
rect 2507 336 2567 362
rect 2625 336 2685 362
rect 2743 336 2803 362
rect 2861 336 2921 362
rect -2921 -295 -2861 -264
rect -2803 -295 -2743 -264
rect -2685 -295 -2625 -264
rect -2567 -295 -2507 -264
rect -2449 -295 -2389 -264
rect -2331 -295 -2271 -264
rect -2213 -295 -2153 -264
rect -2095 -295 -2035 -264
rect -1977 -295 -1917 -264
rect -1859 -295 -1799 -264
rect -1741 -295 -1681 -264
rect -1623 -295 -1563 -264
rect -1505 -295 -1445 -264
rect -1387 -295 -1327 -264
rect -1269 -295 -1209 -264
rect -1151 -295 -1091 -264
rect -1033 -295 -973 -264
rect -915 -295 -855 -264
rect -797 -295 -737 -264
rect -679 -295 -619 -264
rect -561 -295 -501 -264
rect -443 -295 -383 -264
rect -325 -295 -265 -264
rect -207 -295 -147 -264
rect -89 -295 -29 -264
rect 29 -295 89 -264
rect 147 -295 207 -264
rect 265 -295 325 -264
rect 383 -295 443 -264
rect 501 -295 561 -264
rect 619 -295 679 -264
rect 737 -295 797 -264
rect 855 -295 915 -264
rect 973 -295 1033 -264
rect 1091 -295 1151 -264
rect 1209 -295 1269 -264
rect 1327 -295 1387 -264
rect 1445 -295 1505 -264
rect 1563 -295 1623 -264
rect 1681 -295 1741 -264
rect 1799 -295 1859 -264
rect 1917 -295 1977 -264
rect 2035 -295 2095 -264
rect 2153 -295 2213 -264
rect 2271 -295 2331 -264
rect 2389 -295 2449 -264
rect 2507 -295 2567 -264
rect 2625 -295 2685 -264
rect 2743 -295 2803 -264
rect 2861 -295 2921 -264
rect -2924 -311 -2858 -295
rect -2924 -345 -2908 -311
rect -2874 -345 -2858 -311
rect -2924 -361 -2858 -345
rect -2806 -311 -2740 -295
rect -2806 -345 -2790 -311
rect -2756 -345 -2740 -311
rect -2806 -361 -2740 -345
rect -2688 -311 -2622 -295
rect -2688 -345 -2672 -311
rect -2638 -345 -2622 -311
rect -2688 -361 -2622 -345
rect -2570 -311 -2504 -295
rect -2570 -345 -2554 -311
rect -2520 -345 -2504 -311
rect -2570 -361 -2504 -345
rect -2452 -311 -2386 -295
rect -2452 -345 -2436 -311
rect -2402 -345 -2386 -311
rect -2452 -361 -2386 -345
rect -2334 -311 -2268 -295
rect -2334 -345 -2318 -311
rect -2284 -345 -2268 -311
rect -2334 -361 -2268 -345
rect -2216 -311 -2150 -295
rect -2216 -345 -2200 -311
rect -2166 -345 -2150 -311
rect -2216 -361 -2150 -345
rect -2098 -311 -2032 -295
rect -2098 -345 -2082 -311
rect -2048 -345 -2032 -311
rect -2098 -361 -2032 -345
rect -1980 -311 -1914 -295
rect -1980 -345 -1964 -311
rect -1930 -345 -1914 -311
rect -1980 -361 -1914 -345
rect -1862 -311 -1796 -295
rect -1862 -345 -1846 -311
rect -1812 -345 -1796 -311
rect -1862 -361 -1796 -345
rect -1744 -311 -1678 -295
rect -1744 -345 -1728 -311
rect -1694 -345 -1678 -311
rect -1744 -361 -1678 -345
rect -1626 -311 -1560 -295
rect -1626 -345 -1610 -311
rect -1576 -345 -1560 -311
rect -1626 -361 -1560 -345
rect -1508 -311 -1442 -295
rect -1508 -345 -1492 -311
rect -1458 -345 -1442 -311
rect -1508 -361 -1442 -345
rect -1390 -311 -1324 -295
rect -1390 -345 -1374 -311
rect -1340 -345 -1324 -311
rect -1390 -361 -1324 -345
rect -1272 -311 -1206 -295
rect -1272 -345 -1256 -311
rect -1222 -345 -1206 -311
rect -1272 -361 -1206 -345
rect -1154 -311 -1088 -295
rect -1154 -345 -1138 -311
rect -1104 -345 -1088 -311
rect -1154 -361 -1088 -345
rect -1036 -311 -970 -295
rect -1036 -345 -1020 -311
rect -986 -345 -970 -311
rect -1036 -361 -970 -345
rect -918 -311 -852 -295
rect -918 -345 -902 -311
rect -868 -345 -852 -311
rect -918 -361 -852 -345
rect -800 -311 -734 -295
rect -800 -345 -784 -311
rect -750 -345 -734 -311
rect -800 -361 -734 -345
rect -682 -311 -616 -295
rect -682 -345 -666 -311
rect -632 -345 -616 -311
rect -682 -361 -616 -345
rect -564 -311 -498 -295
rect -564 -345 -548 -311
rect -514 -345 -498 -311
rect -564 -361 -498 -345
rect -446 -311 -380 -295
rect -446 -345 -430 -311
rect -396 -345 -380 -311
rect -446 -361 -380 -345
rect -328 -311 -262 -295
rect -328 -345 -312 -311
rect -278 -345 -262 -311
rect -328 -361 -262 -345
rect -210 -311 -144 -295
rect -210 -345 -194 -311
rect -160 -345 -144 -311
rect -210 -361 -144 -345
rect -92 -311 -26 -295
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect -92 -361 -26 -345
rect 26 -311 92 -295
rect 26 -345 42 -311
rect 76 -345 92 -311
rect 26 -361 92 -345
rect 144 -311 210 -295
rect 144 -345 160 -311
rect 194 -345 210 -311
rect 144 -361 210 -345
rect 262 -311 328 -295
rect 262 -345 278 -311
rect 312 -345 328 -311
rect 262 -361 328 -345
rect 380 -311 446 -295
rect 380 -345 396 -311
rect 430 -345 446 -311
rect 380 -361 446 -345
rect 498 -311 564 -295
rect 498 -345 514 -311
rect 548 -345 564 -311
rect 498 -361 564 -345
rect 616 -311 682 -295
rect 616 -345 632 -311
rect 666 -345 682 -311
rect 616 -361 682 -345
rect 734 -311 800 -295
rect 734 -345 750 -311
rect 784 -345 800 -311
rect 734 -361 800 -345
rect 852 -311 918 -295
rect 852 -345 868 -311
rect 902 -345 918 -311
rect 852 -361 918 -345
rect 970 -311 1036 -295
rect 970 -345 986 -311
rect 1020 -345 1036 -311
rect 970 -361 1036 -345
rect 1088 -311 1154 -295
rect 1088 -345 1104 -311
rect 1138 -345 1154 -311
rect 1088 -361 1154 -345
rect 1206 -311 1272 -295
rect 1206 -345 1222 -311
rect 1256 -345 1272 -311
rect 1206 -361 1272 -345
rect 1324 -311 1390 -295
rect 1324 -345 1340 -311
rect 1374 -345 1390 -311
rect 1324 -361 1390 -345
rect 1442 -311 1508 -295
rect 1442 -345 1458 -311
rect 1492 -345 1508 -311
rect 1442 -361 1508 -345
rect 1560 -311 1626 -295
rect 1560 -345 1576 -311
rect 1610 -345 1626 -311
rect 1560 -361 1626 -345
rect 1678 -311 1744 -295
rect 1678 -345 1694 -311
rect 1728 -345 1744 -311
rect 1678 -361 1744 -345
rect 1796 -311 1862 -295
rect 1796 -345 1812 -311
rect 1846 -345 1862 -311
rect 1796 -361 1862 -345
rect 1914 -311 1980 -295
rect 1914 -345 1930 -311
rect 1964 -345 1980 -311
rect 1914 -361 1980 -345
rect 2032 -311 2098 -295
rect 2032 -345 2048 -311
rect 2082 -345 2098 -311
rect 2032 -361 2098 -345
rect 2150 -311 2216 -295
rect 2150 -345 2166 -311
rect 2200 -345 2216 -311
rect 2150 -361 2216 -345
rect 2268 -311 2334 -295
rect 2268 -345 2284 -311
rect 2318 -345 2334 -311
rect 2268 -361 2334 -345
rect 2386 -311 2452 -295
rect 2386 -345 2402 -311
rect 2436 -345 2452 -311
rect 2386 -361 2452 -345
rect 2504 -311 2570 -295
rect 2504 -345 2520 -311
rect 2554 -345 2570 -311
rect 2504 -361 2570 -345
rect 2622 -311 2688 -295
rect 2622 -345 2638 -311
rect 2672 -345 2688 -311
rect 2622 -361 2688 -345
rect 2740 -311 2806 -295
rect 2740 -345 2756 -311
rect 2790 -345 2806 -311
rect 2740 -361 2806 -345
rect 2858 -311 2924 -295
rect 2858 -345 2874 -311
rect 2908 -345 2924 -311
rect 2858 -361 2924 -345
<< polycont >>
rect -2908 -345 -2874 -311
rect -2790 -345 -2756 -311
rect -2672 -345 -2638 -311
rect -2554 -345 -2520 -311
rect -2436 -345 -2402 -311
rect -2318 -345 -2284 -311
rect -2200 -345 -2166 -311
rect -2082 -345 -2048 -311
rect -1964 -345 -1930 -311
rect -1846 -345 -1812 -311
rect -1728 -345 -1694 -311
rect -1610 -345 -1576 -311
rect -1492 -345 -1458 -311
rect -1374 -345 -1340 -311
rect -1256 -345 -1222 -311
rect -1138 -345 -1104 -311
rect -1020 -345 -986 -311
rect -902 -345 -868 -311
rect -784 -345 -750 -311
rect -666 -345 -632 -311
rect -548 -345 -514 -311
rect -430 -345 -396 -311
rect -312 -345 -278 -311
rect -194 -345 -160 -311
rect -76 -345 -42 -311
rect 42 -345 76 -311
rect 160 -345 194 -311
rect 278 -345 312 -311
rect 396 -345 430 -311
rect 514 -345 548 -311
rect 632 -345 666 -311
rect 750 -345 784 -311
rect 868 -345 902 -311
rect 986 -345 1020 -311
rect 1104 -345 1138 -311
rect 1222 -345 1256 -311
rect 1340 -345 1374 -311
rect 1458 -345 1492 -311
rect 1576 -345 1610 -311
rect 1694 -345 1728 -311
rect 1812 -345 1846 -311
rect 1930 -345 1964 -311
rect 2048 -345 2082 -311
rect 2166 -345 2200 -311
rect 2284 -345 2318 -311
rect 2402 -345 2436 -311
rect 2520 -345 2554 -311
rect 2638 -345 2672 -311
rect 2756 -345 2790 -311
rect 2874 -345 2908 -311
<< locali >>
rect -3081 414 -2985 448
rect 2985 414 3081 448
rect -3081 351 -3047 414
rect 3047 351 3081 414
rect -2967 324 -2933 340
rect -2967 -268 -2933 -252
rect -2849 324 -2815 340
rect -2849 -268 -2815 -252
rect -2731 324 -2697 340
rect -2731 -268 -2697 -252
rect -2613 324 -2579 340
rect -2613 -268 -2579 -252
rect -2495 324 -2461 340
rect -2495 -268 -2461 -252
rect -2377 324 -2343 340
rect -2377 -268 -2343 -252
rect -2259 324 -2225 340
rect -2259 -268 -2225 -252
rect -2141 324 -2107 340
rect -2141 -268 -2107 -252
rect -2023 324 -1989 340
rect -2023 -268 -1989 -252
rect -1905 324 -1871 340
rect -1905 -268 -1871 -252
rect -1787 324 -1753 340
rect -1787 -268 -1753 -252
rect -1669 324 -1635 340
rect -1669 -268 -1635 -252
rect -1551 324 -1517 340
rect -1551 -268 -1517 -252
rect -1433 324 -1399 340
rect -1433 -268 -1399 -252
rect -1315 324 -1281 340
rect -1315 -268 -1281 -252
rect -1197 324 -1163 340
rect -1197 -268 -1163 -252
rect -1079 324 -1045 340
rect -1079 -268 -1045 -252
rect -961 324 -927 340
rect -961 -268 -927 -252
rect -843 324 -809 340
rect -843 -268 -809 -252
rect -725 324 -691 340
rect -725 -268 -691 -252
rect -607 324 -573 340
rect -607 -268 -573 -252
rect -489 324 -455 340
rect -489 -268 -455 -252
rect -371 324 -337 340
rect -371 -268 -337 -252
rect -253 324 -219 340
rect -253 -268 -219 -252
rect -135 324 -101 340
rect -135 -268 -101 -252
rect -17 324 17 340
rect -17 -268 17 -252
rect 101 324 135 340
rect 101 -268 135 -252
rect 219 324 253 340
rect 219 -268 253 -252
rect 337 324 371 340
rect 337 -268 371 -252
rect 455 324 489 340
rect 455 -268 489 -252
rect 573 324 607 340
rect 573 -268 607 -252
rect 691 324 725 340
rect 691 -268 725 -252
rect 809 324 843 340
rect 809 -268 843 -252
rect 927 324 961 340
rect 927 -268 961 -252
rect 1045 324 1079 340
rect 1045 -268 1079 -252
rect 1163 324 1197 340
rect 1163 -268 1197 -252
rect 1281 324 1315 340
rect 1281 -268 1315 -252
rect 1399 324 1433 340
rect 1399 -268 1433 -252
rect 1517 324 1551 340
rect 1517 -268 1551 -252
rect 1635 324 1669 340
rect 1635 -268 1669 -252
rect 1753 324 1787 340
rect 1753 -268 1787 -252
rect 1871 324 1905 340
rect 1871 -268 1905 -252
rect 1989 324 2023 340
rect 1989 -268 2023 -252
rect 2107 324 2141 340
rect 2107 -268 2141 -252
rect 2225 324 2259 340
rect 2225 -268 2259 -252
rect 2343 324 2377 340
rect 2343 -268 2377 -252
rect 2461 324 2495 340
rect 2461 -268 2495 -252
rect 2579 324 2613 340
rect 2579 -268 2613 -252
rect 2697 324 2731 340
rect 2697 -268 2731 -252
rect 2815 324 2849 340
rect 2815 -268 2849 -252
rect 2933 324 2967 340
rect 2933 -268 2967 -252
rect -2924 -345 -2908 -311
rect -2874 -345 -2858 -311
rect -2806 -345 -2790 -311
rect -2756 -345 -2740 -311
rect -2688 -345 -2672 -311
rect -2638 -345 -2622 -311
rect -2570 -345 -2554 -311
rect -2520 -345 -2504 -311
rect -2452 -345 -2436 -311
rect -2402 -345 -2386 -311
rect -2334 -345 -2318 -311
rect -2284 -345 -2268 -311
rect -2216 -345 -2200 -311
rect -2166 -345 -2150 -311
rect -2098 -345 -2082 -311
rect -2048 -345 -2032 -311
rect -1980 -345 -1964 -311
rect -1930 -345 -1914 -311
rect -1862 -345 -1846 -311
rect -1812 -345 -1796 -311
rect -1744 -345 -1728 -311
rect -1694 -345 -1678 -311
rect -1626 -345 -1610 -311
rect -1576 -345 -1560 -311
rect -1508 -345 -1492 -311
rect -1458 -345 -1442 -311
rect -1390 -345 -1374 -311
rect -1340 -345 -1324 -311
rect -1272 -345 -1256 -311
rect -1222 -345 -1206 -311
rect -1154 -345 -1138 -311
rect -1104 -345 -1088 -311
rect -1036 -345 -1020 -311
rect -986 -345 -970 -311
rect -918 -345 -902 -311
rect -868 -345 -852 -311
rect -800 -345 -784 -311
rect -750 -345 -734 -311
rect -682 -345 -666 -311
rect -632 -345 -616 -311
rect -564 -345 -548 -311
rect -514 -345 -498 -311
rect -446 -345 -430 -311
rect -396 -345 -380 -311
rect -328 -345 -312 -311
rect -278 -345 -262 -311
rect -210 -345 -194 -311
rect -160 -345 -144 -311
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect 26 -345 42 -311
rect 76 -345 92 -311
rect 144 -345 160 -311
rect 194 -345 210 -311
rect 262 -345 278 -311
rect 312 -345 328 -311
rect 380 -345 396 -311
rect 430 -345 446 -311
rect 498 -345 514 -311
rect 548 -345 564 -311
rect 616 -345 632 -311
rect 666 -345 682 -311
rect 734 -345 750 -311
rect 784 -345 800 -311
rect 852 -345 868 -311
rect 902 -345 918 -311
rect 970 -345 986 -311
rect 1020 -345 1036 -311
rect 1088 -345 1104 -311
rect 1138 -345 1154 -311
rect 1206 -345 1222 -311
rect 1256 -345 1272 -311
rect 1324 -345 1340 -311
rect 1374 -345 1390 -311
rect 1442 -345 1458 -311
rect 1492 -345 1508 -311
rect 1560 -345 1576 -311
rect 1610 -345 1626 -311
rect 1678 -345 1694 -311
rect 1728 -345 1744 -311
rect 1796 -345 1812 -311
rect 1846 -345 1862 -311
rect 1914 -345 1930 -311
rect 1964 -345 1980 -311
rect 2032 -345 2048 -311
rect 2082 -345 2098 -311
rect 2150 -345 2166 -311
rect 2200 -345 2216 -311
rect 2268 -345 2284 -311
rect 2318 -345 2334 -311
rect 2386 -345 2402 -311
rect 2436 -345 2452 -311
rect 2504 -345 2520 -311
rect 2554 -345 2570 -311
rect 2622 -345 2638 -311
rect 2672 -345 2688 -311
rect 2740 -345 2756 -311
rect 2790 -345 2806 -311
rect 2858 -345 2874 -311
rect 2908 -345 2924 -311
rect -3081 -414 -3047 -351
rect 3047 -414 3081 -351
rect -3081 -448 -2985 -414
rect 2985 -448 3081 -414
<< viali >>
rect -2967 -252 -2933 324
rect -2849 -252 -2815 324
rect -2731 -252 -2697 324
rect -2613 -252 -2579 324
rect -2495 -252 -2461 324
rect -2377 -252 -2343 324
rect -2259 -252 -2225 324
rect -2141 -252 -2107 324
rect -2023 -252 -1989 324
rect -1905 -252 -1871 324
rect -1787 -252 -1753 324
rect -1669 -252 -1635 324
rect -1551 -252 -1517 324
rect -1433 -252 -1399 324
rect -1315 -252 -1281 324
rect -1197 -252 -1163 324
rect -1079 -252 -1045 324
rect -961 -252 -927 324
rect -843 -252 -809 324
rect -725 -252 -691 324
rect -607 -252 -573 324
rect -489 -252 -455 324
rect -371 -252 -337 324
rect -253 -252 -219 324
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
rect 219 -252 253 324
rect 337 -252 371 324
rect 455 -252 489 324
rect 573 -252 607 324
rect 691 -252 725 324
rect 809 -252 843 324
rect 927 -252 961 324
rect 1045 -252 1079 324
rect 1163 -252 1197 324
rect 1281 -252 1315 324
rect 1399 -252 1433 324
rect 1517 -252 1551 324
rect 1635 -252 1669 324
rect 1753 -252 1787 324
rect 1871 -252 1905 324
rect 1989 -252 2023 324
rect 2107 -252 2141 324
rect 2225 -252 2259 324
rect 2343 -252 2377 324
rect 2461 -252 2495 324
rect 2579 -252 2613 324
rect 2697 -252 2731 324
rect 2815 -252 2849 324
rect 2933 -252 2967 324
rect -2908 -345 -2874 -311
rect -2790 -345 -2756 -311
rect -2672 -345 -2638 -311
rect -2554 -345 -2520 -311
rect -2436 -345 -2402 -311
rect -2318 -345 -2284 -311
rect -2200 -345 -2166 -311
rect -2082 -345 -2048 -311
rect -1964 -345 -1930 -311
rect -1846 -345 -1812 -311
rect -1728 -345 -1694 -311
rect -1610 -345 -1576 -311
rect -1492 -345 -1458 -311
rect -1374 -345 -1340 -311
rect -1256 -345 -1222 -311
rect -1138 -345 -1104 -311
rect -1020 -345 -986 -311
rect -902 -345 -868 -311
rect -784 -345 -750 -311
rect -666 -345 -632 -311
rect -548 -345 -514 -311
rect -430 -345 -396 -311
rect -312 -345 -278 -311
rect -194 -345 -160 -311
rect -76 -345 -42 -311
rect 42 -345 76 -311
rect 160 -345 194 -311
rect 278 -345 312 -311
rect 396 -345 430 -311
rect 514 -345 548 -311
rect 632 -345 666 -311
rect 750 -345 784 -311
rect 868 -345 902 -311
rect 986 -345 1020 -311
rect 1104 -345 1138 -311
rect 1222 -345 1256 -311
rect 1340 -345 1374 -311
rect 1458 -345 1492 -311
rect 1576 -345 1610 -311
rect 1694 -345 1728 -311
rect 1812 -345 1846 -311
rect 1930 -345 1964 -311
rect 2048 -345 2082 -311
rect 2166 -345 2200 -311
rect 2284 -345 2318 -311
rect 2402 -345 2436 -311
rect 2520 -345 2554 -311
rect 2638 -345 2672 -311
rect 2756 -345 2790 -311
rect 2874 -345 2908 -311
<< metal1 >>
rect -2973 324 -2927 336
rect -2973 -252 -2967 324
rect -2933 -252 -2927 324
rect -2973 -264 -2927 -252
rect -2855 324 -2809 336
rect -2855 -252 -2849 324
rect -2815 -252 -2809 324
rect -2855 -264 -2809 -252
rect -2737 324 -2691 336
rect -2737 -252 -2731 324
rect -2697 -252 -2691 324
rect -2737 -264 -2691 -252
rect -2619 324 -2573 336
rect -2619 -252 -2613 324
rect -2579 -252 -2573 324
rect -2619 -264 -2573 -252
rect -2501 324 -2455 336
rect -2501 -252 -2495 324
rect -2461 -252 -2455 324
rect -2501 -264 -2455 -252
rect -2383 324 -2337 336
rect -2383 -252 -2377 324
rect -2343 -252 -2337 324
rect -2383 -264 -2337 -252
rect -2265 324 -2219 336
rect -2265 -252 -2259 324
rect -2225 -252 -2219 324
rect -2265 -264 -2219 -252
rect -2147 324 -2101 336
rect -2147 -252 -2141 324
rect -2107 -252 -2101 324
rect -2147 -264 -2101 -252
rect -2029 324 -1983 336
rect -2029 -252 -2023 324
rect -1989 -252 -1983 324
rect -2029 -264 -1983 -252
rect -1911 324 -1865 336
rect -1911 -252 -1905 324
rect -1871 -252 -1865 324
rect -1911 -264 -1865 -252
rect -1793 324 -1747 336
rect -1793 -252 -1787 324
rect -1753 -252 -1747 324
rect -1793 -264 -1747 -252
rect -1675 324 -1629 336
rect -1675 -252 -1669 324
rect -1635 -252 -1629 324
rect -1675 -264 -1629 -252
rect -1557 324 -1511 336
rect -1557 -252 -1551 324
rect -1517 -252 -1511 324
rect -1557 -264 -1511 -252
rect -1439 324 -1393 336
rect -1439 -252 -1433 324
rect -1399 -252 -1393 324
rect -1439 -264 -1393 -252
rect -1321 324 -1275 336
rect -1321 -252 -1315 324
rect -1281 -252 -1275 324
rect -1321 -264 -1275 -252
rect -1203 324 -1157 336
rect -1203 -252 -1197 324
rect -1163 -252 -1157 324
rect -1203 -264 -1157 -252
rect -1085 324 -1039 336
rect -1085 -252 -1079 324
rect -1045 -252 -1039 324
rect -1085 -264 -1039 -252
rect -967 324 -921 336
rect -967 -252 -961 324
rect -927 -252 -921 324
rect -967 -264 -921 -252
rect -849 324 -803 336
rect -849 -252 -843 324
rect -809 -252 -803 324
rect -849 -264 -803 -252
rect -731 324 -685 336
rect -731 -252 -725 324
rect -691 -252 -685 324
rect -731 -264 -685 -252
rect -613 324 -567 336
rect -613 -252 -607 324
rect -573 -252 -567 324
rect -613 -264 -567 -252
rect -495 324 -449 336
rect -495 -252 -489 324
rect -455 -252 -449 324
rect -495 -264 -449 -252
rect -377 324 -331 336
rect -377 -252 -371 324
rect -337 -252 -331 324
rect -377 -264 -331 -252
rect -259 324 -213 336
rect -259 -252 -253 324
rect -219 -252 -213 324
rect -259 -264 -213 -252
rect -141 324 -95 336
rect -141 -252 -135 324
rect -101 -252 -95 324
rect -141 -264 -95 -252
rect -23 324 23 336
rect -23 -252 -17 324
rect 17 -252 23 324
rect -23 -264 23 -252
rect 95 324 141 336
rect 95 -252 101 324
rect 135 -252 141 324
rect 95 -264 141 -252
rect 213 324 259 336
rect 213 -252 219 324
rect 253 -252 259 324
rect 213 -264 259 -252
rect 331 324 377 336
rect 331 -252 337 324
rect 371 -252 377 324
rect 331 -264 377 -252
rect 449 324 495 336
rect 449 -252 455 324
rect 489 -252 495 324
rect 449 -264 495 -252
rect 567 324 613 336
rect 567 -252 573 324
rect 607 -252 613 324
rect 567 -264 613 -252
rect 685 324 731 336
rect 685 -252 691 324
rect 725 -252 731 324
rect 685 -264 731 -252
rect 803 324 849 336
rect 803 -252 809 324
rect 843 -252 849 324
rect 803 -264 849 -252
rect 921 324 967 336
rect 921 -252 927 324
rect 961 -252 967 324
rect 921 -264 967 -252
rect 1039 324 1085 336
rect 1039 -252 1045 324
rect 1079 -252 1085 324
rect 1039 -264 1085 -252
rect 1157 324 1203 336
rect 1157 -252 1163 324
rect 1197 -252 1203 324
rect 1157 -264 1203 -252
rect 1275 324 1321 336
rect 1275 -252 1281 324
rect 1315 -252 1321 324
rect 1275 -264 1321 -252
rect 1393 324 1439 336
rect 1393 -252 1399 324
rect 1433 -252 1439 324
rect 1393 -264 1439 -252
rect 1511 324 1557 336
rect 1511 -252 1517 324
rect 1551 -252 1557 324
rect 1511 -264 1557 -252
rect 1629 324 1675 336
rect 1629 -252 1635 324
rect 1669 -252 1675 324
rect 1629 -264 1675 -252
rect 1747 324 1793 336
rect 1747 -252 1753 324
rect 1787 -252 1793 324
rect 1747 -264 1793 -252
rect 1865 324 1911 336
rect 1865 -252 1871 324
rect 1905 -252 1911 324
rect 1865 -264 1911 -252
rect 1983 324 2029 336
rect 1983 -252 1989 324
rect 2023 -252 2029 324
rect 1983 -264 2029 -252
rect 2101 324 2147 336
rect 2101 -252 2107 324
rect 2141 -252 2147 324
rect 2101 -264 2147 -252
rect 2219 324 2265 336
rect 2219 -252 2225 324
rect 2259 -252 2265 324
rect 2219 -264 2265 -252
rect 2337 324 2383 336
rect 2337 -252 2343 324
rect 2377 -252 2383 324
rect 2337 -264 2383 -252
rect 2455 324 2501 336
rect 2455 -252 2461 324
rect 2495 -252 2501 324
rect 2455 -264 2501 -252
rect 2573 324 2619 336
rect 2573 -252 2579 324
rect 2613 -252 2619 324
rect 2573 -264 2619 -252
rect 2691 324 2737 336
rect 2691 -252 2697 324
rect 2731 -252 2737 324
rect 2691 -264 2737 -252
rect 2809 324 2855 336
rect 2809 -252 2815 324
rect 2849 -252 2855 324
rect 2809 -264 2855 -252
rect 2927 324 2973 336
rect 2927 -252 2933 324
rect 2967 -252 2973 324
rect 2927 -264 2973 -252
rect -2920 -311 -2862 -305
rect -2920 -345 -2908 -311
rect -2874 -345 -2862 -311
rect -2920 -351 -2862 -345
rect -2802 -311 -2744 -305
rect -2802 -345 -2790 -311
rect -2756 -345 -2744 -311
rect -2802 -351 -2744 -345
rect -2684 -311 -2626 -305
rect -2684 -345 -2672 -311
rect -2638 -345 -2626 -311
rect -2684 -351 -2626 -345
rect -2566 -311 -2508 -305
rect -2566 -345 -2554 -311
rect -2520 -345 -2508 -311
rect -2566 -351 -2508 -345
rect -2448 -311 -2390 -305
rect -2448 -345 -2436 -311
rect -2402 -345 -2390 -311
rect -2448 -351 -2390 -345
rect -2330 -311 -2272 -305
rect -2330 -345 -2318 -311
rect -2284 -345 -2272 -311
rect -2330 -351 -2272 -345
rect -2212 -311 -2154 -305
rect -2212 -345 -2200 -311
rect -2166 -345 -2154 -311
rect -2212 -351 -2154 -345
rect -2094 -311 -2036 -305
rect -2094 -345 -2082 -311
rect -2048 -345 -2036 -311
rect -2094 -351 -2036 -345
rect -1976 -311 -1918 -305
rect -1976 -345 -1964 -311
rect -1930 -345 -1918 -311
rect -1976 -351 -1918 -345
rect -1858 -311 -1800 -305
rect -1858 -345 -1846 -311
rect -1812 -345 -1800 -311
rect -1858 -351 -1800 -345
rect -1740 -311 -1682 -305
rect -1740 -345 -1728 -311
rect -1694 -345 -1682 -311
rect -1740 -351 -1682 -345
rect -1622 -311 -1564 -305
rect -1622 -345 -1610 -311
rect -1576 -345 -1564 -311
rect -1622 -351 -1564 -345
rect -1504 -311 -1446 -305
rect -1504 -345 -1492 -311
rect -1458 -345 -1446 -311
rect -1504 -351 -1446 -345
rect -1386 -311 -1328 -305
rect -1386 -345 -1374 -311
rect -1340 -345 -1328 -311
rect -1386 -351 -1328 -345
rect -1268 -311 -1210 -305
rect -1268 -345 -1256 -311
rect -1222 -345 -1210 -311
rect -1268 -351 -1210 -345
rect -1150 -311 -1092 -305
rect -1150 -345 -1138 -311
rect -1104 -345 -1092 -311
rect -1150 -351 -1092 -345
rect -1032 -311 -974 -305
rect -1032 -345 -1020 -311
rect -986 -345 -974 -311
rect -1032 -351 -974 -345
rect -914 -311 -856 -305
rect -914 -345 -902 -311
rect -868 -345 -856 -311
rect -914 -351 -856 -345
rect -796 -311 -738 -305
rect -796 -345 -784 -311
rect -750 -345 -738 -311
rect -796 -351 -738 -345
rect -678 -311 -620 -305
rect -678 -345 -666 -311
rect -632 -345 -620 -311
rect -678 -351 -620 -345
rect -560 -311 -502 -305
rect -560 -345 -548 -311
rect -514 -345 -502 -311
rect -560 -351 -502 -345
rect -442 -311 -384 -305
rect -442 -345 -430 -311
rect -396 -345 -384 -311
rect -442 -351 -384 -345
rect -324 -311 -266 -305
rect -324 -345 -312 -311
rect -278 -345 -266 -311
rect -324 -351 -266 -345
rect -206 -311 -148 -305
rect -206 -345 -194 -311
rect -160 -345 -148 -311
rect -206 -351 -148 -345
rect -88 -311 -30 -305
rect -88 -345 -76 -311
rect -42 -345 -30 -311
rect -88 -351 -30 -345
rect 30 -311 88 -305
rect 30 -345 42 -311
rect 76 -345 88 -311
rect 30 -351 88 -345
rect 148 -311 206 -305
rect 148 -345 160 -311
rect 194 -345 206 -311
rect 148 -351 206 -345
rect 266 -311 324 -305
rect 266 -345 278 -311
rect 312 -345 324 -311
rect 266 -351 324 -345
rect 384 -311 442 -305
rect 384 -345 396 -311
rect 430 -345 442 -311
rect 384 -351 442 -345
rect 502 -311 560 -305
rect 502 -345 514 -311
rect 548 -345 560 -311
rect 502 -351 560 -345
rect 620 -311 678 -305
rect 620 -345 632 -311
rect 666 -345 678 -311
rect 620 -351 678 -345
rect 738 -311 796 -305
rect 738 -345 750 -311
rect 784 -345 796 -311
rect 738 -351 796 -345
rect 856 -311 914 -305
rect 856 -345 868 -311
rect 902 -345 914 -311
rect 856 -351 914 -345
rect 974 -311 1032 -305
rect 974 -345 986 -311
rect 1020 -345 1032 -311
rect 974 -351 1032 -345
rect 1092 -311 1150 -305
rect 1092 -345 1104 -311
rect 1138 -345 1150 -311
rect 1092 -351 1150 -345
rect 1210 -311 1268 -305
rect 1210 -345 1222 -311
rect 1256 -345 1268 -311
rect 1210 -351 1268 -345
rect 1328 -311 1386 -305
rect 1328 -345 1340 -311
rect 1374 -345 1386 -311
rect 1328 -351 1386 -345
rect 1446 -311 1504 -305
rect 1446 -345 1458 -311
rect 1492 -345 1504 -311
rect 1446 -351 1504 -345
rect 1564 -311 1622 -305
rect 1564 -345 1576 -311
rect 1610 -345 1622 -311
rect 1564 -351 1622 -345
rect 1682 -311 1740 -305
rect 1682 -345 1694 -311
rect 1728 -345 1740 -311
rect 1682 -351 1740 -345
rect 1800 -311 1858 -305
rect 1800 -345 1812 -311
rect 1846 -345 1858 -311
rect 1800 -351 1858 -345
rect 1918 -311 1976 -305
rect 1918 -345 1930 -311
rect 1964 -345 1976 -311
rect 1918 -351 1976 -345
rect 2036 -311 2094 -305
rect 2036 -345 2048 -311
rect 2082 -345 2094 -311
rect 2036 -351 2094 -345
rect 2154 -311 2212 -305
rect 2154 -345 2166 -311
rect 2200 -345 2212 -311
rect 2154 -351 2212 -345
rect 2272 -311 2330 -305
rect 2272 -345 2284 -311
rect 2318 -345 2330 -311
rect 2272 -351 2330 -345
rect 2390 -311 2448 -305
rect 2390 -345 2402 -311
rect 2436 -345 2448 -311
rect 2390 -351 2448 -345
rect 2508 -311 2566 -305
rect 2508 -345 2520 -311
rect 2554 -345 2566 -311
rect 2508 -351 2566 -345
rect 2626 -311 2684 -305
rect 2626 -345 2638 -311
rect 2672 -345 2684 -311
rect 2626 -351 2684 -345
rect 2744 -311 2802 -305
rect 2744 -345 2756 -311
rect 2790 -345 2802 -311
rect 2744 -351 2802 -345
rect 2862 -311 2920 -305
rect 2862 -345 2874 -311
rect 2908 -345 2920 -311
rect 2862 -351 2920 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -431 3064 431
string parameters w 3 l 0.3 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
