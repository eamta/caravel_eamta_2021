magic
tech sky130A
magscale 1 2
timestamp 1623248045
<< pwell >>
rect -1127 -1110 1127 1110
<< nmoslvt >>
rect -927 -900 -897 900
rect -831 -900 -801 900
rect -735 -900 -705 900
rect -639 -900 -609 900
rect -543 -900 -513 900
rect -447 -900 -417 900
rect -351 -900 -321 900
rect -255 -900 -225 900
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
rect 225 -900 255 900
rect 321 -900 351 900
rect 417 -900 447 900
rect 513 -900 543 900
rect 609 -900 639 900
rect 705 -900 735 900
rect 801 -900 831 900
rect 897 -900 927 900
<< ndiff >>
rect -989 888 -927 900
rect -989 -888 -977 888
rect -943 -888 -927 888
rect -989 -900 -927 -888
rect -897 888 -831 900
rect -897 -888 -881 888
rect -847 -888 -831 888
rect -897 -900 -831 -888
rect -801 888 -735 900
rect -801 -888 -785 888
rect -751 -888 -735 888
rect -801 -900 -735 -888
rect -705 888 -639 900
rect -705 -888 -689 888
rect -655 -888 -639 888
rect -705 -900 -639 -888
rect -609 888 -543 900
rect -609 -888 -593 888
rect -559 -888 -543 888
rect -609 -900 -543 -888
rect -513 888 -447 900
rect -513 -888 -497 888
rect -463 -888 -447 888
rect -513 -900 -447 -888
rect -417 888 -351 900
rect -417 -888 -401 888
rect -367 -888 -351 888
rect -417 -900 -351 -888
rect -321 888 -255 900
rect -321 -888 -305 888
rect -271 -888 -255 888
rect -321 -900 -255 -888
rect -225 888 -159 900
rect -225 -888 -209 888
rect -175 -888 -159 888
rect -225 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 225 900
rect 159 -888 175 888
rect 209 -888 225 888
rect 159 -900 225 -888
rect 255 888 321 900
rect 255 -888 271 888
rect 305 -888 321 888
rect 255 -900 321 -888
rect 351 888 417 900
rect 351 -888 367 888
rect 401 -888 417 888
rect 351 -900 417 -888
rect 447 888 513 900
rect 447 -888 463 888
rect 497 -888 513 888
rect 447 -900 513 -888
rect 543 888 609 900
rect 543 -888 559 888
rect 593 -888 609 888
rect 543 -900 609 -888
rect 639 888 705 900
rect 639 -888 655 888
rect 689 -888 705 888
rect 639 -900 705 -888
rect 735 888 801 900
rect 735 -888 751 888
rect 785 -888 801 888
rect 735 -900 801 -888
rect 831 888 897 900
rect 831 -888 847 888
rect 881 -888 897 888
rect 831 -900 897 -888
rect 927 888 989 900
rect 927 -888 943 888
rect 977 -888 989 888
rect 927 -900 989 -888
<< ndiffc >>
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
<< psubdiff >>
rect -1091 1041 -995 1075
rect 995 1041 1091 1075
rect -1091 978 -1057 1041
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1041
rect -1091 -1074 1091 -1040
<< psubdiffcont >>
rect -995 1041 995 1075
rect -1091 -978 -1057 978
<< poly >>
rect -927 990 945 1019
rect -927 956 -906 990
rect 924 956 945 990
rect -927 922 945 956
rect -927 900 -897 922
rect -831 900 -801 922
rect -735 900 -705 922
rect -639 900 -609 922
rect -543 900 -513 922
rect -447 900 -417 922
rect -351 900 -321 922
rect -255 900 -225 922
rect -159 900 -129 922
rect -63 900 -33 922
rect 33 900 63 922
rect 129 900 159 922
rect 225 900 255 922
rect 321 900 351 922
rect 417 900 447 922
rect 513 900 543 922
rect 609 900 639 922
rect 705 900 735 922
rect 801 900 831 922
rect 897 900 927 922
rect -927 -926 -897 -900
rect -831 -926 -801 -900
rect -735 -926 -705 -900
rect -639 -926 -609 -900
rect -543 -926 -513 -900
rect -447 -926 -417 -900
rect -351 -926 -321 -900
rect -255 -926 -225 -900
rect -159 -926 -129 -900
rect -63 -926 -33 -900
rect 33 -926 63 -900
rect 129 -926 159 -900
rect 225 -926 255 -900
rect 321 -926 351 -900
rect 417 -926 447 -900
rect 513 -926 543 -900
rect 609 -926 639 -900
rect 705 -926 735 -900
rect 801 -926 831 -900
rect 897 -926 927 -900
<< polycont >>
rect -906 956 924 990
<< locali >>
rect -1091 1041 -995 1075
rect 995 1041 1091 1075
rect -1091 978 -1057 1041
rect -922 1001 940 1006
rect -922 949 -906 1001
rect 924 949 940 1001
rect -922 940 940 949
rect -977 888 -943 904
rect -977 -904 -943 -888
rect -881 888 -847 904
rect -881 -904 -847 -888
rect -785 888 -751 904
rect -785 -904 -751 -888
rect -689 888 -655 904
rect -689 -904 -655 -888
rect -593 888 -559 904
rect -593 -904 -559 -888
rect -497 888 -463 904
rect -497 -904 -463 -888
rect -401 888 -367 904
rect -401 -904 -367 -888
rect -305 888 -271 904
rect -305 -904 -271 -888
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect 271 888 305 904
rect 271 -904 305 -888
rect 367 888 401 904
rect 367 -904 401 -888
rect 463 888 497 904
rect 463 -904 497 -888
rect 559 888 593 904
rect 559 -904 593 -888
rect 655 888 689 904
rect 655 -904 689 -888
rect 751 888 785 904
rect 751 -904 785 -888
rect 847 888 881 904
rect 847 -904 881 -888
rect 943 888 977 904
rect 943 -904 977 -888
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1041
rect -1091 -1074 1091 -1040
<< viali >>
rect -906 990 924 1001
rect -906 956 924 990
rect -906 949 924 956
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
<< metal1 >>
rect -918 1001 936 1007
rect -918 949 -906 1001
rect 924 949 936 1001
rect -918 943 936 949
rect -983 888 -937 900
rect -983 -888 -977 888
rect -943 -888 -937 888
rect -983 -900 -937 -888
rect -887 888 -841 900
rect -887 -888 -881 888
rect -847 -888 -841 888
rect -887 -900 -841 -888
rect -791 888 -745 900
rect -791 -888 -785 888
rect -751 -888 -745 888
rect -791 -900 -745 -888
rect -695 888 -649 900
rect -695 -888 -689 888
rect -655 -888 -649 888
rect -695 -900 -649 -888
rect -599 888 -553 900
rect -599 -888 -593 888
rect -559 -888 -553 888
rect -599 -900 -553 -888
rect -503 888 -457 900
rect -503 -888 -497 888
rect -463 -888 -457 888
rect -503 -900 -457 -888
rect -407 888 -361 900
rect -407 -888 -401 888
rect -367 -888 -361 888
rect -407 -900 -361 -888
rect -311 888 -265 900
rect -311 -888 -305 888
rect -271 -888 -265 888
rect -311 -900 -265 -888
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect 265 888 311 900
rect 265 -888 271 888
rect 305 -888 311 888
rect 265 -900 311 -888
rect 361 888 407 900
rect 361 -888 367 888
rect 401 -888 407 888
rect 361 -900 407 -888
rect 457 888 503 900
rect 457 -888 463 888
rect 497 -888 503 888
rect 457 -900 503 -888
rect 553 888 599 900
rect 553 -888 559 888
rect 593 -888 599 888
rect 553 -900 599 -888
rect 649 888 695 900
rect 649 -888 655 888
rect 689 -888 695 888
rect 649 -900 695 -888
rect 745 888 791 900
rect 745 -888 751 888
rect 785 -888 791 888
rect 745 -900 791 -888
rect 841 888 887 900
rect 841 -888 847 888
rect 881 -888 887 888
rect 841 -900 887 -888
rect 937 888 983 900
rect 937 -888 943 888
rect 977 -888 983 888
rect 937 -900 983 -888
<< via1 >>
rect -906 949 924 1001
<< metal2 >>
rect -906 1001 924 1011
rect -906 939 924 949
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string FIXED_BBOX -1074 -1057 1074 1057
string parameters w 9 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
