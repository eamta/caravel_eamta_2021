magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 380 1729 415 1747
rect 344 1714 415 1729
rect 18 1578 45 1596
rect 157 1591 215 1597
rect 157 1580 169 1591
rect 157 1578 203 1580
rect 344 1578 414 1714
rect 526 1646 584 1652
rect 526 1612 538 1646
rect 696 1623 730 1641
rect 1118 1623 1153 1641
rect 526 1606 584 1612
rect 696 1587 766 1623
rect 1082 1608 1153 1623
rect 1433 1608 1468 1642
rect 0 1542 414 1578
rect 713 1578 845 1587
rect 494 1542 528 1576
rect 582 1542 616 1576
rect 0 1508 650 1542
rect 0 1236 414 1508
rect 613 1470 628 1485
rect 570 1440 628 1470
rect 482 1385 540 1418
rect 548 1385 556 1426
rect 570 1418 598 1440
rect 613 1425 628 1440
rect 696 1470 707 1481
rect 713 1470 892 1578
rect 696 1440 892 1470
rect 895 1485 953 1491
rect 895 1451 920 1485
rect 895 1445 953 1451
rect 696 1429 707 1440
rect 568 1385 628 1418
rect 494 1381 528 1385
rect 540 1372 556 1385
rect 582 1381 616 1385
rect 434 1236 448 1368
rect 460 1364 468 1368
rect 504 1364 556 1372
rect 610 1364 644 1368
rect 460 1357 474 1364
rect 460 1352 468 1357
rect 504 1338 568 1364
rect 572 1347 644 1364
rect 696 1366 710 1418
rect 713 1366 892 1440
rect 572 1338 622 1347
rect 522 1304 622 1338
rect 522 1288 568 1304
rect 576 1298 584 1304
rect 604 1270 622 1304
rect 696 1236 892 1366
rect 895 1285 953 1291
rect 895 1251 907 1285
rect 895 1245 953 1251
rect 0 1219 656 1236
rect 380 1202 656 1219
rect 710 1202 892 1236
rect 346 1196 392 1202
rect 334 1184 392 1196
rect 422 1184 480 1202
rect 510 1184 656 1202
rect 346 1180 380 1182
rect 434 1180 468 1182
rect 522 1180 556 1184
rect 610 1180 644 1182
rect 713 1148 892 1202
rect 380 1146 892 1148
rect 380 1137 433 1146
rect 469 1137 521 1146
rect 663 1137 892 1146
rect 380 1129 422 1137
rect 0 1125 422 1129
rect 480 1125 510 1137
rect 674 1134 892 1137
rect 0 1114 433 1125
rect 469 1122 521 1125
rect 530 1122 634 1126
rect 674 1125 704 1134
rect 469 1114 652 1122
rect 663 1114 704 1125
rect 0 1038 414 1114
rect 480 1088 552 1104
rect 480 1074 618 1088
rect 552 1054 618 1074
rect 696 1056 704 1114
rect 713 1113 892 1134
rect 1082 1149 1152 1608
rect 1434 1589 1468 1608
rect 1264 1540 1322 1546
rect 1264 1506 1276 1540
rect 1264 1500 1322 1506
rect 1264 1232 1322 1238
rect 1264 1198 1276 1232
rect 1264 1192 1322 1198
rect 1082 1113 1135 1149
rect 719 1056 730 1067
rect 11 978 45 1038
rect 111 1026 261 1038
rect 327 1026 414 1038
rect 111 1007 134 1026
rect 153 984 176 1007
rect 327 1002 480 1026
rect 522 1020 588 1046
rect 696 1026 730 1056
rect 1082 1042 1146 1113
rect 1453 1096 1468 1589
rect 1487 1555 1522 1589
rect 1802 1555 1837 1589
rect 1487 1129 1521 1555
rect 1803 1536 1837 1555
rect 1633 1487 1691 1493
rect 1633 1453 1645 1487
rect 1633 1447 1691 1453
rect 1633 1179 1691 1185
rect 1633 1145 1645 1179
rect 1633 1139 1691 1145
rect 1822 1129 1837 1536
rect 1856 1502 1891 1536
rect 2171 1502 2206 1536
rect 1856 1129 1890 1502
rect 2172 1483 2206 1502
rect 2191 1440 2206 1483
rect 2002 1434 2060 1440
rect 2002 1400 2014 1434
rect 2002 1394 2060 1400
rect 1958 1173 2016 1202
rect 2046 1173 2104 1202
rect 1970 1169 2004 1173
rect 2058 1169 2092 1173
rect 2016 1148 2082 1160
rect 2172 1148 2206 1440
rect 1920 1135 2206 1148
rect 1920 1129 1955 1135
rect 1487 1114 1955 1129
rect 1976 1126 2206 1135
rect 1998 1125 2206 1126
rect 1987 1114 2206 1125
rect 1487 1093 1954 1114
rect 2002 1098 2014 1114
rect 2020 1098 2064 1104
rect 1487 1056 1502 1093
rect 1515 1056 1954 1093
rect 1998 1076 2064 1098
rect 2172 1086 2206 1114
rect 1487 1043 1954 1056
rect 2172 1056 2183 1067
rect 2191 1056 2206 1086
rect 1082 1038 1468 1042
rect 522 1006 584 1020
rect 522 1004 552 1006
rect 510 1002 552 1004
rect 169 978 203 980
rect 327 978 414 1002
rect 490 996 552 1002
rect 490 978 612 996
rect 696 984 704 1026
rect 712 1023 730 1026
rect 1118 1026 1468 1038
rect 1118 1023 1153 1026
rect 712 1010 766 1023
rect 712 987 768 1010
rect 1082 1008 1153 1023
rect 1433 1008 1468 1026
rect 712 984 845 987
rect 902 984 1065 987
rect 1082 984 1152 1008
rect 696 978 1152 984
rect 0 956 414 978
rect 468 965 488 978
rect 490 965 576 978
rect 582 965 616 976
rect 622 965 1152 978
rect 1434 989 1468 1008
rect 1515 1024 1954 1043
rect 2066 1046 2124 1052
rect 2066 1026 2078 1046
rect 2172 1026 2206 1056
rect 2062 1024 2080 1026
rect 2110 1024 2128 1026
rect 2172 1024 2183 1026
rect 1515 1015 2183 1024
rect 1515 1012 2150 1015
rect 1515 1004 2128 1012
rect 1515 1003 2160 1004
rect 1515 996 2190 1003
rect 2191 996 2206 1026
rect 1515 990 2206 996
rect 2225 1449 2260 1483
rect 2540 1449 2575 1466
rect 2225 1148 2259 1449
rect 2541 1448 2575 1449
rect 2541 1412 2611 1448
rect 2558 1387 2629 1412
rect 2371 1381 2429 1387
rect 2371 1347 2383 1381
rect 2541 1378 2629 1387
rect 2909 1378 2944 1412
rect 2371 1341 2429 1347
rect 1515 989 1954 990
rect 1434 984 1445 989
rect 1453 984 1468 989
rect 468 962 1152 965
rect 460 956 468 962
rect 482 956 540 962
rect 570 956 628 962
rect 0 950 628 956
rect 696 954 1152 962
rect 696 950 704 954
rect 712 950 1152 954
rect 0 942 1152 950
rect 1242 942 1344 974
rect 1434 954 1468 984
rect 1434 946 1445 954
rect 1453 946 1468 954
rect 1434 942 1468 946
rect 1487 942 1954 989
rect 2030 965 2080 990
rect 2022 954 2080 965
rect 2110 965 2160 990
rect 2225 971 2270 1148
rect 2327 1120 2385 1149
rect 2415 1120 2473 1149
rect 2541 1131 2628 1378
rect 2910 1359 2944 1378
rect 2740 1310 2798 1316
rect 2740 1276 2752 1310
rect 2740 1270 2798 1276
rect 2339 1116 2373 1120
rect 2427 1116 2461 1120
rect 2385 1095 2451 1107
rect 2541 1095 2675 1131
rect 2289 1082 2675 1095
rect 2289 1067 2324 1082
rect 2345 1073 2675 1082
rect 2367 1072 2675 1073
rect 2356 1067 2675 1072
rect 2289 1061 2675 1067
rect 2289 971 2323 1061
rect 2371 1039 2383 1061
rect 2389 1039 2539 1051
rect 2371 1033 2539 1039
rect 2389 1026 2539 1033
rect 2367 1023 2433 1026
rect 2435 993 2493 999
rect 2435 980 2447 993
rect 2435 978 2481 980
rect 2541 978 2675 1061
rect 2696 1058 2754 1071
rect 2784 1058 2842 1071
rect 2910 1056 2921 1067
rect 2929 1056 2944 1359
rect 2910 1026 2944 1056
rect 2740 1020 2798 1026
rect 2740 986 2752 1020
rect 2910 1015 2921 1026
rect 2740 980 2798 986
rect 2910 984 2921 995
rect 2910 978 2924 984
rect 2929 978 2944 1026
rect 2963 1325 2998 1359
rect 3278 1325 3313 1359
rect 2963 1025 2997 1325
rect 3279 1306 3313 1325
rect 3109 1257 3167 1263
rect 3109 1223 3121 1257
rect 3109 1217 3167 1223
rect 3095 1177 3233 1207
rect 2999 1143 3051 1177
rect 3065 1143 3211 1177
rect 3279 1143 3287 1211
rect 3298 1177 3313 1306
rect 3332 1272 3367 1306
rect 3647 1272 3682 1306
rect 3332 1178 3366 1272
rect 3648 1253 3682 1272
rect 4034 1253 4087 1254
rect 3478 1204 3536 1210
rect 3478 1180 3490 1204
rect 3478 1178 3492 1180
rect 3522 1178 3524 1180
rect 3667 1178 3682 1253
rect 3701 1219 3736 1253
rect 4016 1219 4087 1253
rect 3701 1178 3735 1219
rect 4017 1218 4087 1219
rect 4034 1184 4105 1218
rect 3332 1177 3754 1178
rect 3314 1143 3754 1177
rect 2999 1025 3033 1143
rect 3065 1057 3087 1143
rect 3165 1109 3203 1113
rect 3107 1057 3111 1109
rect 3165 1091 3225 1109
rect 3065 1025 3123 1057
rect 3141 1041 3145 1075
rect 3153 1041 3225 1091
rect 3281 1057 3313 1143
rect 3153 1025 3211 1041
rect 3279 1025 3313 1057
rect 3315 1099 3754 1143
rect 3847 1151 3905 1157
rect 3847 1117 3859 1151
rect 3847 1111 3905 1117
rect 4034 1107 4104 1184
rect 4216 1116 4274 1122
rect 3833 1099 3971 1101
rect 4017 1099 4025 1105
rect 4034 1099 4123 1107
rect 3315 1025 4123 1099
rect 4216 1082 4228 1116
rect 4216 1076 4274 1082
rect 4202 1036 4340 1057
rect 4202 1035 4271 1036
rect 2963 978 4123 1025
rect 2435 971 2493 978
rect 2541 971 4123 978
rect 4172 1010 4360 1035
rect 4386 1010 4420 1122
rect 4172 976 4420 1010
rect 2110 954 2168 965
rect 2022 942 2068 954
rect 2122 942 2168 954
rect 2225 954 4123 971
rect 2225 943 2270 954
rect 2236 942 2270 943
rect 2289 950 2497 954
rect 2289 942 2521 950
rect 2558 942 4123 954
rect 0 940 4123 942
rect 0 934 4140 940
rect 0 922 656 934
rect 663 931 704 934
rect 0 908 660 922
rect 674 919 704 931
rect 663 908 704 919
rect 713 914 4140 934
rect 4147 914 4168 976
rect 713 908 4168 914
rect 0 764 414 908
rect 434 854 468 908
rect 482 885 650 908
rect 656 885 1152 908
rect 482 870 1152 885
rect 434 826 474 854
rect 482 840 656 870
rect 696 840 1152 870
rect 1278 859 1294 860
rect 1220 845 1278 859
rect 1308 845 1366 859
rect 1220 844 1266 845
rect 434 792 468 826
rect 482 825 1152 840
rect 482 797 650 825
rect 434 766 474 792
rect 482 790 628 797
rect 482 785 644 790
rect 494 781 502 785
rect 522 772 568 785
rect 582 781 590 785
rect 434 764 448 766
rect 460 764 474 766
rect 504 764 568 772
rect 572 766 598 776
rect 610 766 644 785
rect 572 764 622 766
rect 656 764 1152 825
rect 0 754 656 764
rect 0 640 414 754
rect 434 752 448 754
rect 460 752 468 754
rect 434 728 468 752
rect 504 738 568 754
rect 572 752 622 754
rect 572 738 644 752
rect 522 728 644 738
rect 434 686 448 728
rect 522 704 622 728
rect 522 698 584 704
rect 522 688 568 698
rect 604 688 622 704
rect 562 686 622 688
rect 641 686 656 701
rect 422 670 480 686
rect 510 670 656 686
rect 422 666 656 670
rect 696 666 1152 764
rect 1176 762 1186 766
rect 1198 762 1210 766
rect 1222 762 1266 844
rect 1320 833 1354 845
rect 1320 818 1366 833
rect 422 656 1152 666
rect 434 641 1152 656
rect 434 640 644 641
rect 656 640 1152 641
rect 0 619 1152 640
rect 70 606 1152 619
rect 380 602 656 606
rect 710 602 1152 606
rect 522 580 556 602
rect 713 530 1152 602
rect 1164 651 1216 762
rect 1226 750 1266 762
rect 1286 762 1298 790
rect 1310 773 1366 818
rect 1286 761 1304 762
rect 1278 750 1304 761
rect 1226 691 1304 750
rect 1226 679 1244 691
rect 1232 675 1244 679
rect 1264 679 1304 691
rect 1310 750 1354 773
rect 1310 691 1386 750
rect 1310 679 1340 691
rect 1352 679 1386 691
rect 1264 666 1308 679
rect 1164 641 1210 651
rect 1242 648 1308 666
rect 1310 648 1386 679
rect 1164 584 1206 641
rect 1242 632 1386 648
rect 1260 598 1386 632
rect 1260 584 1310 598
rect 1318 592 1322 598
rect 1346 584 1350 598
rect 1352 594 1386 598
rect 1352 584 1360 594
rect 1164 582 1222 584
rect 1252 582 1374 584
rect 1434 582 1468 908
rect 1176 578 1186 582
rect 1352 578 1360 582
rect 713 513 1170 530
rect 1211 519 1263 530
rect 1299 525 1415 530
rect 1363 519 1415 525
rect 1118 506 1170 513
rect 1222 507 1252 519
rect 1374 507 1404 519
rect 1118 496 1159 506
rect 1211 503 1263 507
rect 1211 496 1343 503
rect 1363 496 1415 507
rect 1452 496 1468 582
rect 1487 902 2168 908
rect 2191 902 2206 908
rect 1487 636 1954 902
rect 2022 890 2037 902
rect 2138 890 2168 902
rect 1956 868 2018 890
rect 2022 881 2080 890
rect 2022 868 2081 881
rect 1956 860 2082 868
rect 2110 860 2168 890
rect 1974 854 2082 860
rect 2022 840 2082 854
rect 2002 828 2082 840
rect 1998 816 2082 828
rect 2138 816 2168 860
rect 1998 800 2168 816
rect 2002 794 2079 800
rect 1956 790 1990 794
rect 1956 769 2002 790
rect 2022 785 2079 794
rect 2080 785 2168 800
rect 1956 766 1996 769
rect 1956 741 1990 766
rect 2001 753 2002 769
rect 2020 781 2068 785
rect 2080 784 2106 785
rect 2020 772 2048 781
rect 2080 772 2090 784
rect 2122 781 2156 785
rect 2020 754 2092 772
rect 2172 766 2206 902
rect 2236 883 2270 908
rect 2289 883 2323 908
rect 2403 883 2437 900
rect 2491 883 2525 900
rect 2558 883 4168 908
rect 2144 762 2206 766
rect 2044 753 2092 754
rect 1956 636 2004 741
rect 2044 738 2104 753
rect 2132 747 2206 762
rect 2046 636 2048 738
rect 2062 688 2104 738
rect 2106 704 2128 738
rect 2110 698 2124 704
rect 2089 673 2104 688
rect 2132 670 2162 747
rect 2058 636 2092 670
rect 2132 636 2158 670
rect 2172 636 2206 747
rect 2225 874 4168 883
rect 2225 849 2537 874
rect 2558 866 4168 874
rect 2540 849 4168 866
rect 4172 907 4222 976
rect 4272 968 4318 976
rect 4259 950 4260 955
rect 4272 950 4332 968
rect 4172 857 4230 907
rect 4248 900 4252 934
rect 4259 908 4332 950
rect 4260 891 4318 908
rect 4326 900 4340 908
rect 4324 891 4340 900
rect 4260 874 4342 891
rect 4260 868 4338 874
rect 4260 857 4318 868
rect 4172 855 4254 857
rect 4260 855 4342 857
rect 4184 853 4218 855
rect 4220 853 4254 855
rect 4266 853 4306 855
rect 4308 853 4342 855
rect 4184 851 4266 853
rect 4272 851 4354 853
rect 2225 636 2270 849
rect 1487 619 2104 636
rect 1487 477 1521 619
rect 1552 477 1555 619
rect 1563 600 1592 619
rect 1640 613 1686 619
rect 1567 598 1592 600
rect 1567 588 1586 598
rect 1611 579 1686 613
rect 1702 579 1732 619
rect 1629 545 1732 579
rect 1629 529 1686 545
rect 1702 529 1732 545
rect 1803 564 1837 619
rect 1856 606 1902 619
rect 1920 610 2104 619
rect 1803 530 1840 564
rect 1856 550 1890 606
rect 1920 602 1955 610
rect 1958 602 2104 610
rect 2132 602 2270 636
rect 2289 750 2323 849
rect 2403 815 2450 828
rect 2343 812 2397 815
rect 2403 812 2451 815
rect 2343 792 2451 812
rect 2476 810 2491 844
rect 2507 826 2537 849
rect 2391 787 2451 792
rect 2371 781 2451 787
rect 2333 762 2354 766
rect 2333 750 2360 762
rect 2289 713 2360 750
rect 2367 761 2451 781
rect 2367 747 2453 761
rect 2494 760 2537 826
rect 2507 747 2537 760
rect 2371 741 2388 747
rect 2396 732 2442 747
rect 2449 732 2453 747
rect 2503 732 2537 747
rect 2396 719 2454 732
rect 2507 728 2539 732
rect 2518 719 2539 728
rect 2289 688 2354 713
rect 2396 700 2461 719
rect 2467 700 2539 719
rect 2366 688 2373 699
rect 1958 573 1959 602
rect 1970 585 2004 602
rect 2046 588 2048 602
rect 2046 585 2058 588
rect 2046 573 2063 585
rect 2132 582 2158 602
rect 2172 582 2206 602
rect 1671 514 1686 529
rect 1803 477 1837 530
rect 1487 443 1686 477
rect 1691 472 1743 477
rect 1822 472 1837 477
rect 1691 466 1837 472
rect 1702 454 1837 466
rect 1691 443 1837 454
rect 1856 514 1874 550
rect 1879 539 1890 550
rect 1856 472 1890 514
rect 1856 409 1871 472
rect 1974 458 1990 560
rect 2002 526 2060 532
rect 2002 492 2018 526
rect 2190 492 2206 582
rect 2002 486 2060 492
rect 1998 476 2064 478
rect 1903 413 2073 424
rect 2105 413 2157 424
rect 1856 401 1870 409
rect 1914 406 2062 413
rect 2032 401 2062 406
rect 2116 401 2146 413
rect 1856 390 1881 401
rect 2021 390 2073 401
rect 2105 390 2157 401
rect 2191 390 2206 492
rect 2225 582 2266 602
rect 2225 492 2240 582
rect 2255 578 2266 582
rect 2289 594 2373 688
rect 2289 583 2323 594
rect 2339 583 2373 594
rect 2374 583 2379 700
rect 2402 583 2407 700
rect 2408 698 2539 700
rect 2408 691 2473 698
rect 2408 685 2493 691
rect 2408 670 2495 685
rect 2408 620 2473 670
rect 2481 651 2495 670
rect 2518 635 2539 698
rect 2541 706 4168 849
rect 4208 842 4266 851
rect 4296 843 4354 851
rect 4296 842 4348 843
rect 4194 840 4348 842
rect 4194 827 4342 840
rect 4194 808 4296 827
rect 4208 774 4296 808
rect 4302 815 4342 827
rect 4352 827 4370 831
rect 4352 815 4382 827
rect 4208 706 4288 774
rect 4302 706 4382 815
rect 4386 706 4420 976
rect 2541 672 4382 706
rect 4388 672 4420 706
rect 4422 914 4474 976
rect 4422 911 4484 914
rect 4844 911 4879 929
rect 2408 594 2461 620
rect 2427 583 2461 594
rect 2541 618 4168 672
rect 4230 642 4248 660
rect 4266 652 4294 672
rect 4264 642 4294 652
rect 4230 626 4294 642
rect 4298 626 4370 672
rect 4248 618 4370 626
rect 2541 586 4382 618
rect 2541 583 4123 586
rect 2289 582 4123 583
rect 2255 515 2259 578
rect 2289 554 2313 582
rect 2327 560 4123 582
rect 2327 554 3457 560
rect 2289 549 3457 554
rect 2339 532 2385 549
rect 2541 536 3457 549
rect 3496 554 3540 560
rect 3556 554 3582 560
rect 3496 542 3522 554
rect 3554 542 3602 554
rect 3538 536 3602 542
rect 2351 525 2385 532
rect 2327 520 2385 525
rect 2444 520 2467 536
rect 2541 532 3464 536
rect 3534 532 3602 536
rect 2225 390 2259 492
rect 2343 458 2354 507
rect 2472 492 2495 508
rect 2367 450 2368 480
rect 2371 473 2429 479
rect 2371 450 2383 473
rect 2367 423 2433 450
rect 2541 426 3484 532
rect 3516 526 3602 532
rect 3523 517 3580 526
rect 3538 476 3580 517
rect 3588 492 3602 526
rect 3565 461 3580 476
rect 2541 416 2944 426
rect 2368 405 2434 408
rect 2225 380 2240 390
rect 224 126 228 362
rect 1906 354 2452 380
rect 2541 371 2548 416
rect 2507 360 2548 371
rect 252 154 256 334
rect 2189 312 2452 354
rect 2518 348 2548 360
rect 2558 386 2944 416
rect 2558 348 2628 386
rect 2740 380 2798 386
rect 2910 380 2944 386
rect 2507 337 2628 348
rect 2250 303 2284 312
rect 2338 303 2372 312
rect 2384 308 2452 312
rect 2558 318 2628 337
rect 2910 337 2924 380
rect 2929 337 2944 380
rect 2910 318 2944 337
rect 2558 308 2647 318
rect 2695 316 2823 318
rect 2384 307 2647 308
rect 2384 301 2636 307
rect 1540 276 1796 300
rect 2594 295 2636 301
rect 2692 298 2826 316
rect 2849 298 2944 318
rect 2594 294 2647 295
rect 2692 294 2944 298
rect 2594 290 2944 294
rect 2963 424 3484 426
rect 3534 424 3568 458
rect 3648 424 3682 560
rect 2963 407 3682 424
rect 2963 306 2997 407
rect 3065 405 3115 407
rect 3153 405 3211 407
rect 3070 383 3100 405
rect 3123 383 3142 405
rect 3158 383 3188 405
rect 3105 380 3142 383
rect 3024 358 3031 362
rect 3105 358 3180 380
rect 2594 284 2946 290
rect 1568 248 1768 272
rect 2726 250 2792 282
rect 2929 256 2946 284
rect 1744 126 1768 248
rect 1772 154 1796 244
rect 2963 231 2980 306
rect 2987 265 2997 306
rect 3012 265 3051 358
rect 3100 343 3193 358
rect 3105 333 3193 343
rect 3105 317 3158 333
rect 3166 327 3167 333
rect 3194 299 3195 358
rect 3200 299 3205 362
rect 3279 277 3313 407
rect 3279 273 3300 277
rect 3279 265 3313 273
rect 3012 231 3246 265
rect 3300 231 3313 265
rect 3112 174 3146 231
rect 3332 212 3366 407
rect 3396 390 3400 407
rect 3412 390 3682 407
rect 3412 324 3434 390
rect 3440 352 3462 390
rect 3478 314 3536 320
rect 3478 280 3490 314
rect 3478 274 3536 280
rect 3648 274 3682 390
rect 3332 183 3446 212
rect 3332 178 3399 183
rect 3667 178 3682 274
rect 3701 507 4123 560
rect 4134 584 4382 586
rect 4388 584 4420 618
rect 3701 337 4115 507
rect 3701 301 4104 337
rect 3701 178 3735 301
rect 3847 261 3905 267
rect 3847 227 3859 261
rect 3847 221 3905 227
rect 1750 88 1768 126
rect 1778 88 1796 154
rect 3701 144 3716 178
rect 4034 125 4104 301
rect 4134 318 4168 584
rect 4248 576 4294 584
rect 4248 550 4282 576
rect 4330 558 4382 584
rect 4194 524 4282 550
rect 4336 524 4382 558
rect 4386 524 4420 584
rect 4422 573 4520 911
rect 4808 896 4879 911
rect 4808 779 4878 896
rect 4990 828 5048 834
rect 4990 794 5002 828
rect 4990 788 5048 794
rect 4621 773 4679 779
rect 4621 739 4633 773
rect 4621 733 4679 739
rect 4791 705 4878 779
rect 6294 711 6329 745
rect 4565 689 4623 703
rect 4565 669 4589 689
rect 4677 669 4711 703
rect 4577 635 4723 669
rect 4791 652 4889 705
rect 6295 692 6329 711
rect 4577 611 4591 635
rect 4422 524 4537 573
rect 4633 539 4695 573
rect 4661 533 4695 539
rect 4791 533 5230 652
rect 5610 599 5645 617
rect 5574 584 5645 599
rect 4190 490 4382 524
rect 4236 482 4296 490
rect 4236 467 4293 482
rect 4352 467 4382 490
rect 4234 463 4282 467
rect 4294 466 4320 467
rect 4234 454 4260 463
rect 4294 454 4302 466
rect 4352 463 4370 467
rect 4184 435 4202 439
rect 4234 436 4306 454
rect 4258 435 4306 436
rect 4172 318 4222 435
rect 4258 420 4318 435
rect 4276 370 4318 420
rect 4326 386 4340 420
rect 4303 355 4318 370
rect 4272 318 4306 352
rect 4386 318 4420 522
rect 4439 401 4537 524
rect 4617 471 4651 499
rect 4791 471 4805 533
rect 4605 437 4751 471
rect 4617 401 4651 437
rect 4450 318 4537 401
rect 4649 367 4707 373
rect 4649 333 4661 367
rect 4808 348 5230 533
rect 5241 529 5276 563
rect 4649 327 4707 333
rect 4134 284 4158 318
rect 4172 284 4420 318
rect 4216 208 4274 214
rect 4216 174 4228 208
rect 4216 168 4274 174
rect 4386 168 4420 284
rect 4467 284 4537 318
rect 4467 248 4520 284
rect 4838 231 4853 348
rect 4872 231 4906 348
rect 5018 314 5076 320
rect 5018 280 5030 314
rect 5018 274 5076 280
rect 4872 197 4887 231
rect 5207 178 5222 348
rect 5241 178 5275 529
rect 5387 461 5445 467
rect 5387 427 5399 461
rect 5387 421 5445 427
rect 5387 261 5445 267
rect 5387 227 5399 261
rect 5387 221 5445 227
rect 5241 144 5256 178
rect 5574 125 5644 584
rect 5756 516 5814 522
rect 5756 482 5768 516
rect 5756 476 5814 482
rect 5756 208 5814 214
rect 5756 174 5768 208
rect 5756 168 5814 174
rect 4034 89 4087 125
rect 5574 89 5627 125
rect 5945 72 5960 618
rect 5979 72 6013 672
rect 6125 643 6183 649
rect 6125 609 6137 643
rect 6125 603 6183 609
rect 6125 155 6183 161
rect 6125 121 6137 155
rect 6125 115 6183 121
rect 5979 38 5994 72
rect 6314 19 6329 692
rect 6348 658 6383 692
rect 6348 19 6382 658
rect 6348 -15 6363 19
rect 6681 0 6734 387
rect 7788 0 7841 281
rect 8157 0 8210 175
rect 8526 0 8579 175
rect 8895 0 8948 69
rect 9264 0 9317 69
rect 6681 -34 6751 0
rect 6681 -70 6734 -34
rect 7052 -87 7067 0
rect 7086 -87 7120 0
rect 7232 -4 7290 0
rect 7232 -38 7244 -4
rect 7232 -44 7290 -38
rect 7086 -121 7101 -87
rect 7421 -140 7436 0
rect 7455 -140 7489 0
rect 7601 -57 7659 -51
rect 7601 -91 7613 -57
rect 7601 -97 7659 -91
rect 7455 -174 7470 -140
rect 7788 -193 7858 0
rect 7970 -110 8028 -104
rect 7970 -144 7982 -110
rect 7970 -150 8028 -144
rect 7788 -229 7841 -193
rect 8157 -246 8227 0
rect 8339 -3 8397 0
rect 8339 -163 8397 -157
rect 8339 -197 8351 -163
rect 8339 -203 8397 -197
rect 8157 -282 8210 -246
rect 8526 -299 8596 0
rect 8895 -1 8966 0
rect 8708 -216 8766 -210
rect 8708 -250 8720 -216
rect 8708 -256 8766 -250
rect 8526 -335 8579 -299
rect 8895 -352 8965 -1
rect 9077 -69 9135 -63
rect 9077 -103 9089 -69
rect 9077 -109 9135 -103
rect 9077 -269 9135 -263
rect 9077 -303 9089 -269
rect 9077 -309 9135 -303
rect 8895 -388 8948 -352
rect 9264 -405 9334 0
rect 9446 -14 9504 -8
rect 9446 -48 9458 -14
rect 9446 -54 9504 -48
rect 9446 -322 9504 -316
rect 9446 -356 9458 -322
rect 9446 -362 9504 -356
rect 9264 -441 9317 -405
rect 284 -1623 337 -1622
rect 266 -1657 337 -1623
rect 267 -1658 337 -1657
rect 284 -1692 355 -1658
rect 1447 -1671 1482 -1653
rect 635 -1692 670 -1675
rect -43 -1822 -15 -1804
rect 284 -1822 354 -1692
rect 636 -1693 670 -1692
rect 1411 -1686 1482 -1671
rect 1762 -1686 1797 -1652
rect 636 -1729 706 -1693
rect 1078 -1728 1093 -1707
rect 1112 -1728 1394 -1710
rect 1411 -1728 1481 -1686
rect 1763 -1705 1797 -1686
rect 1022 -1729 1481 -1728
rect 653 -1754 724 -1729
rect 466 -1760 524 -1754
rect 466 -1794 478 -1760
rect 636 -1763 724 -1754
rect 1004 -1763 1481 -1729
rect 1782 -1748 1797 -1705
rect 466 -1800 524 -1794
rect -72 -2136 354 -1822
rect 636 -1822 723 -1763
rect 1005 -1764 1481 -1763
rect 1022 -1822 1481 -1764
rect 428 -1850 437 -1841
rect 391 -1946 409 -1850
rect 419 -1853 437 -1850
rect 419 -1858 468 -1853
rect 522 -1858 556 -1853
rect 636 -1858 1481 -1822
rect 1561 -1858 1595 -1824
rect 1649 -1858 1683 -1824
rect 1763 -1858 1797 -1748
rect 1816 -1739 1851 -1705
rect 1816 -1858 1850 -1739
rect 3607 -1771 3642 -1737
rect 1962 -1807 2020 -1801
rect 1962 -1820 1974 -1807
rect 1962 -1822 2008 -1820
rect 1962 -1824 2020 -1822
rect 1958 -1841 2024 -1824
rect 2132 -1830 2166 -1801
rect 2518 -1830 2729 -1775
rect 3608 -1790 3642 -1771
rect 1962 -1847 2020 -1841
rect 1934 -1858 2048 -1850
rect 2132 -1858 2475 -1830
rect 419 -1892 2475 -1858
rect 419 -1946 468 -1892
rect 428 -1948 468 -1946
rect 522 -1935 556 -1892
rect 636 -1910 1813 -1892
rect 1816 -1910 1850 -1892
rect 1892 -1904 2064 -1892
rect 428 -1974 474 -1948
rect 434 -2009 474 -1974
rect 495 -1975 502 -1972
rect 522 -1975 568 -1935
rect 495 -1976 568 -1975
rect 583 -1976 590 -1946
rect 489 -1977 562 -1976
rect 484 -1988 562 -1977
rect 461 -2021 474 -2009
rect 489 -2009 562 -1988
rect 489 -2021 529 -2009
rect 549 -2021 562 -2009
rect 577 -1988 590 -1976
rect 602 -1976 617 -1972
rect 461 -2025 468 -2021
rect 483 -2034 542 -2021
rect 549 -2025 556 -2021
rect 483 -2102 546 -2034
rect 577 -2047 594 -1988
rect 577 -2049 590 -2047
rect 583 -2059 590 -2049
rect 483 -2116 528 -2102
rect 602 -2116 629 -1976
rect -72 -2165 386 -2136
rect 483 -2156 541 -2116
rect 571 -2156 629 -2116
rect 636 -2155 1850 -1910
rect 1930 -1930 1964 -1904
rect 2018 -1925 2052 -1904
rect 1988 -1930 2052 -1925
rect 2112 -1920 2118 -1904
rect 2132 -1920 2475 -1892
rect 1988 -1938 2035 -1930
rect 1920 -1972 1930 -1938
rect 1970 -1946 2038 -1938
rect 1938 -1966 1976 -1956
rect 1988 -1966 2038 -1946
rect 1938 -1974 2038 -1966
rect 2049 -1974 2064 -1959
rect 1918 -2006 1933 -1997
rect 1938 -2006 2064 -1974
rect 1918 -2010 1976 -2006
rect 2018 -2008 2064 -2006
rect 1984 -2010 2000 -2008
rect 1918 -2012 2000 -2010
rect 1876 -2038 1881 -2034
rect 1918 -2038 1976 -2012
rect 2012 -2038 2064 -2008
rect 2071 -2024 2087 -1990
rect 1876 -2050 1887 -2038
rect 495 -2160 529 -2156
rect 583 -2160 617 -2156
rect -72 -2170 354 -2165
rect 636 -2170 1864 -2155
rect -72 -2181 420 -2170
rect -72 -2187 340 -2181
rect 16 -2200 28 -2194
rect 320 -2204 340 -2187
rect 354 -2199 420 -2181
rect 461 -2181 1864 -2170
rect 461 -2194 1092 -2181
rect 510 -2202 571 -2194
rect 510 -2204 562 -2202
rect 634 -2204 1092 -2194
rect 653 -2240 1092 -2204
rect 419 -2276 1092 -2240
rect 1178 -2239 1213 -2181
rect 1216 -2208 1239 -2181
rect 1259 -2220 1266 -2181
rect 1374 -2206 1864 -2181
rect 1872 -2183 1887 -2050
rect 1910 -2053 1915 -2049
rect 1904 -2054 1915 -2053
rect 1930 -2053 1976 -2038
rect 1998 -2049 2064 -2038
rect 1998 -2053 2003 -2049
rect 1899 -2065 1923 -2054
rect 1930 -2056 1975 -2053
rect 1992 -2054 2003 -2053
rect 1935 -2065 1975 -2056
rect 1987 -2065 2006 -2054
rect 2018 -2056 2064 -2049
rect 2030 -2065 2064 -2056
rect 1904 -2068 1975 -2065
rect 1992 -2068 2064 -2065
rect 1904 -2099 1969 -2068
rect 1976 -2081 1981 -2068
rect 1986 -2081 2044 -2068
rect 1975 -2099 2044 -2081
rect 1904 -2102 2044 -2099
rect 1904 -2109 1981 -2102
rect 1986 -2109 2044 -2102
rect 1904 -2149 2044 -2109
rect 1904 -2165 1981 -2149
rect 1986 -2165 2024 -2149
rect 1904 -2183 1975 -2165
rect 1872 -2206 1975 -2183
rect 1374 -2217 1850 -2206
rect 1876 -2217 1944 -2206
rect 1964 -2217 1975 -2206
rect 1992 -2183 2007 -2165
rect 2030 -2183 2044 -2149
rect 1992 -2217 2044 -2183
rect 1374 -2218 2086 -2217
rect 1301 -2224 1308 -2220
rect 1178 -2246 1201 -2239
rect 1340 -2242 1367 -2236
rect 1301 -2270 1367 -2242
rect 1374 -2246 1835 -2218
rect 1374 -2251 1831 -2246
rect 1374 -2276 1830 -2251
rect 1876 -2261 1881 -2218
rect 1893 -2228 2086 -2218
rect 1893 -2233 2044 -2228
rect 1893 -2240 1923 -2233
rect 1956 -2240 1986 -2233
rect 2045 -2240 2075 -2228
rect 1882 -2242 1934 -2240
rect 1945 -2242 1997 -2240
rect 1882 -2246 2026 -2242
rect 2034 -2246 2086 -2240
rect 1882 -2251 2086 -2246
rect 2112 -2251 2475 -1920
rect 1896 -2264 1923 -2251
rect 1956 -2264 1965 -2251
rect 419 -2293 1213 -2276
rect 1218 -2287 1830 -2276
rect 177 -2352 200 -2323
rect 205 -2324 228 -2323
rect 186 -2396 200 -2352
rect 123 -2400 200 -2396
rect 214 -2424 228 -2324
rect 419 -2362 663 -2293
rect 1024 -2344 1025 -2293
rect 1058 -2310 1213 -2293
rect 1229 -2299 1259 -2287
rect 1267 -2299 1830 -2287
rect 1218 -2304 1830 -2299
rect 1218 -2310 1270 -2304
rect 1391 -2363 1830 -2304
rect 1938 -2280 1965 -2264
rect 1938 -2285 2004 -2280
rect 1938 -2320 1965 -2285
rect 2045 -2330 2046 -2251
rect 2112 -2320 2146 -2251
rect 1391 -2399 1813 -2363
rect 1823 -2382 1830 -2363
rect 2112 -2350 2123 -2339
rect 2135 -2350 2146 -2339
rect 2149 -2340 2475 -2251
rect 2518 -1845 2589 -1830
rect 3438 -1839 3496 -1833
rect 2518 -2304 2588 -1845
rect 3438 -1873 3450 -1839
rect 3438 -1879 3496 -1873
rect 2700 -1913 2758 -1907
rect 2700 -1947 2712 -1913
rect 2870 -1936 2904 -1918
rect 3292 -1936 3326 -1918
rect 2700 -1953 2758 -1947
rect 2870 -1972 2940 -1936
rect 2887 -2006 2958 -1972
rect 2700 -2221 2758 -2215
rect 2700 -2255 2712 -2221
rect 2700 -2261 2758 -2255
rect 2518 -2340 2571 -2304
rect 2112 -2382 2146 -2350
rect 1823 -2393 1864 -2382
rect 2034 -2384 2146 -2382
rect 1823 -2405 1853 -2393
rect 1812 -2406 1853 -2405
rect 1895 -2405 1961 -2392
rect 2034 -2393 2075 -2384
rect 2045 -2405 2075 -2393
rect 2135 -2395 2146 -2384
rect 2518 -2374 2729 -2340
rect 2887 -2357 2957 -2006
rect 3069 -2074 3127 -2068
rect 3069 -2108 3081 -2074
rect 3069 -2114 3127 -2108
rect 3069 -2274 3127 -2268
rect 3069 -2308 3081 -2274
rect 3069 -2314 3127 -2308
rect 2518 -2393 2695 -2374
rect 2887 -2393 2940 -2357
rect 1895 -2406 1972 -2405
rect 1812 -2416 1972 -2406
rect 2034 -2416 2086 -2405
rect 3256 -2410 3326 -1936
rect 3438 -2327 3496 -2321
rect 3438 -2361 3450 -2327
rect 3438 -2367 3496 -2361
rect 2122 -2416 2146 -2415
rect 151 -2428 228 -2424
rect 1760 -2452 1979 -2420
rect 3256 -2446 3309 -2410
rect 3627 -2463 3642 -1790
rect 3661 -1824 3696 -1790
rect 3661 -2463 3695 -1824
rect 3807 -1892 3865 -1886
rect 3807 -1926 3819 -1892
rect 3807 -1932 3865 -1926
rect 3977 -2095 4011 -2077
rect 5821 -2089 5856 -2055
rect 3977 -2131 4047 -2095
rect 5822 -2108 5856 -2089
rect 3994 -2165 4065 -2131
rect 4345 -2165 4380 -2131
rect 3807 -2380 3865 -2374
rect 3807 -2414 3819 -2380
rect 3807 -2420 3865 -2414
rect 3661 -2497 3676 -2463
rect 1067 -2524 1323 -2500
rect 3994 -2516 4064 -2165
rect 4346 -2184 4380 -2165
rect 4176 -2233 4234 -2227
rect 4176 -2267 4188 -2233
rect 4176 -2273 4234 -2267
rect 4176 -2433 4234 -2427
rect 4176 -2467 4188 -2433
rect 4176 -2473 4234 -2467
rect 389 -2594 398 -2540
rect 1095 -2552 1295 -2528
rect 3994 -2552 4047 -2516
rect 443 -2617 452 -2594
rect 1271 -2674 1295 -2552
rect 1299 -2646 1323 -2556
rect 4365 -2569 4380 -2184
rect 4399 -2218 4434 -2184
rect 4714 -2218 4749 -2184
rect 5137 -2201 5172 -2183
rect 4399 -2569 4433 -2218
rect 4715 -2237 4749 -2218
rect 5101 -2216 5172 -2201
rect 4545 -2286 4603 -2280
rect 4545 -2320 4557 -2286
rect 4545 -2326 4603 -2320
rect 4545 -2486 4603 -2480
rect 4545 -2520 4557 -2486
rect 4545 -2526 4603 -2520
rect 4399 -2603 4414 -2569
rect 4734 -2622 4749 -2237
rect 4768 -2271 4803 -2237
rect 4768 -2622 4802 -2271
rect 4914 -2339 4972 -2333
rect 4914 -2373 4926 -2339
rect 4914 -2379 4972 -2373
rect 4914 -2539 4972 -2533
rect 4914 -2573 4926 -2539
rect 4914 -2579 4972 -2573
rect 1277 -2712 1295 -2674
rect 1305 -2712 1323 -2646
rect 4768 -2656 4783 -2622
rect 5101 -2675 5171 -2216
rect 5283 -2284 5341 -2278
rect 5283 -2318 5295 -2284
rect 5283 -2324 5341 -2318
rect 5283 -2592 5341 -2586
rect 5283 -2626 5295 -2592
rect 5283 -2632 5341 -2626
rect 5101 -2711 5154 -2675
rect 391 -2718 409 -2712
rect 419 -2718 437 -2712
rect 5472 -2728 5487 -2182
rect 5506 -2728 5540 -2128
rect 5652 -2157 5710 -2151
rect 5652 -2191 5664 -2157
rect 5652 -2197 5710 -2191
rect 5652 -2645 5710 -2639
rect 5652 -2679 5664 -2645
rect 5652 -2685 5710 -2679
rect 391 -2800 409 -2748
rect 419 -2800 437 -2748
rect 5506 -2762 5521 -2728
rect 5841 -2781 5856 -2108
rect 5875 -2142 5910 -2108
rect 5875 -2781 5909 -2142
rect 6021 -2210 6079 -2204
rect 6021 -2244 6033 -2210
rect 6021 -2250 6079 -2244
rect 6191 -2413 6225 -2395
rect 6191 -2449 6261 -2413
rect 6208 -2483 6279 -2449
rect 6559 -2483 6594 -2449
rect 6021 -2698 6079 -2692
rect 6021 -2732 6033 -2698
rect 6021 -2738 6079 -2732
rect 5875 -2815 5890 -2781
rect 6208 -2834 6278 -2483
rect 6560 -2502 6594 -2483
rect 6390 -2551 6448 -2545
rect 6390 -2585 6402 -2551
rect 6390 -2591 6448 -2585
rect 6390 -2751 6448 -2745
rect 6390 -2785 6402 -2751
rect 6390 -2791 6448 -2785
rect 6208 -2870 6261 -2834
rect 6579 -2887 6594 -2502
rect 6613 -2536 6648 -2502
rect 6928 -2536 6963 -2502
rect 7351 -2519 7386 -2501
rect 6613 -2887 6647 -2536
rect 6929 -2555 6963 -2536
rect 7315 -2534 7386 -2519
rect 6759 -2604 6817 -2598
rect 6759 -2638 6771 -2604
rect 6759 -2644 6817 -2638
rect 6759 -2804 6817 -2798
rect 6759 -2838 6771 -2804
rect 6759 -2844 6817 -2838
rect 6613 -2921 6628 -2887
rect 6948 -2940 6963 -2555
rect 6982 -2589 7017 -2555
rect 6982 -2940 7016 -2589
rect 7128 -2657 7186 -2651
rect 7128 -2691 7140 -2657
rect 7128 -2697 7186 -2691
rect 7128 -2857 7186 -2851
rect 7128 -2891 7140 -2857
rect 7128 -2897 7186 -2891
rect 6982 -2974 6997 -2940
rect 7315 -2993 7385 -2534
rect 7497 -2602 7555 -2596
rect 7497 -2636 7509 -2602
rect 7667 -2625 7701 -2607
rect 8089 -2625 8124 -2607
rect 7497 -2642 7555 -2636
rect 7667 -2661 7737 -2625
rect 8053 -2640 8124 -2625
rect 7684 -2695 7755 -2661
rect 7497 -2910 7555 -2904
rect 7497 -2944 7509 -2910
rect 7497 -2950 7555 -2944
rect 7315 -3029 7368 -2993
rect 7684 -3046 7754 -2695
rect 7866 -2763 7924 -2757
rect 7866 -2797 7878 -2763
rect 7866 -2803 7924 -2797
rect 7866 -2963 7924 -2957
rect 7866 -2997 7878 -2963
rect 7866 -3003 7924 -2997
rect 7684 -3082 7737 -3046
rect 8053 -3099 8123 -2640
rect 8235 -2708 8293 -2702
rect 8235 -2742 8247 -2708
rect 8405 -2731 8439 -2713
rect 8827 -2731 8862 -2713
rect 8235 -2748 8293 -2742
rect 8405 -2767 8475 -2731
rect 8791 -2746 8862 -2731
rect 8422 -2801 8493 -2767
rect 8235 -3016 8293 -3010
rect 8235 -3050 8247 -3016
rect 8235 -3056 8293 -3050
rect 8053 -3135 8106 -3099
rect 8422 -3152 8492 -2801
rect 8604 -2869 8662 -2863
rect 8604 -2903 8616 -2869
rect 8604 -2909 8662 -2903
rect 8604 -3069 8662 -3063
rect 8604 -3103 8616 -3069
rect 8604 -3109 8662 -3103
rect 8422 -3188 8475 -3152
rect 8791 -3205 8861 -2746
rect 8973 -2814 9031 -2808
rect 8973 -2848 8985 -2814
rect 8973 -2854 9031 -2848
rect 8973 -3122 9031 -3116
rect 8973 -3156 8985 -3122
rect 8973 -3162 9031 -3156
rect 8791 -3241 8844 -3205
<< nwell >>
rect 2948 474 2978 978
rect 2948 426 2976 474
<< poly >>
rect -72 1026 2996 1056
rect -72 314 -42 1026
rect 0 954 2924 984
rect 0 464 30 954
rect -72 278 2 314
rect 2894 306 2924 954
rect 2966 548 2996 1026
rect 3442 635 3457 669
rect 2966 496 3070 548
rect 2880 298 2946 306
rect 2780 290 2946 298
rect 2780 268 2896 290
rect 2880 256 2896 268
rect 2930 256 2946 290
rect 11 178 21 250
rect 2880 240 2946 256
rect 2942 132 2988 162
rect 882 -6 912 82
rect 1059 62 1119 78
rect 1661 58 1721 74
rect 0 -36 912 -6
rect 2874 -78 2904 52
rect 0 -108 2904 -78
<< polycont >>
rect 2896 256 2930 290
<< locali >>
rect 2880 256 2896 290
rect 2930 256 2946 290
<< viali >>
rect 2896 256 2930 290
<< metal1 >>
rect 635 880 679 902
rect 2948 854 2978 950
rect 3351 644 3365 656
rect 2880 298 2946 306
rect 2878 246 2888 298
rect 2940 246 2950 298
rect 2880 240 2946 246
rect 0 0 200 200
rect 1431 50 1493 76
rect 2946 0 2976 88
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
<< via1 >>
rect 2888 290 2940 298
rect 2888 256 2896 290
rect 2896 256 2930 290
rect 2930 256 2940 290
rect 2888 246 2940 256
<< metal2 >>
rect 2888 298 2940 308
rect 2888 236 2940 246
use flipflop  flipflop_0
timestamp 1624053917
transform 1 0 1568 0 1 72
box -686 -2400 8118 1112
use flipflop  x1
timestamp 1624053917
transform 1 0 1095 0 1 -2728
box -686 -2400 8118 1112
use and_masa  and_masa_0
timestamp 1624053917
transform 1 0 3016 0 1 66
box -53 -2000 2214 1147
use and_masa  x4
timestamp 1624053917
transform 1 0 -32 0 1 -2734
box -53 -2000 2214 1147
use xor_masa  xor_masa_0
timestamp 1624053917
transform 1 0 28 0 1 72
box -53 -2000 4428 1112
use xor_masa  xor_masa_1
timestamp 1624053917
transform 1 0 28 0 1 672
box -53 -2000 4428 1112
<< labels >>
rlabel space -28 278 30 314 1 ce
rlabel poly 2880 240 2946 306 1 Q
rlabel space 3418 635 3457 669 1 out
rlabel poly 1059 62 1119 78 1 clk
rlabel poly 1661 58 1721 74 1 clr
rlabel metal1 635 880 679 902 1 vdd
rlabel poly 11 178 21 250 1 ce
rlabel metal1 3351 644 3365 656 1 out
rlabel metal1 1431 50 1493 76 1 vss
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 ce
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 clr
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Q
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 out
port 7 nsew
<< end >>
