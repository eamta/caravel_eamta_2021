magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 3217 1639 3639 1658
rect 3639 1631 3665 1639
rect 3639 1623 4034 1631
rect 3568 1622 4034 1623
rect -196 1588 -161 1622
rect 3253 1619 4034 1622
rect -195 1569 -161 1588
rect 3217 1605 4034 1619
rect -365 1520 -307 1526
rect -365 1486 -353 1520
rect -365 1480 -307 1486
rect -365 1212 -307 1218
rect -365 1178 -353 1212
rect -365 1172 -307 1178
rect -176 1129 -161 1569
rect -142 1535 -107 1569
rect 173 1535 208 1569
rect 604 1549 613 1552
rect 3217 1551 3253 1605
rect 3287 1588 3622 1605
rect 3281 1569 3622 1588
rect 3281 1551 3586 1569
rect 3588 1555 3657 1569
rect 3745 1558 3797 1569
rect 3603 1551 3657 1555
rect 3756 1551 3786 1558
rect -142 1129 -108 1535
rect 174 1516 208 1535
rect 193 1473 208 1516
rect 4 1467 62 1473
rect 4 1433 16 1467
rect 4 1427 62 1433
rect 4 1159 62 1165
rect 4 1129 16 1159
rect 41 1152 66 1159
rect 174 1152 208 1473
rect 227 1482 262 1516
rect 542 1499 577 1516
rect 672 1499 681 1549
rect 3217 1499 3230 1551
rect 3234 1499 3235 1551
rect 542 1482 613 1499
rect 227 1152 261 1482
rect 543 1463 613 1482
rect 684 1471 718 1497
rect 772 1471 806 1497
rect 860 1471 884 1497
rect 560 1429 631 1463
rect 672 1459 906 1463
rect 730 1440 760 1459
rect 818 1440 848 1459
rect 719 1429 771 1440
rect 807 1429 859 1440
rect 911 1429 946 1463
rect 373 1414 431 1420
rect 373 1380 385 1414
rect 373 1374 431 1380
rect 560 1222 630 1429
rect 714 1390 720 1395
rect 818 1390 846 1419
rect 912 1410 946 1429
rect 1110 1418 1144 1444
rect 1226 1418 1253 1444
rect 1281 1411 1314 1436
rect 1351 1411 1448 1461
rect 1281 1410 1448 1411
rect 931 1390 946 1410
rect 636 1252 946 1390
rect 965 1376 1000 1410
rect 1010 1406 1156 1410
rect 1214 1406 1448 1410
rect 1603 1406 1749 1461
rect 1964 1406 2110 1408
rect 1068 1387 1098 1406
rect 1272 1393 1315 1406
rect 1272 1387 1351 1393
rect 1057 1376 1109 1387
rect 1261 1376 1351 1387
rect 965 1252 999 1376
rect 1068 1324 1098 1366
rect 1281 1357 1351 1376
rect 1491 1363 1558 1391
rect 3217 1372 3252 1499
rect 3253 1372 3287 1551
rect 3361 1461 3368 1551
rect 3371 1543 3485 1551
rect 3422 1537 3483 1543
rect 3333 1439 3368 1461
rect 3371 1452 3374 1515
rect 3388 1503 3483 1537
rect 3395 1486 3402 1503
rect 3399 1480 3402 1486
rect 3410 1486 3479 1503
rect 3410 1470 3461 1486
rect 3413 1461 3443 1470
rect 3510 1467 3523 1477
rect 3504 1465 3523 1467
rect 3388 1439 3401 1443
rect 3413 1439 3456 1461
rect 3476 1439 3489 1443
rect 3333 1427 3501 1439
rect 3355 1417 3501 1427
rect 3334 1383 3501 1417
rect 3355 1372 3501 1383
rect 3504 1383 3527 1465
rect 3504 1372 3523 1383
rect 3535 1372 3544 1551
rect 3569 1372 3603 1551
rect 3622 1372 3644 1551
rect 3698 1535 3844 1551
rect 3876 1535 3881 1578
rect 3972 1569 4008 1605
rect 3945 1558 4008 1569
rect 3956 1552 4008 1558
rect 4158 1552 4178 1578
rect 3956 1550 4377 1552
rect 3898 1535 3972 1550
rect 3698 1462 3710 1535
rect 3844 1507 3912 1535
rect 3938 1507 3972 1535
rect 3998 1516 4006 1550
rect 4044 1516 4150 1550
rect 4158 1516 4178 1550
rect 4198 1516 4232 1538
rect 4332 1516 4377 1550
rect 3844 1505 3972 1507
rect 3742 1501 3744 1505
rect 3730 1462 3744 1501
rect 3798 1491 3972 1505
rect 3796 1483 3972 1491
rect 3786 1473 3972 1483
rect 3991 1482 4044 1516
rect 4087 1499 4341 1516
rect 4436 1499 4445 1549
rect 4087 1482 4377 1499
rect 3786 1472 3978 1473
rect 3786 1467 3912 1472
rect 3764 1462 3778 1467
rect 3780 1462 3912 1467
rect 3698 1461 3912 1462
rect 3938 1461 3972 1472
rect 3991 1461 4025 1482
rect 4044 1461 4112 1482
rect 3730 1457 3744 1461
rect 3764 1433 3778 1461
rect 3780 1435 3836 1461
rect 3786 1433 3836 1435
rect 3876 1433 3881 1461
rect 3898 1460 4112 1461
rect 3217 1371 3644 1372
rect 3741 1371 3782 1386
rect 1281 1352 1592 1357
rect 1107 1264 1140 1324
rect 1281 1323 1369 1352
rect 1457 1329 1592 1352
rect 1649 1323 1684 1357
rect 1107 1258 1141 1264
rect 636 1222 999 1252
rect 1125 1236 1141 1258
rect 560 1210 999 1222
rect 1067 1221 1113 1236
rect 1067 1210 1098 1221
rect 1133 1210 1141 1236
rect 1161 1210 1169 1236
rect 329 1153 387 1206
rect 417 1183 475 1206
rect 395 1153 475 1183
rect 560 1202 1192 1210
rect 1281 1202 1368 1323
rect 1434 1280 1584 1310
rect 1492 1221 1556 1255
rect 1522 1212 1556 1221
rect 1506 1202 1573 1212
rect 395 1152 429 1153
rect -254 1125 43 1129
rect 45 1125 66 1152
rect -254 1119 62 1125
rect -254 1057 43 1119
rect 79 1091 100 1152
rect 174 1128 429 1152
rect 174 1119 333 1128
rect 175 1118 333 1119
rect 335 1118 429 1128
rect 193 1084 208 1118
rect -254 1056 112 1057
rect -254 1040 113 1056
rect -178 1023 113 1040
rect 187 1023 208 1084
rect 227 1056 261 1118
rect 395 1117 429 1118
rect 560 1117 1368 1202
rect 1414 1144 1433 1202
rect 1505 1199 1604 1202
rect 1505 1186 1573 1199
rect 1448 1174 1470 1178
rect 1442 1162 1470 1174
rect 1472 1174 1482 1178
rect 1536 1174 1570 1178
rect 1472 1162 1488 1174
rect 1524 1169 1582 1174
rect 1414 1128 1436 1144
rect 1442 1140 1474 1162
rect 1530 1158 1576 1169
rect 395 1112 1368 1117
rect 373 1106 1368 1112
rect 369 1084 1368 1106
rect 373 1072 385 1084
rect 395 1072 1368 1084
rect 373 1066 1368 1072
rect 225 1050 283 1056
rect 221 1038 261 1050
rect -178 987 43 1023
rect 79 702 113 1023
rect 221 1016 287 1038
rect 225 1010 283 1016
rect 395 1011 1368 1066
rect 1410 1011 1436 1128
rect 1448 1049 1474 1140
rect 1479 1049 1482 1129
rect 1518 1095 1524 1106
rect 1536 1095 1570 1158
rect 1650 1107 1684 1323
rect 1703 1300 2053 1304
rect 1703 1270 1718 1300
rect 1727 1293 2053 1300
rect 1738 1287 2053 1293
rect 1738 1281 2089 1287
rect 1727 1280 2089 1281
rect 1727 1270 1826 1280
rect 2018 1270 2089 1280
rect 2214 1279 2476 1304
rect 2495 1287 2530 1304
rect 2495 1279 2566 1287
rect 2214 1270 2566 1279
rect 1703 1232 1737 1270
rect 1738 1266 1775 1270
rect 2019 1258 2089 1270
rect 2496 1261 2566 1270
rect 2272 1258 2566 1261
rect 2019 1251 2566 1258
rect 2036 1247 2584 1251
rect 2694 1247 2803 1251
rect 2036 1240 2803 1247
rect 2863 1240 2899 1251
rect 2036 1234 2792 1240
rect 2794 1234 2803 1240
rect 1703 1164 1718 1232
rect 2036 1228 2827 1234
rect 2874 1228 2899 1240
rect 3217 1234 3252 1371
rect 1726 1164 1737 1175
rect 1821 1164 1845 1182
rect 1650 1095 1697 1107
rect 1513 1061 1516 1095
rect 1529 1061 1701 1095
rect 1523 1049 1524 1050
rect 1448 1020 1494 1049
rect 1524 1048 1525 1049
rect 1442 1011 1494 1020
rect 1524 1019 1525 1020
rect 1523 1018 1524 1019
rect 1518 1011 1524 1018
rect 1536 1011 1570 1061
rect 1650 1049 1697 1061
rect 1650 1019 1684 1049
rect 227 1004 261 1010
rect 395 1007 1572 1011
rect 1650 1007 1697 1019
rect 395 1004 1701 1007
rect 193 973 1701 1004
rect 227 970 1573 973
rect 227 945 239 969
rect 269 945 327 969
rect 395 961 1573 970
rect 1637 961 1697 973
rect 395 958 1572 961
rect 1650 958 1684 961
rect 1703 958 1737 1164
rect 1894 1162 1907 1208
rect 1863 1149 1893 1152
rect 1783 1121 1805 1149
rect 1863 1134 1894 1149
rect 1922 1134 1935 1222
rect 2036 1217 2899 1228
rect 2036 1181 2827 1217
rect 2831 1181 2862 1217
rect 2865 1181 2899 1217
rect 2916 1198 2933 1232
rect 3219 1198 3250 1225
rect 3253 1198 3287 1371
rect 3380 1274 3410 1371
rect 3422 1367 3435 1371
rect 3367 1271 3413 1274
rect 3365 1259 3413 1271
rect 3422 1259 3435 1343
rect 3468 1279 3498 1371
rect 3510 1343 3523 1371
rect 3535 1367 3544 1371
rect 3569 1352 3586 1371
rect 3588 1352 3603 1367
rect 3468 1274 3501 1279
rect 3455 1271 3501 1274
rect 3453 1259 3501 1271
rect 3569 1264 3603 1352
rect 3622 1280 3656 1371
rect 3724 1352 3739 1367
rect 3756 1352 3782 1371
rect 3724 1322 3782 1352
rect 3724 1307 3739 1322
rect 3413 1228 3443 1259
rect 3468 1229 3503 1259
rect 3539 1230 3555 1264
rect 3569 1230 3606 1264
rect 2916 1191 3287 1198
rect 2916 1181 3250 1191
rect 2036 1175 3250 1181
rect 3276 1180 3287 1191
rect 3411 1179 3445 1183
rect 3395 1178 3461 1179
rect 2036 1172 3214 1175
rect 1980 1160 2005 1172
rect 1821 1121 1943 1134
rect 1976 1126 2005 1160
rect 1783 1119 1863 1121
rect 1783 1073 1805 1119
rect 1806 1106 1863 1119
rect 1811 1084 1863 1106
rect 1866 1114 1894 1121
rect 1899 1114 1922 1121
rect 1936 1114 1951 1121
rect 1980 1114 2005 1126
rect 2019 1164 3214 1172
rect 3468 1170 3498 1229
rect 3569 1170 3603 1230
rect 3622 1214 3640 1280
rect 3756 1221 3782 1322
rect 3852 1284 3864 1386
rect 3880 1312 3892 1366
rect 3622 1172 3656 1214
rect 3741 1206 3782 1221
rect 3938 1275 3972 1460
rect 3991 1275 4006 1460
rect 4098 1387 4099 1460
rect 4130 1452 4150 1482
rect 4111 1430 4150 1452
rect 4158 1448 4178 1482
rect 4198 1452 4232 1482
rect 4306 1463 4377 1482
rect 4448 1471 4482 1497
rect 4536 1471 4570 1497
rect 4624 1471 4648 1497
rect 4307 1454 4395 1463
rect 4436 1459 4670 1463
rect 4183 1448 4232 1452
rect 4111 1420 4156 1430
rect 4158 1422 4232 1448
rect 4183 1420 4232 1422
rect 4273 1429 4395 1454
rect 4494 1440 4524 1459
rect 4582 1440 4612 1459
rect 4483 1429 4535 1440
rect 4571 1429 4623 1440
rect 4675 1429 4710 1463
rect 4273 1420 4394 1429
rect 4111 1387 4232 1420
rect 4307 1416 4394 1420
rect 4098 1382 4274 1387
rect 4286 1382 4394 1416
rect 4478 1390 4484 1395
rect 4582 1390 4610 1419
rect 4676 1410 4710 1429
rect 4874 1418 4908 1444
rect 4990 1418 5017 1444
rect 5045 1411 5078 1436
rect 5115 1411 5212 1461
rect 5045 1410 5212 1411
rect 4695 1390 4710 1410
rect 4098 1380 4293 1382
rect 4098 1371 4181 1380
rect 4186 1371 4293 1380
rect 4307 1371 4394 1382
rect 4098 1370 4394 1371
rect 4110 1366 4151 1370
rect 4198 1366 4232 1370
rect 4133 1364 4151 1366
rect 4105 1333 4139 1337
rect 4193 1333 4227 1337
rect 4105 1332 4151 1333
rect 4121 1321 4151 1332
rect 3938 1263 4006 1275
rect 4113 1310 4151 1321
rect 4181 1310 4239 1333
rect 4113 1276 4239 1310
rect 4014 1263 4025 1274
rect 3938 1241 4025 1263
rect 4113 1254 4151 1276
rect 4181 1261 4223 1276
rect 3622 1170 3640 1172
rect 3740 1170 3744 1193
rect 2019 1128 3196 1164
rect 3330 1145 3752 1170
rect 3322 1144 3752 1145
rect 3234 1133 3245 1144
rect 3321 1133 3752 1144
rect 3234 1128 3752 1133
rect 3768 1159 3826 1165
rect 3768 1128 3780 1159
rect 3805 1152 3830 1159
rect 3938 1152 3972 1241
rect 3986 1207 4025 1241
rect 4036 1207 4059 1241
rect 4113 1238 4139 1254
rect 3991 1152 4025 1207
rect 4181 1206 4186 1261
rect 4193 1256 4223 1261
rect 4229 1256 4239 1276
rect 4193 1238 4239 1256
rect 4324 1247 4394 1370
rect 4209 1223 4239 1238
rect 4244 1223 4261 1226
rect 4209 1209 4261 1223
rect 4307 1222 4394 1247
rect 4400 1252 4710 1390
rect 4729 1376 4764 1410
rect 4774 1406 4920 1410
rect 4978 1406 5212 1410
rect 5367 1406 5513 1461
rect 5728 1406 5874 1408
rect 4832 1387 4862 1406
rect 5036 1393 5079 1406
rect 5036 1387 5115 1393
rect 4821 1376 4873 1387
rect 5025 1376 5115 1387
rect 4729 1252 4763 1376
rect 4832 1324 4862 1366
rect 5045 1357 5115 1376
rect 5255 1363 5322 1391
rect 5045 1352 5356 1357
rect 4871 1264 4904 1324
rect 5045 1323 5133 1352
rect 5221 1329 5356 1352
rect 5413 1323 5448 1357
rect 4871 1258 4905 1264
rect 4400 1222 4763 1252
rect 4889 1236 4905 1258
rect 4307 1210 4763 1222
rect 4831 1221 4877 1236
rect 4831 1210 4862 1221
rect 4897 1210 4905 1236
rect 4925 1210 4933 1236
rect 4209 1206 4286 1209
rect 4093 1153 4151 1206
rect 4181 1183 4286 1206
rect 4159 1175 4286 1183
rect 4307 1202 4956 1210
rect 5045 1202 5132 1323
rect 5198 1280 5348 1310
rect 5256 1221 5320 1255
rect 5286 1212 5320 1221
rect 5270 1202 5337 1212
rect 4307 1175 5132 1202
rect 4159 1163 4261 1175
rect 4159 1153 4239 1163
rect 4244 1160 4261 1163
rect 4307 1160 4310 1175
rect 4159 1152 4193 1153
rect 3809 1139 3830 1152
rect 3786 1128 3830 1139
rect 3843 1128 3864 1152
rect 3938 1146 4193 1152
rect 4209 1149 4227 1153
rect 4307 1149 4318 1160
rect 3877 1130 4193 1146
rect 3877 1128 4261 1130
rect 2019 1125 4261 1128
rect 2019 1118 4193 1125
rect 2019 1117 4042 1118
rect 4159 1117 4193 1118
rect 4324 1117 5132 1175
rect 5178 1144 5197 1202
rect 5269 1199 5368 1202
rect 5269 1186 5337 1199
rect 5212 1174 5234 1178
rect 5206 1162 5234 1174
rect 5236 1174 5246 1178
rect 5300 1174 5334 1178
rect 5236 1162 5252 1174
rect 5288 1169 5346 1174
rect 5178 1128 5200 1144
rect 5206 1140 5238 1162
rect 5294 1158 5340 1169
rect 1866 1084 1951 1114
rect 2019 1106 4121 1117
rect 4159 1106 5132 1117
rect 1811 1073 1833 1084
rect 1838 1073 1857 1084
rect 1783 1043 1864 1073
rect 1805 992 1864 1043
rect 1866 1026 1894 1084
rect 1899 1026 1922 1084
rect 1936 1069 1951 1084
rect 1980 1072 2005 1084
rect 1936 1026 1951 1041
rect 1976 1038 2005 1072
rect 1980 1026 2005 1038
rect 1866 996 1951 1026
rect 2019 1011 5132 1106
rect 5174 1011 5200 1128
rect 5212 1049 5238 1140
rect 5243 1049 5246 1129
rect 5282 1095 5288 1106
rect 5300 1095 5334 1158
rect 5414 1107 5448 1323
rect 5467 1300 5817 1304
rect 5467 1270 5482 1300
rect 5491 1293 5817 1300
rect 5502 1287 5817 1293
rect 5502 1281 5853 1287
rect 5491 1280 5853 1281
rect 5491 1270 5590 1280
rect 5782 1270 5853 1280
rect 5467 1232 5501 1270
rect 5502 1266 5539 1270
rect 5783 1258 5853 1270
rect 6036 1258 6222 1261
rect 5783 1251 6222 1258
rect 5800 1234 6222 1251
rect 5467 1164 5482 1232
rect 5490 1164 5501 1175
rect 5585 1164 5609 1182
rect 5414 1095 5461 1107
rect 5277 1061 5280 1095
rect 5293 1061 5465 1095
rect 5287 1049 5288 1050
rect 5212 1020 5258 1049
rect 5288 1048 5289 1049
rect 5206 1011 5258 1020
rect 5288 1019 5289 1020
rect 5287 1018 5288 1019
rect 5282 1011 5288 1018
rect 5300 1011 5334 1061
rect 5414 1049 5461 1061
rect 5414 1019 5448 1049
rect 2019 1007 5336 1011
rect 5414 1007 5461 1019
rect 1805 976 1857 992
rect 1866 990 1894 996
rect 1899 990 1922 996
rect 1805 958 1863 976
rect 1866 962 1885 990
rect 1936 981 1951 996
rect 1980 984 2005 996
rect 1893 958 1951 976
rect 395 941 1951 958
rect 1976 950 2005 984
rect 1980 941 2005 950
rect 2019 973 5465 1007
rect 2019 961 5337 973
rect 5401 961 5461 973
rect 2019 958 5336 961
rect 5414 958 5448 961
rect 5467 958 5501 1164
rect 5658 1162 5671 1208
rect 5627 1149 5657 1152
rect 5547 1121 5569 1149
rect 5627 1134 5658 1149
rect 5686 1134 5699 1222
rect 5800 1181 6591 1234
rect 5800 1172 6762 1181
rect 5744 1160 5769 1172
rect 5585 1121 5707 1134
rect 5740 1126 5769 1160
rect 5547 1119 5627 1121
rect 5547 1073 5569 1119
rect 5570 1106 5627 1119
rect 5575 1084 5627 1106
rect 5630 1114 5658 1121
rect 5663 1114 5686 1121
rect 5700 1114 5715 1121
rect 5744 1114 5769 1126
rect 5783 1137 6762 1172
rect 6827 1137 6879 1145
rect 6889 1137 6924 1145
rect 5783 1128 6960 1137
rect 7094 1128 7516 1137
rect 5783 1117 7516 1128
rect 5630 1084 5715 1114
rect 5575 1073 5597 1084
rect 5602 1073 5621 1084
rect 5547 1043 5628 1073
rect 5569 992 5628 1043
rect 5630 1026 5658 1084
rect 5663 1026 5686 1084
rect 5700 1069 5715 1084
rect 5744 1072 5769 1084
rect 5700 1026 5715 1041
rect 5740 1038 5769 1072
rect 5744 1026 5769 1038
rect 5630 996 5715 1026
rect 5569 976 5621 992
rect 5630 990 5658 996
rect 5663 990 5686 996
rect 5569 958 5627 976
rect 5630 962 5649 990
rect 5700 981 5715 996
rect 5744 984 5769 996
rect 5657 958 5715 976
rect 2019 941 5715 958
rect 5740 950 5769 984
rect 5744 941 5769 950
rect 395 934 1941 941
rect 395 875 482 934
rect 553 887 1941 934
rect 2019 887 5705 941
rect 5783 887 7741 1117
rect 7832 1081 7885 1082
rect 7814 1047 7885 1081
rect 7815 1046 7885 1047
rect 553 875 7741 887
rect 395 866 7741 875
rect 395 844 1945 866
rect 1958 854 5709 866
rect 1958 853 2019 854
rect 2020 853 5709 854
rect 5722 854 7741 866
rect 5722 853 5783 854
rect 5784 853 7741 854
rect 2036 844 5709 853
rect 395 840 1958 844
rect 2036 840 5722 844
rect 181 805 327 839
rect 395 826 1945 840
rect 395 805 1941 826
rect 1958 805 2019 840
rect 2036 826 5709 840
rect 2036 819 5705 826
rect 2032 805 5705 819
rect 5722 805 5783 840
rect 5800 819 7741 853
rect 159 761 179 799
rect 181 791 221 804
rect 181 789 236 791
rect 199 785 227 788
rect 239 772 263 805
rect 315 801 327 804
rect 279 789 327 801
rect 237 754 301 772
rect 339 761 349 799
rect 395 792 1958 805
rect 2032 792 5722 805
rect 395 791 1957 792
rect 1958 791 2019 792
rect 395 779 2019 791
rect 2032 791 5721 792
rect 5722 791 5783 792
rect 2032 779 5783 791
rect 5796 779 7741 819
rect 395 770 7741 779
rect 7832 1012 7903 1046
rect 8183 1012 8218 1046
rect 395 758 7731 770
rect 145 750 147 754
rect 233 751 301 754
rect 237 750 301 751
rect 108 640 113 702
rect 133 640 167 750
rect 190 742 301 750
rect 221 708 301 742
rect 221 692 279 708
rect 264 677 279 692
rect 361 674 379 754
rect 345 640 379 674
rect 395 640 1958 758
rect 1972 704 1997 707
rect 2036 704 5722 758
rect 5736 704 5761 707
rect 5800 704 7731 758
rect 133 606 279 640
rect 333 606 1958 640
rect 233 566 267 606
rect 412 517 1958 606
rect 2026 687 5722 704
rect 2026 649 2051 687
rect 2092 655 2111 683
rect 2055 649 2078 655
rect 2083 649 2111 655
rect 2113 653 2172 687
rect 2240 684 2274 687
rect 2293 684 2327 687
rect 2242 680 2274 684
rect 2120 649 2172 653
rect 2026 619 2111 649
rect 2114 619 2172 649
rect 2181 619 2194 653
rect 2026 561 2051 619
rect 2055 561 2078 619
rect 2083 561 2111 619
rect 2120 603 2172 619
rect 2120 561 2139 603
rect 2157 602 2172 603
rect 2144 588 2194 602
rect 2144 561 2166 588
rect 2026 531 2111 561
rect 2026 524 2051 531
rect 2055 524 2078 531
rect 2083 524 2111 531
rect 781 508 1958 517
rect 2034 511 2111 524
rect 817 500 914 508
rect 979 464 1958 508
rect 1150 411 1958 464
rect 2042 423 2055 511
rect 2083 496 2111 511
rect 2114 539 2166 561
rect 2114 526 2171 539
rect 2172 526 2194 588
rect 2114 524 2194 526
rect 2114 493 2156 524
rect 2172 496 2194 524
rect 2070 437 2083 483
rect 2240 481 2274 680
rect 2280 672 2328 684
rect 2405 672 5722 687
rect 2276 638 5722 672
rect 2280 626 2328 638
rect 2405 634 5722 638
rect 2293 596 2327 626
rect 2280 584 2328 596
rect 2407 584 2441 634
rect 2453 626 2454 627
rect 2484 626 2535 634
rect 2452 625 2453 626
rect 2483 625 2535 626
rect 2452 596 2453 597
rect 2483 596 2529 625
rect 2453 595 2454 596
rect 2276 550 2448 584
rect 2453 550 2459 595
rect 2461 550 2464 584
rect 2280 538 2328 550
rect 2240 470 2251 481
rect 2259 417 2274 481
rect 1519 394 1958 411
rect 1519 387 1941 394
rect 1519 384 1705 387
rect 1888 365 1941 387
rect 2206 375 2239 379
rect 2240 375 2274 417
rect 2161 365 2274 375
rect 1888 358 2274 365
rect 1924 345 2274 358
rect 1924 341 2250 345
rect 2259 341 2274 345
rect 2293 511 2327 538
rect 2293 481 2316 511
rect 2407 498 2441 550
rect 2495 516 2498 596
rect 2503 505 2529 596
rect 2541 517 2567 634
rect 2609 539 5722 634
rect 2609 528 3582 539
rect 3620 528 5722 539
rect 2395 483 2495 498
rect 2503 483 2535 505
rect 2541 501 2563 517
rect 2293 324 2327 481
rect 2395 471 2505 483
rect 2407 467 2441 471
rect 2495 467 2505 471
rect 2507 471 2535 483
rect 2507 467 2529 471
rect 2404 451 2472 459
rect 2404 446 2485 451
rect 2373 443 2485 446
rect 2544 443 2563 501
rect 2609 505 3434 528
rect 3548 527 3582 528
rect 3699 527 5722 528
rect 3514 520 5722 527
rect 5790 687 7731 704
rect 5790 649 5815 687
rect 5856 655 5875 683
rect 5819 649 5842 655
rect 5847 649 5875 655
rect 5877 653 5936 687
rect 6004 684 6038 687
rect 6057 684 6091 687
rect 6006 680 6038 684
rect 5884 649 5936 653
rect 5790 619 5875 649
rect 5878 619 5936 649
rect 5945 619 5958 653
rect 5790 561 5815 619
rect 5819 561 5842 619
rect 5847 561 5875 619
rect 5884 603 5936 619
rect 5884 561 5903 603
rect 5921 602 5936 603
rect 5908 588 5958 602
rect 5908 561 5930 588
rect 5790 531 5875 561
rect 5790 524 5815 531
rect 5819 524 5842 531
rect 5847 524 5875 531
rect 3480 517 5722 520
rect 3480 515 3803 517
rect 2609 479 2617 505
rect 2626 479 3434 505
rect 3514 496 3803 515
rect 3514 492 3532 496
rect 3548 493 3803 496
rect 3877 493 3898 517
rect 3911 493 3936 517
rect 3502 487 3560 492
rect 2609 443 3434 479
rect 3480 482 3497 485
rect 3502 482 3532 487
rect 3480 470 3532 482
rect 3540 477 3560 487
rect 2404 433 2485 443
rect 2421 417 2485 433
rect 2451 407 2485 417
rect 2435 374 2501 407
rect 2609 335 2696 443
rect 2785 435 3434 443
rect 3476 436 3532 470
rect 3548 468 3560 477
rect 3590 468 3648 492
rect 3716 472 3750 493
rect 3769 472 3803 493
rect 3911 486 3932 493
rect 3969 486 3973 517
rect 3915 480 3973 486
rect 3989 512 4507 517
rect 3989 501 4420 512
rect 4496 501 4507 512
rect 3989 475 4411 501
rect 4470 481 4507 492
rect 4545 481 5722 517
rect 5798 511 5875 524
rect 2808 409 2816 435
rect 2836 381 2844 435
rect 2879 424 2910 435
rect 2864 409 2910 424
rect 2609 324 2620 335
rect 2293 307 2316 324
rect 2397 316 2507 320
rect 2385 307 2520 316
rect 2626 307 2696 335
rect 2879 321 2909 409
rect 2978 393 3021 435
rect 3031 423 3434 435
rect 2978 382 2989 393
rect 1888 305 2081 307
rect 2160 305 2696 307
rect 2257 288 2696 305
rect 2257 282 2442 288
rect 2461 282 2696 288
rect 2257 269 2696 282
rect 2257 258 2716 269
rect 2868 261 2920 269
rect 2257 254 2705 258
rect 2257 252 2442 254
rect 2461 252 2705 254
rect 2629 243 2705 252
rect 2662 239 2705 243
rect 2758 239 2785 261
rect 2662 235 2785 239
rect 2799 258 2920 261
rect 2799 239 2916 258
rect 2799 235 2967 239
rect 2997 235 3012 393
rect 3031 255 3341 423
rect 3347 317 3359 423
rect 3364 343 3434 423
rect 3480 422 3532 436
rect 3480 419 3497 422
rect 3502 407 3532 422
rect 3502 391 3548 407
rect 3502 343 3512 391
rect 3518 384 3548 391
rect 3555 384 3560 468
rect 3518 369 3560 384
rect 3590 369 3637 416
rect 3716 404 3803 472
rect 3997 452 4001 475
rect 4101 455 4119 475
rect 4104 449 4119 455
rect 4138 449 4172 475
rect 3716 382 3750 404
rect 3716 371 3727 382
rect 3518 343 3637 369
rect 3364 335 3711 343
rect 3364 312 3585 335
rect 3364 308 3548 312
rect 3364 279 3542 308
rect 3364 275 3543 279
rect 3555 275 3585 312
rect 3590 311 3711 335
rect 3602 308 3711 311
rect 3608 279 3711 308
rect 3597 275 3711 279
rect 3364 263 3435 275
rect 3509 274 3555 275
rect 3527 263 3555 274
rect 3585 274 3631 275
rect 3585 265 3630 274
rect 3031 235 3065 255
rect 3257 250 3263 255
rect 3031 201 3046 235
rect 3364 225 3468 263
rect 3509 251 3555 263
rect 3558 253 3630 265
rect 3643 253 3711 275
rect 3735 253 3750 382
rect 3769 253 3803 404
rect 3959 424 4000 439
rect 3849 279 3861 333
rect 3877 259 3889 361
rect 3959 323 3985 424
rect 4101 415 4172 449
rect 4280 467 4315 475
rect 4280 466 4346 467
rect 4280 417 4315 466
rect 4454 454 4465 465
rect 4470 464 5722 481
rect 4470 458 4580 464
rect 4637 458 4667 464
rect 4470 454 4590 458
rect 4454 447 4590 454
rect 4626 447 4678 458
rect 4779 447 4825 464
rect 4101 347 4119 415
rect 4135 381 4172 415
rect 4186 381 4206 415
rect 4298 414 4315 417
rect 4298 386 4319 414
rect 4331 386 4361 417
rect 4104 342 4119 347
rect 4138 342 4172 381
rect 4240 374 4288 386
rect 4240 371 4286 374
rect 4240 366 4273 371
rect 4002 323 4017 338
rect 3959 293 4017 323
rect 4085 323 4096 334
rect 4104 323 4240 342
rect 4085 296 4240 323
rect 3959 274 3985 293
rect 4002 278 4017 293
rect 4075 274 4240 296
rect 4243 274 4273 366
rect 4306 302 4319 386
rect 4328 374 4376 386
rect 4328 371 4374 374
rect 4306 274 4319 278
rect 4331 274 4361 371
rect 4454 342 4488 447
rect 4491 420 4522 447
rect 4808 413 4825 447
rect 4842 428 4876 464
rect 4879 462 4910 464
rect 4879 429 4913 462
rect 4879 428 4910 429
rect 4914 428 5722 464
rect 4842 417 5722 428
rect 5806 423 5819 511
rect 5847 496 5875 511
rect 5878 539 5930 561
rect 5878 526 5935 539
rect 5936 526 5958 588
rect 5878 524 5958 526
rect 5878 493 5920 524
rect 5936 496 5958 524
rect 5834 437 5847 483
rect 6004 481 6038 680
rect 6044 672 6092 684
rect 6169 672 7731 687
rect 6040 658 7731 672
rect 7832 658 7902 1012
rect 8184 993 8218 1012
rect 8014 944 8072 950
rect 8014 910 8026 944
rect 8014 904 8072 910
rect 6040 638 7902 658
rect 6044 626 6092 638
rect 6169 634 7902 638
rect 6057 596 6091 626
rect 6044 584 6092 596
rect 6171 584 6205 634
rect 6217 626 6218 627
rect 6248 626 6299 634
rect 6216 625 6217 626
rect 6247 625 6299 626
rect 6216 596 6217 597
rect 6247 596 6293 625
rect 6217 595 6218 596
rect 6040 550 6212 584
rect 6217 550 6223 595
rect 6225 550 6228 584
rect 6044 538 6092 550
rect 6004 470 6015 481
rect 6023 417 6038 481
rect 4743 355 4778 411
rect 4842 405 4867 417
rect 4914 411 5722 417
rect 4949 405 4979 411
rect 4842 394 4878 405
rect 4938 394 4990 405
rect 5009 398 5158 411
rect 5175 394 5722 411
rect 5175 387 5705 394
rect 5175 384 5469 387
rect 5175 358 5228 384
rect 5285 360 5527 375
rect 5652 365 5705 387
rect 5970 375 6003 379
rect 6004 375 6038 417
rect 5925 365 6038 375
rect 5433 352 5463 360
rect 5652 358 6038 365
rect 4386 328 4524 342
rect 5422 341 5474 352
rect 5688 345 6038 358
rect 5688 341 6014 345
rect 6023 341 6038 345
rect 6057 511 6091 538
rect 6057 481 6080 511
rect 6171 498 6205 550
rect 6259 516 6262 596
rect 6267 505 6293 596
rect 6305 517 6331 634
rect 6373 622 7902 634
rect 8014 636 8072 642
rect 6373 570 7885 622
rect 8014 607 8026 636
rect 8014 603 8060 607
rect 8010 602 8076 603
rect 8014 596 8072 602
rect 6373 539 7399 570
rect 6373 528 7346 539
rect 6159 483 6259 498
rect 6267 483 6299 505
rect 6305 501 6327 517
rect 4365 274 4524 328
rect 6057 324 6091 481
rect 6159 471 6269 483
rect 6171 467 6205 471
rect 6259 467 6269 471
rect 6271 471 6299 483
rect 6271 467 6293 471
rect 6168 451 6236 459
rect 6168 446 6249 451
rect 6137 443 6249 446
rect 6308 443 6327 501
rect 6373 505 7198 528
rect 7312 527 7346 528
rect 7463 527 7885 570
rect 8203 569 8218 993
rect 8237 959 8272 993
rect 8552 959 8587 993
rect 8237 569 8271 959
rect 8553 940 8587 959
rect 8383 891 8441 897
rect 8383 857 8395 891
rect 8383 851 8441 857
rect 8383 583 8441 589
rect 7936 535 8184 569
rect 8383 549 8395 583
rect 8383 543 8441 549
rect 7278 520 7885 527
rect 7244 517 7885 520
rect 7244 515 7567 517
rect 6373 479 6381 505
rect 6390 479 7198 505
rect 7278 496 7567 515
rect 7278 492 7296 496
rect 7312 493 7567 496
rect 7641 493 7662 517
rect 7675 493 7700 517
rect 7266 487 7324 492
rect 6373 443 7198 479
rect 7244 482 7261 485
rect 7266 482 7296 487
rect 7244 470 7296 482
rect 7304 477 7324 487
rect 6168 433 6249 443
rect 6185 417 6249 433
rect 6215 407 6249 417
rect 6199 374 6265 407
rect 6373 335 6460 443
rect 6549 435 7198 443
rect 7240 436 7296 470
rect 7312 468 7324 477
rect 7354 468 7412 492
rect 7480 472 7514 493
rect 7533 472 7567 493
rect 7675 486 7696 493
rect 6572 409 6580 435
rect 6600 381 6608 435
rect 6643 424 6674 435
rect 6628 409 6674 424
rect 6373 324 6384 335
rect 6057 307 6080 324
rect 6161 316 6271 320
rect 6149 307 6284 316
rect 6390 307 6460 335
rect 6643 321 6673 409
rect 6742 393 6785 435
rect 6795 423 7198 435
rect 6742 382 6753 393
rect 5652 305 5845 307
rect 5924 305 6460 307
rect 3959 259 4000 274
rect 4075 262 4119 274
rect 4138 262 4177 274
rect 3558 251 3716 253
rect 3509 225 3716 251
rect 3118 208 3170 216
rect 3206 208 3258 216
rect 3118 205 3285 208
rect 3127 186 3285 205
rect 3071 182 3305 186
rect 3364 182 3435 225
rect 3509 223 3555 225
rect 3509 215 3583 223
rect 3585 215 3716 225
rect 3364 163 3434 182
rect 3509 163 3543 215
rect 3549 197 3583 215
rect 3563 163 3583 197
rect 3591 185 3716 215
rect 3735 212 3911 253
rect 4097 252 4177 262
rect 3735 210 3955 212
rect 3961 210 4177 252
rect 3735 185 4177 210
rect 3591 163 3631 185
rect 3643 163 3711 185
rect 3716 163 3750 185
rect 3763 173 3803 185
rect 3829 184 4177 185
rect 3832 173 3837 184
rect 3364 146 3643 163
rect 3364 96 3373 146
rect 3409 129 3643 146
rect 3654 129 3665 163
rect 3697 129 3750 163
rect 3769 172 3837 173
rect 3409 96 3410 129
rect 3509 107 3543 129
rect 3563 96 3583 129
rect 3591 96 3611 129
rect 3643 96 3711 129
rect 3735 96 3743 129
rect 3769 110 3803 172
rect 3832 110 3837 172
rect 3843 178 4011 184
rect 3843 162 3955 178
rect 3843 110 3943 162
rect 3997 144 4011 178
rect 4043 172 4177 184
rect 4043 144 4119 172
rect 3997 110 4119 144
rect 3769 96 3843 110
rect 3409 95 3843 96
rect 3563 67 3583 95
rect 3735 91 3743 95
rect 3769 94 3785 95
rect 3860 94 3865 110
rect 3897 106 4057 110
rect 3897 94 4043 106
rect 4097 95 4119 110
rect 4138 119 4177 172
rect 4138 111 4172 119
rect 4197 111 4206 274
rect 4218 262 4237 274
rect 4214 180 4237 262
rect 4240 262 4386 274
rect 4427 262 4488 274
rect 4507 262 4524 274
rect 4240 206 4407 262
rect 4252 202 4265 206
rect 4218 178 4237 180
rect 4218 168 4231 178
rect 4285 175 4328 206
rect 4340 202 4353 206
rect 4330 193 4368 197
rect 4330 175 4370 193
rect 4280 130 4370 175
rect 4373 142 4407 206
rect 4280 125 4368 130
rect 4280 119 4342 125
rect 4280 111 4331 119
rect 4373 111 4380 142
rect 4454 119 4524 262
rect 6021 288 6460 305
rect 6021 282 6206 288
rect 6225 282 6460 288
rect 6021 269 6460 282
rect 6021 258 6480 269
rect 6632 261 6684 269
rect 6021 254 6469 258
rect 6021 252 6206 254
rect 6225 252 6469 254
rect 6393 243 6469 252
rect 6426 239 6469 243
rect 6522 239 6549 261
rect 6426 235 6549 239
rect 6563 258 6684 261
rect 6563 239 6680 258
rect 6563 235 6731 239
rect 6761 235 6776 393
rect 6795 255 7105 423
rect 7111 317 7123 423
rect 7128 343 7198 423
rect 7244 422 7296 436
rect 7244 419 7261 422
rect 7266 407 7296 422
rect 7266 391 7312 407
rect 7266 343 7276 391
rect 7282 384 7312 391
rect 7319 384 7324 468
rect 7282 369 7324 384
rect 7354 369 7401 416
rect 7480 404 7567 472
rect 7480 382 7514 404
rect 7480 371 7491 382
rect 7282 343 7401 369
rect 7128 335 7475 343
rect 7128 312 7349 335
rect 7128 308 7312 312
rect 7128 279 7306 308
rect 7128 275 7307 279
rect 7319 275 7349 312
rect 7354 311 7475 335
rect 7366 308 7475 311
rect 7372 279 7475 308
rect 7361 275 7475 279
rect 7128 263 7199 275
rect 7273 274 7319 275
rect 7291 263 7319 274
rect 7349 274 7395 275
rect 7349 265 7394 274
rect 6795 235 6829 255
rect 7021 250 7027 255
rect 6795 201 6810 235
rect 7128 225 7232 263
rect 7273 251 7319 263
rect 7322 253 7394 265
rect 7407 253 7475 275
rect 7499 253 7514 382
rect 7533 253 7567 404
rect 7613 279 7625 333
rect 7641 259 7653 361
rect 7322 251 7480 253
rect 7273 225 7480 251
rect 6882 208 6934 216
rect 6970 208 7022 216
rect 6882 205 7049 208
rect 6891 186 7049 205
rect 4454 111 4488 119
rect 4138 95 4488 111
rect 4507 95 4524 119
rect 4097 94 4524 95
rect 4579 94 4592 184
rect 6835 182 7069 186
rect 7128 182 7199 225
rect 7273 223 7319 225
rect 7273 215 7347 223
rect 7349 215 7480 225
rect 7128 163 7198 182
rect 7273 163 7307 215
rect 7313 197 7347 215
rect 7327 163 7347 197
rect 7355 185 7480 215
rect 7499 185 7675 253
rect 7701 231 7703 467
rect 7729 259 7731 439
rect 7355 163 7395 185
rect 7407 163 7475 185
rect 7480 163 7514 185
rect 7527 173 7567 185
rect 7128 146 7407 163
rect 7128 96 7137 146
rect 7173 129 7407 146
rect 7418 129 7429 163
rect 7461 129 7514 163
rect 7533 172 7601 173
rect 7173 96 7174 129
rect 7273 107 7307 129
rect 7327 96 7347 129
rect 7355 96 7375 129
rect 7407 96 7475 129
rect 7499 96 7507 129
rect 7533 110 7567 172
rect 7607 110 7675 185
rect 7533 96 7607 110
rect 7173 95 7607 96
rect 3769 76 4119 94
rect 4138 76 4172 94
rect 4197 91 4206 94
rect 4256 91 4370 94
rect 4373 91 4380 94
rect 4197 90 4231 91
rect 4285 90 4319 91
rect 4373 90 4407 91
rect 3860 67 3865 76
rect 4138 66 4153 76
rect 4155 68 4172 76
rect 3733 42 4153 66
rect 4161 57 4172 68
rect 4234 57 4392 74
rect 4454 57 4460 94
rect 7327 67 7347 95
rect 7499 91 7507 95
rect 7533 94 7549 95
rect 7533 76 7749 94
rect 7868 76 7883 507
rect 7936 501 8184 534
rect 8010 500 8122 501
rect 7902 76 7936 500
rect 8048 467 8106 473
rect 8044 466 8110 467
rect 8048 433 8060 466
rect 8572 447 8587 940
rect 8606 906 8641 940
rect 8606 447 8640 906
rect 8752 838 8810 844
rect 8752 804 8764 838
rect 8922 815 8956 833
rect 8752 798 8810 804
rect 8922 779 8992 815
rect 8939 745 9010 779
rect 8752 530 8810 536
rect 8752 496 8764 530
rect 8752 490 8810 496
rect 8048 427 8106 433
rect 8606 413 8621 447
rect 8939 394 9009 745
rect 9121 677 9179 683
rect 9121 643 9133 677
rect 9121 637 9179 643
rect 9121 477 9179 483
rect 9121 443 9133 477
rect 9121 437 9179 443
rect 8939 358 8992 394
rect 8048 159 8106 165
rect 8048 125 8060 159
rect 8048 119 8106 125
rect 4163 56 4441 57
rect 3733 40 4138 42
rect 4234 40 4392 56
rect 4488 40 4524 66
rect 7497 40 7721 66
rect 7902 42 7917 76
rect 4138 23 4488 40
rect 4524 7 4550 40
rect 4102 6 4550 7
rect 43 -2483 450 -2430
rect 43 -2519 465 -2483
rect 766 -2519 834 -2518
rect 43 -2553 483 -2519
rect 529 -2553 702 -2519
rect 748 -2536 834 -2519
rect 748 -2553 1188 -2536
rect 43 -2725 482 -2553
rect 749 -2554 1188 -2553
rect 766 -2571 1188 -2554
rect 766 -2589 1203 -2571
rect 766 -2615 1557 -2589
rect 591 -2655 640 -2621
rect 749 -2624 1557 -2615
rect 749 -2642 1572 -2624
rect 749 -2677 1926 -2642
rect 535 -2725 536 -2693
rect 593 -2705 596 -2694
rect 547 -2725 596 -2705
rect 601 -2725 602 -2693
rect 629 -2694 630 -2693
rect 624 -2705 638 -2694
rect 629 -2725 630 -2705
rect 635 -2725 684 -2705
rect 749 -2713 1941 -2677
rect 749 -2725 1959 -2713
rect 28 -2747 1959 -2725
rect 2239 -2747 2274 -2713
rect 28 -2785 1958 -2747
rect 2240 -2766 2274 -2747
rect 2259 -2785 2274 -2766
rect 2293 -2785 2328 -2766
rect 28 -2800 2328 -2785
rect 28 -3030 2327 -2800
rect 2439 -2868 2497 -2862
rect 2439 -2902 2451 -2868
rect 2609 -2891 2643 -2873
rect 2439 -2908 2497 -2902
rect 2609 -2927 2679 -2891
rect 173 -3057 200 -3030
rect 207 -3033 213 -3030
rect 253 -3057 267 -3030
rect 295 -3057 301 -3030
rect 311 -3033 329 -3030
rect 345 -3034 363 -3030
rect 373 -3034 379 -3030
rect 199 -3058 233 -3057
rect 253 -3075 263 -3057
rect 267 -3058 301 -3057
rect 397 -3083 2327 -3030
rect 195 -3216 221 -3174
rect 253 -3216 263 -3109
rect 371 -3124 437 -3110
rect 366 -3127 447 -3124
rect 453 -3127 479 -3083
rect 781 -3136 2327 -3083
rect 366 -3155 453 -3152
rect 237 -3277 263 -3216
rect 388 -3196 437 -3162
rect 1150 -3189 2327 -3136
rect 2626 -2961 2697 -2927
rect 2977 -2961 3012 -2927
rect 3400 -2944 3435 -2926
rect 388 -3219 422 -3196
rect 343 -3263 366 -3219
rect 371 -3235 394 -3219
rect 453 -3235 479 -3219
rect 261 -3307 267 -3297
rect 253 -3325 267 -3307
rect 453 -3298 463 -3235
rect 1519 -3242 2327 -3189
rect 2439 -3176 2497 -3170
rect 2439 -3210 2451 -3176
rect 2439 -3216 2497 -3210
rect 1888 -3259 2327 -3242
rect 1888 -3293 2308 -3259
rect 1888 -3295 2295 -3293
rect 195 -3337 236 -3325
rect 119 -3428 153 -3337
rect 173 -3417 179 -3412
rect 195 -3416 241 -3337
rect 261 -3377 267 -3325
rect 289 -3377 295 -3325
rect 311 -3337 329 -3321
rect 307 -3354 329 -3337
rect 345 -3338 363 -3322
rect 453 -3326 467 -3298
rect 485 -3321 501 -3298
rect 526 -3321 559 -3298
rect 2626 -3312 2696 -2961
rect 2978 -2980 3012 -2961
rect 3364 -2959 3435 -2944
rect 3715 -2959 3750 -2925
rect 2808 -3029 2866 -3023
rect 2808 -3063 2820 -3029
rect 2808 -3069 2866 -3063
rect 2808 -3229 2866 -3223
rect 2808 -3263 2820 -3229
rect 2808 -3269 2866 -3263
rect 438 -3338 479 -3326
rect 345 -3354 367 -3338
rect 295 -3390 301 -3378
rect 165 -3428 179 -3417
rect 119 -3493 179 -3428
rect 145 -3494 179 -3493
rect 150 -3505 165 -3494
rect 173 -3505 179 -3494
rect 207 -3428 241 -3416
rect 261 -3417 267 -3412
rect 253 -3428 267 -3417
rect 207 -3493 267 -3428
rect 150 -3506 191 -3505
rect 173 -3510 179 -3506
rect 207 -3509 213 -3493
rect 233 -3494 267 -3493
rect 238 -3505 267 -3494
rect 295 -3493 305 -3390
rect 307 -3493 335 -3354
rect 238 -3506 279 -3505
rect 253 -3510 267 -3506
rect 295 -3509 301 -3493
rect 311 -3505 335 -3493
rect 339 -3494 367 -3354
rect 373 -3387 379 -3377
rect 373 -3389 385 -3387
rect 369 -3494 385 -3389
rect 407 -3415 413 -3411
rect 401 -3416 413 -3415
rect 433 -3415 479 -3338
rect 498 -3411 501 -3321
rect 526 -3338 561 -3326
rect 495 -3415 501 -3411
rect 396 -3424 421 -3416
rect 433 -3424 473 -3415
rect 489 -3416 501 -3415
rect 521 -3349 561 -3338
rect 2626 -3348 2679 -3312
rect 396 -3427 473 -3424
rect 484 -3424 509 -3416
rect 521 -3424 555 -3349
rect 2997 -3365 3012 -2980
rect 3031 -3014 3066 -2980
rect 3031 -3365 3065 -3014
rect 3177 -3082 3235 -3076
rect 3177 -3116 3189 -3082
rect 3177 -3122 3235 -3116
rect 3177 -3282 3235 -3276
rect 3177 -3316 3189 -3282
rect 3177 -3322 3235 -3316
rect 3031 -3399 3046 -3365
rect 484 -3427 555 -3424
rect 311 -3509 329 -3505
rect 253 -3531 263 -3510
rect 339 -3526 363 -3494
rect 373 -3498 385 -3494
rect 401 -3458 473 -3427
rect 401 -3491 441 -3458
rect 461 -3470 473 -3458
rect 489 -3458 555 -3427
rect 3364 -3418 3434 -2959
rect 3716 -2978 3750 -2959
rect 3546 -3027 3604 -3021
rect 3546 -3061 3558 -3027
rect 3546 -3067 3604 -3061
rect 3546 -3335 3604 -3329
rect 3546 -3369 3558 -3335
rect 3546 -3375 3604 -3369
rect 3364 -3454 3417 -3418
rect 401 -3493 453 -3491
rect 461 -3493 467 -3470
rect 489 -3493 529 -3458
rect 3735 -3471 3750 -2978
rect 3769 -3012 3804 -2978
rect 4084 -3012 4119 -2978
rect 3769 -3471 3803 -3012
rect 4085 -3031 4119 -3012
rect 3915 -3080 3973 -3074
rect 3915 -3114 3927 -3080
rect 3915 -3120 3973 -3114
rect 3915 -3388 3973 -3382
rect 3915 -3422 3927 -3388
rect 3915 -3428 3973 -3422
rect 401 -3498 413 -3493
rect 373 -3510 379 -3498
rect 407 -3509 413 -3498
rect 438 -3505 467 -3493
rect 438 -3506 479 -3505
rect 453 -3510 467 -3506
rect 495 -3509 501 -3493
rect 3769 -3505 3784 -3471
rect 453 -3531 463 -3510
rect 4104 -3524 4119 -3031
rect 4138 -3065 4173 -3031
rect 4138 -3524 4172 -3065
rect 4284 -3133 4342 -3127
rect 4284 -3167 4296 -3133
rect 4284 -3173 4342 -3167
rect 4284 -3441 4342 -3435
rect 4284 -3475 4296 -3441
rect 4284 -3481 4342 -3475
rect 4138 -3558 4153 -3524
rect 144 -3594 920 -3560
<< metal1 >>
rect 7647 1599 7703 1645
rect 0 0 200 200
rect 7675 46 7703 1599
rect 7586 0 7703 46
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
<< metal2 >>
rect 355 1571 7727 1599
rect 2267 1567 2335 1571
rect 6031 1567 6099 1571
rect 356 1418 7671 1446
rect 3013 1291 3944 1319
rect 4139 1291 7615 1319
rect 947 1177 3606 1205
rect 4247 1177 7370 1205
rect 2104 947 3466 975
rect 5859 947 7221 975
rect 520 676 1882 704
rect 4275 676 5637 704
rect 371 446 3494 474
rect 4135 446 7258 474
rect 142 328 3602 356
rect 3797 328 7313 356
rect 7587 333 7615 1291
rect 7643 233 7671 1418
rect 116 205 7671 233
rect 1642 74 1710 78
rect 5406 74 5474 78
rect 7699 74 7727 1571
rect 1642 46 7727 74
use dffc_2  dffc_2_3
timestamp 1624053917
transform -1 0 2989 0 -1 1622
box -67 -23 2436 852
use dffc_2  dffc_2_0
timestamp 1624053917
transform 1 0 988 0 1 23
box -67 -23 2436 852
use dffc_2  dffc_2_2
timestamp 1624053917
transform -1 0 6753 0 -1 1622
box -67 -23 2436 852
use dffc_2  dffc_2_1
timestamp 1624053917
transform 1 0 4752 0 1 23
box -67 -23 2436 852
use xor_somo  xor_somo_0
timestamp 1624053917
transform 1 0 96 0 1 23
box -96 -2000 4428 1165
use xor_somo  xor_somo_3
timestamp 1624053917
transform -1 0 3881 0 -1 1622
box -96 -2000 4428 1165
use xor_somo  xor_somo_1
timestamp 1624053917
transform 1 0 3860 0 1 23
box -96 -2000 4428 1165
use xor_somo  xor_somo_2
timestamp 1624053917
transform -1 0 7645 0 -1 1622
box -96 -2000 4428 1165
use xor_somo  xor_somo_4
timestamp 1624053917
transform 1 0 96 0 1 -3577
box -96 -2000 4428 1165
use and_somo  and_somo_2
timestamp 1624053917
transform -1 0 4358 0 -1 1622
box -81 -2000 2214 1147
use and_somo  and_somo_0
timestamp 1624053917
transform 1 0 3383 0 1 23
box -81 -2000 2214 1147
use and_somo  and_somo_1
timestamp 1624053917
transform 1 0 7147 0 1 23
box -81 -2000 2214 1147
use and_somo  and_somo_3
timestamp 1624053917
transform 1 0 81 0 1 -3577
box -81 -2000 2214 1147
<< labels >>
rlabel space 3797 279 3851 333 1 D0
rlabel metal2 355 1571 434 1599 1 CLR
rlabel metal2 356 1418 451 1446 1 CLK
rlabel space 948 1191 1000 1246 1 D3
rlabel space 4247 1163 4307 1223 1 D2
rlabel space 6741 399 6793 454 1 D1
rlabel space 2977 399 3029 454 1 D0
rlabel space 111 805 163 841 1 vdd
rlabel space 578 1602 623 1638 1 vss
rlabel metal2 142 328 185 356 1 CE
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 D0
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 CE
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLR
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLK
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 vdd
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 D1
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 D2
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 D3
port 9 nsew
<< end >>
