magic
tech sky130A
magscale 1 2
timestamp 1615944125
<< error_p >>
rect -1202 292 -1144 298
rect -998 292 -940 298
rect -794 292 -736 298
rect -590 292 -532 298
rect -386 292 -328 298
rect -182 292 -124 298
rect 22 292 80 298
rect 226 292 284 298
rect 430 292 488 298
rect 634 292 692 298
rect 838 292 896 298
rect 1042 292 1100 298
rect 1246 292 1304 298
rect -1202 258 -1190 292
rect -998 258 -986 292
rect -794 258 -782 292
rect -590 258 -578 292
rect -386 258 -374 292
rect -182 258 -170 292
rect 22 258 34 292
rect 226 258 238 292
rect 430 258 442 292
rect 634 258 646 292
rect 838 258 850 292
rect 1042 258 1054 292
rect 1246 258 1258 292
rect -1202 252 -1144 258
rect -998 252 -940 258
rect -794 252 -736 258
rect -590 252 -532 258
rect -386 252 -328 258
rect -182 252 -124 258
rect 22 252 80 258
rect 226 252 284 258
rect 430 252 488 258
rect 634 252 692 258
rect 838 252 896 258
rect 1042 252 1100 258
rect 1246 252 1304 258
rect -1304 -258 -1246 -252
rect -1100 -258 -1042 -252
rect -896 -258 -838 -252
rect -692 -258 -634 -252
rect -488 -258 -430 -252
rect -284 -258 -226 -252
rect -80 -258 -22 -252
rect 124 -258 182 -252
rect 328 -258 386 -252
rect 532 -258 590 -252
rect 736 -258 794 -252
rect 940 -258 998 -252
rect 1144 -258 1202 -252
rect -1304 -292 -1292 -258
rect -1100 -292 -1088 -258
rect -896 -292 -884 -258
rect -692 -292 -680 -258
rect -488 -292 -476 -258
rect -284 -292 -272 -258
rect -80 -292 -68 -258
rect 124 -292 136 -258
rect 328 -292 340 -258
rect 532 -292 544 -258
rect 736 -292 748 -258
rect 940 -292 952 -258
rect 1144 -292 1156 -258
rect -1304 -298 -1246 -292
rect -1100 -298 -1042 -292
rect -896 -298 -838 -292
rect -692 -298 -634 -292
rect -488 -298 -430 -292
rect -284 -298 -226 -292
rect -80 -298 -22 -292
rect 124 -298 182 -292
rect 328 -298 386 -292
rect 532 -298 590 -292
rect 736 -298 794 -292
rect 940 -298 998 -292
rect 1144 -298 1202 -292
<< pwell >>
rect -1493 -430 1493 430
<< nmos >>
rect -1297 -220 -1253 220
rect -1195 -220 -1151 220
rect -1093 -220 -1049 220
rect -991 -220 -947 220
rect -889 -220 -845 220
rect -787 -220 -743 220
rect -685 -220 -641 220
rect -583 -220 -539 220
rect -481 -220 -437 220
rect -379 -220 -335 220
rect -277 -220 -233 220
rect -175 -220 -131 220
rect -73 -220 -29 220
rect 29 -220 73 220
rect 131 -220 175 220
rect 233 -220 277 220
rect 335 -220 379 220
rect 437 -220 481 220
rect 539 -220 583 220
rect 641 -220 685 220
rect 743 -220 787 220
rect 845 -220 889 220
rect 947 -220 991 220
rect 1049 -220 1093 220
rect 1151 -220 1195 220
rect 1253 -220 1297 220
<< ndiff >>
rect -1355 208 -1297 220
rect -1355 -208 -1343 208
rect -1309 -208 -1297 208
rect -1355 -220 -1297 -208
rect -1253 208 -1195 220
rect -1253 -208 -1241 208
rect -1207 -208 -1195 208
rect -1253 -220 -1195 -208
rect -1151 208 -1093 220
rect -1151 -208 -1139 208
rect -1105 -208 -1093 208
rect -1151 -220 -1093 -208
rect -1049 208 -991 220
rect -1049 -208 -1037 208
rect -1003 -208 -991 208
rect -1049 -220 -991 -208
rect -947 208 -889 220
rect -947 -208 -935 208
rect -901 -208 -889 208
rect -947 -220 -889 -208
rect -845 208 -787 220
rect -845 -208 -833 208
rect -799 -208 -787 208
rect -845 -220 -787 -208
rect -743 208 -685 220
rect -743 -208 -731 208
rect -697 -208 -685 208
rect -743 -220 -685 -208
rect -641 208 -583 220
rect -641 -208 -629 208
rect -595 -208 -583 208
rect -641 -220 -583 -208
rect -539 208 -481 220
rect -539 -208 -527 208
rect -493 -208 -481 208
rect -539 -220 -481 -208
rect -437 208 -379 220
rect -437 -208 -425 208
rect -391 -208 -379 208
rect -437 -220 -379 -208
rect -335 208 -277 220
rect -335 -208 -323 208
rect -289 -208 -277 208
rect -335 -220 -277 -208
rect -233 208 -175 220
rect -233 -208 -221 208
rect -187 -208 -175 208
rect -233 -220 -175 -208
rect -131 208 -73 220
rect -131 -208 -119 208
rect -85 -208 -73 208
rect -131 -220 -73 -208
rect -29 208 29 220
rect -29 -208 -17 208
rect 17 -208 29 208
rect -29 -220 29 -208
rect 73 208 131 220
rect 73 -208 85 208
rect 119 -208 131 208
rect 73 -220 131 -208
rect 175 208 233 220
rect 175 -208 187 208
rect 221 -208 233 208
rect 175 -220 233 -208
rect 277 208 335 220
rect 277 -208 289 208
rect 323 -208 335 208
rect 277 -220 335 -208
rect 379 208 437 220
rect 379 -208 391 208
rect 425 -208 437 208
rect 379 -220 437 -208
rect 481 208 539 220
rect 481 -208 493 208
rect 527 -208 539 208
rect 481 -220 539 -208
rect 583 208 641 220
rect 583 -208 595 208
rect 629 -208 641 208
rect 583 -220 641 -208
rect 685 208 743 220
rect 685 -208 697 208
rect 731 -208 743 208
rect 685 -220 743 -208
rect 787 208 845 220
rect 787 -208 799 208
rect 833 -208 845 208
rect 787 -220 845 -208
rect 889 208 947 220
rect 889 -208 901 208
rect 935 -208 947 208
rect 889 -220 947 -208
rect 991 208 1049 220
rect 991 -208 1003 208
rect 1037 -208 1049 208
rect 991 -220 1049 -208
rect 1093 208 1151 220
rect 1093 -208 1105 208
rect 1139 -208 1151 208
rect 1093 -220 1151 -208
rect 1195 208 1253 220
rect 1195 -208 1207 208
rect 1241 -208 1253 208
rect 1195 -220 1253 -208
rect 1297 208 1355 220
rect 1297 -208 1309 208
rect 1343 -208 1355 208
rect 1297 -220 1355 -208
<< ndiffc >>
rect -1343 -208 -1309 208
rect -1241 -208 -1207 208
rect -1139 -208 -1105 208
rect -1037 -208 -1003 208
rect -935 -208 -901 208
rect -833 -208 -799 208
rect -731 -208 -697 208
rect -629 -208 -595 208
rect -527 -208 -493 208
rect -425 -208 -391 208
rect -323 -208 -289 208
rect -221 -208 -187 208
rect -119 -208 -85 208
rect -17 -208 17 208
rect 85 -208 119 208
rect 187 -208 221 208
rect 289 -208 323 208
rect 391 -208 425 208
rect 493 -208 527 208
rect 595 -208 629 208
rect 697 -208 731 208
rect 799 -208 833 208
rect 901 -208 935 208
rect 1003 -208 1037 208
rect 1105 -208 1139 208
rect 1207 -208 1241 208
rect 1309 -208 1343 208
<< psubdiff >>
rect -1457 360 -1361 394
rect 1361 360 1457 394
rect -1457 298 -1423 360
rect 1423 298 1457 360
rect -1457 -360 -1423 -298
rect 1423 -360 1457 -298
rect -1457 -394 -1361 -360
rect 1361 -394 1457 -360
<< psubdiffcont >>
rect -1361 360 1361 394
rect -1457 -298 -1423 298
rect 1423 -298 1457 298
rect -1361 -394 1361 -360
<< poly >>
rect -1206 292 -1140 308
rect -1206 258 -1190 292
rect -1156 258 -1140 292
rect -1297 220 -1253 246
rect -1206 242 -1140 258
rect -1002 292 -936 308
rect -1002 258 -986 292
rect -952 258 -936 292
rect -1195 220 -1151 242
rect -1093 220 -1049 246
rect -1002 242 -936 258
rect -798 292 -732 308
rect -798 258 -782 292
rect -748 258 -732 292
rect -991 220 -947 242
rect -889 220 -845 246
rect -798 242 -732 258
rect -594 292 -528 308
rect -594 258 -578 292
rect -544 258 -528 292
rect -787 220 -743 242
rect -685 220 -641 246
rect -594 242 -528 258
rect -390 292 -324 308
rect -390 258 -374 292
rect -340 258 -324 292
rect -583 220 -539 242
rect -481 220 -437 246
rect -390 242 -324 258
rect -186 292 -120 308
rect -186 258 -170 292
rect -136 258 -120 292
rect -379 220 -335 242
rect -277 220 -233 246
rect -186 242 -120 258
rect 18 292 84 308
rect 18 258 34 292
rect 68 258 84 292
rect -175 220 -131 242
rect -73 220 -29 246
rect 18 242 84 258
rect 222 292 288 308
rect 222 258 238 292
rect 272 258 288 292
rect 29 220 73 242
rect 131 220 175 246
rect 222 242 288 258
rect 426 292 492 308
rect 426 258 442 292
rect 476 258 492 292
rect 233 220 277 242
rect 335 220 379 246
rect 426 242 492 258
rect 630 292 696 308
rect 630 258 646 292
rect 680 258 696 292
rect 437 220 481 242
rect 539 220 583 246
rect 630 242 696 258
rect 834 292 900 308
rect 834 258 850 292
rect 884 258 900 292
rect 641 220 685 242
rect 743 220 787 246
rect 834 242 900 258
rect 1038 292 1104 308
rect 1038 258 1054 292
rect 1088 258 1104 292
rect 845 220 889 242
rect 947 220 991 246
rect 1038 242 1104 258
rect 1242 292 1308 308
rect 1242 258 1258 292
rect 1292 258 1308 292
rect 1049 220 1093 242
rect 1151 220 1195 246
rect 1242 242 1308 258
rect 1253 220 1297 242
rect -1297 -242 -1253 -220
rect -1308 -258 -1242 -242
rect -1195 -246 -1151 -220
rect -1093 -242 -1049 -220
rect -1308 -292 -1292 -258
rect -1258 -292 -1242 -258
rect -1308 -308 -1242 -292
rect -1104 -258 -1038 -242
rect -991 -246 -947 -220
rect -889 -242 -845 -220
rect -1104 -292 -1088 -258
rect -1054 -292 -1038 -258
rect -1104 -308 -1038 -292
rect -900 -258 -834 -242
rect -787 -246 -743 -220
rect -685 -242 -641 -220
rect -900 -292 -884 -258
rect -850 -292 -834 -258
rect -900 -308 -834 -292
rect -696 -258 -630 -242
rect -583 -246 -539 -220
rect -481 -242 -437 -220
rect -696 -292 -680 -258
rect -646 -292 -630 -258
rect -696 -308 -630 -292
rect -492 -258 -426 -242
rect -379 -246 -335 -220
rect -277 -242 -233 -220
rect -492 -292 -476 -258
rect -442 -292 -426 -258
rect -492 -308 -426 -292
rect -288 -258 -222 -242
rect -175 -246 -131 -220
rect -73 -242 -29 -220
rect -288 -292 -272 -258
rect -238 -292 -222 -258
rect -288 -308 -222 -292
rect -84 -258 -18 -242
rect 29 -246 73 -220
rect 131 -242 175 -220
rect -84 -292 -68 -258
rect -34 -292 -18 -258
rect -84 -308 -18 -292
rect 120 -258 186 -242
rect 233 -246 277 -220
rect 335 -242 379 -220
rect 120 -292 136 -258
rect 170 -292 186 -258
rect 120 -308 186 -292
rect 324 -258 390 -242
rect 437 -246 481 -220
rect 539 -242 583 -220
rect 324 -292 340 -258
rect 374 -292 390 -258
rect 324 -308 390 -292
rect 528 -258 594 -242
rect 641 -246 685 -220
rect 743 -242 787 -220
rect 528 -292 544 -258
rect 578 -292 594 -258
rect 528 -308 594 -292
rect 732 -258 798 -242
rect 845 -246 889 -220
rect 947 -242 991 -220
rect 732 -292 748 -258
rect 782 -292 798 -258
rect 732 -308 798 -292
rect 936 -258 1002 -242
rect 1049 -246 1093 -220
rect 1151 -242 1195 -220
rect 936 -292 952 -258
rect 986 -292 1002 -258
rect 936 -308 1002 -292
rect 1140 -258 1206 -242
rect 1253 -246 1297 -220
rect 1140 -292 1156 -258
rect 1190 -292 1206 -258
rect 1140 -308 1206 -292
<< polycont >>
rect -1190 258 -1156 292
rect -986 258 -952 292
rect -782 258 -748 292
rect -578 258 -544 292
rect -374 258 -340 292
rect -170 258 -136 292
rect 34 258 68 292
rect 238 258 272 292
rect 442 258 476 292
rect 646 258 680 292
rect 850 258 884 292
rect 1054 258 1088 292
rect 1258 258 1292 292
rect -1292 -292 -1258 -258
rect -1088 -292 -1054 -258
rect -884 -292 -850 -258
rect -680 -292 -646 -258
rect -476 -292 -442 -258
rect -272 -292 -238 -258
rect -68 -292 -34 -258
rect 136 -292 170 -258
rect 340 -292 374 -258
rect 544 -292 578 -258
rect 748 -292 782 -258
rect 952 -292 986 -258
rect 1156 -292 1190 -258
<< locali >>
rect -1457 360 -1361 394
rect 1361 360 1457 394
rect -1457 298 -1423 360
rect 1423 298 1457 360
rect -1206 258 -1190 292
rect -1156 258 -1140 292
rect -1002 258 -986 292
rect -952 258 -936 292
rect -798 258 -782 292
rect -748 258 -732 292
rect -594 258 -578 292
rect -544 258 -528 292
rect -390 258 -374 292
rect -340 258 -324 292
rect -186 258 -170 292
rect -136 258 -120 292
rect 18 258 34 292
rect 68 258 84 292
rect 222 258 238 292
rect 272 258 288 292
rect 426 258 442 292
rect 476 258 492 292
rect 630 258 646 292
rect 680 258 696 292
rect 834 258 850 292
rect 884 258 900 292
rect 1038 258 1054 292
rect 1088 258 1104 292
rect 1242 258 1258 292
rect 1292 258 1308 292
rect -1343 208 -1309 224
rect -1343 -224 -1309 -208
rect -1241 208 -1207 224
rect -1241 -224 -1207 -208
rect -1139 208 -1105 224
rect -1139 -224 -1105 -208
rect -1037 208 -1003 224
rect -1037 -224 -1003 -208
rect -935 208 -901 224
rect -935 -224 -901 -208
rect -833 208 -799 224
rect -833 -224 -799 -208
rect -731 208 -697 224
rect -731 -224 -697 -208
rect -629 208 -595 224
rect -629 -224 -595 -208
rect -527 208 -493 224
rect -527 -224 -493 -208
rect -425 208 -391 224
rect -425 -224 -391 -208
rect -323 208 -289 224
rect -323 -224 -289 -208
rect -221 208 -187 224
rect -221 -224 -187 -208
rect -119 208 -85 224
rect -119 -224 -85 -208
rect -17 208 17 224
rect -17 -224 17 -208
rect 85 208 119 224
rect 85 -224 119 -208
rect 187 208 221 224
rect 187 -224 221 -208
rect 289 208 323 224
rect 289 -224 323 -208
rect 391 208 425 224
rect 391 -224 425 -208
rect 493 208 527 224
rect 493 -224 527 -208
rect 595 208 629 224
rect 595 -224 629 -208
rect 697 208 731 224
rect 697 -224 731 -208
rect 799 208 833 224
rect 799 -224 833 -208
rect 901 208 935 224
rect 901 -224 935 -208
rect 1003 208 1037 224
rect 1003 -224 1037 -208
rect 1105 208 1139 224
rect 1105 -224 1139 -208
rect 1207 208 1241 224
rect 1207 -224 1241 -208
rect 1309 208 1343 224
rect 1309 -224 1343 -208
rect -1308 -292 -1292 -258
rect -1258 -292 -1242 -258
rect -1104 -292 -1088 -258
rect -1054 -292 -1038 -258
rect -900 -292 -884 -258
rect -850 -292 -834 -258
rect -696 -292 -680 -258
rect -646 -292 -630 -258
rect -492 -292 -476 -258
rect -442 -292 -426 -258
rect -288 -292 -272 -258
rect -238 -292 -222 -258
rect -84 -292 -68 -258
rect -34 -292 -18 -258
rect 120 -292 136 -258
rect 170 -292 186 -258
rect 324 -292 340 -258
rect 374 -292 390 -258
rect 528 -292 544 -258
rect 578 -292 594 -258
rect 732 -292 748 -258
rect 782 -292 798 -258
rect 936 -292 952 -258
rect 986 -292 1002 -258
rect 1140 -292 1156 -258
rect 1190 -292 1206 -258
rect -1457 -360 -1423 -298
rect 1423 -360 1457 -298
rect -1457 -394 -1361 -360
rect 1361 -394 1457 -360
<< viali >>
rect -1190 258 -1156 292
rect -986 258 -952 292
rect -782 258 -748 292
rect -578 258 -544 292
rect -374 258 -340 292
rect -170 258 -136 292
rect 34 258 68 292
rect 238 258 272 292
rect 442 258 476 292
rect 646 258 680 292
rect 850 258 884 292
rect 1054 258 1088 292
rect 1258 258 1292 292
rect -1343 -208 -1309 208
rect -1241 -208 -1207 208
rect -1139 -208 -1105 208
rect -1037 -208 -1003 208
rect -935 -208 -901 208
rect -833 -208 -799 208
rect -731 -208 -697 208
rect -629 -208 -595 208
rect -527 -208 -493 208
rect -425 -208 -391 208
rect -323 -208 -289 208
rect -221 -208 -187 208
rect -119 -208 -85 208
rect -17 -208 17 208
rect 85 -208 119 208
rect 187 -208 221 208
rect 289 -208 323 208
rect 391 -208 425 208
rect 493 -208 527 208
rect 595 -208 629 208
rect 697 -208 731 208
rect 799 -208 833 208
rect 901 -208 935 208
rect 1003 -208 1037 208
rect 1105 -208 1139 208
rect 1207 -208 1241 208
rect 1309 -208 1343 208
rect -1292 -292 -1258 -258
rect -1088 -292 -1054 -258
rect -884 -292 -850 -258
rect -680 -292 -646 -258
rect -476 -292 -442 -258
rect -272 -292 -238 -258
rect -68 -292 -34 -258
rect 136 -292 170 -258
rect 340 -292 374 -258
rect 544 -292 578 -258
rect 748 -292 782 -258
rect 952 -292 986 -258
rect 1156 -292 1190 -258
<< metal1 >>
rect -1202 292 -1144 298
rect -1202 258 -1190 292
rect -1156 258 -1144 292
rect -1202 252 -1144 258
rect -998 292 -940 298
rect -998 258 -986 292
rect -952 258 -940 292
rect -998 252 -940 258
rect -794 292 -736 298
rect -794 258 -782 292
rect -748 258 -736 292
rect -794 252 -736 258
rect -590 292 -532 298
rect -590 258 -578 292
rect -544 258 -532 292
rect -590 252 -532 258
rect -386 292 -328 298
rect -386 258 -374 292
rect -340 258 -328 292
rect -386 252 -328 258
rect -182 292 -124 298
rect -182 258 -170 292
rect -136 258 -124 292
rect -182 252 -124 258
rect 22 292 80 298
rect 22 258 34 292
rect 68 258 80 292
rect 22 252 80 258
rect 226 292 284 298
rect 226 258 238 292
rect 272 258 284 292
rect 226 252 284 258
rect 430 292 488 298
rect 430 258 442 292
rect 476 258 488 292
rect 430 252 488 258
rect 634 292 692 298
rect 634 258 646 292
rect 680 258 692 292
rect 634 252 692 258
rect 838 292 896 298
rect 838 258 850 292
rect 884 258 896 292
rect 838 252 896 258
rect 1042 292 1100 298
rect 1042 258 1054 292
rect 1088 258 1100 292
rect 1042 252 1100 258
rect 1246 292 1304 298
rect 1246 258 1258 292
rect 1292 258 1304 292
rect 1246 252 1304 258
rect -1349 208 -1303 220
rect -1349 -208 -1343 208
rect -1309 -208 -1303 208
rect -1349 -220 -1303 -208
rect -1247 208 -1201 220
rect -1247 -208 -1241 208
rect -1207 -208 -1201 208
rect -1247 -220 -1201 -208
rect -1145 208 -1099 220
rect -1145 -208 -1139 208
rect -1105 -208 -1099 208
rect -1145 -220 -1099 -208
rect -1043 208 -997 220
rect -1043 -208 -1037 208
rect -1003 -208 -997 208
rect -1043 -220 -997 -208
rect -941 208 -895 220
rect -941 -208 -935 208
rect -901 -208 -895 208
rect -941 -220 -895 -208
rect -839 208 -793 220
rect -839 -208 -833 208
rect -799 -208 -793 208
rect -839 -220 -793 -208
rect -737 208 -691 220
rect -737 -208 -731 208
rect -697 -208 -691 208
rect -737 -220 -691 -208
rect -635 208 -589 220
rect -635 -208 -629 208
rect -595 -208 -589 208
rect -635 -220 -589 -208
rect -533 208 -487 220
rect -533 -208 -527 208
rect -493 -208 -487 208
rect -533 -220 -487 -208
rect -431 208 -385 220
rect -431 -208 -425 208
rect -391 -208 -385 208
rect -431 -220 -385 -208
rect -329 208 -283 220
rect -329 -208 -323 208
rect -289 -208 -283 208
rect -329 -220 -283 -208
rect -227 208 -181 220
rect -227 -208 -221 208
rect -187 -208 -181 208
rect -227 -220 -181 -208
rect -125 208 -79 220
rect -125 -208 -119 208
rect -85 -208 -79 208
rect -125 -220 -79 -208
rect -23 208 23 220
rect -23 -208 -17 208
rect 17 -208 23 208
rect -23 -220 23 -208
rect 79 208 125 220
rect 79 -208 85 208
rect 119 -208 125 208
rect 79 -220 125 -208
rect 181 208 227 220
rect 181 -208 187 208
rect 221 -208 227 208
rect 181 -220 227 -208
rect 283 208 329 220
rect 283 -208 289 208
rect 323 -208 329 208
rect 283 -220 329 -208
rect 385 208 431 220
rect 385 -208 391 208
rect 425 -208 431 208
rect 385 -220 431 -208
rect 487 208 533 220
rect 487 -208 493 208
rect 527 -208 533 208
rect 487 -220 533 -208
rect 589 208 635 220
rect 589 -208 595 208
rect 629 -208 635 208
rect 589 -220 635 -208
rect 691 208 737 220
rect 691 -208 697 208
rect 731 -208 737 208
rect 691 -220 737 -208
rect 793 208 839 220
rect 793 -208 799 208
rect 833 -208 839 208
rect 793 -220 839 -208
rect 895 208 941 220
rect 895 -208 901 208
rect 935 -208 941 208
rect 895 -220 941 -208
rect 997 208 1043 220
rect 997 -208 1003 208
rect 1037 -208 1043 208
rect 997 -220 1043 -208
rect 1099 208 1145 220
rect 1099 -208 1105 208
rect 1139 -208 1145 208
rect 1099 -220 1145 -208
rect 1201 208 1247 220
rect 1201 -208 1207 208
rect 1241 -208 1247 208
rect 1201 -220 1247 -208
rect 1303 208 1349 220
rect 1303 -208 1309 208
rect 1343 -208 1349 208
rect 1303 -220 1349 -208
rect -1304 -258 -1246 -252
rect -1304 -292 -1292 -258
rect -1258 -292 -1246 -258
rect -1304 -298 -1246 -292
rect -1100 -258 -1042 -252
rect -1100 -292 -1088 -258
rect -1054 -292 -1042 -258
rect -1100 -298 -1042 -292
rect -896 -258 -838 -252
rect -896 -292 -884 -258
rect -850 -292 -838 -258
rect -896 -298 -838 -292
rect -692 -258 -634 -252
rect -692 -292 -680 -258
rect -646 -292 -634 -258
rect -692 -298 -634 -292
rect -488 -258 -430 -252
rect -488 -292 -476 -258
rect -442 -292 -430 -258
rect -488 -298 -430 -292
rect -284 -258 -226 -252
rect -284 -292 -272 -258
rect -238 -292 -226 -258
rect -284 -298 -226 -292
rect -80 -258 -22 -252
rect -80 -292 -68 -258
rect -34 -292 -22 -258
rect -80 -298 -22 -292
rect 124 -258 182 -252
rect 124 -292 136 -258
rect 170 -292 182 -258
rect 124 -298 182 -292
rect 328 -258 386 -252
rect 328 -292 340 -258
rect 374 -292 386 -258
rect 328 -298 386 -292
rect 532 -258 590 -252
rect 532 -292 544 -258
rect 578 -292 590 -258
rect 532 -298 590 -292
rect 736 -258 794 -252
rect 736 -292 748 -258
rect 782 -292 794 -258
rect 736 -298 794 -292
rect 940 -258 998 -252
rect 940 -292 952 -258
rect 986 -292 998 -258
rect 940 -298 998 -292
rect 1144 -258 1202 -252
rect 1144 -292 1156 -258
rect 1190 -292 1202 -258
rect 1144 -298 1202 -292
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1440 -377 1440 377
string parameters w 2.2 l 0.22 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
