magic
tech sky130A
magscale 1 2
timestamp 1615909117
<< error_p >>
rect -2920 306 -2862 312
rect -2802 306 -2744 312
rect -2684 306 -2626 312
rect -2566 306 -2508 312
rect -2448 306 -2390 312
rect -2330 306 -2272 312
rect -2212 306 -2154 312
rect -2094 306 -2036 312
rect -1976 306 -1918 312
rect -1858 306 -1800 312
rect -1740 306 -1682 312
rect -1622 306 -1564 312
rect -1504 306 -1446 312
rect -1386 306 -1328 312
rect -1268 306 -1210 312
rect -1150 306 -1092 312
rect -1032 306 -974 312
rect -914 306 -856 312
rect -796 306 -738 312
rect -678 306 -620 312
rect -560 306 -502 312
rect -442 306 -384 312
rect -324 306 -266 312
rect -206 306 -148 312
rect -88 306 -30 312
rect 30 306 88 312
rect 148 306 206 312
rect 266 306 324 312
rect 384 306 442 312
rect 502 306 560 312
rect 620 306 678 312
rect 738 306 796 312
rect 856 306 914 312
rect 974 306 1032 312
rect 1092 306 1150 312
rect 1210 306 1268 312
rect 1328 306 1386 312
rect 1446 306 1504 312
rect 1564 306 1622 312
rect 1682 306 1740 312
rect 1800 306 1858 312
rect 1918 306 1976 312
rect 2036 306 2094 312
rect 2154 306 2212 312
rect 2272 306 2330 312
rect 2390 306 2448 312
rect 2508 306 2566 312
rect 2626 306 2684 312
rect 2744 306 2802 312
rect 2862 306 2920 312
rect -2920 272 -2908 306
rect -2802 272 -2790 306
rect -2684 272 -2672 306
rect -2566 272 -2554 306
rect -2448 272 -2436 306
rect -2330 272 -2318 306
rect -2212 272 -2200 306
rect -2094 272 -2082 306
rect -1976 272 -1964 306
rect -1858 272 -1846 306
rect -1740 272 -1728 306
rect -1622 272 -1610 306
rect -1504 272 -1492 306
rect -1386 272 -1374 306
rect -1268 272 -1256 306
rect -1150 272 -1138 306
rect -1032 272 -1020 306
rect -914 272 -902 306
rect -796 272 -784 306
rect -678 272 -666 306
rect -560 272 -548 306
rect -442 272 -430 306
rect -324 272 -312 306
rect -206 272 -194 306
rect -88 272 -76 306
rect 30 272 42 306
rect 148 272 160 306
rect 266 272 278 306
rect 384 272 396 306
rect 502 272 514 306
rect 620 272 632 306
rect 738 272 750 306
rect 856 272 868 306
rect 974 272 986 306
rect 1092 272 1104 306
rect 1210 272 1222 306
rect 1328 272 1340 306
rect 1446 272 1458 306
rect 1564 272 1576 306
rect 1682 272 1694 306
rect 1800 272 1812 306
rect 1918 272 1930 306
rect 2036 272 2048 306
rect 2154 272 2166 306
rect 2272 272 2284 306
rect 2390 272 2402 306
rect 2508 272 2520 306
rect 2626 272 2638 306
rect 2744 272 2756 306
rect 2862 272 2874 306
rect -2920 266 -2862 272
rect -2802 266 -2744 272
rect -2684 266 -2626 272
rect -2566 266 -2508 272
rect -2448 266 -2390 272
rect -2330 266 -2272 272
rect -2212 266 -2154 272
rect -2094 266 -2036 272
rect -1976 266 -1918 272
rect -1858 266 -1800 272
rect -1740 266 -1682 272
rect -1622 266 -1564 272
rect -1504 266 -1446 272
rect -1386 266 -1328 272
rect -1268 266 -1210 272
rect -1150 266 -1092 272
rect -1032 266 -974 272
rect -914 266 -856 272
rect -796 266 -738 272
rect -678 266 -620 272
rect -560 266 -502 272
rect -442 266 -384 272
rect -324 266 -266 272
rect -206 266 -148 272
rect -88 266 -30 272
rect 30 266 88 272
rect 148 266 206 272
rect 266 266 324 272
rect 384 266 442 272
rect 502 266 560 272
rect 620 266 678 272
rect 738 266 796 272
rect 856 266 914 272
rect 974 266 1032 272
rect 1092 266 1150 272
rect 1210 266 1268 272
rect 1328 266 1386 272
rect 1446 266 1504 272
rect 1564 266 1622 272
rect 1682 266 1740 272
rect 1800 266 1858 272
rect 1918 266 1976 272
rect 2036 266 2094 272
rect 2154 266 2212 272
rect 2272 266 2330 272
rect 2390 266 2448 272
rect 2508 266 2566 272
rect 2626 266 2684 272
rect 2744 266 2802 272
rect 2862 266 2920 272
rect -2920 -272 -2862 -266
rect -2802 -272 -2744 -266
rect -2684 -272 -2626 -266
rect -2566 -272 -2508 -266
rect -2448 -272 -2390 -266
rect -2330 -272 -2272 -266
rect -2212 -272 -2154 -266
rect -2094 -272 -2036 -266
rect -1976 -272 -1918 -266
rect -1858 -272 -1800 -266
rect -1740 -272 -1682 -266
rect -1622 -272 -1564 -266
rect -1504 -272 -1446 -266
rect -1386 -272 -1328 -266
rect -1268 -272 -1210 -266
rect -1150 -272 -1092 -266
rect -1032 -272 -974 -266
rect -914 -272 -856 -266
rect -796 -272 -738 -266
rect -678 -272 -620 -266
rect -560 -272 -502 -266
rect -442 -272 -384 -266
rect -324 -272 -266 -266
rect -206 -272 -148 -266
rect -88 -272 -30 -266
rect 30 -272 88 -266
rect 148 -272 206 -266
rect 266 -272 324 -266
rect 384 -272 442 -266
rect 502 -272 560 -266
rect 620 -272 678 -266
rect 738 -272 796 -266
rect 856 -272 914 -266
rect 974 -272 1032 -266
rect 1092 -272 1150 -266
rect 1210 -272 1268 -266
rect 1328 -272 1386 -266
rect 1446 -272 1504 -266
rect 1564 -272 1622 -266
rect 1682 -272 1740 -266
rect 1800 -272 1858 -266
rect 1918 -272 1976 -266
rect 2036 -272 2094 -266
rect 2154 -272 2212 -266
rect 2272 -272 2330 -266
rect 2390 -272 2448 -266
rect 2508 -272 2566 -266
rect 2626 -272 2684 -266
rect 2744 -272 2802 -266
rect 2862 -272 2920 -266
rect -2920 -306 -2908 -272
rect -2802 -306 -2790 -272
rect -2684 -306 -2672 -272
rect -2566 -306 -2554 -272
rect -2448 -306 -2436 -272
rect -2330 -306 -2318 -272
rect -2212 -306 -2200 -272
rect -2094 -306 -2082 -272
rect -1976 -306 -1964 -272
rect -1858 -306 -1846 -272
rect -1740 -306 -1728 -272
rect -1622 -306 -1610 -272
rect -1504 -306 -1492 -272
rect -1386 -306 -1374 -272
rect -1268 -306 -1256 -272
rect -1150 -306 -1138 -272
rect -1032 -306 -1020 -272
rect -914 -306 -902 -272
rect -796 -306 -784 -272
rect -678 -306 -666 -272
rect -560 -306 -548 -272
rect -442 -306 -430 -272
rect -324 -306 -312 -272
rect -206 -306 -194 -272
rect -88 -306 -76 -272
rect 30 -306 42 -272
rect 148 -306 160 -272
rect 266 -306 278 -272
rect 384 -306 396 -272
rect 502 -306 514 -272
rect 620 -306 632 -272
rect 738 -306 750 -272
rect 856 -306 868 -272
rect 974 -306 986 -272
rect 1092 -306 1104 -272
rect 1210 -306 1222 -272
rect 1328 -306 1340 -272
rect 1446 -306 1458 -272
rect 1564 -306 1576 -272
rect 1682 -306 1694 -272
rect 1800 -306 1812 -272
rect 1918 -306 1930 -272
rect 2036 -306 2048 -272
rect 2154 -306 2166 -272
rect 2272 -306 2284 -272
rect 2390 -306 2402 -272
rect 2508 -306 2520 -272
rect 2626 -306 2638 -272
rect 2744 -306 2756 -272
rect 2862 -306 2874 -272
rect -2920 -312 -2862 -306
rect -2802 -312 -2744 -306
rect -2684 -312 -2626 -306
rect -2566 -312 -2508 -306
rect -2448 -312 -2390 -306
rect -2330 -312 -2272 -306
rect -2212 -312 -2154 -306
rect -2094 -312 -2036 -306
rect -1976 -312 -1918 -306
rect -1858 -312 -1800 -306
rect -1740 -312 -1682 -306
rect -1622 -312 -1564 -306
rect -1504 -312 -1446 -306
rect -1386 -312 -1328 -306
rect -1268 -312 -1210 -306
rect -1150 -312 -1092 -306
rect -1032 -312 -974 -306
rect -914 -312 -856 -306
rect -796 -312 -738 -306
rect -678 -312 -620 -306
rect -560 -312 -502 -306
rect -442 -312 -384 -306
rect -324 -312 -266 -306
rect -206 -312 -148 -306
rect -88 -312 -30 -306
rect 30 -312 88 -306
rect 148 -312 206 -306
rect 266 -312 324 -306
rect 384 -312 442 -306
rect 502 -312 560 -306
rect 620 -312 678 -306
rect 738 -312 796 -306
rect 856 -312 914 -306
rect 974 -312 1032 -306
rect 1092 -312 1150 -306
rect 1210 -312 1268 -306
rect 1328 -312 1386 -306
rect 1446 -312 1504 -306
rect 1564 -312 1622 -306
rect 1682 -312 1740 -306
rect 1800 -312 1858 -306
rect 1918 -312 1976 -306
rect 2036 -312 2094 -306
rect 2154 -312 2212 -306
rect 2272 -312 2330 -306
rect 2390 -312 2448 -306
rect 2508 -312 2566 -306
rect 2626 -312 2684 -306
rect 2744 -312 2802 -306
rect 2862 -312 2920 -306
<< nwell >>
rect -3117 -444 3117 444
<< pmos >>
rect -2921 -225 -2861 225
rect -2803 -225 -2743 225
rect -2685 -225 -2625 225
rect -2567 -225 -2507 225
rect -2449 -225 -2389 225
rect -2331 -225 -2271 225
rect -2213 -225 -2153 225
rect -2095 -225 -2035 225
rect -1977 -225 -1917 225
rect -1859 -225 -1799 225
rect -1741 -225 -1681 225
rect -1623 -225 -1563 225
rect -1505 -225 -1445 225
rect -1387 -225 -1327 225
rect -1269 -225 -1209 225
rect -1151 -225 -1091 225
rect -1033 -225 -973 225
rect -915 -225 -855 225
rect -797 -225 -737 225
rect -679 -225 -619 225
rect -561 -225 -501 225
rect -443 -225 -383 225
rect -325 -225 -265 225
rect -207 -225 -147 225
rect -89 -225 -29 225
rect 29 -225 89 225
rect 147 -225 207 225
rect 265 -225 325 225
rect 383 -225 443 225
rect 501 -225 561 225
rect 619 -225 679 225
rect 737 -225 797 225
rect 855 -225 915 225
rect 973 -225 1033 225
rect 1091 -225 1151 225
rect 1209 -225 1269 225
rect 1327 -225 1387 225
rect 1445 -225 1505 225
rect 1563 -225 1623 225
rect 1681 -225 1741 225
rect 1799 -225 1859 225
rect 1917 -225 1977 225
rect 2035 -225 2095 225
rect 2153 -225 2213 225
rect 2271 -225 2331 225
rect 2389 -225 2449 225
rect 2507 -225 2567 225
rect 2625 -225 2685 225
rect 2743 -225 2803 225
rect 2861 -225 2921 225
<< pdiff >>
rect -2979 213 -2921 225
rect -2979 -213 -2967 213
rect -2933 -213 -2921 213
rect -2979 -225 -2921 -213
rect -2861 213 -2803 225
rect -2861 -213 -2849 213
rect -2815 -213 -2803 213
rect -2861 -225 -2803 -213
rect -2743 213 -2685 225
rect -2743 -213 -2731 213
rect -2697 -213 -2685 213
rect -2743 -225 -2685 -213
rect -2625 213 -2567 225
rect -2625 -213 -2613 213
rect -2579 -213 -2567 213
rect -2625 -225 -2567 -213
rect -2507 213 -2449 225
rect -2507 -213 -2495 213
rect -2461 -213 -2449 213
rect -2507 -225 -2449 -213
rect -2389 213 -2331 225
rect -2389 -213 -2377 213
rect -2343 -213 -2331 213
rect -2389 -225 -2331 -213
rect -2271 213 -2213 225
rect -2271 -213 -2259 213
rect -2225 -213 -2213 213
rect -2271 -225 -2213 -213
rect -2153 213 -2095 225
rect -2153 -213 -2141 213
rect -2107 -213 -2095 213
rect -2153 -225 -2095 -213
rect -2035 213 -1977 225
rect -2035 -213 -2023 213
rect -1989 -213 -1977 213
rect -2035 -225 -1977 -213
rect -1917 213 -1859 225
rect -1917 -213 -1905 213
rect -1871 -213 -1859 213
rect -1917 -225 -1859 -213
rect -1799 213 -1741 225
rect -1799 -213 -1787 213
rect -1753 -213 -1741 213
rect -1799 -225 -1741 -213
rect -1681 213 -1623 225
rect -1681 -213 -1669 213
rect -1635 -213 -1623 213
rect -1681 -225 -1623 -213
rect -1563 213 -1505 225
rect -1563 -213 -1551 213
rect -1517 -213 -1505 213
rect -1563 -225 -1505 -213
rect -1445 213 -1387 225
rect -1445 -213 -1433 213
rect -1399 -213 -1387 213
rect -1445 -225 -1387 -213
rect -1327 213 -1269 225
rect -1327 -213 -1315 213
rect -1281 -213 -1269 213
rect -1327 -225 -1269 -213
rect -1209 213 -1151 225
rect -1209 -213 -1197 213
rect -1163 -213 -1151 213
rect -1209 -225 -1151 -213
rect -1091 213 -1033 225
rect -1091 -213 -1079 213
rect -1045 -213 -1033 213
rect -1091 -225 -1033 -213
rect -973 213 -915 225
rect -973 -213 -961 213
rect -927 -213 -915 213
rect -973 -225 -915 -213
rect -855 213 -797 225
rect -855 -213 -843 213
rect -809 -213 -797 213
rect -855 -225 -797 -213
rect -737 213 -679 225
rect -737 -213 -725 213
rect -691 -213 -679 213
rect -737 -225 -679 -213
rect -619 213 -561 225
rect -619 -213 -607 213
rect -573 -213 -561 213
rect -619 -225 -561 -213
rect -501 213 -443 225
rect -501 -213 -489 213
rect -455 -213 -443 213
rect -501 -225 -443 -213
rect -383 213 -325 225
rect -383 -213 -371 213
rect -337 -213 -325 213
rect -383 -225 -325 -213
rect -265 213 -207 225
rect -265 -213 -253 213
rect -219 -213 -207 213
rect -265 -225 -207 -213
rect -147 213 -89 225
rect -147 -213 -135 213
rect -101 -213 -89 213
rect -147 -225 -89 -213
rect -29 213 29 225
rect -29 -213 -17 213
rect 17 -213 29 213
rect -29 -225 29 -213
rect 89 213 147 225
rect 89 -213 101 213
rect 135 -213 147 213
rect 89 -225 147 -213
rect 207 213 265 225
rect 207 -213 219 213
rect 253 -213 265 213
rect 207 -225 265 -213
rect 325 213 383 225
rect 325 -213 337 213
rect 371 -213 383 213
rect 325 -225 383 -213
rect 443 213 501 225
rect 443 -213 455 213
rect 489 -213 501 213
rect 443 -225 501 -213
rect 561 213 619 225
rect 561 -213 573 213
rect 607 -213 619 213
rect 561 -225 619 -213
rect 679 213 737 225
rect 679 -213 691 213
rect 725 -213 737 213
rect 679 -225 737 -213
rect 797 213 855 225
rect 797 -213 809 213
rect 843 -213 855 213
rect 797 -225 855 -213
rect 915 213 973 225
rect 915 -213 927 213
rect 961 -213 973 213
rect 915 -225 973 -213
rect 1033 213 1091 225
rect 1033 -213 1045 213
rect 1079 -213 1091 213
rect 1033 -225 1091 -213
rect 1151 213 1209 225
rect 1151 -213 1163 213
rect 1197 -213 1209 213
rect 1151 -225 1209 -213
rect 1269 213 1327 225
rect 1269 -213 1281 213
rect 1315 -213 1327 213
rect 1269 -225 1327 -213
rect 1387 213 1445 225
rect 1387 -213 1399 213
rect 1433 -213 1445 213
rect 1387 -225 1445 -213
rect 1505 213 1563 225
rect 1505 -213 1517 213
rect 1551 -213 1563 213
rect 1505 -225 1563 -213
rect 1623 213 1681 225
rect 1623 -213 1635 213
rect 1669 -213 1681 213
rect 1623 -225 1681 -213
rect 1741 213 1799 225
rect 1741 -213 1753 213
rect 1787 -213 1799 213
rect 1741 -225 1799 -213
rect 1859 213 1917 225
rect 1859 -213 1871 213
rect 1905 -213 1917 213
rect 1859 -225 1917 -213
rect 1977 213 2035 225
rect 1977 -213 1989 213
rect 2023 -213 2035 213
rect 1977 -225 2035 -213
rect 2095 213 2153 225
rect 2095 -213 2107 213
rect 2141 -213 2153 213
rect 2095 -225 2153 -213
rect 2213 213 2271 225
rect 2213 -213 2225 213
rect 2259 -213 2271 213
rect 2213 -225 2271 -213
rect 2331 213 2389 225
rect 2331 -213 2343 213
rect 2377 -213 2389 213
rect 2331 -225 2389 -213
rect 2449 213 2507 225
rect 2449 -213 2461 213
rect 2495 -213 2507 213
rect 2449 -225 2507 -213
rect 2567 213 2625 225
rect 2567 -213 2579 213
rect 2613 -213 2625 213
rect 2567 -225 2625 -213
rect 2685 213 2743 225
rect 2685 -213 2697 213
rect 2731 -213 2743 213
rect 2685 -225 2743 -213
rect 2803 213 2861 225
rect 2803 -213 2815 213
rect 2849 -213 2861 213
rect 2803 -225 2861 -213
rect 2921 213 2979 225
rect 2921 -213 2933 213
rect 2967 -213 2979 213
rect 2921 -225 2979 -213
<< pdiffc >>
rect -2967 -213 -2933 213
rect -2849 -213 -2815 213
rect -2731 -213 -2697 213
rect -2613 -213 -2579 213
rect -2495 -213 -2461 213
rect -2377 -213 -2343 213
rect -2259 -213 -2225 213
rect -2141 -213 -2107 213
rect -2023 -213 -1989 213
rect -1905 -213 -1871 213
rect -1787 -213 -1753 213
rect -1669 -213 -1635 213
rect -1551 -213 -1517 213
rect -1433 -213 -1399 213
rect -1315 -213 -1281 213
rect -1197 -213 -1163 213
rect -1079 -213 -1045 213
rect -961 -213 -927 213
rect -843 -213 -809 213
rect -725 -213 -691 213
rect -607 -213 -573 213
rect -489 -213 -455 213
rect -371 -213 -337 213
rect -253 -213 -219 213
rect -135 -213 -101 213
rect -17 -213 17 213
rect 101 -213 135 213
rect 219 -213 253 213
rect 337 -213 371 213
rect 455 -213 489 213
rect 573 -213 607 213
rect 691 -213 725 213
rect 809 -213 843 213
rect 927 -213 961 213
rect 1045 -213 1079 213
rect 1163 -213 1197 213
rect 1281 -213 1315 213
rect 1399 -213 1433 213
rect 1517 -213 1551 213
rect 1635 -213 1669 213
rect 1753 -213 1787 213
rect 1871 -213 1905 213
rect 1989 -213 2023 213
rect 2107 -213 2141 213
rect 2225 -213 2259 213
rect 2343 -213 2377 213
rect 2461 -213 2495 213
rect 2579 -213 2613 213
rect 2697 -213 2731 213
rect 2815 -213 2849 213
rect 2933 -213 2967 213
<< nsubdiff >>
rect -3081 374 -2985 408
rect 2985 374 3081 408
rect -3081 312 -3047 374
rect 3047 312 3081 374
rect -3081 -374 -3047 -312
rect 3047 -374 3081 -312
rect -3081 -408 -2985 -374
rect 2985 -408 3081 -374
<< nsubdiffcont >>
rect -2985 374 2985 408
rect -3081 -312 -3047 312
rect 3047 -312 3081 312
rect -2985 -408 2985 -374
<< poly >>
rect -2924 306 -2858 322
rect -2924 272 -2908 306
rect -2874 272 -2858 306
rect -2924 256 -2858 272
rect -2806 306 -2740 322
rect -2806 272 -2790 306
rect -2756 272 -2740 306
rect -2806 256 -2740 272
rect -2688 306 -2622 322
rect -2688 272 -2672 306
rect -2638 272 -2622 306
rect -2688 256 -2622 272
rect -2570 306 -2504 322
rect -2570 272 -2554 306
rect -2520 272 -2504 306
rect -2570 256 -2504 272
rect -2452 306 -2386 322
rect -2452 272 -2436 306
rect -2402 272 -2386 306
rect -2452 256 -2386 272
rect -2334 306 -2268 322
rect -2334 272 -2318 306
rect -2284 272 -2268 306
rect -2334 256 -2268 272
rect -2216 306 -2150 322
rect -2216 272 -2200 306
rect -2166 272 -2150 306
rect -2216 256 -2150 272
rect -2098 306 -2032 322
rect -2098 272 -2082 306
rect -2048 272 -2032 306
rect -2098 256 -2032 272
rect -1980 306 -1914 322
rect -1980 272 -1964 306
rect -1930 272 -1914 306
rect -1980 256 -1914 272
rect -1862 306 -1796 322
rect -1862 272 -1846 306
rect -1812 272 -1796 306
rect -1862 256 -1796 272
rect -1744 306 -1678 322
rect -1744 272 -1728 306
rect -1694 272 -1678 306
rect -1744 256 -1678 272
rect -1626 306 -1560 322
rect -1626 272 -1610 306
rect -1576 272 -1560 306
rect -1626 256 -1560 272
rect -1508 306 -1442 322
rect -1508 272 -1492 306
rect -1458 272 -1442 306
rect -1508 256 -1442 272
rect -1390 306 -1324 322
rect -1390 272 -1374 306
rect -1340 272 -1324 306
rect -1390 256 -1324 272
rect -1272 306 -1206 322
rect -1272 272 -1256 306
rect -1222 272 -1206 306
rect -1272 256 -1206 272
rect -1154 306 -1088 322
rect -1154 272 -1138 306
rect -1104 272 -1088 306
rect -1154 256 -1088 272
rect -1036 306 -970 322
rect -1036 272 -1020 306
rect -986 272 -970 306
rect -1036 256 -970 272
rect -918 306 -852 322
rect -918 272 -902 306
rect -868 272 -852 306
rect -918 256 -852 272
rect -800 306 -734 322
rect -800 272 -784 306
rect -750 272 -734 306
rect -800 256 -734 272
rect -682 306 -616 322
rect -682 272 -666 306
rect -632 272 -616 306
rect -682 256 -616 272
rect -564 306 -498 322
rect -564 272 -548 306
rect -514 272 -498 306
rect -564 256 -498 272
rect -446 306 -380 322
rect -446 272 -430 306
rect -396 272 -380 306
rect -446 256 -380 272
rect -328 306 -262 322
rect -328 272 -312 306
rect -278 272 -262 306
rect -328 256 -262 272
rect -210 306 -144 322
rect -210 272 -194 306
rect -160 272 -144 306
rect -210 256 -144 272
rect -92 306 -26 322
rect -92 272 -76 306
rect -42 272 -26 306
rect -92 256 -26 272
rect 26 306 92 322
rect 26 272 42 306
rect 76 272 92 306
rect 26 256 92 272
rect 144 306 210 322
rect 144 272 160 306
rect 194 272 210 306
rect 144 256 210 272
rect 262 306 328 322
rect 262 272 278 306
rect 312 272 328 306
rect 262 256 328 272
rect 380 306 446 322
rect 380 272 396 306
rect 430 272 446 306
rect 380 256 446 272
rect 498 306 564 322
rect 498 272 514 306
rect 548 272 564 306
rect 498 256 564 272
rect 616 306 682 322
rect 616 272 632 306
rect 666 272 682 306
rect 616 256 682 272
rect 734 306 800 322
rect 734 272 750 306
rect 784 272 800 306
rect 734 256 800 272
rect 852 306 918 322
rect 852 272 868 306
rect 902 272 918 306
rect 852 256 918 272
rect 970 306 1036 322
rect 970 272 986 306
rect 1020 272 1036 306
rect 970 256 1036 272
rect 1088 306 1154 322
rect 1088 272 1104 306
rect 1138 272 1154 306
rect 1088 256 1154 272
rect 1206 306 1272 322
rect 1206 272 1222 306
rect 1256 272 1272 306
rect 1206 256 1272 272
rect 1324 306 1390 322
rect 1324 272 1340 306
rect 1374 272 1390 306
rect 1324 256 1390 272
rect 1442 306 1508 322
rect 1442 272 1458 306
rect 1492 272 1508 306
rect 1442 256 1508 272
rect 1560 306 1626 322
rect 1560 272 1576 306
rect 1610 272 1626 306
rect 1560 256 1626 272
rect 1678 306 1744 322
rect 1678 272 1694 306
rect 1728 272 1744 306
rect 1678 256 1744 272
rect 1796 306 1862 322
rect 1796 272 1812 306
rect 1846 272 1862 306
rect 1796 256 1862 272
rect 1914 306 1980 322
rect 1914 272 1930 306
rect 1964 272 1980 306
rect 1914 256 1980 272
rect 2032 306 2098 322
rect 2032 272 2048 306
rect 2082 272 2098 306
rect 2032 256 2098 272
rect 2150 306 2216 322
rect 2150 272 2166 306
rect 2200 272 2216 306
rect 2150 256 2216 272
rect 2268 306 2334 322
rect 2268 272 2284 306
rect 2318 272 2334 306
rect 2268 256 2334 272
rect 2386 306 2452 322
rect 2386 272 2402 306
rect 2436 272 2452 306
rect 2386 256 2452 272
rect 2504 306 2570 322
rect 2504 272 2520 306
rect 2554 272 2570 306
rect 2504 256 2570 272
rect 2622 306 2688 322
rect 2622 272 2638 306
rect 2672 272 2688 306
rect 2622 256 2688 272
rect 2740 306 2806 322
rect 2740 272 2756 306
rect 2790 272 2806 306
rect 2740 256 2806 272
rect 2858 306 2924 322
rect 2858 272 2874 306
rect 2908 272 2924 306
rect 2858 256 2924 272
rect -2921 225 -2861 256
rect -2803 225 -2743 256
rect -2685 225 -2625 256
rect -2567 225 -2507 256
rect -2449 225 -2389 256
rect -2331 225 -2271 256
rect -2213 225 -2153 256
rect -2095 225 -2035 256
rect -1977 225 -1917 256
rect -1859 225 -1799 256
rect -1741 225 -1681 256
rect -1623 225 -1563 256
rect -1505 225 -1445 256
rect -1387 225 -1327 256
rect -1269 225 -1209 256
rect -1151 225 -1091 256
rect -1033 225 -973 256
rect -915 225 -855 256
rect -797 225 -737 256
rect -679 225 -619 256
rect -561 225 -501 256
rect -443 225 -383 256
rect -325 225 -265 256
rect -207 225 -147 256
rect -89 225 -29 256
rect 29 225 89 256
rect 147 225 207 256
rect 265 225 325 256
rect 383 225 443 256
rect 501 225 561 256
rect 619 225 679 256
rect 737 225 797 256
rect 855 225 915 256
rect 973 225 1033 256
rect 1091 225 1151 256
rect 1209 225 1269 256
rect 1327 225 1387 256
rect 1445 225 1505 256
rect 1563 225 1623 256
rect 1681 225 1741 256
rect 1799 225 1859 256
rect 1917 225 1977 256
rect 2035 225 2095 256
rect 2153 225 2213 256
rect 2271 225 2331 256
rect 2389 225 2449 256
rect 2507 225 2567 256
rect 2625 225 2685 256
rect 2743 225 2803 256
rect 2861 225 2921 256
rect -2921 -256 -2861 -225
rect -2803 -256 -2743 -225
rect -2685 -256 -2625 -225
rect -2567 -256 -2507 -225
rect -2449 -256 -2389 -225
rect -2331 -256 -2271 -225
rect -2213 -256 -2153 -225
rect -2095 -256 -2035 -225
rect -1977 -256 -1917 -225
rect -1859 -256 -1799 -225
rect -1741 -256 -1681 -225
rect -1623 -256 -1563 -225
rect -1505 -256 -1445 -225
rect -1387 -256 -1327 -225
rect -1269 -256 -1209 -225
rect -1151 -256 -1091 -225
rect -1033 -256 -973 -225
rect -915 -256 -855 -225
rect -797 -256 -737 -225
rect -679 -256 -619 -225
rect -561 -256 -501 -225
rect -443 -256 -383 -225
rect -325 -256 -265 -225
rect -207 -256 -147 -225
rect -89 -256 -29 -225
rect 29 -256 89 -225
rect 147 -256 207 -225
rect 265 -256 325 -225
rect 383 -256 443 -225
rect 501 -256 561 -225
rect 619 -256 679 -225
rect 737 -256 797 -225
rect 855 -256 915 -225
rect 973 -256 1033 -225
rect 1091 -256 1151 -225
rect 1209 -256 1269 -225
rect 1327 -256 1387 -225
rect 1445 -256 1505 -225
rect 1563 -256 1623 -225
rect 1681 -256 1741 -225
rect 1799 -256 1859 -225
rect 1917 -256 1977 -225
rect 2035 -256 2095 -225
rect 2153 -256 2213 -225
rect 2271 -256 2331 -225
rect 2389 -256 2449 -225
rect 2507 -256 2567 -225
rect 2625 -256 2685 -225
rect 2743 -256 2803 -225
rect 2861 -256 2921 -225
rect -2924 -272 -2858 -256
rect -2924 -306 -2908 -272
rect -2874 -306 -2858 -272
rect -2924 -322 -2858 -306
rect -2806 -272 -2740 -256
rect -2806 -306 -2790 -272
rect -2756 -306 -2740 -272
rect -2806 -322 -2740 -306
rect -2688 -272 -2622 -256
rect -2688 -306 -2672 -272
rect -2638 -306 -2622 -272
rect -2688 -322 -2622 -306
rect -2570 -272 -2504 -256
rect -2570 -306 -2554 -272
rect -2520 -306 -2504 -272
rect -2570 -322 -2504 -306
rect -2452 -272 -2386 -256
rect -2452 -306 -2436 -272
rect -2402 -306 -2386 -272
rect -2452 -322 -2386 -306
rect -2334 -272 -2268 -256
rect -2334 -306 -2318 -272
rect -2284 -306 -2268 -272
rect -2334 -322 -2268 -306
rect -2216 -272 -2150 -256
rect -2216 -306 -2200 -272
rect -2166 -306 -2150 -272
rect -2216 -322 -2150 -306
rect -2098 -272 -2032 -256
rect -2098 -306 -2082 -272
rect -2048 -306 -2032 -272
rect -2098 -322 -2032 -306
rect -1980 -272 -1914 -256
rect -1980 -306 -1964 -272
rect -1930 -306 -1914 -272
rect -1980 -322 -1914 -306
rect -1862 -272 -1796 -256
rect -1862 -306 -1846 -272
rect -1812 -306 -1796 -272
rect -1862 -322 -1796 -306
rect -1744 -272 -1678 -256
rect -1744 -306 -1728 -272
rect -1694 -306 -1678 -272
rect -1744 -322 -1678 -306
rect -1626 -272 -1560 -256
rect -1626 -306 -1610 -272
rect -1576 -306 -1560 -272
rect -1626 -322 -1560 -306
rect -1508 -272 -1442 -256
rect -1508 -306 -1492 -272
rect -1458 -306 -1442 -272
rect -1508 -322 -1442 -306
rect -1390 -272 -1324 -256
rect -1390 -306 -1374 -272
rect -1340 -306 -1324 -272
rect -1390 -322 -1324 -306
rect -1272 -272 -1206 -256
rect -1272 -306 -1256 -272
rect -1222 -306 -1206 -272
rect -1272 -322 -1206 -306
rect -1154 -272 -1088 -256
rect -1154 -306 -1138 -272
rect -1104 -306 -1088 -272
rect -1154 -322 -1088 -306
rect -1036 -272 -970 -256
rect -1036 -306 -1020 -272
rect -986 -306 -970 -272
rect -1036 -322 -970 -306
rect -918 -272 -852 -256
rect -918 -306 -902 -272
rect -868 -306 -852 -272
rect -918 -322 -852 -306
rect -800 -272 -734 -256
rect -800 -306 -784 -272
rect -750 -306 -734 -272
rect -800 -322 -734 -306
rect -682 -272 -616 -256
rect -682 -306 -666 -272
rect -632 -306 -616 -272
rect -682 -322 -616 -306
rect -564 -272 -498 -256
rect -564 -306 -548 -272
rect -514 -306 -498 -272
rect -564 -322 -498 -306
rect -446 -272 -380 -256
rect -446 -306 -430 -272
rect -396 -306 -380 -272
rect -446 -322 -380 -306
rect -328 -272 -262 -256
rect -328 -306 -312 -272
rect -278 -306 -262 -272
rect -328 -322 -262 -306
rect -210 -272 -144 -256
rect -210 -306 -194 -272
rect -160 -306 -144 -272
rect -210 -322 -144 -306
rect -92 -272 -26 -256
rect -92 -306 -76 -272
rect -42 -306 -26 -272
rect -92 -322 -26 -306
rect 26 -272 92 -256
rect 26 -306 42 -272
rect 76 -306 92 -272
rect 26 -322 92 -306
rect 144 -272 210 -256
rect 144 -306 160 -272
rect 194 -306 210 -272
rect 144 -322 210 -306
rect 262 -272 328 -256
rect 262 -306 278 -272
rect 312 -306 328 -272
rect 262 -322 328 -306
rect 380 -272 446 -256
rect 380 -306 396 -272
rect 430 -306 446 -272
rect 380 -322 446 -306
rect 498 -272 564 -256
rect 498 -306 514 -272
rect 548 -306 564 -272
rect 498 -322 564 -306
rect 616 -272 682 -256
rect 616 -306 632 -272
rect 666 -306 682 -272
rect 616 -322 682 -306
rect 734 -272 800 -256
rect 734 -306 750 -272
rect 784 -306 800 -272
rect 734 -322 800 -306
rect 852 -272 918 -256
rect 852 -306 868 -272
rect 902 -306 918 -272
rect 852 -322 918 -306
rect 970 -272 1036 -256
rect 970 -306 986 -272
rect 1020 -306 1036 -272
rect 970 -322 1036 -306
rect 1088 -272 1154 -256
rect 1088 -306 1104 -272
rect 1138 -306 1154 -272
rect 1088 -322 1154 -306
rect 1206 -272 1272 -256
rect 1206 -306 1222 -272
rect 1256 -306 1272 -272
rect 1206 -322 1272 -306
rect 1324 -272 1390 -256
rect 1324 -306 1340 -272
rect 1374 -306 1390 -272
rect 1324 -322 1390 -306
rect 1442 -272 1508 -256
rect 1442 -306 1458 -272
rect 1492 -306 1508 -272
rect 1442 -322 1508 -306
rect 1560 -272 1626 -256
rect 1560 -306 1576 -272
rect 1610 -306 1626 -272
rect 1560 -322 1626 -306
rect 1678 -272 1744 -256
rect 1678 -306 1694 -272
rect 1728 -306 1744 -272
rect 1678 -322 1744 -306
rect 1796 -272 1862 -256
rect 1796 -306 1812 -272
rect 1846 -306 1862 -272
rect 1796 -322 1862 -306
rect 1914 -272 1980 -256
rect 1914 -306 1930 -272
rect 1964 -306 1980 -272
rect 1914 -322 1980 -306
rect 2032 -272 2098 -256
rect 2032 -306 2048 -272
rect 2082 -306 2098 -272
rect 2032 -322 2098 -306
rect 2150 -272 2216 -256
rect 2150 -306 2166 -272
rect 2200 -306 2216 -272
rect 2150 -322 2216 -306
rect 2268 -272 2334 -256
rect 2268 -306 2284 -272
rect 2318 -306 2334 -272
rect 2268 -322 2334 -306
rect 2386 -272 2452 -256
rect 2386 -306 2402 -272
rect 2436 -306 2452 -272
rect 2386 -322 2452 -306
rect 2504 -272 2570 -256
rect 2504 -306 2520 -272
rect 2554 -306 2570 -272
rect 2504 -322 2570 -306
rect 2622 -272 2688 -256
rect 2622 -306 2638 -272
rect 2672 -306 2688 -272
rect 2622 -322 2688 -306
rect 2740 -272 2806 -256
rect 2740 -306 2756 -272
rect 2790 -306 2806 -272
rect 2740 -322 2806 -306
rect 2858 -272 2924 -256
rect 2858 -306 2874 -272
rect 2908 -306 2924 -272
rect 2858 -322 2924 -306
<< polycont >>
rect -2908 272 -2874 306
rect -2790 272 -2756 306
rect -2672 272 -2638 306
rect -2554 272 -2520 306
rect -2436 272 -2402 306
rect -2318 272 -2284 306
rect -2200 272 -2166 306
rect -2082 272 -2048 306
rect -1964 272 -1930 306
rect -1846 272 -1812 306
rect -1728 272 -1694 306
rect -1610 272 -1576 306
rect -1492 272 -1458 306
rect -1374 272 -1340 306
rect -1256 272 -1222 306
rect -1138 272 -1104 306
rect -1020 272 -986 306
rect -902 272 -868 306
rect -784 272 -750 306
rect -666 272 -632 306
rect -548 272 -514 306
rect -430 272 -396 306
rect -312 272 -278 306
rect -194 272 -160 306
rect -76 272 -42 306
rect 42 272 76 306
rect 160 272 194 306
rect 278 272 312 306
rect 396 272 430 306
rect 514 272 548 306
rect 632 272 666 306
rect 750 272 784 306
rect 868 272 902 306
rect 986 272 1020 306
rect 1104 272 1138 306
rect 1222 272 1256 306
rect 1340 272 1374 306
rect 1458 272 1492 306
rect 1576 272 1610 306
rect 1694 272 1728 306
rect 1812 272 1846 306
rect 1930 272 1964 306
rect 2048 272 2082 306
rect 2166 272 2200 306
rect 2284 272 2318 306
rect 2402 272 2436 306
rect 2520 272 2554 306
rect 2638 272 2672 306
rect 2756 272 2790 306
rect 2874 272 2908 306
rect -2908 -306 -2874 -272
rect -2790 -306 -2756 -272
rect -2672 -306 -2638 -272
rect -2554 -306 -2520 -272
rect -2436 -306 -2402 -272
rect -2318 -306 -2284 -272
rect -2200 -306 -2166 -272
rect -2082 -306 -2048 -272
rect -1964 -306 -1930 -272
rect -1846 -306 -1812 -272
rect -1728 -306 -1694 -272
rect -1610 -306 -1576 -272
rect -1492 -306 -1458 -272
rect -1374 -306 -1340 -272
rect -1256 -306 -1222 -272
rect -1138 -306 -1104 -272
rect -1020 -306 -986 -272
rect -902 -306 -868 -272
rect -784 -306 -750 -272
rect -666 -306 -632 -272
rect -548 -306 -514 -272
rect -430 -306 -396 -272
rect -312 -306 -278 -272
rect -194 -306 -160 -272
rect -76 -306 -42 -272
rect 42 -306 76 -272
rect 160 -306 194 -272
rect 278 -306 312 -272
rect 396 -306 430 -272
rect 514 -306 548 -272
rect 632 -306 666 -272
rect 750 -306 784 -272
rect 868 -306 902 -272
rect 986 -306 1020 -272
rect 1104 -306 1138 -272
rect 1222 -306 1256 -272
rect 1340 -306 1374 -272
rect 1458 -306 1492 -272
rect 1576 -306 1610 -272
rect 1694 -306 1728 -272
rect 1812 -306 1846 -272
rect 1930 -306 1964 -272
rect 2048 -306 2082 -272
rect 2166 -306 2200 -272
rect 2284 -306 2318 -272
rect 2402 -306 2436 -272
rect 2520 -306 2554 -272
rect 2638 -306 2672 -272
rect 2756 -306 2790 -272
rect 2874 -306 2908 -272
<< locali >>
rect -3081 374 -2985 408
rect 2985 374 3081 408
rect -3081 312 -3047 374
rect 3047 312 3081 374
rect -2924 272 -2908 306
rect -2874 272 -2858 306
rect -2806 272 -2790 306
rect -2756 272 -2740 306
rect -2688 272 -2672 306
rect -2638 272 -2622 306
rect -2570 272 -2554 306
rect -2520 272 -2504 306
rect -2452 272 -2436 306
rect -2402 272 -2386 306
rect -2334 272 -2318 306
rect -2284 272 -2268 306
rect -2216 272 -2200 306
rect -2166 272 -2150 306
rect -2098 272 -2082 306
rect -2048 272 -2032 306
rect -1980 272 -1964 306
rect -1930 272 -1914 306
rect -1862 272 -1846 306
rect -1812 272 -1796 306
rect -1744 272 -1728 306
rect -1694 272 -1678 306
rect -1626 272 -1610 306
rect -1576 272 -1560 306
rect -1508 272 -1492 306
rect -1458 272 -1442 306
rect -1390 272 -1374 306
rect -1340 272 -1324 306
rect -1272 272 -1256 306
rect -1222 272 -1206 306
rect -1154 272 -1138 306
rect -1104 272 -1088 306
rect -1036 272 -1020 306
rect -986 272 -970 306
rect -918 272 -902 306
rect -868 272 -852 306
rect -800 272 -784 306
rect -750 272 -734 306
rect -682 272 -666 306
rect -632 272 -616 306
rect -564 272 -548 306
rect -514 272 -498 306
rect -446 272 -430 306
rect -396 272 -380 306
rect -328 272 -312 306
rect -278 272 -262 306
rect -210 272 -194 306
rect -160 272 -144 306
rect -92 272 -76 306
rect -42 272 -26 306
rect 26 272 42 306
rect 76 272 92 306
rect 144 272 160 306
rect 194 272 210 306
rect 262 272 278 306
rect 312 272 328 306
rect 380 272 396 306
rect 430 272 446 306
rect 498 272 514 306
rect 548 272 564 306
rect 616 272 632 306
rect 666 272 682 306
rect 734 272 750 306
rect 784 272 800 306
rect 852 272 868 306
rect 902 272 918 306
rect 970 272 986 306
rect 1020 272 1036 306
rect 1088 272 1104 306
rect 1138 272 1154 306
rect 1206 272 1222 306
rect 1256 272 1272 306
rect 1324 272 1340 306
rect 1374 272 1390 306
rect 1442 272 1458 306
rect 1492 272 1508 306
rect 1560 272 1576 306
rect 1610 272 1626 306
rect 1678 272 1694 306
rect 1728 272 1744 306
rect 1796 272 1812 306
rect 1846 272 1862 306
rect 1914 272 1930 306
rect 1964 272 1980 306
rect 2032 272 2048 306
rect 2082 272 2098 306
rect 2150 272 2166 306
rect 2200 272 2216 306
rect 2268 272 2284 306
rect 2318 272 2334 306
rect 2386 272 2402 306
rect 2436 272 2452 306
rect 2504 272 2520 306
rect 2554 272 2570 306
rect 2622 272 2638 306
rect 2672 272 2688 306
rect 2740 272 2756 306
rect 2790 272 2806 306
rect 2858 272 2874 306
rect 2908 272 2924 306
rect -2967 213 -2933 229
rect -2967 -229 -2933 -213
rect -2849 213 -2815 229
rect -2849 -229 -2815 -213
rect -2731 213 -2697 229
rect -2731 -229 -2697 -213
rect -2613 213 -2579 229
rect -2613 -229 -2579 -213
rect -2495 213 -2461 229
rect -2495 -229 -2461 -213
rect -2377 213 -2343 229
rect -2377 -229 -2343 -213
rect -2259 213 -2225 229
rect -2259 -229 -2225 -213
rect -2141 213 -2107 229
rect -2141 -229 -2107 -213
rect -2023 213 -1989 229
rect -2023 -229 -1989 -213
rect -1905 213 -1871 229
rect -1905 -229 -1871 -213
rect -1787 213 -1753 229
rect -1787 -229 -1753 -213
rect -1669 213 -1635 229
rect -1669 -229 -1635 -213
rect -1551 213 -1517 229
rect -1551 -229 -1517 -213
rect -1433 213 -1399 229
rect -1433 -229 -1399 -213
rect -1315 213 -1281 229
rect -1315 -229 -1281 -213
rect -1197 213 -1163 229
rect -1197 -229 -1163 -213
rect -1079 213 -1045 229
rect -1079 -229 -1045 -213
rect -961 213 -927 229
rect -961 -229 -927 -213
rect -843 213 -809 229
rect -843 -229 -809 -213
rect -725 213 -691 229
rect -725 -229 -691 -213
rect -607 213 -573 229
rect -607 -229 -573 -213
rect -489 213 -455 229
rect -489 -229 -455 -213
rect -371 213 -337 229
rect -371 -229 -337 -213
rect -253 213 -219 229
rect -253 -229 -219 -213
rect -135 213 -101 229
rect -135 -229 -101 -213
rect -17 213 17 229
rect -17 -229 17 -213
rect 101 213 135 229
rect 101 -229 135 -213
rect 219 213 253 229
rect 219 -229 253 -213
rect 337 213 371 229
rect 337 -229 371 -213
rect 455 213 489 229
rect 455 -229 489 -213
rect 573 213 607 229
rect 573 -229 607 -213
rect 691 213 725 229
rect 691 -229 725 -213
rect 809 213 843 229
rect 809 -229 843 -213
rect 927 213 961 229
rect 927 -229 961 -213
rect 1045 213 1079 229
rect 1045 -229 1079 -213
rect 1163 213 1197 229
rect 1163 -229 1197 -213
rect 1281 213 1315 229
rect 1281 -229 1315 -213
rect 1399 213 1433 229
rect 1399 -229 1433 -213
rect 1517 213 1551 229
rect 1517 -229 1551 -213
rect 1635 213 1669 229
rect 1635 -229 1669 -213
rect 1753 213 1787 229
rect 1753 -229 1787 -213
rect 1871 213 1905 229
rect 1871 -229 1905 -213
rect 1989 213 2023 229
rect 1989 -229 2023 -213
rect 2107 213 2141 229
rect 2107 -229 2141 -213
rect 2225 213 2259 229
rect 2225 -229 2259 -213
rect 2343 213 2377 229
rect 2343 -229 2377 -213
rect 2461 213 2495 229
rect 2461 -229 2495 -213
rect 2579 213 2613 229
rect 2579 -229 2613 -213
rect 2697 213 2731 229
rect 2697 -229 2731 -213
rect 2815 213 2849 229
rect 2815 -229 2849 -213
rect 2933 213 2967 229
rect 2933 -229 2967 -213
rect -2924 -306 -2908 -272
rect -2874 -306 -2858 -272
rect -2806 -306 -2790 -272
rect -2756 -306 -2740 -272
rect -2688 -306 -2672 -272
rect -2638 -306 -2622 -272
rect -2570 -306 -2554 -272
rect -2520 -306 -2504 -272
rect -2452 -306 -2436 -272
rect -2402 -306 -2386 -272
rect -2334 -306 -2318 -272
rect -2284 -306 -2268 -272
rect -2216 -306 -2200 -272
rect -2166 -306 -2150 -272
rect -2098 -306 -2082 -272
rect -2048 -306 -2032 -272
rect -1980 -306 -1964 -272
rect -1930 -306 -1914 -272
rect -1862 -306 -1846 -272
rect -1812 -306 -1796 -272
rect -1744 -306 -1728 -272
rect -1694 -306 -1678 -272
rect -1626 -306 -1610 -272
rect -1576 -306 -1560 -272
rect -1508 -306 -1492 -272
rect -1458 -306 -1442 -272
rect -1390 -306 -1374 -272
rect -1340 -306 -1324 -272
rect -1272 -306 -1256 -272
rect -1222 -306 -1206 -272
rect -1154 -306 -1138 -272
rect -1104 -306 -1088 -272
rect -1036 -306 -1020 -272
rect -986 -306 -970 -272
rect -918 -306 -902 -272
rect -868 -306 -852 -272
rect -800 -306 -784 -272
rect -750 -306 -734 -272
rect -682 -306 -666 -272
rect -632 -306 -616 -272
rect -564 -306 -548 -272
rect -514 -306 -498 -272
rect -446 -306 -430 -272
rect -396 -306 -380 -272
rect -328 -306 -312 -272
rect -278 -306 -262 -272
rect -210 -306 -194 -272
rect -160 -306 -144 -272
rect -92 -306 -76 -272
rect -42 -306 -26 -272
rect 26 -306 42 -272
rect 76 -306 92 -272
rect 144 -306 160 -272
rect 194 -306 210 -272
rect 262 -306 278 -272
rect 312 -306 328 -272
rect 380 -306 396 -272
rect 430 -306 446 -272
rect 498 -306 514 -272
rect 548 -306 564 -272
rect 616 -306 632 -272
rect 666 -306 682 -272
rect 734 -306 750 -272
rect 784 -306 800 -272
rect 852 -306 868 -272
rect 902 -306 918 -272
rect 970 -306 986 -272
rect 1020 -306 1036 -272
rect 1088 -306 1104 -272
rect 1138 -306 1154 -272
rect 1206 -306 1222 -272
rect 1256 -306 1272 -272
rect 1324 -306 1340 -272
rect 1374 -306 1390 -272
rect 1442 -306 1458 -272
rect 1492 -306 1508 -272
rect 1560 -306 1576 -272
rect 1610 -306 1626 -272
rect 1678 -306 1694 -272
rect 1728 -306 1744 -272
rect 1796 -306 1812 -272
rect 1846 -306 1862 -272
rect 1914 -306 1930 -272
rect 1964 -306 1980 -272
rect 2032 -306 2048 -272
rect 2082 -306 2098 -272
rect 2150 -306 2166 -272
rect 2200 -306 2216 -272
rect 2268 -306 2284 -272
rect 2318 -306 2334 -272
rect 2386 -306 2402 -272
rect 2436 -306 2452 -272
rect 2504 -306 2520 -272
rect 2554 -306 2570 -272
rect 2622 -306 2638 -272
rect 2672 -306 2688 -272
rect 2740 -306 2756 -272
rect 2790 -306 2806 -272
rect 2858 -306 2874 -272
rect 2908 -306 2924 -272
rect -3081 -374 -3047 -312
rect 3047 -374 3081 -312
rect -3081 -408 -2985 -374
rect 2985 -408 3081 -374
<< viali >>
rect -2908 272 -2874 306
rect -2790 272 -2756 306
rect -2672 272 -2638 306
rect -2554 272 -2520 306
rect -2436 272 -2402 306
rect -2318 272 -2284 306
rect -2200 272 -2166 306
rect -2082 272 -2048 306
rect -1964 272 -1930 306
rect -1846 272 -1812 306
rect -1728 272 -1694 306
rect -1610 272 -1576 306
rect -1492 272 -1458 306
rect -1374 272 -1340 306
rect -1256 272 -1222 306
rect -1138 272 -1104 306
rect -1020 272 -986 306
rect -902 272 -868 306
rect -784 272 -750 306
rect -666 272 -632 306
rect -548 272 -514 306
rect -430 272 -396 306
rect -312 272 -278 306
rect -194 272 -160 306
rect -76 272 -42 306
rect 42 272 76 306
rect 160 272 194 306
rect 278 272 312 306
rect 396 272 430 306
rect 514 272 548 306
rect 632 272 666 306
rect 750 272 784 306
rect 868 272 902 306
rect 986 272 1020 306
rect 1104 272 1138 306
rect 1222 272 1256 306
rect 1340 272 1374 306
rect 1458 272 1492 306
rect 1576 272 1610 306
rect 1694 272 1728 306
rect 1812 272 1846 306
rect 1930 272 1964 306
rect 2048 272 2082 306
rect 2166 272 2200 306
rect 2284 272 2318 306
rect 2402 272 2436 306
rect 2520 272 2554 306
rect 2638 272 2672 306
rect 2756 272 2790 306
rect 2874 272 2908 306
rect -2967 -213 -2933 213
rect -2849 -213 -2815 213
rect -2731 -213 -2697 213
rect -2613 -213 -2579 213
rect -2495 -213 -2461 213
rect -2377 -213 -2343 213
rect -2259 -213 -2225 213
rect -2141 -213 -2107 213
rect -2023 -213 -1989 213
rect -1905 -213 -1871 213
rect -1787 -213 -1753 213
rect -1669 -213 -1635 213
rect -1551 -213 -1517 213
rect -1433 -213 -1399 213
rect -1315 -213 -1281 213
rect -1197 -213 -1163 213
rect -1079 -213 -1045 213
rect -961 -213 -927 213
rect -843 -213 -809 213
rect -725 -213 -691 213
rect -607 -213 -573 213
rect -489 -213 -455 213
rect -371 -213 -337 213
rect -253 -213 -219 213
rect -135 -213 -101 213
rect -17 -213 17 213
rect 101 -213 135 213
rect 219 -213 253 213
rect 337 -213 371 213
rect 455 -213 489 213
rect 573 -213 607 213
rect 691 -213 725 213
rect 809 -213 843 213
rect 927 -213 961 213
rect 1045 -213 1079 213
rect 1163 -213 1197 213
rect 1281 -213 1315 213
rect 1399 -213 1433 213
rect 1517 -213 1551 213
rect 1635 -213 1669 213
rect 1753 -213 1787 213
rect 1871 -213 1905 213
rect 1989 -213 2023 213
rect 2107 -213 2141 213
rect 2225 -213 2259 213
rect 2343 -213 2377 213
rect 2461 -213 2495 213
rect 2579 -213 2613 213
rect 2697 -213 2731 213
rect 2815 -213 2849 213
rect 2933 -213 2967 213
rect -2908 -306 -2874 -272
rect -2790 -306 -2756 -272
rect -2672 -306 -2638 -272
rect -2554 -306 -2520 -272
rect -2436 -306 -2402 -272
rect -2318 -306 -2284 -272
rect -2200 -306 -2166 -272
rect -2082 -306 -2048 -272
rect -1964 -306 -1930 -272
rect -1846 -306 -1812 -272
rect -1728 -306 -1694 -272
rect -1610 -306 -1576 -272
rect -1492 -306 -1458 -272
rect -1374 -306 -1340 -272
rect -1256 -306 -1222 -272
rect -1138 -306 -1104 -272
rect -1020 -306 -986 -272
rect -902 -306 -868 -272
rect -784 -306 -750 -272
rect -666 -306 -632 -272
rect -548 -306 -514 -272
rect -430 -306 -396 -272
rect -312 -306 -278 -272
rect -194 -306 -160 -272
rect -76 -306 -42 -272
rect 42 -306 76 -272
rect 160 -306 194 -272
rect 278 -306 312 -272
rect 396 -306 430 -272
rect 514 -306 548 -272
rect 632 -306 666 -272
rect 750 -306 784 -272
rect 868 -306 902 -272
rect 986 -306 1020 -272
rect 1104 -306 1138 -272
rect 1222 -306 1256 -272
rect 1340 -306 1374 -272
rect 1458 -306 1492 -272
rect 1576 -306 1610 -272
rect 1694 -306 1728 -272
rect 1812 -306 1846 -272
rect 1930 -306 1964 -272
rect 2048 -306 2082 -272
rect 2166 -306 2200 -272
rect 2284 -306 2318 -272
rect 2402 -306 2436 -272
rect 2520 -306 2554 -272
rect 2638 -306 2672 -272
rect 2756 -306 2790 -272
rect 2874 -306 2908 -272
<< metal1 >>
rect -2920 306 -2862 312
rect -2920 272 -2908 306
rect -2874 272 -2862 306
rect -2920 266 -2862 272
rect -2802 306 -2744 312
rect -2802 272 -2790 306
rect -2756 272 -2744 306
rect -2802 266 -2744 272
rect -2684 306 -2626 312
rect -2684 272 -2672 306
rect -2638 272 -2626 306
rect -2684 266 -2626 272
rect -2566 306 -2508 312
rect -2566 272 -2554 306
rect -2520 272 -2508 306
rect -2566 266 -2508 272
rect -2448 306 -2390 312
rect -2448 272 -2436 306
rect -2402 272 -2390 306
rect -2448 266 -2390 272
rect -2330 306 -2272 312
rect -2330 272 -2318 306
rect -2284 272 -2272 306
rect -2330 266 -2272 272
rect -2212 306 -2154 312
rect -2212 272 -2200 306
rect -2166 272 -2154 306
rect -2212 266 -2154 272
rect -2094 306 -2036 312
rect -2094 272 -2082 306
rect -2048 272 -2036 306
rect -2094 266 -2036 272
rect -1976 306 -1918 312
rect -1976 272 -1964 306
rect -1930 272 -1918 306
rect -1976 266 -1918 272
rect -1858 306 -1800 312
rect -1858 272 -1846 306
rect -1812 272 -1800 306
rect -1858 266 -1800 272
rect -1740 306 -1682 312
rect -1740 272 -1728 306
rect -1694 272 -1682 306
rect -1740 266 -1682 272
rect -1622 306 -1564 312
rect -1622 272 -1610 306
rect -1576 272 -1564 306
rect -1622 266 -1564 272
rect -1504 306 -1446 312
rect -1504 272 -1492 306
rect -1458 272 -1446 306
rect -1504 266 -1446 272
rect -1386 306 -1328 312
rect -1386 272 -1374 306
rect -1340 272 -1328 306
rect -1386 266 -1328 272
rect -1268 306 -1210 312
rect -1268 272 -1256 306
rect -1222 272 -1210 306
rect -1268 266 -1210 272
rect -1150 306 -1092 312
rect -1150 272 -1138 306
rect -1104 272 -1092 306
rect -1150 266 -1092 272
rect -1032 306 -974 312
rect -1032 272 -1020 306
rect -986 272 -974 306
rect -1032 266 -974 272
rect -914 306 -856 312
rect -914 272 -902 306
rect -868 272 -856 306
rect -914 266 -856 272
rect -796 306 -738 312
rect -796 272 -784 306
rect -750 272 -738 306
rect -796 266 -738 272
rect -678 306 -620 312
rect -678 272 -666 306
rect -632 272 -620 306
rect -678 266 -620 272
rect -560 306 -502 312
rect -560 272 -548 306
rect -514 272 -502 306
rect -560 266 -502 272
rect -442 306 -384 312
rect -442 272 -430 306
rect -396 272 -384 306
rect -442 266 -384 272
rect -324 306 -266 312
rect -324 272 -312 306
rect -278 272 -266 306
rect -324 266 -266 272
rect -206 306 -148 312
rect -206 272 -194 306
rect -160 272 -148 306
rect -206 266 -148 272
rect -88 306 -30 312
rect -88 272 -76 306
rect -42 272 -30 306
rect -88 266 -30 272
rect 30 306 88 312
rect 30 272 42 306
rect 76 272 88 306
rect 30 266 88 272
rect 148 306 206 312
rect 148 272 160 306
rect 194 272 206 306
rect 148 266 206 272
rect 266 306 324 312
rect 266 272 278 306
rect 312 272 324 306
rect 266 266 324 272
rect 384 306 442 312
rect 384 272 396 306
rect 430 272 442 306
rect 384 266 442 272
rect 502 306 560 312
rect 502 272 514 306
rect 548 272 560 306
rect 502 266 560 272
rect 620 306 678 312
rect 620 272 632 306
rect 666 272 678 306
rect 620 266 678 272
rect 738 306 796 312
rect 738 272 750 306
rect 784 272 796 306
rect 738 266 796 272
rect 856 306 914 312
rect 856 272 868 306
rect 902 272 914 306
rect 856 266 914 272
rect 974 306 1032 312
rect 974 272 986 306
rect 1020 272 1032 306
rect 974 266 1032 272
rect 1092 306 1150 312
rect 1092 272 1104 306
rect 1138 272 1150 306
rect 1092 266 1150 272
rect 1210 306 1268 312
rect 1210 272 1222 306
rect 1256 272 1268 306
rect 1210 266 1268 272
rect 1328 306 1386 312
rect 1328 272 1340 306
rect 1374 272 1386 306
rect 1328 266 1386 272
rect 1446 306 1504 312
rect 1446 272 1458 306
rect 1492 272 1504 306
rect 1446 266 1504 272
rect 1564 306 1622 312
rect 1564 272 1576 306
rect 1610 272 1622 306
rect 1564 266 1622 272
rect 1682 306 1740 312
rect 1682 272 1694 306
rect 1728 272 1740 306
rect 1682 266 1740 272
rect 1800 306 1858 312
rect 1800 272 1812 306
rect 1846 272 1858 306
rect 1800 266 1858 272
rect 1918 306 1976 312
rect 1918 272 1930 306
rect 1964 272 1976 306
rect 1918 266 1976 272
rect 2036 306 2094 312
rect 2036 272 2048 306
rect 2082 272 2094 306
rect 2036 266 2094 272
rect 2154 306 2212 312
rect 2154 272 2166 306
rect 2200 272 2212 306
rect 2154 266 2212 272
rect 2272 306 2330 312
rect 2272 272 2284 306
rect 2318 272 2330 306
rect 2272 266 2330 272
rect 2390 306 2448 312
rect 2390 272 2402 306
rect 2436 272 2448 306
rect 2390 266 2448 272
rect 2508 306 2566 312
rect 2508 272 2520 306
rect 2554 272 2566 306
rect 2508 266 2566 272
rect 2626 306 2684 312
rect 2626 272 2638 306
rect 2672 272 2684 306
rect 2626 266 2684 272
rect 2744 306 2802 312
rect 2744 272 2756 306
rect 2790 272 2802 306
rect 2744 266 2802 272
rect 2862 306 2920 312
rect 2862 272 2874 306
rect 2908 272 2920 306
rect 2862 266 2920 272
rect -2973 213 -2927 225
rect -2973 -213 -2967 213
rect -2933 -213 -2927 213
rect -2973 -225 -2927 -213
rect -2855 213 -2809 225
rect -2855 -213 -2849 213
rect -2815 -213 -2809 213
rect -2855 -225 -2809 -213
rect -2737 213 -2691 225
rect -2737 -213 -2731 213
rect -2697 -213 -2691 213
rect -2737 -225 -2691 -213
rect -2619 213 -2573 225
rect -2619 -213 -2613 213
rect -2579 -213 -2573 213
rect -2619 -225 -2573 -213
rect -2501 213 -2455 225
rect -2501 -213 -2495 213
rect -2461 -213 -2455 213
rect -2501 -225 -2455 -213
rect -2383 213 -2337 225
rect -2383 -213 -2377 213
rect -2343 -213 -2337 213
rect -2383 -225 -2337 -213
rect -2265 213 -2219 225
rect -2265 -213 -2259 213
rect -2225 -213 -2219 213
rect -2265 -225 -2219 -213
rect -2147 213 -2101 225
rect -2147 -213 -2141 213
rect -2107 -213 -2101 213
rect -2147 -225 -2101 -213
rect -2029 213 -1983 225
rect -2029 -213 -2023 213
rect -1989 -213 -1983 213
rect -2029 -225 -1983 -213
rect -1911 213 -1865 225
rect -1911 -213 -1905 213
rect -1871 -213 -1865 213
rect -1911 -225 -1865 -213
rect -1793 213 -1747 225
rect -1793 -213 -1787 213
rect -1753 -213 -1747 213
rect -1793 -225 -1747 -213
rect -1675 213 -1629 225
rect -1675 -213 -1669 213
rect -1635 -213 -1629 213
rect -1675 -225 -1629 -213
rect -1557 213 -1511 225
rect -1557 -213 -1551 213
rect -1517 -213 -1511 213
rect -1557 -225 -1511 -213
rect -1439 213 -1393 225
rect -1439 -213 -1433 213
rect -1399 -213 -1393 213
rect -1439 -225 -1393 -213
rect -1321 213 -1275 225
rect -1321 -213 -1315 213
rect -1281 -213 -1275 213
rect -1321 -225 -1275 -213
rect -1203 213 -1157 225
rect -1203 -213 -1197 213
rect -1163 -213 -1157 213
rect -1203 -225 -1157 -213
rect -1085 213 -1039 225
rect -1085 -213 -1079 213
rect -1045 -213 -1039 213
rect -1085 -225 -1039 -213
rect -967 213 -921 225
rect -967 -213 -961 213
rect -927 -213 -921 213
rect -967 -225 -921 -213
rect -849 213 -803 225
rect -849 -213 -843 213
rect -809 -213 -803 213
rect -849 -225 -803 -213
rect -731 213 -685 225
rect -731 -213 -725 213
rect -691 -213 -685 213
rect -731 -225 -685 -213
rect -613 213 -567 225
rect -613 -213 -607 213
rect -573 -213 -567 213
rect -613 -225 -567 -213
rect -495 213 -449 225
rect -495 -213 -489 213
rect -455 -213 -449 213
rect -495 -225 -449 -213
rect -377 213 -331 225
rect -377 -213 -371 213
rect -337 -213 -331 213
rect -377 -225 -331 -213
rect -259 213 -213 225
rect -259 -213 -253 213
rect -219 -213 -213 213
rect -259 -225 -213 -213
rect -141 213 -95 225
rect -141 -213 -135 213
rect -101 -213 -95 213
rect -141 -225 -95 -213
rect -23 213 23 225
rect -23 -213 -17 213
rect 17 -213 23 213
rect -23 -225 23 -213
rect 95 213 141 225
rect 95 -213 101 213
rect 135 -213 141 213
rect 95 -225 141 -213
rect 213 213 259 225
rect 213 -213 219 213
rect 253 -213 259 213
rect 213 -225 259 -213
rect 331 213 377 225
rect 331 -213 337 213
rect 371 -213 377 213
rect 331 -225 377 -213
rect 449 213 495 225
rect 449 -213 455 213
rect 489 -213 495 213
rect 449 -225 495 -213
rect 567 213 613 225
rect 567 -213 573 213
rect 607 -213 613 213
rect 567 -225 613 -213
rect 685 213 731 225
rect 685 -213 691 213
rect 725 -213 731 213
rect 685 -225 731 -213
rect 803 213 849 225
rect 803 -213 809 213
rect 843 -213 849 213
rect 803 -225 849 -213
rect 921 213 967 225
rect 921 -213 927 213
rect 961 -213 967 213
rect 921 -225 967 -213
rect 1039 213 1085 225
rect 1039 -213 1045 213
rect 1079 -213 1085 213
rect 1039 -225 1085 -213
rect 1157 213 1203 225
rect 1157 -213 1163 213
rect 1197 -213 1203 213
rect 1157 -225 1203 -213
rect 1275 213 1321 225
rect 1275 -213 1281 213
rect 1315 -213 1321 213
rect 1275 -225 1321 -213
rect 1393 213 1439 225
rect 1393 -213 1399 213
rect 1433 -213 1439 213
rect 1393 -225 1439 -213
rect 1511 213 1557 225
rect 1511 -213 1517 213
rect 1551 -213 1557 213
rect 1511 -225 1557 -213
rect 1629 213 1675 225
rect 1629 -213 1635 213
rect 1669 -213 1675 213
rect 1629 -225 1675 -213
rect 1747 213 1793 225
rect 1747 -213 1753 213
rect 1787 -213 1793 213
rect 1747 -225 1793 -213
rect 1865 213 1911 225
rect 1865 -213 1871 213
rect 1905 -213 1911 213
rect 1865 -225 1911 -213
rect 1983 213 2029 225
rect 1983 -213 1989 213
rect 2023 -213 2029 213
rect 1983 -225 2029 -213
rect 2101 213 2147 225
rect 2101 -213 2107 213
rect 2141 -213 2147 213
rect 2101 -225 2147 -213
rect 2219 213 2265 225
rect 2219 -213 2225 213
rect 2259 -213 2265 213
rect 2219 -225 2265 -213
rect 2337 213 2383 225
rect 2337 -213 2343 213
rect 2377 -213 2383 213
rect 2337 -225 2383 -213
rect 2455 213 2501 225
rect 2455 -213 2461 213
rect 2495 -213 2501 213
rect 2455 -225 2501 -213
rect 2573 213 2619 225
rect 2573 -213 2579 213
rect 2613 -213 2619 213
rect 2573 -225 2619 -213
rect 2691 213 2737 225
rect 2691 -213 2697 213
rect 2731 -213 2737 213
rect 2691 -225 2737 -213
rect 2809 213 2855 225
rect 2809 -213 2815 213
rect 2849 -213 2855 213
rect 2809 -225 2855 -213
rect 2927 213 2973 225
rect 2927 -213 2933 213
rect 2967 -213 2973 213
rect 2927 -225 2973 -213
rect -2920 -272 -2862 -266
rect -2920 -306 -2908 -272
rect -2874 -306 -2862 -272
rect -2920 -312 -2862 -306
rect -2802 -272 -2744 -266
rect -2802 -306 -2790 -272
rect -2756 -306 -2744 -272
rect -2802 -312 -2744 -306
rect -2684 -272 -2626 -266
rect -2684 -306 -2672 -272
rect -2638 -306 -2626 -272
rect -2684 -312 -2626 -306
rect -2566 -272 -2508 -266
rect -2566 -306 -2554 -272
rect -2520 -306 -2508 -272
rect -2566 -312 -2508 -306
rect -2448 -272 -2390 -266
rect -2448 -306 -2436 -272
rect -2402 -306 -2390 -272
rect -2448 -312 -2390 -306
rect -2330 -272 -2272 -266
rect -2330 -306 -2318 -272
rect -2284 -306 -2272 -272
rect -2330 -312 -2272 -306
rect -2212 -272 -2154 -266
rect -2212 -306 -2200 -272
rect -2166 -306 -2154 -272
rect -2212 -312 -2154 -306
rect -2094 -272 -2036 -266
rect -2094 -306 -2082 -272
rect -2048 -306 -2036 -272
rect -2094 -312 -2036 -306
rect -1976 -272 -1918 -266
rect -1976 -306 -1964 -272
rect -1930 -306 -1918 -272
rect -1976 -312 -1918 -306
rect -1858 -272 -1800 -266
rect -1858 -306 -1846 -272
rect -1812 -306 -1800 -272
rect -1858 -312 -1800 -306
rect -1740 -272 -1682 -266
rect -1740 -306 -1728 -272
rect -1694 -306 -1682 -272
rect -1740 -312 -1682 -306
rect -1622 -272 -1564 -266
rect -1622 -306 -1610 -272
rect -1576 -306 -1564 -272
rect -1622 -312 -1564 -306
rect -1504 -272 -1446 -266
rect -1504 -306 -1492 -272
rect -1458 -306 -1446 -272
rect -1504 -312 -1446 -306
rect -1386 -272 -1328 -266
rect -1386 -306 -1374 -272
rect -1340 -306 -1328 -272
rect -1386 -312 -1328 -306
rect -1268 -272 -1210 -266
rect -1268 -306 -1256 -272
rect -1222 -306 -1210 -272
rect -1268 -312 -1210 -306
rect -1150 -272 -1092 -266
rect -1150 -306 -1138 -272
rect -1104 -306 -1092 -272
rect -1150 -312 -1092 -306
rect -1032 -272 -974 -266
rect -1032 -306 -1020 -272
rect -986 -306 -974 -272
rect -1032 -312 -974 -306
rect -914 -272 -856 -266
rect -914 -306 -902 -272
rect -868 -306 -856 -272
rect -914 -312 -856 -306
rect -796 -272 -738 -266
rect -796 -306 -784 -272
rect -750 -306 -738 -272
rect -796 -312 -738 -306
rect -678 -272 -620 -266
rect -678 -306 -666 -272
rect -632 -306 -620 -272
rect -678 -312 -620 -306
rect -560 -272 -502 -266
rect -560 -306 -548 -272
rect -514 -306 -502 -272
rect -560 -312 -502 -306
rect -442 -272 -384 -266
rect -442 -306 -430 -272
rect -396 -306 -384 -272
rect -442 -312 -384 -306
rect -324 -272 -266 -266
rect -324 -306 -312 -272
rect -278 -306 -266 -272
rect -324 -312 -266 -306
rect -206 -272 -148 -266
rect -206 -306 -194 -272
rect -160 -306 -148 -272
rect -206 -312 -148 -306
rect -88 -272 -30 -266
rect -88 -306 -76 -272
rect -42 -306 -30 -272
rect -88 -312 -30 -306
rect 30 -272 88 -266
rect 30 -306 42 -272
rect 76 -306 88 -272
rect 30 -312 88 -306
rect 148 -272 206 -266
rect 148 -306 160 -272
rect 194 -306 206 -272
rect 148 -312 206 -306
rect 266 -272 324 -266
rect 266 -306 278 -272
rect 312 -306 324 -272
rect 266 -312 324 -306
rect 384 -272 442 -266
rect 384 -306 396 -272
rect 430 -306 442 -272
rect 384 -312 442 -306
rect 502 -272 560 -266
rect 502 -306 514 -272
rect 548 -306 560 -272
rect 502 -312 560 -306
rect 620 -272 678 -266
rect 620 -306 632 -272
rect 666 -306 678 -272
rect 620 -312 678 -306
rect 738 -272 796 -266
rect 738 -306 750 -272
rect 784 -306 796 -272
rect 738 -312 796 -306
rect 856 -272 914 -266
rect 856 -306 868 -272
rect 902 -306 914 -272
rect 856 -312 914 -306
rect 974 -272 1032 -266
rect 974 -306 986 -272
rect 1020 -306 1032 -272
rect 974 -312 1032 -306
rect 1092 -272 1150 -266
rect 1092 -306 1104 -272
rect 1138 -306 1150 -272
rect 1092 -312 1150 -306
rect 1210 -272 1268 -266
rect 1210 -306 1222 -272
rect 1256 -306 1268 -272
rect 1210 -312 1268 -306
rect 1328 -272 1386 -266
rect 1328 -306 1340 -272
rect 1374 -306 1386 -272
rect 1328 -312 1386 -306
rect 1446 -272 1504 -266
rect 1446 -306 1458 -272
rect 1492 -306 1504 -272
rect 1446 -312 1504 -306
rect 1564 -272 1622 -266
rect 1564 -306 1576 -272
rect 1610 -306 1622 -272
rect 1564 -312 1622 -306
rect 1682 -272 1740 -266
rect 1682 -306 1694 -272
rect 1728 -306 1740 -272
rect 1682 -312 1740 -306
rect 1800 -272 1858 -266
rect 1800 -306 1812 -272
rect 1846 -306 1858 -272
rect 1800 -312 1858 -306
rect 1918 -272 1976 -266
rect 1918 -306 1930 -272
rect 1964 -306 1976 -272
rect 1918 -312 1976 -306
rect 2036 -272 2094 -266
rect 2036 -306 2048 -272
rect 2082 -306 2094 -272
rect 2036 -312 2094 -306
rect 2154 -272 2212 -266
rect 2154 -306 2166 -272
rect 2200 -306 2212 -272
rect 2154 -312 2212 -306
rect 2272 -272 2330 -266
rect 2272 -306 2284 -272
rect 2318 -306 2330 -272
rect 2272 -312 2330 -306
rect 2390 -272 2448 -266
rect 2390 -306 2402 -272
rect 2436 -306 2448 -272
rect 2390 -312 2448 -306
rect 2508 -272 2566 -266
rect 2508 -306 2520 -272
rect 2554 -306 2566 -272
rect 2508 -312 2566 -306
rect 2626 -272 2684 -266
rect 2626 -306 2638 -272
rect 2672 -306 2684 -272
rect 2626 -312 2684 -306
rect 2744 -272 2802 -266
rect 2744 -306 2756 -272
rect 2790 -306 2802 -272
rect 2744 -312 2802 -306
rect 2862 -272 2920 -266
rect 2862 -306 2874 -272
rect 2908 -306 2920 -272
rect 2862 -312 2920 -306
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -391 3064 391
string parameters w 2.25 l 0.3 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
