magic
tech sky130A
magscale 1 2
timestamp 1619358404
<< error_p >>
rect -1730 1700 -1670 4900
rect -1650 1700 -1590 4900
rect 1589 1700 1649 4900
rect 1669 1700 1729 4900
rect -1730 -1600 -1670 1600
rect -1650 -1600 -1590 1600
rect 1589 -1600 1649 1600
rect 1669 -1600 1729 1600
rect -1730 -4900 -1670 -1700
rect -1650 -4900 -1590 -1700
rect 1589 -4900 1649 -1700
rect 1669 -4900 1729 -1700
<< metal3 >>
rect -4969 4872 -1670 4900
rect -4969 1728 -1754 4872
rect -1690 1728 -1670 4872
rect -4969 1700 -1670 1728
rect -1650 4872 1649 4900
rect -1650 1728 1565 4872
rect 1629 1728 1649 4872
rect -1650 1700 1649 1728
rect 1669 4872 4968 4900
rect 1669 1728 4884 4872
rect 4948 1728 4968 4872
rect 1669 1700 4968 1728
rect -4969 1572 -1670 1600
rect -4969 -1572 -1754 1572
rect -1690 -1572 -1670 1572
rect -4969 -1600 -1670 -1572
rect -1650 1572 1649 1600
rect -1650 -1572 1565 1572
rect 1629 -1572 1649 1572
rect -1650 -1600 1649 -1572
rect 1669 1572 4968 1600
rect 1669 -1572 4884 1572
rect 4948 -1572 4968 1572
rect 1669 -1600 4968 -1572
rect -4969 -1728 -1670 -1700
rect -4969 -4872 -1754 -1728
rect -1690 -4872 -1670 -1728
rect -4969 -4900 -1670 -4872
rect -1650 -1728 1649 -1700
rect -1650 -4872 1565 -1728
rect 1629 -4872 1649 -1728
rect -1650 -4900 1649 -4872
rect 1669 -1728 4968 -1700
rect 1669 -4872 4884 -1728
rect 4948 -4872 4968 -1728
rect 1669 -4900 4968 -4872
<< via3 >>
rect -1754 1728 -1690 4872
rect 1565 1728 1629 4872
rect 4884 1728 4948 4872
rect -1754 -1572 -1690 1572
rect 1565 -1572 1629 1572
rect 4884 -1572 4948 1572
rect -1754 -4872 -1690 -1728
rect 1565 -4872 1629 -1728
rect 4884 -4872 4948 -1728
<< mimcap >>
rect -4869 4760 -1869 4800
rect -4869 1840 -4829 4760
rect -1909 1840 -1869 4760
rect -4869 1800 -1869 1840
rect -1550 4760 1450 4800
rect -1550 1840 -1510 4760
rect 1410 1840 1450 4760
rect -1550 1800 1450 1840
rect 1769 4760 4769 4800
rect 1769 1840 1809 4760
rect 4729 1840 4769 4760
rect 1769 1800 4769 1840
rect -4869 1460 -1869 1500
rect -4869 -1460 -4829 1460
rect -1909 -1460 -1869 1460
rect -4869 -1500 -1869 -1460
rect -1550 1460 1450 1500
rect -1550 -1460 -1510 1460
rect 1410 -1460 1450 1460
rect -1550 -1500 1450 -1460
rect 1769 1460 4769 1500
rect 1769 -1460 1809 1460
rect 4729 -1460 4769 1460
rect 1769 -1500 4769 -1460
rect -4869 -1840 -1869 -1800
rect -4869 -4760 -4829 -1840
rect -1909 -4760 -1869 -1840
rect -4869 -4800 -1869 -4760
rect -1550 -1840 1450 -1800
rect -1550 -4760 -1510 -1840
rect 1410 -4760 1450 -1840
rect -1550 -4800 1450 -4760
rect 1769 -1840 4769 -1800
rect 1769 -4760 1809 -1840
rect 4729 -4760 4769 -1840
rect 1769 -4800 4769 -4760
<< mimcapcontact >>
rect -4829 1840 -1909 4760
rect -1510 1840 1410 4760
rect 1809 1840 4729 4760
rect -4829 -1460 -1909 1460
rect -1510 -1460 1410 1460
rect 1809 -1460 4729 1460
rect -4829 -4760 -1909 -1840
rect -1510 -4760 1410 -1840
rect 1809 -4760 4729 -1840
<< metal4 >>
rect -1770 4872 -1674 4888
rect -4830 4760 -1908 4761
rect -4830 1840 -4829 4760
rect -1909 1840 -1908 4760
rect -4830 1839 -1908 1840
rect -1770 1728 -1754 4872
rect -1690 1728 -1674 4872
rect 1549 4872 1645 4888
rect -1511 4760 1411 4761
rect -1511 1840 -1510 4760
rect 1410 1840 1411 4760
rect -1511 1839 1411 1840
rect -1770 1712 -1674 1728
rect 1549 1728 1565 4872
rect 1629 1728 1645 4872
rect 4868 4872 4964 4888
rect 1808 4760 4730 4761
rect 1808 1840 1809 4760
rect 4729 1840 4730 4760
rect 1808 1839 4730 1840
rect 1549 1712 1645 1728
rect 4868 1728 4884 4872
rect 4948 1728 4964 4872
rect 4868 1712 4964 1728
rect -1770 1572 -1674 1588
rect -4830 1460 -1908 1461
rect -4830 -1460 -4829 1460
rect -1909 -1460 -1908 1460
rect -4830 -1461 -1908 -1460
rect -1770 -1572 -1754 1572
rect -1690 -1572 -1674 1572
rect 1549 1572 1645 1588
rect -1511 1460 1411 1461
rect -1511 -1460 -1510 1460
rect 1410 -1460 1411 1460
rect -1511 -1461 1411 -1460
rect -1770 -1588 -1674 -1572
rect 1549 -1572 1565 1572
rect 1629 -1572 1645 1572
rect 4868 1572 4964 1588
rect 1808 1460 4730 1461
rect 1808 -1460 1809 1460
rect 4729 -1460 4730 1460
rect 1808 -1461 4730 -1460
rect 1549 -1588 1645 -1572
rect 4868 -1572 4884 1572
rect 4948 -1572 4964 1572
rect 4868 -1588 4964 -1572
rect -1770 -1728 -1674 -1712
rect -4830 -1840 -1908 -1839
rect -4830 -4760 -4829 -1840
rect -1909 -4760 -1908 -1840
rect -4830 -4761 -1908 -4760
rect -1770 -4872 -1754 -1728
rect -1690 -4872 -1674 -1728
rect 1549 -1728 1645 -1712
rect -1511 -1840 1411 -1839
rect -1511 -4760 -1510 -1840
rect 1410 -4760 1411 -1840
rect -1511 -4761 1411 -4760
rect -1770 -4888 -1674 -4872
rect 1549 -4872 1565 -1728
rect 1629 -4872 1645 -1728
rect 4868 -1728 4964 -1712
rect 1808 -1840 4730 -1839
rect 1808 -4760 1809 -1840
rect 4729 -4760 4730 -1840
rect 1808 -4761 4730 -4760
rect 1549 -4888 1645 -4872
rect 4868 -4872 4884 -1728
rect 4948 -4872 4964 -1728
rect 4868 -4888 4964 -4872
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1669 1700 4869 4900
string parameters w 15 l 15 val 235.2 carea 1.00 cperi 0.17 nx 3 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>
