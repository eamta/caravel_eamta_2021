magic
tech sky130A
magscale 1 2
timestamp 1616003964
<< nwell >>
rect -109 -242 109 242
<< pmos >>
rect -15 -180 15 180
<< pdiff >>
rect -73 168 -15 180
rect -73 -168 -61 168
rect -27 -168 -15 168
rect -73 -180 -15 -168
rect 15 168 73 180
rect 15 -168 27 168
rect 61 -168 73 168
rect 15 -180 73 -168
<< pdiffc >>
rect -61 -168 -27 168
rect 27 -168 61 168
<< poly >>
rect -15 180 15 206
rect -15 -206 15 -180
<< locali >>
rect -61 168 -27 184
rect -61 -184 -27 -168
rect 27 168 61 184
rect 27 -184 61 -168
<< viali >>
rect -61 -168 -27 168
rect 27 -168 61 168
<< metal1 >>
rect -67 168 -21 180
rect -67 -168 -61 168
rect -27 -168 -21 168
rect -67 -180 -21 -168
rect 21 168 67 180
rect 21 -168 27 168
rect 61 -168 67 168
rect 21 -180 67 -168
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
