magic
tech sky130A
magscale 1 2
timestamp 1621207460
<< metal1 >>
rect 4000 21800 22400 22100
rect 4000 21500 20440 21800
rect 20840 21500 22400 21800
rect 4020 21140 21940 21380
rect 22340 21140 22350 21380
rect 21450 12060 21460 12180
rect 21440 11920 21460 12060
rect 21820 12060 21830 12180
rect 21820 11920 21840 12060
rect 21440 11900 21840 11920
rect 11090 11760 12010 11770
rect 11090 10940 11100 11760
rect 11470 10940 12010 11760
rect 11090 10930 12010 10940
rect 2720 10810 3530 10910
rect 2720 10610 3530 10710
rect 10530 10210 11490 10310
rect 11090 9710 11490 10210
rect 11090 9700 16850 9710
rect 11090 9620 16570 9700
rect 16940 9620 16950 9700
rect 11090 9610 16850 9620
rect 10720 260 11480 270
rect 10720 180 11100 260
rect 2020 20 11100 180
rect 11470 180 11480 260
rect 11470 20 26790 180
rect 2020 -80 26790 20
<< via1 >>
rect 20440 21500 20840 21800
rect 21940 21140 22340 21380
rect 21460 11920 21820 12180
rect 11100 10940 11470 11760
rect 16570 9620 16940 9700
rect 11100 20 11470 260
<< metal2 >>
rect 20440 21800 20840 21810
rect 20440 20580 20840 21500
rect 21940 21380 22340 21390
rect 21940 20860 22340 21140
rect 9440 12070 9810 12080
rect 9440 11910 9450 12070
rect 9800 11910 9810 12070
rect 9440 10410 9810 11910
rect 11090 11760 11480 11770
rect 11090 10940 11100 11760
rect 11470 10940 11480 11760
rect 11090 260 11480 10940
rect 11540 11750 11930 11770
rect 11540 10940 11550 11750
rect 11920 10940 11930 11750
rect 11540 5500 11930 10940
rect 20440 11750 20840 12090
rect 20440 10940 20450 11750
rect 20830 10940 20840 11750
rect 20440 10930 20840 10940
rect 20940 10760 21340 12240
rect 21460 12180 21820 12190
rect 21460 11910 21820 11920
rect 20940 10230 20950 10760
rect 21330 10230 21340 10760
rect 20940 10220 21340 10230
rect 16560 9700 16950 9710
rect 16560 9620 16570 9700
rect 16940 9620 16950 9700
rect 16560 9310 16950 9620
rect 11540 5090 12200 5500
rect 11090 20 11100 260
rect 11470 20 11480 260
rect 11090 10 11480 20
<< via2 >>
rect 9450 11910 9800 12070
rect 11550 10940 11920 11750
rect 20450 10940 20830 11750
rect 21460 11920 21820 12180
rect 20950 10230 21330 10760
<< metal3 >>
rect 9440 12180 21840 12200
rect 9440 12070 21460 12180
rect 9440 11910 9450 12070
rect 9800 11920 21460 12070
rect 21820 11920 21840 12180
rect 9800 11910 21840 11920
rect 9440 11900 21840 11910
rect 11090 11750 20840 11760
rect 11090 10940 11550 11750
rect 11920 10940 20450 11750
rect 20830 10940 20840 11750
rect 11090 10930 20840 10940
rect 20940 10760 21340 10765
rect 20940 10230 20950 10760
rect 21330 10230 21340 10760
rect 20940 10225 21340 10230
<< via3 >>
rect 20950 10230 21330 10760
<< metal4 >>
rect 20949 10760 21331 10761
rect 20949 10230 20950 10760
rect 21330 10230 21331 10760
rect 20949 10229 21331 10230
use mirror  mirror_0
timestamp 1619550847
transform 1 0 4040 0 1 12065
box -40 -65 18300 9043
use input  input_0
timestamp 1619394249
transform 1 0 3626 0 1 410
box -1626 -410 7400 10510
use output  output_0
timestamp 1619566814
transform 1 0 23490 0 1 6790
box -11490 -6790 3299 4990
<< labels >>
rlabel metal2 11090 260 11480 10940 1 vss
rlabel metal1 2720 10810 3530 10910 1 vin_p
rlabel metal1 2720 10610 3530 10710 1 vin_n
rlabel metal1 4020 21140 4520 21380 1 iref
rlabel space 25470 10220 26070 10770 1 vout
rlabel metal1 4000 21500 22400 21800 1 vdd
rlabel metal1 2020 -80 26790 180 1 vss
rlabel metal1 4000 21500 22400 22100 1 vdd
<< end >>
