magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 298 1095 333 1129
rect 299 1076 333 1095
rect -17 871 0 1033
rect 129 1027 187 1033
rect 129 993 141 1027
rect 129 987 187 993
rect -105 837 0 871
rect -17 826 0 837
rect 6 826 17 837
rect -17 796 17 826
rect -17 782 0 796
rect 6 785 17 796
rect 85 826 100 841
rect 118 826 137 831
rect 85 796 143 826
rect 146 796 165 831
rect 216 826 231 841
rect 173 796 231 826
rect -51 560 -50 732
rect -42 583 -38 728
rect -17 682 16 782
rect 85 781 100 796
rect 118 766 137 796
rect 112 762 131 766
rect 146 754 173 796
rect 206 782 231 796
rect 191 769 231 782
rect 177 766 231 769
rect 185 762 219 766
rect 146 750 165 754
rect 112 732 175 750
rect 112 728 180 732
rect 192 728 222 754
rect 234 738 253 790
rect 234 728 253 732
rect 112 716 222 728
rect 134 685 209 716
rect -17 617 17 682
rect 134 669 191 685
rect 134 654 149 669
rect 265 617 268 732
rect 299 728 310 837
rect 318 732 333 1076
rect 352 1042 387 1076
rect 667 1042 702 1076
rect 299 617 333 728
rect -17 610 99 617
rect -17 606 88 610
rect -17 594 77 606
rect -17 583 16 594
rect 36 583 88 594
rect 134 583 333 617
rect 146 544 180 583
rect 352 564 386 1042
rect 668 1023 702 1042
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect 454 826 469 841
rect 454 796 512 826
rect 410 564 420 732
rect 432 728 444 790
rect 454 781 472 796
rect 460 766 472 781
rect 460 754 478 766
rect 456 743 500 754
rect 520 743 532 831
rect 548 826 560 831
rect 585 826 600 841
rect 542 796 600 826
rect 456 732 532 743
rect 456 728 500 732
rect 432 716 450 728
rect 428 687 450 716
rect 460 725 500 728
rect 520 728 532 732
rect 548 771 600 796
rect 668 826 679 837
rect 687 826 702 1023
rect 548 755 622 771
rect 548 728 588 755
rect 593 728 626 755
rect 520 727 538 728
rect 460 713 478 725
rect 512 716 538 727
rect 466 709 478 713
rect 498 713 538 716
rect 548 721 626 728
rect 548 713 622 721
rect 498 700 542 713
rect 554 709 588 713
rect 593 705 622 713
rect 634 705 659 771
rect 432 685 450 687
rect 476 697 542 700
rect 476 687 544 697
rect 432 675 444 685
rect 476 682 498 687
rect 512 682 544 687
rect 476 666 544 682
rect 559 666 560 682
rect 494 632 566 666
rect 494 616 544 632
rect 601 616 602 663
rect 529 601 544 616
rect 634 598 667 663
rect 601 596 667 598
rect 668 564 702 826
rect 721 989 756 1023
rect 1036 989 1071 1023
rect 721 732 755 989
rect 1037 970 1071 989
rect 867 921 925 927
rect 867 905 879 921
rect 867 887 908 905
rect 867 881 925 887
rect 839 853 880 877
rect 835 754 866 766
rect 352 548 544 564
rect 567 562 702 564
rect 590 553 642 562
rect 352 541 398 548
rect 456 541 486 548
rect 352 530 409 541
rect 445 533 486 541
rect 601 541 631 553
rect 601 533 642 541
rect 445 530 642 533
rect 676 530 702 562
rect 710 565 755 732
rect 801 716 832 732
rect 798 660 832 716
rect 835 672 869 754
rect 835 660 866 672
rect 798 656 866 660
rect 798 634 844 656
rect 801 622 844 634
rect 829 613 844 622
rect 867 613 925 619
rect 829 565 832 613
rect 863 579 866 613
rect 867 579 891 613
rect 867 573 925 579
rect 710 548 756 565
rect 786 548 844 565
rect 710 544 755 548
rect 798 544 832 545
rect 721 511 755 544
rect 721 510 866 511
rect 721 500 797 510
rect 721 488 786 500
rect 721 477 797 488
rect 1056 477 1071 970
rect 1090 936 1125 970
rect 1405 936 1440 970
rect 1090 477 1124 936
rect 1406 917 1440 936
rect 1236 868 1294 874
rect 1236 834 1248 868
rect 1236 828 1294 834
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1054 428 1134 441
rect 1425 424 1440 917
rect 1459 883 1494 917
rect 1774 883 1809 917
rect 1459 424 1493 883
rect 1775 864 1809 883
rect 1605 815 1663 821
rect 1605 781 1617 815
rect 1605 775 1663 781
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1794 371 1809 864
rect 1828 830 1863 864
rect 2143 830 2178 847
rect 1828 371 1862 830
rect 2144 829 2178 830
rect 2144 793 2214 829
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 2161 759 2232 793
rect 2512 759 2547 793
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1828 337 1843 371
rect 2161 318 2231 759
rect 2513 740 2547 759
rect 2343 691 2401 697
rect 2343 657 2355 691
rect 2343 651 2401 657
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2161 282 2214 318
rect 2532 265 2547 740
rect 2566 706 2601 740
rect 2566 265 2600 706
rect 2712 638 2770 644
rect 2712 604 2724 638
rect 2712 598 2770 604
rect 2882 597 2916 651
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect 2901 212 2916 597
rect 2935 563 2970 597
rect 3250 563 3285 597
rect 2935 212 2969 563
rect 3251 544 3285 563
rect 3673 547 3708 581
rect 3988 547 4023 581
rect 3081 495 3139 501
rect 3081 461 3093 495
rect 3081 455 3139 461
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3270 159 3285 544
rect 3304 510 3339 544
rect 3304 159 3338 510
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 544
rect 3673 106 3707 547
rect 3989 528 4023 547
rect 3819 479 3877 485
rect 3819 445 3831 479
rect 3819 439 3877 445
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4008 53 4023 528
rect 4042 494 4077 528
rect 4042 53 4076 494
rect 4188 426 4246 432
rect 4188 392 4200 426
rect 4188 386 4246 392
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
<< nwell >>
rect -219 539 880 917
rect -219 486 -96 539
rect -95 534 880 539
rect -95 526 172 534
rect 192 526 222 534
rect 242 526 880 534
rect -95 486 880 526
rect -219 428 880 486
<< psubdiff >>
rect -180 37 -156 71
rect 21 37 45 71
<< nsubdiff >>
rect -150 837 -105 871
rect -13 837 27 871
<< psubdiffcont >>
rect -156 37 21 71
<< nsubdiffcont >>
rect -105 837 -13 871
<< poly >>
rect -126 796 310 826
rect -126 748 -96 796
rect 280 752 310 796
rect 368 796 786 826
rect 368 728 398 796
rect 593 755 659 796
rect 593 721 609 755
rect 643 721 659 755
rect 756 745 786 796
rect 593 705 659 721
rect 11 644 77 660
rect 11 610 27 644
rect 61 610 77 644
rect 11 594 77 610
rect -126 499 -96 539
rect 47 533 77 594
rect 601 647 667 663
rect 601 613 617 647
rect 651 613 667 647
rect 601 597 667 613
rect 601 533 631 597
rect 47 503 222 533
rect -192 483 -96 499
rect -192 449 -176 483
rect -142 449 -96 483
rect -192 433 -96 449
rect -126 296 -96 433
rect 280 458 310 530
rect 456 503 631 533
rect 280 428 398 458
rect 46 389 222 405
rect 46 355 62 389
rect 96 375 222 389
rect 368 386 398 428
rect 96 355 112 375
rect 46 339 112 355
rect 756 284 786 533
rect -16 232 50 248
rect -16 198 0 232
rect 34 198 50 232
rect -16 182 50 198
rect 20 112 50 182
rect 280 112 310 168
rect 20 82 310 112
rect 456 112 486 180
rect 756 112 786 162
rect 456 82 786 112
<< polycont >>
rect 609 721 643 755
rect 27 610 61 644
rect 617 613 651 647
rect -176 449 -142 483
rect 62 355 96 389
rect 0 198 34 232
<< locali >>
rect 593 755 659 771
rect 593 721 609 755
rect 643 721 659 755
rect 593 705 659 721
rect 11 644 77 660
rect 11 610 27 644
rect 61 610 77 644
rect 11 594 77 610
rect 601 647 667 663
rect 601 613 617 647
rect 651 613 667 647
rect 601 596 667 613
rect -192 483 -126 499
rect -192 449 -176 483
rect -142 449 -126 483
rect -192 433 -126 449
rect 46 389 112 405
rect 46 355 62 389
rect 96 355 112 389
rect 46 339 112 355
rect -16 232 50 248
rect -16 198 0 232
rect 34 198 50 232
rect -16 182 50 198
<< viali >>
rect -150 837 -105 871
rect -105 837 -13 871
rect -13 837 27 871
rect 609 721 643 755
rect 27 610 61 644
rect 617 613 651 647
rect -176 449 -142 483
rect 62 355 96 389
rect 0 198 34 232
rect -180 37 -156 71
rect -156 37 21 71
rect 21 37 45 71
<< metal1 >>
rect -219 871 880 877
rect -219 837 -150 871
rect 27 837 880 871
rect -219 831 880 837
rect -172 548 -138 831
rect 11 644 77 660
rect -65 610 27 644
rect 61 610 77 644
rect 11 594 77 610
rect -192 483 -126 499
rect -192 449 -176 483
rect -142 449 -126 483
rect -192 433 -126 449
rect -178 77 -132 270
rect -84 246 -50 557
rect 146 548 180 831
rect 234 756 444 790
rect 234 725 268 756
rect 410 727 444 756
rect 322 422 356 559
rect 498 548 532 831
rect 593 757 659 771
rect 590 705 600 757
rect 652 705 662 757
rect 601 647 667 663
rect 601 613 617 647
rect 651 613 733 647
rect 601 596 667 613
rect 576 422 586 427
rect 46 398 112 405
rect 39 346 49 398
rect 101 346 112 398
rect 322 388 586 422
rect 46 339 112 346
rect -16 232 50 248
rect -57 198 0 232
rect 34 200 50 232
rect 140 200 186 360
rect 322 349 356 388
rect 576 375 586 388
rect 638 375 648 427
rect 34 198 200 200
rect -16 182 200 198
rect 0 77 200 182
rect 492 77 538 360
rect 710 261 744 579
rect 798 548 832 831
rect 594 176 604 228
rect 656 210 666 228
rect 656 176 744 210
rect 792 77 838 270
rect -197 71 880 77
rect -197 37 -180 71
rect 45 37 880 71
rect -197 31 880 37
rect 0 0 200 31
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
<< via1 >>
rect 600 755 652 757
rect 600 721 609 755
rect 609 721 643 755
rect 643 721 652 755
rect 600 705 652 721
rect 49 389 101 398
rect 49 355 62 389
rect 62 355 96 389
rect 96 355 101 389
rect 49 346 101 355
rect 586 375 638 427
rect 604 176 656 228
<< metal2 >>
rect 600 757 652 767
rect 600 695 652 705
rect 586 428 638 437
rect 586 427 881 428
rect 49 398 101 408
rect 638 375 881 427
rect 586 365 638 375
rect 49 336 101 346
rect 64 230 97 336
rect 604 230 656 238
rect 64 228 656 230
rect 64 195 604 228
rect 594 176 604 195
rect 656 176 662 228
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615150785
transform 1 0 -111 0 1 225
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_1
timestamp 1615077590
transform 1 0 207 0 1 270
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_2
timestamp 1615077590
transform 1 0 295 0 1 270
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_3
timestamp 1615077590
transform 1 0 383 0 1 270
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_4
timestamp 1615077590
transform 1 0 471 0 1 270
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_1
timestamp 1615150785
transform 1 0 771 0 1 225
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_XSLFBL  XM4
timestamp 1624053917
transform 1 0 1265 0 1 697
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_L9ESED  XM7
timestamp 1624053917
transform 1 0 2372 0 1 529
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_XSLFBL  XM6
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 1634 0 1 644
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3110 0 1 378
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_L9ESED  XM8
timestamp 1624053917
transform 1 0 2741 0 1 476
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM11
timestamp 1624053917
transform 1 0 3848 0 1 317
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_HVW3BE  XM10
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_L9ESED  XM12
timestamp 1624053917
transform 1 0 4217 0 1 264
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_0
timestamp 1614978561
transform 1 0 -111 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_1
timestamp 1614978561
transform 1 0 207 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_2
timestamp 1614978561
transform 1 0 295 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_5
timestamp 1614978561
transform 1 0 383 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_4
timestamp 1614978561
transform 1 0 471 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 158 0 1 856
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_3
timestamp 1614978561
transform 1 0 771 0 1 638
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_XSLFBL  XM3
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
<< labels >>
rlabel metal1 -142 433 -126 499 1 a
rlabel metal2 600 695 652 705 1 b
rlabel metal2 638 375 881 428 1 z
rlabel nwell -150 837 27 871 1 vdd!
rlabel metal1 -156 37 21 71 1 vss!
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 b
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 z
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
<< end >>
