magic
tech sky130A
magscale 1 2
timestamp 1624338677
<< nwell >>
rect -263 -330 263 330
<< pmos >>
rect -63 -111 -33 111
rect 33 -111 63 111
<< pdiff >>
rect -125 99 -63 111
rect -125 -99 -113 99
rect -79 -99 -63 99
rect -125 -111 -63 -99
rect -33 99 33 111
rect -33 -99 -17 99
rect 17 -99 33 99
rect -33 -111 33 -99
rect 63 99 125 111
rect 63 -99 79 99
rect 113 -99 125 99
rect 63 -111 125 -99
<< pdiffc >>
rect -113 -99 -79 99
rect -17 -99 17 99
rect 79 -99 113 99
<< nsubdiff >>
rect -227 260 227 294
rect -227 198 -193 260
rect 193 198 227 260
rect -227 -260 -193 -198
rect 193 -260 227 -198
rect -227 -294 -131 -260
rect 131 -294 227 -260
<< nsubdiffcont >>
rect -227 -198 -193 198
rect 193 -198 227 198
rect -131 -294 131 -260
<< poly >>
rect -87 192 -21 208
rect -87 158 -71 192
rect -37 158 -21 192
rect -87 142 -21 158
rect 21 192 87 208
rect 21 158 37 192
rect 71 158 87 192
rect 21 142 87 158
rect -63 111 -33 142
rect 33 111 63 142
rect -63 -137 -33 -111
rect 33 -137 63 -111
<< polycont >>
rect -71 158 -37 192
rect 37 158 71 192
<< locali >>
rect -227 260 227 294
rect -227 198 -193 260
rect 193 198 227 260
rect -87 158 -71 192
rect -37 158 -21 192
rect 21 158 37 192
rect 71 158 87 192
rect -113 99 -79 115
rect -113 -115 -79 -99
rect -17 99 17 115
rect -17 -115 17 -99
rect 79 99 113 115
rect 79 -115 113 -99
rect -227 -260 -193 -198
rect 193 -260 227 -198
rect -227 -294 -131 -260
rect 131 -294 227 -260
<< viali >>
rect -71 158 -37 192
rect 37 158 71 192
rect -113 -99 -79 99
rect -17 -99 17 99
rect 79 -99 113 99
<< metal1 >>
rect -87 192 -21 204
rect -87 158 -71 192
rect -37 158 -21 192
rect -87 146 -21 158
rect 21 192 87 204
rect 21 158 37 192
rect 71 158 87 192
rect 21 146 87 158
rect -119 99 -73 111
rect -119 -99 -113 99
rect -79 -99 -73 99
rect -119 -111 -73 -99
rect -23 99 23 111
rect -23 -99 -17 99
rect 17 -99 23 99
rect -23 -111 23 -99
rect 73 99 119 111
rect 73 -99 79 99
rect 113 -99 119 99
rect 73 -111 119 -99
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -210 -277 210 277
string parameters w 1.11 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
