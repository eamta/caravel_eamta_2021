magic
tech sky130A
magscale 1 2
timestamp 1615997521
<< nwell >>
rect -13567 -569 13567 569
<< pmoslvt >>
rect -13371 -350 -13161 350
rect -13103 -350 -12893 350
rect -12835 -350 -12625 350
rect -12567 -350 -12357 350
rect -12299 -350 -12089 350
rect -12031 -350 -11821 350
rect -11763 -350 -11553 350
rect -11495 -350 -11285 350
rect -11227 -350 -11017 350
rect -10959 -350 -10749 350
rect -10691 -350 -10481 350
rect -10423 -350 -10213 350
rect -10155 -350 -9945 350
rect -9887 -350 -9677 350
rect -9619 -350 -9409 350
rect -9351 -350 -9141 350
rect -9083 -350 -8873 350
rect -8815 -350 -8605 350
rect -8547 -350 -8337 350
rect -8279 -350 -8069 350
rect -8011 -350 -7801 350
rect -7743 -350 -7533 350
rect -7475 -350 -7265 350
rect -7207 -350 -6997 350
rect -6939 -350 -6729 350
rect -6671 -350 -6461 350
rect -6403 -350 -6193 350
rect -6135 -350 -5925 350
rect -5867 -350 -5657 350
rect -5599 -350 -5389 350
rect -5331 -350 -5121 350
rect -5063 -350 -4853 350
rect -4795 -350 -4585 350
rect -4527 -350 -4317 350
rect -4259 -350 -4049 350
rect -3991 -350 -3781 350
rect -3723 -350 -3513 350
rect -3455 -350 -3245 350
rect -3187 -350 -2977 350
rect -2919 -350 -2709 350
rect -2651 -350 -2441 350
rect -2383 -350 -2173 350
rect -2115 -350 -1905 350
rect -1847 -350 -1637 350
rect -1579 -350 -1369 350
rect -1311 -350 -1101 350
rect -1043 -350 -833 350
rect -775 -350 -565 350
rect -507 -350 -297 350
rect -239 -350 -29 350
rect 29 -350 239 350
rect 297 -350 507 350
rect 565 -350 775 350
rect 833 -350 1043 350
rect 1101 -350 1311 350
rect 1369 -350 1579 350
rect 1637 -350 1847 350
rect 1905 -350 2115 350
rect 2173 -350 2383 350
rect 2441 -350 2651 350
rect 2709 -350 2919 350
rect 2977 -350 3187 350
rect 3245 -350 3455 350
rect 3513 -350 3723 350
rect 3781 -350 3991 350
rect 4049 -350 4259 350
rect 4317 -350 4527 350
rect 4585 -350 4795 350
rect 4853 -350 5063 350
rect 5121 -350 5331 350
rect 5389 -350 5599 350
rect 5657 -350 5867 350
rect 5925 -350 6135 350
rect 6193 -350 6403 350
rect 6461 -350 6671 350
rect 6729 -350 6939 350
rect 6997 -350 7207 350
rect 7265 -350 7475 350
rect 7533 -350 7743 350
rect 7801 -350 8011 350
rect 8069 -350 8279 350
rect 8337 -350 8547 350
rect 8605 -350 8815 350
rect 8873 -350 9083 350
rect 9141 -350 9351 350
rect 9409 -350 9619 350
rect 9677 -350 9887 350
rect 9945 -350 10155 350
rect 10213 -350 10423 350
rect 10481 -350 10691 350
rect 10749 -350 10959 350
rect 11017 -350 11227 350
rect 11285 -350 11495 350
rect 11553 -350 11763 350
rect 11821 -350 12031 350
rect 12089 -350 12299 350
rect 12357 -350 12567 350
rect 12625 -350 12835 350
rect 12893 -350 13103 350
rect 13161 -350 13371 350
<< pdiff >>
rect -13429 338 -13371 350
rect -13429 -338 -13417 338
rect -13383 -338 -13371 338
rect -13429 -350 -13371 -338
rect -13161 338 -13103 350
rect -13161 -338 -13149 338
rect -13115 -338 -13103 338
rect -13161 -350 -13103 -338
rect -12893 338 -12835 350
rect -12893 -338 -12881 338
rect -12847 -338 -12835 338
rect -12893 -350 -12835 -338
rect -12625 338 -12567 350
rect -12625 -338 -12613 338
rect -12579 -338 -12567 338
rect -12625 -350 -12567 -338
rect -12357 338 -12299 350
rect -12357 -338 -12345 338
rect -12311 -338 -12299 338
rect -12357 -350 -12299 -338
rect -12089 338 -12031 350
rect -12089 -338 -12077 338
rect -12043 -338 -12031 338
rect -12089 -350 -12031 -338
rect -11821 338 -11763 350
rect -11821 -338 -11809 338
rect -11775 -338 -11763 338
rect -11821 -350 -11763 -338
rect -11553 338 -11495 350
rect -11553 -338 -11541 338
rect -11507 -338 -11495 338
rect -11553 -350 -11495 -338
rect -11285 338 -11227 350
rect -11285 -338 -11273 338
rect -11239 -338 -11227 338
rect -11285 -350 -11227 -338
rect -11017 338 -10959 350
rect -11017 -338 -11005 338
rect -10971 -338 -10959 338
rect -11017 -350 -10959 -338
rect -10749 338 -10691 350
rect -10749 -338 -10737 338
rect -10703 -338 -10691 338
rect -10749 -350 -10691 -338
rect -10481 338 -10423 350
rect -10481 -338 -10469 338
rect -10435 -338 -10423 338
rect -10481 -350 -10423 -338
rect -10213 338 -10155 350
rect -10213 -338 -10201 338
rect -10167 -338 -10155 338
rect -10213 -350 -10155 -338
rect -9945 338 -9887 350
rect -9945 -338 -9933 338
rect -9899 -338 -9887 338
rect -9945 -350 -9887 -338
rect -9677 338 -9619 350
rect -9677 -338 -9665 338
rect -9631 -338 -9619 338
rect -9677 -350 -9619 -338
rect -9409 338 -9351 350
rect -9409 -338 -9397 338
rect -9363 -338 -9351 338
rect -9409 -350 -9351 -338
rect -9141 338 -9083 350
rect -9141 -338 -9129 338
rect -9095 -338 -9083 338
rect -9141 -350 -9083 -338
rect -8873 338 -8815 350
rect -8873 -338 -8861 338
rect -8827 -338 -8815 338
rect -8873 -350 -8815 -338
rect -8605 338 -8547 350
rect -8605 -338 -8593 338
rect -8559 -338 -8547 338
rect -8605 -350 -8547 -338
rect -8337 338 -8279 350
rect -8337 -338 -8325 338
rect -8291 -338 -8279 338
rect -8337 -350 -8279 -338
rect -8069 338 -8011 350
rect -8069 -338 -8057 338
rect -8023 -338 -8011 338
rect -8069 -350 -8011 -338
rect -7801 338 -7743 350
rect -7801 -338 -7789 338
rect -7755 -338 -7743 338
rect -7801 -350 -7743 -338
rect -7533 338 -7475 350
rect -7533 -338 -7521 338
rect -7487 -338 -7475 338
rect -7533 -350 -7475 -338
rect -7265 338 -7207 350
rect -7265 -338 -7253 338
rect -7219 -338 -7207 338
rect -7265 -350 -7207 -338
rect -6997 338 -6939 350
rect -6997 -338 -6985 338
rect -6951 -338 -6939 338
rect -6997 -350 -6939 -338
rect -6729 338 -6671 350
rect -6729 -338 -6717 338
rect -6683 -338 -6671 338
rect -6729 -350 -6671 -338
rect -6461 338 -6403 350
rect -6461 -338 -6449 338
rect -6415 -338 -6403 338
rect -6461 -350 -6403 -338
rect -6193 338 -6135 350
rect -6193 -338 -6181 338
rect -6147 -338 -6135 338
rect -6193 -350 -6135 -338
rect -5925 338 -5867 350
rect -5925 -338 -5913 338
rect -5879 -338 -5867 338
rect -5925 -350 -5867 -338
rect -5657 338 -5599 350
rect -5657 -338 -5645 338
rect -5611 -338 -5599 338
rect -5657 -350 -5599 -338
rect -5389 338 -5331 350
rect -5389 -338 -5377 338
rect -5343 -338 -5331 338
rect -5389 -350 -5331 -338
rect -5121 338 -5063 350
rect -5121 -338 -5109 338
rect -5075 -338 -5063 338
rect -5121 -350 -5063 -338
rect -4853 338 -4795 350
rect -4853 -338 -4841 338
rect -4807 -338 -4795 338
rect -4853 -350 -4795 -338
rect -4585 338 -4527 350
rect -4585 -338 -4573 338
rect -4539 -338 -4527 338
rect -4585 -350 -4527 -338
rect -4317 338 -4259 350
rect -4317 -338 -4305 338
rect -4271 -338 -4259 338
rect -4317 -350 -4259 -338
rect -4049 338 -3991 350
rect -4049 -338 -4037 338
rect -4003 -338 -3991 338
rect -4049 -350 -3991 -338
rect -3781 338 -3723 350
rect -3781 -338 -3769 338
rect -3735 -338 -3723 338
rect -3781 -350 -3723 -338
rect -3513 338 -3455 350
rect -3513 -338 -3501 338
rect -3467 -338 -3455 338
rect -3513 -350 -3455 -338
rect -3245 338 -3187 350
rect -3245 -338 -3233 338
rect -3199 -338 -3187 338
rect -3245 -350 -3187 -338
rect -2977 338 -2919 350
rect -2977 -338 -2965 338
rect -2931 -338 -2919 338
rect -2977 -350 -2919 -338
rect -2709 338 -2651 350
rect -2709 -338 -2697 338
rect -2663 -338 -2651 338
rect -2709 -350 -2651 -338
rect -2441 338 -2383 350
rect -2441 -338 -2429 338
rect -2395 -338 -2383 338
rect -2441 -350 -2383 -338
rect -2173 338 -2115 350
rect -2173 -338 -2161 338
rect -2127 -338 -2115 338
rect -2173 -350 -2115 -338
rect -1905 338 -1847 350
rect -1905 -338 -1893 338
rect -1859 -338 -1847 338
rect -1905 -350 -1847 -338
rect -1637 338 -1579 350
rect -1637 -338 -1625 338
rect -1591 -338 -1579 338
rect -1637 -350 -1579 -338
rect -1369 338 -1311 350
rect -1369 -338 -1357 338
rect -1323 -338 -1311 338
rect -1369 -350 -1311 -338
rect -1101 338 -1043 350
rect -1101 -338 -1089 338
rect -1055 -338 -1043 338
rect -1101 -350 -1043 -338
rect -833 338 -775 350
rect -833 -338 -821 338
rect -787 -338 -775 338
rect -833 -350 -775 -338
rect -565 338 -507 350
rect -565 -338 -553 338
rect -519 -338 -507 338
rect -565 -350 -507 -338
rect -297 338 -239 350
rect -297 -338 -285 338
rect -251 -338 -239 338
rect -297 -350 -239 -338
rect -29 338 29 350
rect -29 -338 -17 338
rect 17 -338 29 338
rect -29 -350 29 -338
rect 239 338 297 350
rect 239 -338 251 338
rect 285 -338 297 338
rect 239 -350 297 -338
rect 507 338 565 350
rect 507 -338 519 338
rect 553 -338 565 338
rect 507 -350 565 -338
rect 775 338 833 350
rect 775 -338 787 338
rect 821 -338 833 338
rect 775 -350 833 -338
rect 1043 338 1101 350
rect 1043 -338 1055 338
rect 1089 -338 1101 338
rect 1043 -350 1101 -338
rect 1311 338 1369 350
rect 1311 -338 1323 338
rect 1357 -338 1369 338
rect 1311 -350 1369 -338
rect 1579 338 1637 350
rect 1579 -338 1591 338
rect 1625 -338 1637 338
rect 1579 -350 1637 -338
rect 1847 338 1905 350
rect 1847 -338 1859 338
rect 1893 -338 1905 338
rect 1847 -350 1905 -338
rect 2115 338 2173 350
rect 2115 -338 2127 338
rect 2161 -338 2173 338
rect 2115 -350 2173 -338
rect 2383 338 2441 350
rect 2383 -338 2395 338
rect 2429 -338 2441 338
rect 2383 -350 2441 -338
rect 2651 338 2709 350
rect 2651 -338 2663 338
rect 2697 -338 2709 338
rect 2651 -350 2709 -338
rect 2919 338 2977 350
rect 2919 -338 2931 338
rect 2965 -338 2977 338
rect 2919 -350 2977 -338
rect 3187 338 3245 350
rect 3187 -338 3199 338
rect 3233 -338 3245 338
rect 3187 -350 3245 -338
rect 3455 338 3513 350
rect 3455 -338 3467 338
rect 3501 -338 3513 338
rect 3455 -350 3513 -338
rect 3723 338 3781 350
rect 3723 -338 3735 338
rect 3769 -338 3781 338
rect 3723 -350 3781 -338
rect 3991 338 4049 350
rect 3991 -338 4003 338
rect 4037 -338 4049 338
rect 3991 -350 4049 -338
rect 4259 338 4317 350
rect 4259 -338 4271 338
rect 4305 -338 4317 338
rect 4259 -350 4317 -338
rect 4527 338 4585 350
rect 4527 -338 4539 338
rect 4573 -338 4585 338
rect 4527 -350 4585 -338
rect 4795 338 4853 350
rect 4795 -338 4807 338
rect 4841 -338 4853 338
rect 4795 -350 4853 -338
rect 5063 338 5121 350
rect 5063 -338 5075 338
rect 5109 -338 5121 338
rect 5063 -350 5121 -338
rect 5331 338 5389 350
rect 5331 -338 5343 338
rect 5377 -338 5389 338
rect 5331 -350 5389 -338
rect 5599 338 5657 350
rect 5599 -338 5611 338
rect 5645 -338 5657 338
rect 5599 -350 5657 -338
rect 5867 338 5925 350
rect 5867 -338 5879 338
rect 5913 -338 5925 338
rect 5867 -350 5925 -338
rect 6135 338 6193 350
rect 6135 -338 6147 338
rect 6181 -338 6193 338
rect 6135 -350 6193 -338
rect 6403 338 6461 350
rect 6403 -338 6415 338
rect 6449 -338 6461 338
rect 6403 -350 6461 -338
rect 6671 338 6729 350
rect 6671 -338 6683 338
rect 6717 -338 6729 338
rect 6671 -350 6729 -338
rect 6939 338 6997 350
rect 6939 -338 6951 338
rect 6985 -338 6997 338
rect 6939 -350 6997 -338
rect 7207 338 7265 350
rect 7207 -338 7219 338
rect 7253 -338 7265 338
rect 7207 -350 7265 -338
rect 7475 338 7533 350
rect 7475 -338 7487 338
rect 7521 -338 7533 338
rect 7475 -350 7533 -338
rect 7743 338 7801 350
rect 7743 -338 7755 338
rect 7789 -338 7801 338
rect 7743 -350 7801 -338
rect 8011 338 8069 350
rect 8011 -338 8023 338
rect 8057 -338 8069 338
rect 8011 -350 8069 -338
rect 8279 338 8337 350
rect 8279 -338 8291 338
rect 8325 -338 8337 338
rect 8279 -350 8337 -338
rect 8547 338 8605 350
rect 8547 -338 8559 338
rect 8593 -338 8605 338
rect 8547 -350 8605 -338
rect 8815 338 8873 350
rect 8815 -338 8827 338
rect 8861 -338 8873 338
rect 8815 -350 8873 -338
rect 9083 338 9141 350
rect 9083 -338 9095 338
rect 9129 -338 9141 338
rect 9083 -350 9141 -338
rect 9351 338 9409 350
rect 9351 -338 9363 338
rect 9397 -338 9409 338
rect 9351 -350 9409 -338
rect 9619 338 9677 350
rect 9619 -338 9631 338
rect 9665 -338 9677 338
rect 9619 -350 9677 -338
rect 9887 338 9945 350
rect 9887 -338 9899 338
rect 9933 -338 9945 338
rect 9887 -350 9945 -338
rect 10155 338 10213 350
rect 10155 -338 10167 338
rect 10201 -338 10213 338
rect 10155 -350 10213 -338
rect 10423 338 10481 350
rect 10423 -338 10435 338
rect 10469 -338 10481 338
rect 10423 -350 10481 -338
rect 10691 338 10749 350
rect 10691 -338 10703 338
rect 10737 -338 10749 338
rect 10691 -350 10749 -338
rect 10959 338 11017 350
rect 10959 -338 10971 338
rect 11005 -338 11017 338
rect 10959 -350 11017 -338
rect 11227 338 11285 350
rect 11227 -338 11239 338
rect 11273 -338 11285 338
rect 11227 -350 11285 -338
rect 11495 338 11553 350
rect 11495 -338 11507 338
rect 11541 -338 11553 338
rect 11495 -350 11553 -338
rect 11763 338 11821 350
rect 11763 -338 11775 338
rect 11809 -338 11821 338
rect 11763 -350 11821 -338
rect 12031 338 12089 350
rect 12031 -338 12043 338
rect 12077 -338 12089 338
rect 12031 -350 12089 -338
rect 12299 338 12357 350
rect 12299 -338 12311 338
rect 12345 -338 12357 338
rect 12299 -350 12357 -338
rect 12567 338 12625 350
rect 12567 -338 12579 338
rect 12613 -338 12625 338
rect 12567 -350 12625 -338
rect 12835 338 12893 350
rect 12835 -338 12847 338
rect 12881 -338 12893 338
rect 12835 -350 12893 -338
rect 13103 338 13161 350
rect 13103 -338 13115 338
rect 13149 -338 13161 338
rect 13103 -350 13161 -338
rect 13371 338 13429 350
rect 13371 -338 13383 338
rect 13417 -338 13429 338
rect 13371 -350 13429 -338
<< pdiffc >>
rect -13417 -338 -13383 338
rect -13149 -338 -13115 338
rect -12881 -338 -12847 338
rect -12613 -338 -12579 338
rect -12345 -338 -12311 338
rect -12077 -338 -12043 338
rect -11809 -338 -11775 338
rect -11541 -338 -11507 338
rect -11273 -338 -11239 338
rect -11005 -338 -10971 338
rect -10737 -338 -10703 338
rect -10469 -338 -10435 338
rect -10201 -338 -10167 338
rect -9933 -338 -9899 338
rect -9665 -338 -9631 338
rect -9397 -338 -9363 338
rect -9129 -338 -9095 338
rect -8861 -338 -8827 338
rect -8593 -338 -8559 338
rect -8325 -338 -8291 338
rect -8057 -338 -8023 338
rect -7789 -338 -7755 338
rect -7521 -338 -7487 338
rect -7253 -338 -7219 338
rect -6985 -338 -6951 338
rect -6717 -338 -6683 338
rect -6449 -338 -6415 338
rect -6181 -338 -6147 338
rect -5913 -338 -5879 338
rect -5645 -338 -5611 338
rect -5377 -338 -5343 338
rect -5109 -338 -5075 338
rect -4841 -338 -4807 338
rect -4573 -338 -4539 338
rect -4305 -338 -4271 338
rect -4037 -338 -4003 338
rect -3769 -338 -3735 338
rect -3501 -338 -3467 338
rect -3233 -338 -3199 338
rect -2965 -338 -2931 338
rect -2697 -338 -2663 338
rect -2429 -338 -2395 338
rect -2161 -338 -2127 338
rect -1893 -338 -1859 338
rect -1625 -338 -1591 338
rect -1357 -338 -1323 338
rect -1089 -338 -1055 338
rect -821 -338 -787 338
rect -553 -338 -519 338
rect -285 -338 -251 338
rect -17 -338 17 338
rect 251 -338 285 338
rect 519 -338 553 338
rect 787 -338 821 338
rect 1055 -338 1089 338
rect 1323 -338 1357 338
rect 1591 -338 1625 338
rect 1859 -338 1893 338
rect 2127 -338 2161 338
rect 2395 -338 2429 338
rect 2663 -338 2697 338
rect 2931 -338 2965 338
rect 3199 -338 3233 338
rect 3467 -338 3501 338
rect 3735 -338 3769 338
rect 4003 -338 4037 338
rect 4271 -338 4305 338
rect 4539 -338 4573 338
rect 4807 -338 4841 338
rect 5075 -338 5109 338
rect 5343 -338 5377 338
rect 5611 -338 5645 338
rect 5879 -338 5913 338
rect 6147 -338 6181 338
rect 6415 -338 6449 338
rect 6683 -338 6717 338
rect 6951 -338 6985 338
rect 7219 -338 7253 338
rect 7487 -338 7521 338
rect 7755 -338 7789 338
rect 8023 -338 8057 338
rect 8291 -338 8325 338
rect 8559 -338 8593 338
rect 8827 -338 8861 338
rect 9095 -338 9129 338
rect 9363 -338 9397 338
rect 9631 -338 9665 338
rect 9899 -338 9933 338
rect 10167 -338 10201 338
rect 10435 -338 10469 338
rect 10703 -338 10737 338
rect 10971 -338 11005 338
rect 11239 -338 11273 338
rect 11507 -338 11541 338
rect 11775 -338 11809 338
rect 12043 -338 12077 338
rect 12311 -338 12345 338
rect 12579 -338 12613 338
rect 12847 -338 12881 338
rect 13115 -338 13149 338
rect 13383 -338 13417 338
<< nsubdiff >>
rect -13531 499 -13435 533
rect 13435 499 13531 533
rect -13531 437 -13497 499
rect 13497 437 13531 499
rect -13531 -499 -13497 -437
rect 13497 -499 13531 -437
rect -13531 -533 -13435 -499
rect 13435 -533 13531 -499
<< nsubdiffcont >>
rect -13435 499 13435 533
rect -13531 -437 -13497 437
rect 13497 -437 13531 437
rect -13435 -533 13435 -499
<< poly >>
rect -13371 431 -13161 447
rect -13371 397 -13355 431
rect -13177 397 -13161 431
rect -13371 350 -13161 397
rect -13103 431 -12893 447
rect -13103 397 -13087 431
rect -12909 397 -12893 431
rect -13103 350 -12893 397
rect -12835 431 -12625 447
rect -12835 397 -12819 431
rect -12641 397 -12625 431
rect -12835 350 -12625 397
rect -12567 431 -12357 447
rect -12567 397 -12551 431
rect -12373 397 -12357 431
rect -12567 350 -12357 397
rect -12299 431 -12089 447
rect -12299 397 -12283 431
rect -12105 397 -12089 431
rect -12299 350 -12089 397
rect -12031 431 -11821 447
rect -12031 397 -12015 431
rect -11837 397 -11821 431
rect -12031 350 -11821 397
rect -11763 431 -11553 447
rect -11763 397 -11747 431
rect -11569 397 -11553 431
rect -11763 350 -11553 397
rect -11495 431 -11285 447
rect -11495 397 -11479 431
rect -11301 397 -11285 431
rect -11495 350 -11285 397
rect -11227 431 -11017 447
rect -11227 397 -11211 431
rect -11033 397 -11017 431
rect -11227 350 -11017 397
rect -10959 431 -10749 447
rect -10959 397 -10943 431
rect -10765 397 -10749 431
rect -10959 350 -10749 397
rect -10691 431 -10481 447
rect -10691 397 -10675 431
rect -10497 397 -10481 431
rect -10691 350 -10481 397
rect -10423 431 -10213 447
rect -10423 397 -10407 431
rect -10229 397 -10213 431
rect -10423 350 -10213 397
rect -10155 431 -9945 447
rect -10155 397 -10139 431
rect -9961 397 -9945 431
rect -10155 350 -9945 397
rect -9887 431 -9677 447
rect -9887 397 -9871 431
rect -9693 397 -9677 431
rect -9887 350 -9677 397
rect -9619 431 -9409 447
rect -9619 397 -9603 431
rect -9425 397 -9409 431
rect -9619 350 -9409 397
rect -9351 431 -9141 447
rect -9351 397 -9335 431
rect -9157 397 -9141 431
rect -9351 350 -9141 397
rect -9083 431 -8873 447
rect -9083 397 -9067 431
rect -8889 397 -8873 431
rect -9083 350 -8873 397
rect -8815 431 -8605 447
rect -8815 397 -8799 431
rect -8621 397 -8605 431
rect -8815 350 -8605 397
rect -8547 431 -8337 447
rect -8547 397 -8531 431
rect -8353 397 -8337 431
rect -8547 350 -8337 397
rect -8279 431 -8069 447
rect -8279 397 -8263 431
rect -8085 397 -8069 431
rect -8279 350 -8069 397
rect -8011 431 -7801 447
rect -8011 397 -7995 431
rect -7817 397 -7801 431
rect -8011 350 -7801 397
rect -7743 431 -7533 447
rect -7743 397 -7727 431
rect -7549 397 -7533 431
rect -7743 350 -7533 397
rect -7475 431 -7265 447
rect -7475 397 -7459 431
rect -7281 397 -7265 431
rect -7475 350 -7265 397
rect -7207 431 -6997 447
rect -7207 397 -7191 431
rect -7013 397 -6997 431
rect -7207 350 -6997 397
rect -6939 431 -6729 447
rect -6939 397 -6923 431
rect -6745 397 -6729 431
rect -6939 350 -6729 397
rect -6671 431 -6461 447
rect -6671 397 -6655 431
rect -6477 397 -6461 431
rect -6671 350 -6461 397
rect -6403 431 -6193 447
rect -6403 397 -6387 431
rect -6209 397 -6193 431
rect -6403 350 -6193 397
rect -6135 431 -5925 447
rect -6135 397 -6119 431
rect -5941 397 -5925 431
rect -6135 350 -5925 397
rect -5867 431 -5657 447
rect -5867 397 -5851 431
rect -5673 397 -5657 431
rect -5867 350 -5657 397
rect -5599 431 -5389 447
rect -5599 397 -5583 431
rect -5405 397 -5389 431
rect -5599 350 -5389 397
rect -5331 431 -5121 447
rect -5331 397 -5315 431
rect -5137 397 -5121 431
rect -5331 350 -5121 397
rect -5063 431 -4853 447
rect -5063 397 -5047 431
rect -4869 397 -4853 431
rect -5063 350 -4853 397
rect -4795 431 -4585 447
rect -4795 397 -4779 431
rect -4601 397 -4585 431
rect -4795 350 -4585 397
rect -4527 431 -4317 447
rect -4527 397 -4511 431
rect -4333 397 -4317 431
rect -4527 350 -4317 397
rect -4259 431 -4049 447
rect -4259 397 -4243 431
rect -4065 397 -4049 431
rect -4259 350 -4049 397
rect -3991 431 -3781 447
rect -3991 397 -3975 431
rect -3797 397 -3781 431
rect -3991 350 -3781 397
rect -3723 431 -3513 447
rect -3723 397 -3707 431
rect -3529 397 -3513 431
rect -3723 350 -3513 397
rect -3455 431 -3245 447
rect -3455 397 -3439 431
rect -3261 397 -3245 431
rect -3455 350 -3245 397
rect -3187 431 -2977 447
rect -3187 397 -3171 431
rect -2993 397 -2977 431
rect -3187 350 -2977 397
rect -2919 431 -2709 447
rect -2919 397 -2903 431
rect -2725 397 -2709 431
rect -2919 350 -2709 397
rect -2651 431 -2441 447
rect -2651 397 -2635 431
rect -2457 397 -2441 431
rect -2651 350 -2441 397
rect -2383 431 -2173 447
rect -2383 397 -2367 431
rect -2189 397 -2173 431
rect -2383 350 -2173 397
rect -2115 431 -1905 447
rect -2115 397 -2099 431
rect -1921 397 -1905 431
rect -2115 350 -1905 397
rect -1847 431 -1637 447
rect -1847 397 -1831 431
rect -1653 397 -1637 431
rect -1847 350 -1637 397
rect -1579 431 -1369 447
rect -1579 397 -1563 431
rect -1385 397 -1369 431
rect -1579 350 -1369 397
rect -1311 431 -1101 447
rect -1311 397 -1295 431
rect -1117 397 -1101 431
rect -1311 350 -1101 397
rect -1043 431 -833 447
rect -1043 397 -1027 431
rect -849 397 -833 431
rect -1043 350 -833 397
rect -775 431 -565 447
rect -775 397 -759 431
rect -581 397 -565 431
rect -775 350 -565 397
rect -507 431 -297 447
rect -507 397 -491 431
rect -313 397 -297 431
rect -507 350 -297 397
rect -239 431 -29 447
rect -239 397 -223 431
rect -45 397 -29 431
rect -239 350 -29 397
rect 29 431 239 447
rect 29 397 45 431
rect 223 397 239 431
rect 29 350 239 397
rect 297 431 507 447
rect 297 397 313 431
rect 491 397 507 431
rect 297 350 507 397
rect 565 431 775 447
rect 565 397 581 431
rect 759 397 775 431
rect 565 350 775 397
rect 833 431 1043 447
rect 833 397 849 431
rect 1027 397 1043 431
rect 833 350 1043 397
rect 1101 431 1311 447
rect 1101 397 1117 431
rect 1295 397 1311 431
rect 1101 350 1311 397
rect 1369 431 1579 447
rect 1369 397 1385 431
rect 1563 397 1579 431
rect 1369 350 1579 397
rect 1637 431 1847 447
rect 1637 397 1653 431
rect 1831 397 1847 431
rect 1637 350 1847 397
rect 1905 431 2115 447
rect 1905 397 1921 431
rect 2099 397 2115 431
rect 1905 350 2115 397
rect 2173 431 2383 447
rect 2173 397 2189 431
rect 2367 397 2383 431
rect 2173 350 2383 397
rect 2441 431 2651 447
rect 2441 397 2457 431
rect 2635 397 2651 431
rect 2441 350 2651 397
rect 2709 431 2919 447
rect 2709 397 2725 431
rect 2903 397 2919 431
rect 2709 350 2919 397
rect 2977 431 3187 447
rect 2977 397 2993 431
rect 3171 397 3187 431
rect 2977 350 3187 397
rect 3245 431 3455 447
rect 3245 397 3261 431
rect 3439 397 3455 431
rect 3245 350 3455 397
rect 3513 431 3723 447
rect 3513 397 3529 431
rect 3707 397 3723 431
rect 3513 350 3723 397
rect 3781 431 3991 447
rect 3781 397 3797 431
rect 3975 397 3991 431
rect 3781 350 3991 397
rect 4049 431 4259 447
rect 4049 397 4065 431
rect 4243 397 4259 431
rect 4049 350 4259 397
rect 4317 431 4527 447
rect 4317 397 4333 431
rect 4511 397 4527 431
rect 4317 350 4527 397
rect 4585 431 4795 447
rect 4585 397 4601 431
rect 4779 397 4795 431
rect 4585 350 4795 397
rect 4853 431 5063 447
rect 4853 397 4869 431
rect 5047 397 5063 431
rect 4853 350 5063 397
rect 5121 431 5331 447
rect 5121 397 5137 431
rect 5315 397 5331 431
rect 5121 350 5331 397
rect 5389 431 5599 447
rect 5389 397 5405 431
rect 5583 397 5599 431
rect 5389 350 5599 397
rect 5657 431 5867 447
rect 5657 397 5673 431
rect 5851 397 5867 431
rect 5657 350 5867 397
rect 5925 431 6135 447
rect 5925 397 5941 431
rect 6119 397 6135 431
rect 5925 350 6135 397
rect 6193 431 6403 447
rect 6193 397 6209 431
rect 6387 397 6403 431
rect 6193 350 6403 397
rect 6461 431 6671 447
rect 6461 397 6477 431
rect 6655 397 6671 431
rect 6461 350 6671 397
rect 6729 431 6939 447
rect 6729 397 6745 431
rect 6923 397 6939 431
rect 6729 350 6939 397
rect 6997 431 7207 447
rect 6997 397 7013 431
rect 7191 397 7207 431
rect 6997 350 7207 397
rect 7265 431 7475 447
rect 7265 397 7281 431
rect 7459 397 7475 431
rect 7265 350 7475 397
rect 7533 431 7743 447
rect 7533 397 7549 431
rect 7727 397 7743 431
rect 7533 350 7743 397
rect 7801 431 8011 447
rect 7801 397 7817 431
rect 7995 397 8011 431
rect 7801 350 8011 397
rect 8069 431 8279 447
rect 8069 397 8085 431
rect 8263 397 8279 431
rect 8069 350 8279 397
rect 8337 431 8547 447
rect 8337 397 8353 431
rect 8531 397 8547 431
rect 8337 350 8547 397
rect 8605 431 8815 447
rect 8605 397 8621 431
rect 8799 397 8815 431
rect 8605 350 8815 397
rect 8873 431 9083 447
rect 8873 397 8889 431
rect 9067 397 9083 431
rect 8873 350 9083 397
rect 9141 431 9351 447
rect 9141 397 9157 431
rect 9335 397 9351 431
rect 9141 350 9351 397
rect 9409 431 9619 447
rect 9409 397 9425 431
rect 9603 397 9619 431
rect 9409 350 9619 397
rect 9677 431 9887 447
rect 9677 397 9693 431
rect 9871 397 9887 431
rect 9677 350 9887 397
rect 9945 431 10155 447
rect 9945 397 9961 431
rect 10139 397 10155 431
rect 9945 350 10155 397
rect 10213 431 10423 447
rect 10213 397 10229 431
rect 10407 397 10423 431
rect 10213 350 10423 397
rect 10481 431 10691 447
rect 10481 397 10497 431
rect 10675 397 10691 431
rect 10481 350 10691 397
rect 10749 431 10959 447
rect 10749 397 10765 431
rect 10943 397 10959 431
rect 10749 350 10959 397
rect 11017 431 11227 447
rect 11017 397 11033 431
rect 11211 397 11227 431
rect 11017 350 11227 397
rect 11285 431 11495 447
rect 11285 397 11301 431
rect 11479 397 11495 431
rect 11285 350 11495 397
rect 11553 431 11763 447
rect 11553 397 11569 431
rect 11747 397 11763 431
rect 11553 350 11763 397
rect 11821 431 12031 447
rect 11821 397 11837 431
rect 12015 397 12031 431
rect 11821 350 12031 397
rect 12089 431 12299 447
rect 12089 397 12105 431
rect 12283 397 12299 431
rect 12089 350 12299 397
rect 12357 431 12567 447
rect 12357 397 12373 431
rect 12551 397 12567 431
rect 12357 350 12567 397
rect 12625 431 12835 447
rect 12625 397 12641 431
rect 12819 397 12835 431
rect 12625 350 12835 397
rect 12893 431 13103 447
rect 12893 397 12909 431
rect 13087 397 13103 431
rect 12893 350 13103 397
rect 13161 431 13371 447
rect 13161 397 13177 431
rect 13355 397 13371 431
rect 13161 350 13371 397
rect -13371 -397 -13161 -350
rect -13371 -431 -13355 -397
rect -13177 -431 -13161 -397
rect -13371 -447 -13161 -431
rect -13103 -397 -12893 -350
rect -13103 -431 -13087 -397
rect -12909 -431 -12893 -397
rect -13103 -447 -12893 -431
rect -12835 -397 -12625 -350
rect -12835 -431 -12819 -397
rect -12641 -431 -12625 -397
rect -12835 -447 -12625 -431
rect -12567 -397 -12357 -350
rect -12567 -431 -12551 -397
rect -12373 -431 -12357 -397
rect -12567 -447 -12357 -431
rect -12299 -397 -12089 -350
rect -12299 -431 -12283 -397
rect -12105 -431 -12089 -397
rect -12299 -447 -12089 -431
rect -12031 -397 -11821 -350
rect -12031 -431 -12015 -397
rect -11837 -431 -11821 -397
rect -12031 -447 -11821 -431
rect -11763 -397 -11553 -350
rect -11763 -431 -11747 -397
rect -11569 -431 -11553 -397
rect -11763 -447 -11553 -431
rect -11495 -397 -11285 -350
rect -11495 -431 -11479 -397
rect -11301 -431 -11285 -397
rect -11495 -447 -11285 -431
rect -11227 -397 -11017 -350
rect -11227 -431 -11211 -397
rect -11033 -431 -11017 -397
rect -11227 -447 -11017 -431
rect -10959 -397 -10749 -350
rect -10959 -431 -10943 -397
rect -10765 -431 -10749 -397
rect -10959 -447 -10749 -431
rect -10691 -397 -10481 -350
rect -10691 -431 -10675 -397
rect -10497 -431 -10481 -397
rect -10691 -447 -10481 -431
rect -10423 -397 -10213 -350
rect -10423 -431 -10407 -397
rect -10229 -431 -10213 -397
rect -10423 -447 -10213 -431
rect -10155 -397 -9945 -350
rect -10155 -431 -10139 -397
rect -9961 -431 -9945 -397
rect -10155 -447 -9945 -431
rect -9887 -397 -9677 -350
rect -9887 -431 -9871 -397
rect -9693 -431 -9677 -397
rect -9887 -447 -9677 -431
rect -9619 -397 -9409 -350
rect -9619 -431 -9603 -397
rect -9425 -431 -9409 -397
rect -9619 -447 -9409 -431
rect -9351 -397 -9141 -350
rect -9351 -431 -9335 -397
rect -9157 -431 -9141 -397
rect -9351 -447 -9141 -431
rect -9083 -397 -8873 -350
rect -9083 -431 -9067 -397
rect -8889 -431 -8873 -397
rect -9083 -447 -8873 -431
rect -8815 -397 -8605 -350
rect -8815 -431 -8799 -397
rect -8621 -431 -8605 -397
rect -8815 -447 -8605 -431
rect -8547 -397 -8337 -350
rect -8547 -431 -8531 -397
rect -8353 -431 -8337 -397
rect -8547 -447 -8337 -431
rect -8279 -397 -8069 -350
rect -8279 -431 -8263 -397
rect -8085 -431 -8069 -397
rect -8279 -447 -8069 -431
rect -8011 -397 -7801 -350
rect -8011 -431 -7995 -397
rect -7817 -431 -7801 -397
rect -8011 -447 -7801 -431
rect -7743 -397 -7533 -350
rect -7743 -431 -7727 -397
rect -7549 -431 -7533 -397
rect -7743 -447 -7533 -431
rect -7475 -397 -7265 -350
rect -7475 -431 -7459 -397
rect -7281 -431 -7265 -397
rect -7475 -447 -7265 -431
rect -7207 -397 -6997 -350
rect -7207 -431 -7191 -397
rect -7013 -431 -6997 -397
rect -7207 -447 -6997 -431
rect -6939 -397 -6729 -350
rect -6939 -431 -6923 -397
rect -6745 -431 -6729 -397
rect -6939 -447 -6729 -431
rect -6671 -397 -6461 -350
rect -6671 -431 -6655 -397
rect -6477 -431 -6461 -397
rect -6671 -447 -6461 -431
rect -6403 -397 -6193 -350
rect -6403 -431 -6387 -397
rect -6209 -431 -6193 -397
rect -6403 -447 -6193 -431
rect -6135 -397 -5925 -350
rect -6135 -431 -6119 -397
rect -5941 -431 -5925 -397
rect -6135 -447 -5925 -431
rect -5867 -397 -5657 -350
rect -5867 -431 -5851 -397
rect -5673 -431 -5657 -397
rect -5867 -447 -5657 -431
rect -5599 -397 -5389 -350
rect -5599 -431 -5583 -397
rect -5405 -431 -5389 -397
rect -5599 -447 -5389 -431
rect -5331 -397 -5121 -350
rect -5331 -431 -5315 -397
rect -5137 -431 -5121 -397
rect -5331 -447 -5121 -431
rect -5063 -397 -4853 -350
rect -5063 -431 -5047 -397
rect -4869 -431 -4853 -397
rect -5063 -447 -4853 -431
rect -4795 -397 -4585 -350
rect -4795 -431 -4779 -397
rect -4601 -431 -4585 -397
rect -4795 -447 -4585 -431
rect -4527 -397 -4317 -350
rect -4527 -431 -4511 -397
rect -4333 -431 -4317 -397
rect -4527 -447 -4317 -431
rect -4259 -397 -4049 -350
rect -4259 -431 -4243 -397
rect -4065 -431 -4049 -397
rect -4259 -447 -4049 -431
rect -3991 -397 -3781 -350
rect -3991 -431 -3975 -397
rect -3797 -431 -3781 -397
rect -3991 -447 -3781 -431
rect -3723 -397 -3513 -350
rect -3723 -431 -3707 -397
rect -3529 -431 -3513 -397
rect -3723 -447 -3513 -431
rect -3455 -397 -3245 -350
rect -3455 -431 -3439 -397
rect -3261 -431 -3245 -397
rect -3455 -447 -3245 -431
rect -3187 -397 -2977 -350
rect -3187 -431 -3171 -397
rect -2993 -431 -2977 -397
rect -3187 -447 -2977 -431
rect -2919 -397 -2709 -350
rect -2919 -431 -2903 -397
rect -2725 -431 -2709 -397
rect -2919 -447 -2709 -431
rect -2651 -397 -2441 -350
rect -2651 -431 -2635 -397
rect -2457 -431 -2441 -397
rect -2651 -447 -2441 -431
rect -2383 -397 -2173 -350
rect -2383 -431 -2367 -397
rect -2189 -431 -2173 -397
rect -2383 -447 -2173 -431
rect -2115 -397 -1905 -350
rect -2115 -431 -2099 -397
rect -1921 -431 -1905 -397
rect -2115 -447 -1905 -431
rect -1847 -397 -1637 -350
rect -1847 -431 -1831 -397
rect -1653 -431 -1637 -397
rect -1847 -447 -1637 -431
rect -1579 -397 -1369 -350
rect -1579 -431 -1563 -397
rect -1385 -431 -1369 -397
rect -1579 -447 -1369 -431
rect -1311 -397 -1101 -350
rect -1311 -431 -1295 -397
rect -1117 -431 -1101 -397
rect -1311 -447 -1101 -431
rect -1043 -397 -833 -350
rect -1043 -431 -1027 -397
rect -849 -431 -833 -397
rect -1043 -447 -833 -431
rect -775 -397 -565 -350
rect -775 -431 -759 -397
rect -581 -431 -565 -397
rect -775 -447 -565 -431
rect -507 -397 -297 -350
rect -507 -431 -491 -397
rect -313 -431 -297 -397
rect -507 -447 -297 -431
rect -239 -397 -29 -350
rect -239 -431 -223 -397
rect -45 -431 -29 -397
rect -239 -447 -29 -431
rect 29 -397 239 -350
rect 29 -431 45 -397
rect 223 -431 239 -397
rect 29 -447 239 -431
rect 297 -397 507 -350
rect 297 -431 313 -397
rect 491 -431 507 -397
rect 297 -447 507 -431
rect 565 -397 775 -350
rect 565 -431 581 -397
rect 759 -431 775 -397
rect 565 -447 775 -431
rect 833 -397 1043 -350
rect 833 -431 849 -397
rect 1027 -431 1043 -397
rect 833 -447 1043 -431
rect 1101 -397 1311 -350
rect 1101 -431 1117 -397
rect 1295 -431 1311 -397
rect 1101 -447 1311 -431
rect 1369 -397 1579 -350
rect 1369 -431 1385 -397
rect 1563 -431 1579 -397
rect 1369 -447 1579 -431
rect 1637 -397 1847 -350
rect 1637 -431 1653 -397
rect 1831 -431 1847 -397
rect 1637 -447 1847 -431
rect 1905 -397 2115 -350
rect 1905 -431 1921 -397
rect 2099 -431 2115 -397
rect 1905 -447 2115 -431
rect 2173 -397 2383 -350
rect 2173 -431 2189 -397
rect 2367 -431 2383 -397
rect 2173 -447 2383 -431
rect 2441 -397 2651 -350
rect 2441 -431 2457 -397
rect 2635 -431 2651 -397
rect 2441 -447 2651 -431
rect 2709 -397 2919 -350
rect 2709 -431 2725 -397
rect 2903 -431 2919 -397
rect 2709 -447 2919 -431
rect 2977 -397 3187 -350
rect 2977 -431 2993 -397
rect 3171 -431 3187 -397
rect 2977 -447 3187 -431
rect 3245 -397 3455 -350
rect 3245 -431 3261 -397
rect 3439 -431 3455 -397
rect 3245 -447 3455 -431
rect 3513 -397 3723 -350
rect 3513 -431 3529 -397
rect 3707 -431 3723 -397
rect 3513 -447 3723 -431
rect 3781 -397 3991 -350
rect 3781 -431 3797 -397
rect 3975 -431 3991 -397
rect 3781 -447 3991 -431
rect 4049 -397 4259 -350
rect 4049 -431 4065 -397
rect 4243 -431 4259 -397
rect 4049 -447 4259 -431
rect 4317 -397 4527 -350
rect 4317 -431 4333 -397
rect 4511 -431 4527 -397
rect 4317 -447 4527 -431
rect 4585 -397 4795 -350
rect 4585 -431 4601 -397
rect 4779 -431 4795 -397
rect 4585 -447 4795 -431
rect 4853 -397 5063 -350
rect 4853 -431 4869 -397
rect 5047 -431 5063 -397
rect 4853 -447 5063 -431
rect 5121 -397 5331 -350
rect 5121 -431 5137 -397
rect 5315 -431 5331 -397
rect 5121 -447 5331 -431
rect 5389 -397 5599 -350
rect 5389 -431 5405 -397
rect 5583 -431 5599 -397
rect 5389 -447 5599 -431
rect 5657 -397 5867 -350
rect 5657 -431 5673 -397
rect 5851 -431 5867 -397
rect 5657 -447 5867 -431
rect 5925 -397 6135 -350
rect 5925 -431 5941 -397
rect 6119 -431 6135 -397
rect 5925 -447 6135 -431
rect 6193 -397 6403 -350
rect 6193 -431 6209 -397
rect 6387 -431 6403 -397
rect 6193 -447 6403 -431
rect 6461 -397 6671 -350
rect 6461 -431 6477 -397
rect 6655 -431 6671 -397
rect 6461 -447 6671 -431
rect 6729 -397 6939 -350
rect 6729 -431 6745 -397
rect 6923 -431 6939 -397
rect 6729 -447 6939 -431
rect 6997 -397 7207 -350
rect 6997 -431 7013 -397
rect 7191 -431 7207 -397
rect 6997 -447 7207 -431
rect 7265 -397 7475 -350
rect 7265 -431 7281 -397
rect 7459 -431 7475 -397
rect 7265 -447 7475 -431
rect 7533 -397 7743 -350
rect 7533 -431 7549 -397
rect 7727 -431 7743 -397
rect 7533 -447 7743 -431
rect 7801 -397 8011 -350
rect 7801 -431 7817 -397
rect 7995 -431 8011 -397
rect 7801 -447 8011 -431
rect 8069 -397 8279 -350
rect 8069 -431 8085 -397
rect 8263 -431 8279 -397
rect 8069 -447 8279 -431
rect 8337 -397 8547 -350
rect 8337 -431 8353 -397
rect 8531 -431 8547 -397
rect 8337 -447 8547 -431
rect 8605 -397 8815 -350
rect 8605 -431 8621 -397
rect 8799 -431 8815 -397
rect 8605 -447 8815 -431
rect 8873 -397 9083 -350
rect 8873 -431 8889 -397
rect 9067 -431 9083 -397
rect 8873 -447 9083 -431
rect 9141 -397 9351 -350
rect 9141 -431 9157 -397
rect 9335 -431 9351 -397
rect 9141 -447 9351 -431
rect 9409 -397 9619 -350
rect 9409 -431 9425 -397
rect 9603 -431 9619 -397
rect 9409 -447 9619 -431
rect 9677 -397 9887 -350
rect 9677 -431 9693 -397
rect 9871 -431 9887 -397
rect 9677 -447 9887 -431
rect 9945 -397 10155 -350
rect 9945 -431 9961 -397
rect 10139 -431 10155 -397
rect 9945 -447 10155 -431
rect 10213 -397 10423 -350
rect 10213 -431 10229 -397
rect 10407 -431 10423 -397
rect 10213 -447 10423 -431
rect 10481 -397 10691 -350
rect 10481 -431 10497 -397
rect 10675 -431 10691 -397
rect 10481 -447 10691 -431
rect 10749 -397 10959 -350
rect 10749 -431 10765 -397
rect 10943 -431 10959 -397
rect 10749 -447 10959 -431
rect 11017 -397 11227 -350
rect 11017 -431 11033 -397
rect 11211 -431 11227 -397
rect 11017 -447 11227 -431
rect 11285 -397 11495 -350
rect 11285 -431 11301 -397
rect 11479 -431 11495 -397
rect 11285 -447 11495 -431
rect 11553 -397 11763 -350
rect 11553 -431 11569 -397
rect 11747 -431 11763 -397
rect 11553 -447 11763 -431
rect 11821 -397 12031 -350
rect 11821 -431 11837 -397
rect 12015 -431 12031 -397
rect 11821 -447 12031 -431
rect 12089 -397 12299 -350
rect 12089 -431 12105 -397
rect 12283 -431 12299 -397
rect 12089 -447 12299 -431
rect 12357 -397 12567 -350
rect 12357 -431 12373 -397
rect 12551 -431 12567 -397
rect 12357 -447 12567 -431
rect 12625 -397 12835 -350
rect 12625 -431 12641 -397
rect 12819 -431 12835 -397
rect 12625 -447 12835 -431
rect 12893 -397 13103 -350
rect 12893 -431 12909 -397
rect 13087 -431 13103 -397
rect 12893 -447 13103 -431
rect 13161 -397 13371 -350
rect 13161 -431 13177 -397
rect 13355 -431 13371 -397
rect 13161 -447 13371 -431
<< polycont >>
rect -13355 397 -13177 431
rect -13087 397 -12909 431
rect -12819 397 -12641 431
rect -12551 397 -12373 431
rect -12283 397 -12105 431
rect -12015 397 -11837 431
rect -11747 397 -11569 431
rect -11479 397 -11301 431
rect -11211 397 -11033 431
rect -10943 397 -10765 431
rect -10675 397 -10497 431
rect -10407 397 -10229 431
rect -10139 397 -9961 431
rect -9871 397 -9693 431
rect -9603 397 -9425 431
rect -9335 397 -9157 431
rect -9067 397 -8889 431
rect -8799 397 -8621 431
rect -8531 397 -8353 431
rect -8263 397 -8085 431
rect -7995 397 -7817 431
rect -7727 397 -7549 431
rect -7459 397 -7281 431
rect -7191 397 -7013 431
rect -6923 397 -6745 431
rect -6655 397 -6477 431
rect -6387 397 -6209 431
rect -6119 397 -5941 431
rect -5851 397 -5673 431
rect -5583 397 -5405 431
rect -5315 397 -5137 431
rect -5047 397 -4869 431
rect -4779 397 -4601 431
rect -4511 397 -4333 431
rect -4243 397 -4065 431
rect -3975 397 -3797 431
rect -3707 397 -3529 431
rect -3439 397 -3261 431
rect -3171 397 -2993 431
rect -2903 397 -2725 431
rect -2635 397 -2457 431
rect -2367 397 -2189 431
rect -2099 397 -1921 431
rect -1831 397 -1653 431
rect -1563 397 -1385 431
rect -1295 397 -1117 431
rect -1027 397 -849 431
rect -759 397 -581 431
rect -491 397 -313 431
rect -223 397 -45 431
rect 45 397 223 431
rect 313 397 491 431
rect 581 397 759 431
rect 849 397 1027 431
rect 1117 397 1295 431
rect 1385 397 1563 431
rect 1653 397 1831 431
rect 1921 397 2099 431
rect 2189 397 2367 431
rect 2457 397 2635 431
rect 2725 397 2903 431
rect 2993 397 3171 431
rect 3261 397 3439 431
rect 3529 397 3707 431
rect 3797 397 3975 431
rect 4065 397 4243 431
rect 4333 397 4511 431
rect 4601 397 4779 431
rect 4869 397 5047 431
rect 5137 397 5315 431
rect 5405 397 5583 431
rect 5673 397 5851 431
rect 5941 397 6119 431
rect 6209 397 6387 431
rect 6477 397 6655 431
rect 6745 397 6923 431
rect 7013 397 7191 431
rect 7281 397 7459 431
rect 7549 397 7727 431
rect 7817 397 7995 431
rect 8085 397 8263 431
rect 8353 397 8531 431
rect 8621 397 8799 431
rect 8889 397 9067 431
rect 9157 397 9335 431
rect 9425 397 9603 431
rect 9693 397 9871 431
rect 9961 397 10139 431
rect 10229 397 10407 431
rect 10497 397 10675 431
rect 10765 397 10943 431
rect 11033 397 11211 431
rect 11301 397 11479 431
rect 11569 397 11747 431
rect 11837 397 12015 431
rect 12105 397 12283 431
rect 12373 397 12551 431
rect 12641 397 12819 431
rect 12909 397 13087 431
rect 13177 397 13355 431
rect -13355 -431 -13177 -397
rect -13087 -431 -12909 -397
rect -12819 -431 -12641 -397
rect -12551 -431 -12373 -397
rect -12283 -431 -12105 -397
rect -12015 -431 -11837 -397
rect -11747 -431 -11569 -397
rect -11479 -431 -11301 -397
rect -11211 -431 -11033 -397
rect -10943 -431 -10765 -397
rect -10675 -431 -10497 -397
rect -10407 -431 -10229 -397
rect -10139 -431 -9961 -397
rect -9871 -431 -9693 -397
rect -9603 -431 -9425 -397
rect -9335 -431 -9157 -397
rect -9067 -431 -8889 -397
rect -8799 -431 -8621 -397
rect -8531 -431 -8353 -397
rect -8263 -431 -8085 -397
rect -7995 -431 -7817 -397
rect -7727 -431 -7549 -397
rect -7459 -431 -7281 -397
rect -7191 -431 -7013 -397
rect -6923 -431 -6745 -397
rect -6655 -431 -6477 -397
rect -6387 -431 -6209 -397
rect -6119 -431 -5941 -397
rect -5851 -431 -5673 -397
rect -5583 -431 -5405 -397
rect -5315 -431 -5137 -397
rect -5047 -431 -4869 -397
rect -4779 -431 -4601 -397
rect -4511 -431 -4333 -397
rect -4243 -431 -4065 -397
rect -3975 -431 -3797 -397
rect -3707 -431 -3529 -397
rect -3439 -431 -3261 -397
rect -3171 -431 -2993 -397
rect -2903 -431 -2725 -397
rect -2635 -431 -2457 -397
rect -2367 -431 -2189 -397
rect -2099 -431 -1921 -397
rect -1831 -431 -1653 -397
rect -1563 -431 -1385 -397
rect -1295 -431 -1117 -397
rect -1027 -431 -849 -397
rect -759 -431 -581 -397
rect -491 -431 -313 -397
rect -223 -431 -45 -397
rect 45 -431 223 -397
rect 313 -431 491 -397
rect 581 -431 759 -397
rect 849 -431 1027 -397
rect 1117 -431 1295 -397
rect 1385 -431 1563 -397
rect 1653 -431 1831 -397
rect 1921 -431 2099 -397
rect 2189 -431 2367 -397
rect 2457 -431 2635 -397
rect 2725 -431 2903 -397
rect 2993 -431 3171 -397
rect 3261 -431 3439 -397
rect 3529 -431 3707 -397
rect 3797 -431 3975 -397
rect 4065 -431 4243 -397
rect 4333 -431 4511 -397
rect 4601 -431 4779 -397
rect 4869 -431 5047 -397
rect 5137 -431 5315 -397
rect 5405 -431 5583 -397
rect 5673 -431 5851 -397
rect 5941 -431 6119 -397
rect 6209 -431 6387 -397
rect 6477 -431 6655 -397
rect 6745 -431 6923 -397
rect 7013 -431 7191 -397
rect 7281 -431 7459 -397
rect 7549 -431 7727 -397
rect 7817 -431 7995 -397
rect 8085 -431 8263 -397
rect 8353 -431 8531 -397
rect 8621 -431 8799 -397
rect 8889 -431 9067 -397
rect 9157 -431 9335 -397
rect 9425 -431 9603 -397
rect 9693 -431 9871 -397
rect 9961 -431 10139 -397
rect 10229 -431 10407 -397
rect 10497 -431 10675 -397
rect 10765 -431 10943 -397
rect 11033 -431 11211 -397
rect 11301 -431 11479 -397
rect 11569 -431 11747 -397
rect 11837 -431 12015 -397
rect 12105 -431 12283 -397
rect 12373 -431 12551 -397
rect 12641 -431 12819 -397
rect 12909 -431 13087 -397
rect 13177 -431 13355 -397
<< locali >>
rect -13531 499 -13435 533
rect 13435 499 13531 533
rect -13531 437 -13497 499
rect 13497 437 13531 499
rect -13371 397 -13355 431
rect -13177 397 -13161 431
rect -13103 397 -13087 431
rect -12909 397 -12893 431
rect -12835 397 -12819 431
rect -12641 397 -12625 431
rect -12567 397 -12551 431
rect -12373 397 -12357 431
rect -12299 397 -12283 431
rect -12105 397 -12089 431
rect -12031 397 -12015 431
rect -11837 397 -11821 431
rect -11763 397 -11747 431
rect -11569 397 -11553 431
rect -11495 397 -11479 431
rect -11301 397 -11285 431
rect -11227 397 -11211 431
rect -11033 397 -11017 431
rect -10959 397 -10943 431
rect -10765 397 -10749 431
rect -10691 397 -10675 431
rect -10497 397 -10481 431
rect -10423 397 -10407 431
rect -10229 397 -10213 431
rect -10155 397 -10139 431
rect -9961 397 -9945 431
rect -9887 397 -9871 431
rect -9693 397 -9677 431
rect -9619 397 -9603 431
rect -9425 397 -9409 431
rect -9351 397 -9335 431
rect -9157 397 -9141 431
rect -9083 397 -9067 431
rect -8889 397 -8873 431
rect -8815 397 -8799 431
rect -8621 397 -8605 431
rect -8547 397 -8531 431
rect -8353 397 -8337 431
rect -8279 397 -8263 431
rect -8085 397 -8069 431
rect -8011 397 -7995 431
rect -7817 397 -7801 431
rect -7743 397 -7727 431
rect -7549 397 -7533 431
rect -7475 397 -7459 431
rect -7281 397 -7265 431
rect -7207 397 -7191 431
rect -7013 397 -6997 431
rect -6939 397 -6923 431
rect -6745 397 -6729 431
rect -6671 397 -6655 431
rect -6477 397 -6461 431
rect -6403 397 -6387 431
rect -6209 397 -6193 431
rect -6135 397 -6119 431
rect -5941 397 -5925 431
rect -5867 397 -5851 431
rect -5673 397 -5657 431
rect -5599 397 -5583 431
rect -5405 397 -5389 431
rect -5331 397 -5315 431
rect -5137 397 -5121 431
rect -5063 397 -5047 431
rect -4869 397 -4853 431
rect -4795 397 -4779 431
rect -4601 397 -4585 431
rect -4527 397 -4511 431
rect -4333 397 -4317 431
rect -4259 397 -4243 431
rect -4065 397 -4049 431
rect -3991 397 -3975 431
rect -3797 397 -3781 431
rect -3723 397 -3707 431
rect -3529 397 -3513 431
rect -3455 397 -3439 431
rect -3261 397 -3245 431
rect -3187 397 -3171 431
rect -2993 397 -2977 431
rect -2919 397 -2903 431
rect -2725 397 -2709 431
rect -2651 397 -2635 431
rect -2457 397 -2441 431
rect -2383 397 -2367 431
rect -2189 397 -2173 431
rect -2115 397 -2099 431
rect -1921 397 -1905 431
rect -1847 397 -1831 431
rect -1653 397 -1637 431
rect -1579 397 -1563 431
rect -1385 397 -1369 431
rect -1311 397 -1295 431
rect -1117 397 -1101 431
rect -1043 397 -1027 431
rect -849 397 -833 431
rect -775 397 -759 431
rect -581 397 -565 431
rect -507 397 -491 431
rect -313 397 -297 431
rect -239 397 -223 431
rect -45 397 -29 431
rect 29 397 45 431
rect 223 397 239 431
rect 297 397 313 431
rect 491 397 507 431
rect 565 397 581 431
rect 759 397 775 431
rect 833 397 849 431
rect 1027 397 1043 431
rect 1101 397 1117 431
rect 1295 397 1311 431
rect 1369 397 1385 431
rect 1563 397 1579 431
rect 1637 397 1653 431
rect 1831 397 1847 431
rect 1905 397 1921 431
rect 2099 397 2115 431
rect 2173 397 2189 431
rect 2367 397 2383 431
rect 2441 397 2457 431
rect 2635 397 2651 431
rect 2709 397 2725 431
rect 2903 397 2919 431
rect 2977 397 2993 431
rect 3171 397 3187 431
rect 3245 397 3261 431
rect 3439 397 3455 431
rect 3513 397 3529 431
rect 3707 397 3723 431
rect 3781 397 3797 431
rect 3975 397 3991 431
rect 4049 397 4065 431
rect 4243 397 4259 431
rect 4317 397 4333 431
rect 4511 397 4527 431
rect 4585 397 4601 431
rect 4779 397 4795 431
rect 4853 397 4869 431
rect 5047 397 5063 431
rect 5121 397 5137 431
rect 5315 397 5331 431
rect 5389 397 5405 431
rect 5583 397 5599 431
rect 5657 397 5673 431
rect 5851 397 5867 431
rect 5925 397 5941 431
rect 6119 397 6135 431
rect 6193 397 6209 431
rect 6387 397 6403 431
rect 6461 397 6477 431
rect 6655 397 6671 431
rect 6729 397 6745 431
rect 6923 397 6939 431
rect 6997 397 7013 431
rect 7191 397 7207 431
rect 7265 397 7281 431
rect 7459 397 7475 431
rect 7533 397 7549 431
rect 7727 397 7743 431
rect 7801 397 7817 431
rect 7995 397 8011 431
rect 8069 397 8085 431
rect 8263 397 8279 431
rect 8337 397 8353 431
rect 8531 397 8547 431
rect 8605 397 8621 431
rect 8799 397 8815 431
rect 8873 397 8889 431
rect 9067 397 9083 431
rect 9141 397 9157 431
rect 9335 397 9351 431
rect 9409 397 9425 431
rect 9603 397 9619 431
rect 9677 397 9693 431
rect 9871 397 9887 431
rect 9945 397 9961 431
rect 10139 397 10155 431
rect 10213 397 10229 431
rect 10407 397 10423 431
rect 10481 397 10497 431
rect 10675 397 10691 431
rect 10749 397 10765 431
rect 10943 397 10959 431
rect 11017 397 11033 431
rect 11211 397 11227 431
rect 11285 397 11301 431
rect 11479 397 11495 431
rect 11553 397 11569 431
rect 11747 397 11763 431
rect 11821 397 11837 431
rect 12015 397 12031 431
rect 12089 397 12105 431
rect 12283 397 12299 431
rect 12357 397 12373 431
rect 12551 397 12567 431
rect 12625 397 12641 431
rect 12819 397 12835 431
rect 12893 397 12909 431
rect 13087 397 13103 431
rect 13161 397 13177 431
rect 13355 397 13371 431
rect -13417 338 -13383 354
rect -13417 -354 -13383 -338
rect -13149 338 -13115 354
rect -13149 -354 -13115 -338
rect -12881 338 -12847 354
rect -12881 -354 -12847 -338
rect -12613 338 -12579 354
rect -12613 -354 -12579 -338
rect -12345 338 -12311 354
rect -12345 -354 -12311 -338
rect -12077 338 -12043 354
rect -12077 -354 -12043 -338
rect -11809 338 -11775 354
rect -11809 -354 -11775 -338
rect -11541 338 -11507 354
rect -11541 -354 -11507 -338
rect -11273 338 -11239 354
rect -11273 -354 -11239 -338
rect -11005 338 -10971 354
rect -11005 -354 -10971 -338
rect -10737 338 -10703 354
rect -10737 -354 -10703 -338
rect -10469 338 -10435 354
rect -10469 -354 -10435 -338
rect -10201 338 -10167 354
rect -10201 -354 -10167 -338
rect -9933 338 -9899 354
rect -9933 -354 -9899 -338
rect -9665 338 -9631 354
rect -9665 -354 -9631 -338
rect -9397 338 -9363 354
rect -9397 -354 -9363 -338
rect -9129 338 -9095 354
rect -9129 -354 -9095 -338
rect -8861 338 -8827 354
rect -8861 -354 -8827 -338
rect -8593 338 -8559 354
rect -8593 -354 -8559 -338
rect -8325 338 -8291 354
rect -8325 -354 -8291 -338
rect -8057 338 -8023 354
rect -8057 -354 -8023 -338
rect -7789 338 -7755 354
rect -7789 -354 -7755 -338
rect -7521 338 -7487 354
rect -7521 -354 -7487 -338
rect -7253 338 -7219 354
rect -7253 -354 -7219 -338
rect -6985 338 -6951 354
rect -6985 -354 -6951 -338
rect -6717 338 -6683 354
rect -6717 -354 -6683 -338
rect -6449 338 -6415 354
rect -6449 -354 -6415 -338
rect -6181 338 -6147 354
rect -6181 -354 -6147 -338
rect -5913 338 -5879 354
rect -5913 -354 -5879 -338
rect -5645 338 -5611 354
rect -5645 -354 -5611 -338
rect -5377 338 -5343 354
rect -5377 -354 -5343 -338
rect -5109 338 -5075 354
rect -5109 -354 -5075 -338
rect -4841 338 -4807 354
rect -4841 -354 -4807 -338
rect -4573 338 -4539 354
rect -4573 -354 -4539 -338
rect -4305 338 -4271 354
rect -4305 -354 -4271 -338
rect -4037 338 -4003 354
rect -4037 -354 -4003 -338
rect -3769 338 -3735 354
rect -3769 -354 -3735 -338
rect -3501 338 -3467 354
rect -3501 -354 -3467 -338
rect -3233 338 -3199 354
rect -3233 -354 -3199 -338
rect -2965 338 -2931 354
rect -2965 -354 -2931 -338
rect -2697 338 -2663 354
rect -2697 -354 -2663 -338
rect -2429 338 -2395 354
rect -2429 -354 -2395 -338
rect -2161 338 -2127 354
rect -2161 -354 -2127 -338
rect -1893 338 -1859 354
rect -1893 -354 -1859 -338
rect -1625 338 -1591 354
rect -1625 -354 -1591 -338
rect -1357 338 -1323 354
rect -1357 -354 -1323 -338
rect -1089 338 -1055 354
rect -1089 -354 -1055 -338
rect -821 338 -787 354
rect -821 -354 -787 -338
rect -553 338 -519 354
rect -553 -354 -519 -338
rect -285 338 -251 354
rect -285 -354 -251 -338
rect -17 338 17 354
rect -17 -354 17 -338
rect 251 338 285 354
rect 251 -354 285 -338
rect 519 338 553 354
rect 519 -354 553 -338
rect 787 338 821 354
rect 787 -354 821 -338
rect 1055 338 1089 354
rect 1055 -354 1089 -338
rect 1323 338 1357 354
rect 1323 -354 1357 -338
rect 1591 338 1625 354
rect 1591 -354 1625 -338
rect 1859 338 1893 354
rect 1859 -354 1893 -338
rect 2127 338 2161 354
rect 2127 -354 2161 -338
rect 2395 338 2429 354
rect 2395 -354 2429 -338
rect 2663 338 2697 354
rect 2663 -354 2697 -338
rect 2931 338 2965 354
rect 2931 -354 2965 -338
rect 3199 338 3233 354
rect 3199 -354 3233 -338
rect 3467 338 3501 354
rect 3467 -354 3501 -338
rect 3735 338 3769 354
rect 3735 -354 3769 -338
rect 4003 338 4037 354
rect 4003 -354 4037 -338
rect 4271 338 4305 354
rect 4271 -354 4305 -338
rect 4539 338 4573 354
rect 4539 -354 4573 -338
rect 4807 338 4841 354
rect 4807 -354 4841 -338
rect 5075 338 5109 354
rect 5075 -354 5109 -338
rect 5343 338 5377 354
rect 5343 -354 5377 -338
rect 5611 338 5645 354
rect 5611 -354 5645 -338
rect 5879 338 5913 354
rect 5879 -354 5913 -338
rect 6147 338 6181 354
rect 6147 -354 6181 -338
rect 6415 338 6449 354
rect 6415 -354 6449 -338
rect 6683 338 6717 354
rect 6683 -354 6717 -338
rect 6951 338 6985 354
rect 6951 -354 6985 -338
rect 7219 338 7253 354
rect 7219 -354 7253 -338
rect 7487 338 7521 354
rect 7487 -354 7521 -338
rect 7755 338 7789 354
rect 7755 -354 7789 -338
rect 8023 338 8057 354
rect 8023 -354 8057 -338
rect 8291 338 8325 354
rect 8291 -354 8325 -338
rect 8559 338 8593 354
rect 8559 -354 8593 -338
rect 8827 338 8861 354
rect 8827 -354 8861 -338
rect 9095 338 9129 354
rect 9095 -354 9129 -338
rect 9363 338 9397 354
rect 9363 -354 9397 -338
rect 9631 338 9665 354
rect 9631 -354 9665 -338
rect 9899 338 9933 354
rect 9899 -354 9933 -338
rect 10167 338 10201 354
rect 10167 -354 10201 -338
rect 10435 338 10469 354
rect 10435 -354 10469 -338
rect 10703 338 10737 354
rect 10703 -354 10737 -338
rect 10971 338 11005 354
rect 10971 -354 11005 -338
rect 11239 338 11273 354
rect 11239 -354 11273 -338
rect 11507 338 11541 354
rect 11507 -354 11541 -338
rect 11775 338 11809 354
rect 11775 -354 11809 -338
rect 12043 338 12077 354
rect 12043 -354 12077 -338
rect 12311 338 12345 354
rect 12311 -354 12345 -338
rect 12579 338 12613 354
rect 12579 -354 12613 -338
rect 12847 338 12881 354
rect 12847 -354 12881 -338
rect 13115 338 13149 354
rect 13115 -354 13149 -338
rect 13383 338 13417 354
rect 13383 -354 13417 -338
rect -13371 -431 -13355 -397
rect -13177 -431 -13161 -397
rect -13103 -431 -13087 -397
rect -12909 -431 -12893 -397
rect -12835 -431 -12819 -397
rect -12641 -431 -12625 -397
rect -12567 -431 -12551 -397
rect -12373 -431 -12357 -397
rect -12299 -431 -12283 -397
rect -12105 -431 -12089 -397
rect -12031 -431 -12015 -397
rect -11837 -431 -11821 -397
rect -11763 -431 -11747 -397
rect -11569 -431 -11553 -397
rect -11495 -431 -11479 -397
rect -11301 -431 -11285 -397
rect -11227 -431 -11211 -397
rect -11033 -431 -11017 -397
rect -10959 -431 -10943 -397
rect -10765 -431 -10749 -397
rect -10691 -431 -10675 -397
rect -10497 -431 -10481 -397
rect -10423 -431 -10407 -397
rect -10229 -431 -10213 -397
rect -10155 -431 -10139 -397
rect -9961 -431 -9945 -397
rect -9887 -431 -9871 -397
rect -9693 -431 -9677 -397
rect -9619 -431 -9603 -397
rect -9425 -431 -9409 -397
rect -9351 -431 -9335 -397
rect -9157 -431 -9141 -397
rect -9083 -431 -9067 -397
rect -8889 -431 -8873 -397
rect -8815 -431 -8799 -397
rect -8621 -431 -8605 -397
rect -8547 -431 -8531 -397
rect -8353 -431 -8337 -397
rect -8279 -431 -8263 -397
rect -8085 -431 -8069 -397
rect -8011 -431 -7995 -397
rect -7817 -431 -7801 -397
rect -7743 -431 -7727 -397
rect -7549 -431 -7533 -397
rect -7475 -431 -7459 -397
rect -7281 -431 -7265 -397
rect -7207 -431 -7191 -397
rect -7013 -431 -6997 -397
rect -6939 -431 -6923 -397
rect -6745 -431 -6729 -397
rect -6671 -431 -6655 -397
rect -6477 -431 -6461 -397
rect -6403 -431 -6387 -397
rect -6209 -431 -6193 -397
rect -6135 -431 -6119 -397
rect -5941 -431 -5925 -397
rect -5867 -431 -5851 -397
rect -5673 -431 -5657 -397
rect -5599 -431 -5583 -397
rect -5405 -431 -5389 -397
rect -5331 -431 -5315 -397
rect -5137 -431 -5121 -397
rect -5063 -431 -5047 -397
rect -4869 -431 -4853 -397
rect -4795 -431 -4779 -397
rect -4601 -431 -4585 -397
rect -4527 -431 -4511 -397
rect -4333 -431 -4317 -397
rect -4259 -431 -4243 -397
rect -4065 -431 -4049 -397
rect -3991 -431 -3975 -397
rect -3797 -431 -3781 -397
rect -3723 -431 -3707 -397
rect -3529 -431 -3513 -397
rect -3455 -431 -3439 -397
rect -3261 -431 -3245 -397
rect -3187 -431 -3171 -397
rect -2993 -431 -2977 -397
rect -2919 -431 -2903 -397
rect -2725 -431 -2709 -397
rect -2651 -431 -2635 -397
rect -2457 -431 -2441 -397
rect -2383 -431 -2367 -397
rect -2189 -431 -2173 -397
rect -2115 -431 -2099 -397
rect -1921 -431 -1905 -397
rect -1847 -431 -1831 -397
rect -1653 -431 -1637 -397
rect -1579 -431 -1563 -397
rect -1385 -431 -1369 -397
rect -1311 -431 -1295 -397
rect -1117 -431 -1101 -397
rect -1043 -431 -1027 -397
rect -849 -431 -833 -397
rect -775 -431 -759 -397
rect -581 -431 -565 -397
rect -507 -431 -491 -397
rect -313 -431 -297 -397
rect -239 -431 -223 -397
rect -45 -431 -29 -397
rect 29 -431 45 -397
rect 223 -431 239 -397
rect 297 -431 313 -397
rect 491 -431 507 -397
rect 565 -431 581 -397
rect 759 -431 775 -397
rect 833 -431 849 -397
rect 1027 -431 1043 -397
rect 1101 -431 1117 -397
rect 1295 -431 1311 -397
rect 1369 -431 1385 -397
rect 1563 -431 1579 -397
rect 1637 -431 1653 -397
rect 1831 -431 1847 -397
rect 1905 -431 1921 -397
rect 2099 -431 2115 -397
rect 2173 -431 2189 -397
rect 2367 -431 2383 -397
rect 2441 -431 2457 -397
rect 2635 -431 2651 -397
rect 2709 -431 2725 -397
rect 2903 -431 2919 -397
rect 2977 -431 2993 -397
rect 3171 -431 3187 -397
rect 3245 -431 3261 -397
rect 3439 -431 3455 -397
rect 3513 -431 3529 -397
rect 3707 -431 3723 -397
rect 3781 -431 3797 -397
rect 3975 -431 3991 -397
rect 4049 -431 4065 -397
rect 4243 -431 4259 -397
rect 4317 -431 4333 -397
rect 4511 -431 4527 -397
rect 4585 -431 4601 -397
rect 4779 -431 4795 -397
rect 4853 -431 4869 -397
rect 5047 -431 5063 -397
rect 5121 -431 5137 -397
rect 5315 -431 5331 -397
rect 5389 -431 5405 -397
rect 5583 -431 5599 -397
rect 5657 -431 5673 -397
rect 5851 -431 5867 -397
rect 5925 -431 5941 -397
rect 6119 -431 6135 -397
rect 6193 -431 6209 -397
rect 6387 -431 6403 -397
rect 6461 -431 6477 -397
rect 6655 -431 6671 -397
rect 6729 -431 6745 -397
rect 6923 -431 6939 -397
rect 6997 -431 7013 -397
rect 7191 -431 7207 -397
rect 7265 -431 7281 -397
rect 7459 -431 7475 -397
rect 7533 -431 7549 -397
rect 7727 -431 7743 -397
rect 7801 -431 7817 -397
rect 7995 -431 8011 -397
rect 8069 -431 8085 -397
rect 8263 -431 8279 -397
rect 8337 -431 8353 -397
rect 8531 -431 8547 -397
rect 8605 -431 8621 -397
rect 8799 -431 8815 -397
rect 8873 -431 8889 -397
rect 9067 -431 9083 -397
rect 9141 -431 9157 -397
rect 9335 -431 9351 -397
rect 9409 -431 9425 -397
rect 9603 -431 9619 -397
rect 9677 -431 9693 -397
rect 9871 -431 9887 -397
rect 9945 -431 9961 -397
rect 10139 -431 10155 -397
rect 10213 -431 10229 -397
rect 10407 -431 10423 -397
rect 10481 -431 10497 -397
rect 10675 -431 10691 -397
rect 10749 -431 10765 -397
rect 10943 -431 10959 -397
rect 11017 -431 11033 -397
rect 11211 -431 11227 -397
rect 11285 -431 11301 -397
rect 11479 -431 11495 -397
rect 11553 -431 11569 -397
rect 11747 -431 11763 -397
rect 11821 -431 11837 -397
rect 12015 -431 12031 -397
rect 12089 -431 12105 -397
rect 12283 -431 12299 -397
rect 12357 -431 12373 -397
rect 12551 -431 12567 -397
rect 12625 -431 12641 -397
rect 12819 -431 12835 -397
rect 12893 -431 12909 -397
rect 13087 -431 13103 -397
rect 13161 -431 13177 -397
rect 13355 -431 13371 -397
rect -13531 -499 -13497 -437
rect 13497 -499 13531 -437
rect -13531 -533 -13435 -499
rect 13435 -533 13531 -499
<< viali >>
rect -13355 397 -13177 431
rect -13087 397 -12909 431
rect -12819 397 -12641 431
rect -12551 397 -12373 431
rect -12283 397 -12105 431
rect -12015 397 -11837 431
rect -11747 397 -11569 431
rect -11479 397 -11301 431
rect -11211 397 -11033 431
rect -10943 397 -10765 431
rect -10675 397 -10497 431
rect -10407 397 -10229 431
rect -10139 397 -9961 431
rect -9871 397 -9693 431
rect -9603 397 -9425 431
rect -9335 397 -9157 431
rect -9067 397 -8889 431
rect -8799 397 -8621 431
rect -8531 397 -8353 431
rect -8263 397 -8085 431
rect -7995 397 -7817 431
rect -7727 397 -7549 431
rect -7459 397 -7281 431
rect -7191 397 -7013 431
rect -6923 397 -6745 431
rect -6655 397 -6477 431
rect -6387 397 -6209 431
rect -6119 397 -5941 431
rect -5851 397 -5673 431
rect -5583 397 -5405 431
rect -5315 397 -5137 431
rect -5047 397 -4869 431
rect -4779 397 -4601 431
rect -4511 397 -4333 431
rect -4243 397 -4065 431
rect -3975 397 -3797 431
rect -3707 397 -3529 431
rect -3439 397 -3261 431
rect -3171 397 -2993 431
rect -2903 397 -2725 431
rect -2635 397 -2457 431
rect -2367 397 -2189 431
rect -2099 397 -1921 431
rect -1831 397 -1653 431
rect -1563 397 -1385 431
rect -1295 397 -1117 431
rect -1027 397 -849 431
rect -759 397 -581 431
rect -491 397 -313 431
rect -223 397 -45 431
rect 45 397 223 431
rect 313 397 491 431
rect 581 397 759 431
rect 849 397 1027 431
rect 1117 397 1295 431
rect 1385 397 1563 431
rect 1653 397 1831 431
rect 1921 397 2099 431
rect 2189 397 2367 431
rect 2457 397 2635 431
rect 2725 397 2903 431
rect 2993 397 3171 431
rect 3261 397 3439 431
rect 3529 397 3707 431
rect 3797 397 3975 431
rect 4065 397 4243 431
rect 4333 397 4511 431
rect 4601 397 4779 431
rect 4869 397 5047 431
rect 5137 397 5315 431
rect 5405 397 5583 431
rect 5673 397 5851 431
rect 5941 397 6119 431
rect 6209 397 6387 431
rect 6477 397 6655 431
rect 6745 397 6923 431
rect 7013 397 7191 431
rect 7281 397 7459 431
rect 7549 397 7727 431
rect 7817 397 7995 431
rect 8085 397 8263 431
rect 8353 397 8531 431
rect 8621 397 8799 431
rect 8889 397 9067 431
rect 9157 397 9335 431
rect 9425 397 9603 431
rect 9693 397 9871 431
rect 9961 397 10139 431
rect 10229 397 10407 431
rect 10497 397 10675 431
rect 10765 397 10943 431
rect 11033 397 11211 431
rect 11301 397 11479 431
rect 11569 397 11747 431
rect 11837 397 12015 431
rect 12105 397 12283 431
rect 12373 397 12551 431
rect 12641 397 12819 431
rect 12909 397 13087 431
rect 13177 397 13355 431
rect -13417 -338 -13383 338
rect -13149 -338 -13115 338
rect -12881 -338 -12847 338
rect -12613 -338 -12579 338
rect -12345 -338 -12311 338
rect -12077 -338 -12043 338
rect -11809 -338 -11775 338
rect -11541 -338 -11507 338
rect -11273 -338 -11239 338
rect -11005 -338 -10971 338
rect -10737 -338 -10703 338
rect -10469 -338 -10435 338
rect -10201 -338 -10167 338
rect -9933 -338 -9899 338
rect -9665 -338 -9631 338
rect -9397 -338 -9363 338
rect -9129 -338 -9095 338
rect -8861 -338 -8827 338
rect -8593 -338 -8559 338
rect -8325 -338 -8291 338
rect -8057 -338 -8023 338
rect -7789 -338 -7755 338
rect -7521 -338 -7487 338
rect -7253 -338 -7219 338
rect -6985 -338 -6951 338
rect -6717 -338 -6683 338
rect -6449 -338 -6415 338
rect -6181 -338 -6147 338
rect -5913 -338 -5879 338
rect -5645 -338 -5611 338
rect -5377 -338 -5343 338
rect -5109 -338 -5075 338
rect -4841 -338 -4807 338
rect -4573 -338 -4539 338
rect -4305 -338 -4271 338
rect -4037 -338 -4003 338
rect -3769 -338 -3735 338
rect -3501 -338 -3467 338
rect -3233 -338 -3199 338
rect -2965 -338 -2931 338
rect -2697 -338 -2663 338
rect -2429 -338 -2395 338
rect -2161 -338 -2127 338
rect -1893 -338 -1859 338
rect -1625 -338 -1591 338
rect -1357 -338 -1323 338
rect -1089 -338 -1055 338
rect -821 -338 -787 338
rect -553 -338 -519 338
rect -285 -338 -251 338
rect -17 -338 17 338
rect 251 -338 285 338
rect 519 -338 553 338
rect 787 -338 821 338
rect 1055 -338 1089 338
rect 1323 -338 1357 338
rect 1591 -338 1625 338
rect 1859 -338 1893 338
rect 2127 -338 2161 338
rect 2395 -338 2429 338
rect 2663 -338 2697 338
rect 2931 -338 2965 338
rect 3199 -338 3233 338
rect 3467 -338 3501 338
rect 3735 -338 3769 338
rect 4003 -338 4037 338
rect 4271 -338 4305 338
rect 4539 -338 4573 338
rect 4807 -338 4841 338
rect 5075 -338 5109 338
rect 5343 -338 5377 338
rect 5611 -338 5645 338
rect 5879 -338 5913 338
rect 6147 -338 6181 338
rect 6415 -338 6449 338
rect 6683 -338 6717 338
rect 6951 -338 6985 338
rect 7219 -338 7253 338
rect 7487 -338 7521 338
rect 7755 -338 7789 338
rect 8023 -338 8057 338
rect 8291 -338 8325 338
rect 8559 -338 8593 338
rect 8827 -338 8861 338
rect 9095 -338 9129 338
rect 9363 -338 9397 338
rect 9631 -338 9665 338
rect 9899 -338 9933 338
rect 10167 -338 10201 338
rect 10435 -338 10469 338
rect 10703 -338 10737 338
rect 10971 -338 11005 338
rect 11239 -338 11273 338
rect 11507 -338 11541 338
rect 11775 -338 11809 338
rect 12043 -338 12077 338
rect 12311 -338 12345 338
rect 12579 -338 12613 338
rect 12847 -338 12881 338
rect 13115 -338 13149 338
rect 13383 -338 13417 338
rect -13355 -431 -13177 -397
rect -13087 -431 -12909 -397
rect -12819 -431 -12641 -397
rect -12551 -431 -12373 -397
rect -12283 -431 -12105 -397
rect -12015 -431 -11837 -397
rect -11747 -431 -11569 -397
rect -11479 -431 -11301 -397
rect -11211 -431 -11033 -397
rect -10943 -431 -10765 -397
rect -10675 -431 -10497 -397
rect -10407 -431 -10229 -397
rect -10139 -431 -9961 -397
rect -9871 -431 -9693 -397
rect -9603 -431 -9425 -397
rect -9335 -431 -9157 -397
rect -9067 -431 -8889 -397
rect -8799 -431 -8621 -397
rect -8531 -431 -8353 -397
rect -8263 -431 -8085 -397
rect -7995 -431 -7817 -397
rect -7727 -431 -7549 -397
rect -7459 -431 -7281 -397
rect -7191 -431 -7013 -397
rect -6923 -431 -6745 -397
rect -6655 -431 -6477 -397
rect -6387 -431 -6209 -397
rect -6119 -431 -5941 -397
rect -5851 -431 -5673 -397
rect -5583 -431 -5405 -397
rect -5315 -431 -5137 -397
rect -5047 -431 -4869 -397
rect -4779 -431 -4601 -397
rect -4511 -431 -4333 -397
rect -4243 -431 -4065 -397
rect -3975 -431 -3797 -397
rect -3707 -431 -3529 -397
rect -3439 -431 -3261 -397
rect -3171 -431 -2993 -397
rect -2903 -431 -2725 -397
rect -2635 -431 -2457 -397
rect -2367 -431 -2189 -397
rect -2099 -431 -1921 -397
rect -1831 -431 -1653 -397
rect -1563 -431 -1385 -397
rect -1295 -431 -1117 -397
rect -1027 -431 -849 -397
rect -759 -431 -581 -397
rect -491 -431 -313 -397
rect -223 -431 -45 -397
rect 45 -431 223 -397
rect 313 -431 491 -397
rect 581 -431 759 -397
rect 849 -431 1027 -397
rect 1117 -431 1295 -397
rect 1385 -431 1563 -397
rect 1653 -431 1831 -397
rect 1921 -431 2099 -397
rect 2189 -431 2367 -397
rect 2457 -431 2635 -397
rect 2725 -431 2903 -397
rect 2993 -431 3171 -397
rect 3261 -431 3439 -397
rect 3529 -431 3707 -397
rect 3797 -431 3975 -397
rect 4065 -431 4243 -397
rect 4333 -431 4511 -397
rect 4601 -431 4779 -397
rect 4869 -431 5047 -397
rect 5137 -431 5315 -397
rect 5405 -431 5583 -397
rect 5673 -431 5851 -397
rect 5941 -431 6119 -397
rect 6209 -431 6387 -397
rect 6477 -431 6655 -397
rect 6745 -431 6923 -397
rect 7013 -431 7191 -397
rect 7281 -431 7459 -397
rect 7549 -431 7727 -397
rect 7817 -431 7995 -397
rect 8085 -431 8263 -397
rect 8353 -431 8531 -397
rect 8621 -431 8799 -397
rect 8889 -431 9067 -397
rect 9157 -431 9335 -397
rect 9425 -431 9603 -397
rect 9693 -431 9871 -397
rect 9961 -431 10139 -397
rect 10229 -431 10407 -397
rect 10497 -431 10675 -397
rect 10765 -431 10943 -397
rect 11033 -431 11211 -397
rect 11301 -431 11479 -397
rect 11569 -431 11747 -397
rect 11837 -431 12015 -397
rect 12105 -431 12283 -397
rect 12373 -431 12551 -397
rect 12641 -431 12819 -397
rect 12909 -431 13087 -397
rect 13177 -431 13355 -397
<< metal1 >>
rect -13367 431 -13165 437
rect -13367 397 -13355 431
rect -13177 397 -13165 431
rect -13367 391 -13165 397
rect -13099 431 -12897 437
rect -13099 397 -13087 431
rect -12909 397 -12897 431
rect -13099 391 -12897 397
rect -12831 431 -12629 437
rect -12831 397 -12819 431
rect -12641 397 -12629 431
rect -12831 391 -12629 397
rect -12563 431 -12361 437
rect -12563 397 -12551 431
rect -12373 397 -12361 431
rect -12563 391 -12361 397
rect -12295 431 -12093 437
rect -12295 397 -12283 431
rect -12105 397 -12093 431
rect -12295 391 -12093 397
rect -12027 431 -11825 437
rect -12027 397 -12015 431
rect -11837 397 -11825 431
rect -12027 391 -11825 397
rect -11759 431 -11557 437
rect -11759 397 -11747 431
rect -11569 397 -11557 431
rect -11759 391 -11557 397
rect -11491 431 -11289 437
rect -11491 397 -11479 431
rect -11301 397 -11289 431
rect -11491 391 -11289 397
rect -11223 431 -11021 437
rect -11223 397 -11211 431
rect -11033 397 -11021 431
rect -11223 391 -11021 397
rect -10955 431 -10753 437
rect -10955 397 -10943 431
rect -10765 397 -10753 431
rect -10955 391 -10753 397
rect -10687 431 -10485 437
rect -10687 397 -10675 431
rect -10497 397 -10485 431
rect -10687 391 -10485 397
rect -10419 431 -10217 437
rect -10419 397 -10407 431
rect -10229 397 -10217 431
rect -10419 391 -10217 397
rect -10151 431 -9949 437
rect -10151 397 -10139 431
rect -9961 397 -9949 431
rect -10151 391 -9949 397
rect -9883 431 -9681 437
rect -9883 397 -9871 431
rect -9693 397 -9681 431
rect -9883 391 -9681 397
rect -9615 431 -9413 437
rect -9615 397 -9603 431
rect -9425 397 -9413 431
rect -9615 391 -9413 397
rect -9347 431 -9145 437
rect -9347 397 -9335 431
rect -9157 397 -9145 431
rect -9347 391 -9145 397
rect -9079 431 -8877 437
rect -9079 397 -9067 431
rect -8889 397 -8877 431
rect -9079 391 -8877 397
rect -8811 431 -8609 437
rect -8811 397 -8799 431
rect -8621 397 -8609 431
rect -8811 391 -8609 397
rect -8543 431 -8341 437
rect -8543 397 -8531 431
rect -8353 397 -8341 431
rect -8543 391 -8341 397
rect -8275 431 -8073 437
rect -8275 397 -8263 431
rect -8085 397 -8073 431
rect -8275 391 -8073 397
rect -8007 431 -7805 437
rect -8007 397 -7995 431
rect -7817 397 -7805 431
rect -8007 391 -7805 397
rect -7739 431 -7537 437
rect -7739 397 -7727 431
rect -7549 397 -7537 431
rect -7739 391 -7537 397
rect -7471 431 -7269 437
rect -7471 397 -7459 431
rect -7281 397 -7269 431
rect -7471 391 -7269 397
rect -7203 431 -7001 437
rect -7203 397 -7191 431
rect -7013 397 -7001 431
rect -7203 391 -7001 397
rect -6935 431 -6733 437
rect -6935 397 -6923 431
rect -6745 397 -6733 431
rect -6935 391 -6733 397
rect -6667 431 -6465 437
rect -6667 397 -6655 431
rect -6477 397 -6465 431
rect -6667 391 -6465 397
rect -6399 431 -6197 437
rect -6399 397 -6387 431
rect -6209 397 -6197 431
rect -6399 391 -6197 397
rect -6131 431 -5929 437
rect -6131 397 -6119 431
rect -5941 397 -5929 431
rect -6131 391 -5929 397
rect -5863 431 -5661 437
rect -5863 397 -5851 431
rect -5673 397 -5661 431
rect -5863 391 -5661 397
rect -5595 431 -5393 437
rect -5595 397 -5583 431
rect -5405 397 -5393 431
rect -5595 391 -5393 397
rect -5327 431 -5125 437
rect -5327 397 -5315 431
rect -5137 397 -5125 431
rect -5327 391 -5125 397
rect -5059 431 -4857 437
rect -5059 397 -5047 431
rect -4869 397 -4857 431
rect -5059 391 -4857 397
rect -4791 431 -4589 437
rect -4791 397 -4779 431
rect -4601 397 -4589 431
rect -4791 391 -4589 397
rect -4523 431 -4321 437
rect -4523 397 -4511 431
rect -4333 397 -4321 431
rect -4523 391 -4321 397
rect -4255 431 -4053 437
rect -4255 397 -4243 431
rect -4065 397 -4053 431
rect -4255 391 -4053 397
rect -3987 431 -3785 437
rect -3987 397 -3975 431
rect -3797 397 -3785 431
rect -3987 391 -3785 397
rect -3719 431 -3517 437
rect -3719 397 -3707 431
rect -3529 397 -3517 431
rect -3719 391 -3517 397
rect -3451 431 -3249 437
rect -3451 397 -3439 431
rect -3261 397 -3249 431
rect -3451 391 -3249 397
rect -3183 431 -2981 437
rect -3183 397 -3171 431
rect -2993 397 -2981 431
rect -3183 391 -2981 397
rect -2915 431 -2713 437
rect -2915 397 -2903 431
rect -2725 397 -2713 431
rect -2915 391 -2713 397
rect -2647 431 -2445 437
rect -2647 397 -2635 431
rect -2457 397 -2445 431
rect -2647 391 -2445 397
rect -2379 431 -2177 437
rect -2379 397 -2367 431
rect -2189 397 -2177 431
rect -2379 391 -2177 397
rect -2111 431 -1909 437
rect -2111 397 -2099 431
rect -1921 397 -1909 431
rect -2111 391 -1909 397
rect -1843 431 -1641 437
rect -1843 397 -1831 431
rect -1653 397 -1641 431
rect -1843 391 -1641 397
rect -1575 431 -1373 437
rect -1575 397 -1563 431
rect -1385 397 -1373 431
rect -1575 391 -1373 397
rect -1307 431 -1105 437
rect -1307 397 -1295 431
rect -1117 397 -1105 431
rect -1307 391 -1105 397
rect -1039 431 -837 437
rect -1039 397 -1027 431
rect -849 397 -837 431
rect -1039 391 -837 397
rect -771 431 -569 437
rect -771 397 -759 431
rect -581 397 -569 431
rect -771 391 -569 397
rect -503 431 -301 437
rect -503 397 -491 431
rect -313 397 -301 431
rect -503 391 -301 397
rect -235 431 -33 437
rect -235 397 -223 431
rect -45 397 -33 431
rect -235 391 -33 397
rect 33 431 235 437
rect 33 397 45 431
rect 223 397 235 431
rect 33 391 235 397
rect 301 431 503 437
rect 301 397 313 431
rect 491 397 503 431
rect 301 391 503 397
rect 569 431 771 437
rect 569 397 581 431
rect 759 397 771 431
rect 569 391 771 397
rect 837 431 1039 437
rect 837 397 849 431
rect 1027 397 1039 431
rect 837 391 1039 397
rect 1105 431 1307 437
rect 1105 397 1117 431
rect 1295 397 1307 431
rect 1105 391 1307 397
rect 1373 431 1575 437
rect 1373 397 1385 431
rect 1563 397 1575 431
rect 1373 391 1575 397
rect 1641 431 1843 437
rect 1641 397 1653 431
rect 1831 397 1843 431
rect 1641 391 1843 397
rect 1909 431 2111 437
rect 1909 397 1921 431
rect 2099 397 2111 431
rect 1909 391 2111 397
rect 2177 431 2379 437
rect 2177 397 2189 431
rect 2367 397 2379 431
rect 2177 391 2379 397
rect 2445 431 2647 437
rect 2445 397 2457 431
rect 2635 397 2647 431
rect 2445 391 2647 397
rect 2713 431 2915 437
rect 2713 397 2725 431
rect 2903 397 2915 431
rect 2713 391 2915 397
rect 2981 431 3183 437
rect 2981 397 2993 431
rect 3171 397 3183 431
rect 2981 391 3183 397
rect 3249 431 3451 437
rect 3249 397 3261 431
rect 3439 397 3451 431
rect 3249 391 3451 397
rect 3517 431 3719 437
rect 3517 397 3529 431
rect 3707 397 3719 431
rect 3517 391 3719 397
rect 3785 431 3987 437
rect 3785 397 3797 431
rect 3975 397 3987 431
rect 3785 391 3987 397
rect 4053 431 4255 437
rect 4053 397 4065 431
rect 4243 397 4255 431
rect 4053 391 4255 397
rect 4321 431 4523 437
rect 4321 397 4333 431
rect 4511 397 4523 431
rect 4321 391 4523 397
rect 4589 431 4791 437
rect 4589 397 4601 431
rect 4779 397 4791 431
rect 4589 391 4791 397
rect 4857 431 5059 437
rect 4857 397 4869 431
rect 5047 397 5059 431
rect 4857 391 5059 397
rect 5125 431 5327 437
rect 5125 397 5137 431
rect 5315 397 5327 431
rect 5125 391 5327 397
rect 5393 431 5595 437
rect 5393 397 5405 431
rect 5583 397 5595 431
rect 5393 391 5595 397
rect 5661 431 5863 437
rect 5661 397 5673 431
rect 5851 397 5863 431
rect 5661 391 5863 397
rect 5929 431 6131 437
rect 5929 397 5941 431
rect 6119 397 6131 431
rect 5929 391 6131 397
rect 6197 431 6399 437
rect 6197 397 6209 431
rect 6387 397 6399 431
rect 6197 391 6399 397
rect 6465 431 6667 437
rect 6465 397 6477 431
rect 6655 397 6667 431
rect 6465 391 6667 397
rect 6733 431 6935 437
rect 6733 397 6745 431
rect 6923 397 6935 431
rect 6733 391 6935 397
rect 7001 431 7203 437
rect 7001 397 7013 431
rect 7191 397 7203 431
rect 7001 391 7203 397
rect 7269 431 7471 437
rect 7269 397 7281 431
rect 7459 397 7471 431
rect 7269 391 7471 397
rect 7537 431 7739 437
rect 7537 397 7549 431
rect 7727 397 7739 431
rect 7537 391 7739 397
rect 7805 431 8007 437
rect 7805 397 7817 431
rect 7995 397 8007 431
rect 7805 391 8007 397
rect 8073 431 8275 437
rect 8073 397 8085 431
rect 8263 397 8275 431
rect 8073 391 8275 397
rect 8341 431 8543 437
rect 8341 397 8353 431
rect 8531 397 8543 431
rect 8341 391 8543 397
rect 8609 431 8811 437
rect 8609 397 8621 431
rect 8799 397 8811 431
rect 8609 391 8811 397
rect 8877 431 9079 437
rect 8877 397 8889 431
rect 9067 397 9079 431
rect 8877 391 9079 397
rect 9145 431 9347 437
rect 9145 397 9157 431
rect 9335 397 9347 431
rect 9145 391 9347 397
rect 9413 431 9615 437
rect 9413 397 9425 431
rect 9603 397 9615 431
rect 9413 391 9615 397
rect 9681 431 9883 437
rect 9681 397 9693 431
rect 9871 397 9883 431
rect 9681 391 9883 397
rect 9949 431 10151 437
rect 9949 397 9961 431
rect 10139 397 10151 431
rect 9949 391 10151 397
rect 10217 431 10419 437
rect 10217 397 10229 431
rect 10407 397 10419 431
rect 10217 391 10419 397
rect 10485 431 10687 437
rect 10485 397 10497 431
rect 10675 397 10687 431
rect 10485 391 10687 397
rect 10753 431 10955 437
rect 10753 397 10765 431
rect 10943 397 10955 431
rect 10753 391 10955 397
rect 11021 431 11223 437
rect 11021 397 11033 431
rect 11211 397 11223 431
rect 11021 391 11223 397
rect 11289 431 11491 437
rect 11289 397 11301 431
rect 11479 397 11491 431
rect 11289 391 11491 397
rect 11557 431 11759 437
rect 11557 397 11569 431
rect 11747 397 11759 431
rect 11557 391 11759 397
rect 11825 431 12027 437
rect 11825 397 11837 431
rect 12015 397 12027 431
rect 11825 391 12027 397
rect 12093 431 12295 437
rect 12093 397 12105 431
rect 12283 397 12295 431
rect 12093 391 12295 397
rect 12361 431 12563 437
rect 12361 397 12373 431
rect 12551 397 12563 431
rect 12361 391 12563 397
rect 12629 431 12831 437
rect 12629 397 12641 431
rect 12819 397 12831 431
rect 12629 391 12831 397
rect 12897 431 13099 437
rect 12897 397 12909 431
rect 13087 397 13099 431
rect 12897 391 13099 397
rect 13165 431 13367 437
rect 13165 397 13177 431
rect 13355 397 13367 431
rect 13165 391 13367 397
rect -13423 338 -13377 350
rect -13423 -338 -13417 338
rect -13383 -338 -13377 338
rect -13423 -350 -13377 -338
rect -13155 338 -13109 350
rect -13155 -338 -13149 338
rect -13115 -338 -13109 338
rect -13155 -350 -13109 -338
rect -12887 338 -12841 350
rect -12887 -338 -12881 338
rect -12847 -338 -12841 338
rect -12887 -350 -12841 -338
rect -12619 338 -12573 350
rect -12619 -338 -12613 338
rect -12579 -338 -12573 338
rect -12619 -350 -12573 -338
rect -12351 338 -12305 350
rect -12351 -338 -12345 338
rect -12311 -338 -12305 338
rect -12351 -350 -12305 -338
rect -12083 338 -12037 350
rect -12083 -338 -12077 338
rect -12043 -338 -12037 338
rect -12083 -350 -12037 -338
rect -11815 338 -11769 350
rect -11815 -338 -11809 338
rect -11775 -338 -11769 338
rect -11815 -350 -11769 -338
rect -11547 338 -11501 350
rect -11547 -338 -11541 338
rect -11507 -338 -11501 338
rect -11547 -350 -11501 -338
rect -11279 338 -11233 350
rect -11279 -338 -11273 338
rect -11239 -338 -11233 338
rect -11279 -350 -11233 -338
rect -11011 338 -10965 350
rect -11011 -338 -11005 338
rect -10971 -338 -10965 338
rect -11011 -350 -10965 -338
rect -10743 338 -10697 350
rect -10743 -338 -10737 338
rect -10703 -338 -10697 338
rect -10743 -350 -10697 -338
rect -10475 338 -10429 350
rect -10475 -338 -10469 338
rect -10435 -338 -10429 338
rect -10475 -350 -10429 -338
rect -10207 338 -10161 350
rect -10207 -338 -10201 338
rect -10167 -338 -10161 338
rect -10207 -350 -10161 -338
rect -9939 338 -9893 350
rect -9939 -338 -9933 338
rect -9899 -338 -9893 338
rect -9939 -350 -9893 -338
rect -9671 338 -9625 350
rect -9671 -338 -9665 338
rect -9631 -338 -9625 338
rect -9671 -350 -9625 -338
rect -9403 338 -9357 350
rect -9403 -338 -9397 338
rect -9363 -338 -9357 338
rect -9403 -350 -9357 -338
rect -9135 338 -9089 350
rect -9135 -338 -9129 338
rect -9095 -338 -9089 338
rect -9135 -350 -9089 -338
rect -8867 338 -8821 350
rect -8867 -338 -8861 338
rect -8827 -338 -8821 338
rect -8867 -350 -8821 -338
rect -8599 338 -8553 350
rect -8599 -338 -8593 338
rect -8559 -338 -8553 338
rect -8599 -350 -8553 -338
rect -8331 338 -8285 350
rect -8331 -338 -8325 338
rect -8291 -338 -8285 338
rect -8331 -350 -8285 -338
rect -8063 338 -8017 350
rect -8063 -338 -8057 338
rect -8023 -338 -8017 338
rect -8063 -350 -8017 -338
rect -7795 338 -7749 350
rect -7795 -338 -7789 338
rect -7755 -338 -7749 338
rect -7795 -350 -7749 -338
rect -7527 338 -7481 350
rect -7527 -338 -7521 338
rect -7487 -338 -7481 338
rect -7527 -350 -7481 -338
rect -7259 338 -7213 350
rect -7259 -338 -7253 338
rect -7219 -338 -7213 338
rect -7259 -350 -7213 -338
rect -6991 338 -6945 350
rect -6991 -338 -6985 338
rect -6951 -338 -6945 338
rect -6991 -350 -6945 -338
rect -6723 338 -6677 350
rect -6723 -338 -6717 338
rect -6683 -338 -6677 338
rect -6723 -350 -6677 -338
rect -6455 338 -6409 350
rect -6455 -338 -6449 338
rect -6415 -338 -6409 338
rect -6455 -350 -6409 -338
rect -6187 338 -6141 350
rect -6187 -338 -6181 338
rect -6147 -338 -6141 338
rect -6187 -350 -6141 -338
rect -5919 338 -5873 350
rect -5919 -338 -5913 338
rect -5879 -338 -5873 338
rect -5919 -350 -5873 -338
rect -5651 338 -5605 350
rect -5651 -338 -5645 338
rect -5611 -338 -5605 338
rect -5651 -350 -5605 -338
rect -5383 338 -5337 350
rect -5383 -338 -5377 338
rect -5343 -338 -5337 338
rect -5383 -350 -5337 -338
rect -5115 338 -5069 350
rect -5115 -338 -5109 338
rect -5075 -338 -5069 338
rect -5115 -350 -5069 -338
rect -4847 338 -4801 350
rect -4847 -338 -4841 338
rect -4807 -338 -4801 338
rect -4847 -350 -4801 -338
rect -4579 338 -4533 350
rect -4579 -338 -4573 338
rect -4539 -338 -4533 338
rect -4579 -350 -4533 -338
rect -4311 338 -4265 350
rect -4311 -338 -4305 338
rect -4271 -338 -4265 338
rect -4311 -350 -4265 -338
rect -4043 338 -3997 350
rect -4043 -338 -4037 338
rect -4003 -338 -3997 338
rect -4043 -350 -3997 -338
rect -3775 338 -3729 350
rect -3775 -338 -3769 338
rect -3735 -338 -3729 338
rect -3775 -350 -3729 -338
rect -3507 338 -3461 350
rect -3507 -338 -3501 338
rect -3467 -338 -3461 338
rect -3507 -350 -3461 -338
rect -3239 338 -3193 350
rect -3239 -338 -3233 338
rect -3199 -338 -3193 338
rect -3239 -350 -3193 -338
rect -2971 338 -2925 350
rect -2971 -338 -2965 338
rect -2931 -338 -2925 338
rect -2971 -350 -2925 -338
rect -2703 338 -2657 350
rect -2703 -338 -2697 338
rect -2663 -338 -2657 338
rect -2703 -350 -2657 -338
rect -2435 338 -2389 350
rect -2435 -338 -2429 338
rect -2395 -338 -2389 338
rect -2435 -350 -2389 -338
rect -2167 338 -2121 350
rect -2167 -338 -2161 338
rect -2127 -338 -2121 338
rect -2167 -350 -2121 -338
rect -1899 338 -1853 350
rect -1899 -338 -1893 338
rect -1859 -338 -1853 338
rect -1899 -350 -1853 -338
rect -1631 338 -1585 350
rect -1631 -338 -1625 338
rect -1591 -338 -1585 338
rect -1631 -350 -1585 -338
rect -1363 338 -1317 350
rect -1363 -338 -1357 338
rect -1323 -338 -1317 338
rect -1363 -350 -1317 -338
rect -1095 338 -1049 350
rect -1095 -338 -1089 338
rect -1055 -338 -1049 338
rect -1095 -350 -1049 -338
rect -827 338 -781 350
rect -827 -338 -821 338
rect -787 -338 -781 338
rect -827 -350 -781 -338
rect -559 338 -513 350
rect -559 -338 -553 338
rect -519 -338 -513 338
rect -559 -350 -513 -338
rect -291 338 -245 350
rect -291 -338 -285 338
rect -251 -338 -245 338
rect -291 -350 -245 -338
rect -23 338 23 350
rect -23 -338 -17 338
rect 17 -338 23 338
rect -23 -350 23 -338
rect 245 338 291 350
rect 245 -338 251 338
rect 285 -338 291 338
rect 245 -350 291 -338
rect 513 338 559 350
rect 513 -338 519 338
rect 553 -338 559 338
rect 513 -350 559 -338
rect 781 338 827 350
rect 781 -338 787 338
rect 821 -338 827 338
rect 781 -350 827 -338
rect 1049 338 1095 350
rect 1049 -338 1055 338
rect 1089 -338 1095 338
rect 1049 -350 1095 -338
rect 1317 338 1363 350
rect 1317 -338 1323 338
rect 1357 -338 1363 338
rect 1317 -350 1363 -338
rect 1585 338 1631 350
rect 1585 -338 1591 338
rect 1625 -338 1631 338
rect 1585 -350 1631 -338
rect 1853 338 1899 350
rect 1853 -338 1859 338
rect 1893 -338 1899 338
rect 1853 -350 1899 -338
rect 2121 338 2167 350
rect 2121 -338 2127 338
rect 2161 -338 2167 338
rect 2121 -350 2167 -338
rect 2389 338 2435 350
rect 2389 -338 2395 338
rect 2429 -338 2435 338
rect 2389 -350 2435 -338
rect 2657 338 2703 350
rect 2657 -338 2663 338
rect 2697 -338 2703 338
rect 2657 -350 2703 -338
rect 2925 338 2971 350
rect 2925 -338 2931 338
rect 2965 -338 2971 338
rect 2925 -350 2971 -338
rect 3193 338 3239 350
rect 3193 -338 3199 338
rect 3233 -338 3239 338
rect 3193 -350 3239 -338
rect 3461 338 3507 350
rect 3461 -338 3467 338
rect 3501 -338 3507 338
rect 3461 -350 3507 -338
rect 3729 338 3775 350
rect 3729 -338 3735 338
rect 3769 -338 3775 338
rect 3729 -350 3775 -338
rect 3997 338 4043 350
rect 3997 -338 4003 338
rect 4037 -338 4043 338
rect 3997 -350 4043 -338
rect 4265 338 4311 350
rect 4265 -338 4271 338
rect 4305 -338 4311 338
rect 4265 -350 4311 -338
rect 4533 338 4579 350
rect 4533 -338 4539 338
rect 4573 -338 4579 338
rect 4533 -350 4579 -338
rect 4801 338 4847 350
rect 4801 -338 4807 338
rect 4841 -338 4847 338
rect 4801 -350 4847 -338
rect 5069 338 5115 350
rect 5069 -338 5075 338
rect 5109 -338 5115 338
rect 5069 -350 5115 -338
rect 5337 338 5383 350
rect 5337 -338 5343 338
rect 5377 -338 5383 338
rect 5337 -350 5383 -338
rect 5605 338 5651 350
rect 5605 -338 5611 338
rect 5645 -338 5651 338
rect 5605 -350 5651 -338
rect 5873 338 5919 350
rect 5873 -338 5879 338
rect 5913 -338 5919 338
rect 5873 -350 5919 -338
rect 6141 338 6187 350
rect 6141 -338 6147 338
rect 6181 -338 6187 338
rect 6141 -350 6187 -338
rect 6409 338 6455 350
rect 6409 -338 6415 338
rect 6449 -338 6455 338
rect 6409 -350 6455 -338
rect 6677 338 6723 350
rect 6677 -338 6683 338
rect 6717 -338 6723 338
rect 6677 -350 6723 -338
rect 6945 338 6991 350
rect 6945 -338 6951 338
rect 6985 -338 6991 338
rect 6945 -350 6991 -338
rect 7213 338 7259 350
rect 7213 -338 7219 338
rect 7253 -338 7259 338
rect 7213 -350 7259 -338
rect 7481 338 7527 350
rect 7481 -338 7487 338
rect 7521 -338 7527 338
rect 7481 -350 7527 -338
rect 7749 338 7795 350
rect 7749 -338 7755 338
rect 7789 -338 7795 338
rect 7749 -350 7795 -338
rect 8017 338 8063 350
rect 8017 -338 8023 338
rect 8057 -338 8063 338
rect 8017 -350 8063 -338
rect 8285 338 8331 350
rect 8285 -338 8291 338
rect 8325 -338 8331 338
rect 8285 -350 8331 -338
rect 8553 338 8599 350
rect 8553 -338 8559 338
rect 8593 -338 8599 338
rect 8553 -350 8599 -338
rect 8821 338 8867 350
rect 8821 -338 8827 338
rect 8861 -338 8867 338
rect 8821 -350 8867 -338
rect 9089 338 9135 350
rect 9089 -338 9095 338
rect 9129 -338 9135 338
rect 9089 -350 9135 -338
rect 9357 338 9403 350
rect 9357 -338 9363 338
rect 9397 -338 9403 338
rect 9357 -350 9403 -338
rect 9625 338 9671 350
rect 9625 -338 9631 338
rect 9665 -338 9671 338
rect 9625 -350 9671 -338
rect 9893 338 9939 350
rect 9893 -338 9899 338
rect 9933 -338 9939 338
rect 9893 -350 9939 -338
rect 10161 338 10207 350
rect 10161 -338 10167 338
rect 10201 -338 10207 338
rect 10161 -350 10207 -338
rect 10429 338 10475 350
rect 10429 -338 10435 338
rect 10469 -338 10475 338
rect 10429 -350 10475 -338
rect 10697 338 10743 350
rect 10697 -338 10703 338
rect 10737 -338 10743 338
rect 10697 -350 10743 -338
rect 10965 338 11011 350
rect 10965 -338 10971 338
rect 11005 -338 11011 338
rect 10965 -350 11011 -338
rect 11233 338 11279 350
rect 11233 -338 11239 338
rect 11273 -338 11279 338
rect 11233 -350 11279 -338
rect 11501 338 11547 350
rect 11501 -338 11507 338
rect 11541 -338 11547 338
rect 11501 -350 11547 -338
rect 11769 338 11815 350
rect 11769 -338 11775 338
rect 11809 -338 11815 338
rect 11769 -350 11815 -338
rect 12037 338 12083 350
rect 12037 -338 12043 338
rect 12077 -338 12083 338
rect 12037 -350 12083 -338
rect 12305 338 12351 350
rect 12305 -338 12311 338
rect 12345 -338 12351 338
rect 12305 -350 12351 -338
rect 12573 338 12619 350
rect 12573 -338 12579 338
rect 12613 -338 12619 338
rect 12573 -350 12619 -338
rect 12841 338 12887 350
rect 12841 -338 12847 338
rect 12881 -338 12887 338
rect 12841 -350 12887 -338
rect 13109 338 13155 350
rect 13109 -338 13115 338
rect 13149 -338 13155 338
rect 13109 -350 13155 -338
rect 13377 338 13423 350
rect 13377 -338 13383 338
rect 13417 -338 13423 338
rect 13377 -350 13423 -338
rect -13367 -397 -13165 -391
rect -13367 -431 -13355 -397
rect -13177 -431 -13165 -397
rect -13367 -437 -13165 -431
rect -13099 -397 -12897 -391
rect -13099 -431 -13087 -397
rect -12909 -431 -12897 -397
rect -13099 -437 -12897 -431
rect -12831 -397 -12629 -391
rect -12831 -431 -12819 -397
rect -12641 -431 -12629 -397
rect -12831 -437 -12629 -431
rect -12563 -397 -12361 -391
rect -12563 -431 -12551 -397
rect -12373 -431 -12361 -397
rect -12563 -437 -12361 -431
rect -12295 -397 -12093 -391
rect -12295 -431 -12283 -397
rect -12105 -431 -12093 -397
rect -12295 -437 -12093 -431
rect -12027 -397 -11825 -391
rect -12027 -431 -12015 -397
rect -11837 -431 -11825 -397
rect -12027 -437 -11825 -431
rect -11759 -397 -11557 -391
rect -11759 -431 -11747 -397
rect -11569 -431 -11557 -397
rect -11759 -437 -11557 -431
rect -11491 -397 -11289 -391
rect -11491 -431 -11479 -397
rect -11301 -431 -11289 -397
rect -11491 -437 -11289 -431
rect -11223 -397 -11021 -391
rect -11223 -431 -11211 -397
rect -11033 -431 -11021 -397
rect -11223 -437 -11021 -431
rect -10955 -397 -10753 -391
rect -10955 -431 -10943 -397
rect -10765 -431 -10753 -397
rect -10955 -437 -10753 -431
rect -10687 -397 -10485 -391
rect -10687 -431 -10675 -397
rect -10497 -431 -10485 -397
rect -10687 -437 -10485 -431
rect -10419 -397 -10217 -391
rect -10419 -431 -10407 -397
rect -10229 -431 -10217 -397
rect -10419 -437 -10217 -431
rect -10151 -397 -9949 -391
rect -10151 -431 -10139 -397
rect -9961 -431 -9949 -397
rect -10151 -437 -9949 -431
rect -9883 -397 -9681 -391
rect -9883 -431 -9871 -397
rect -9693 -431 -9681 -397
rect -9883 -437 -9681 -431
rect -9615 -397 -9413 -391
rect -9615 -431 -9603 -397
rect -9425 -431 -9413 -397
rect -9615 -437 -9413 -431
rect -9347 -397 -9145 -391
rect -9347 -431 -9335 -397
rect -9157 -431 -9145 -397
rect -9347 -437 -9145 -431
rect -9079 -397 -8877 -391
rect -9079 -431 -9067 -397
rect -8889 -431 -8877 -397
rect -9079 -437 -8877 -431
rect -8811 -397 -8609 -391
rect -8811 -431 -8799 -397
rect -8621 -431 -8609 -397
rect -8811 -437 -8609 -431
rect -8543 -397 -8341 -391
rect -8543 -431 -8531 -397
rect -8353 -431 -8341 -397
rect -8543 -437 -8341 -431
rect -8275 -397 -8073 -391
rect -8275 -431 -8263 -397
rect -8085 -431 -8073 -397
rect -8275 -437 -8073 -431
rect -8007 -397 -7805 -391
rect -8007 -431 -7995 -397
rect -7817 -431 -7805 -397
rect -8007 -437 -7805 -431
rect -7739 -397 -7537 -391
rect -7739 -431 -7727 -397
rect -7549 -431 -7537 -397
rect -7739 -437 -7537 -431
rect -7471 -397 -7269 -391
rect -7471 -431 -7459 -397
rect -7281 -431 -7269 -397
rect -7471 -437 -7269 -431
rect -7203 -397 -7001 -391
rect -7203 -431 -7191 -397
rect -7013 -431 -7001 -397
rect -7203 -437 -7001 -431
rect -6935 -397 -6733 -391
rect -6935 -431 -6923 -397
rect -6745 -431 -6733 -397
rect -6935 -437 -6733 -431
rect -6667 -397 -6465 -391
rect -6667 -431 -6655 -397
rect -6477 -431 -6465 -397
rect -6667 -437 -6465 -431
rect -6399 -397 -6197 -391
rect -6399 -431 -6387 -397
rect -6209 -431 -6197 -397
rect -6399 -437 -6197 -431
rect -6131 -397 -5929 -391
rect -6131 -431 -6119 -397
rect -5941 -431 -5929 -397
rect -6131 -437 -5929 -431
rect -5863 -397 -5661 -391
rect -5863 -431 -5851 -397
rect -5673 -431 -5661 -397
rect -5863 -437 -5661 -431
rect -5595 -397 -5393 -391
rect -5595 -431 -5583 -397
rect -5405 -431 -5393 -397
rect -5595 -437 -5393 -431
rect -5327 -397 -5125 -391
rect -5327 -431 -5315 -397
rect -5137 -431 -5125 -397
rect -5327 -437 -5125 -431
rect -5059 -397 -4857 -391
rect -5059 -431 -5047 -397
rect -4869 -431 -4857 -397
rect -5059 -437 -4857 -431
rect -4791 -397 -4589 -391
rect -4791 -431 -4779 -397
rect -4601 -431 -4589 -397
rect -4791 -437 -4589 -431
rect -4523 -397 -4321 -391
rect -4523 -431 -4511 -397
rect -4333 -431 -4321 -397
rect -4523 -437 -4321 -431
rect -4255 -397 -4053 -391
rect -4255 -431 -4243 -397
rect -4065 -431 -4053 -397
rect -4255 -437 -4053 -431
rect -3987 -397 -3785 -391
rect -3987 -431 -3975 -397
rect -3797 -431 -3785 -397
rect -3987 -437 -3785 -431
rect -3719 -397 -3517 -391
rect -3719 -431 -3707 -397
rect -3529 -431 -3517 -397
rect -3719 -437 -3517 -431
rect -3451 -397 -3249 -391
rect -3451 -431 -3439 -397
rect -3261 -431 -3249 -397
rect -3451 -437 -3249 -431
rect -3183 -397 -2981 -391
rect -3183 -431 -3171 -397
rect -2993 -431 -2981 -397
rect -3183 -437 -2981 -431
rect -2915 -397 -2713 -391
rect -2915 -431 -2903 -397
rect -2725 -431 -2713 -397
rect -2915 -437 -2713 -431
rect -2647 -397 -2445 -391
rect -2647 -431 -2635 -397
rect -2457 -431 -2445 -397
rect -2647 -437 -2445 -431
rect -2379 -397 -2177 -391
rect -2379 -431 -2367 -397
rect -2189 -431 -2177 -397
rect -2379 -437 -2177 -431
rect -2111 -397 -1909 -391
rect -2111 -431 -2099 -397
rect -1921 -431 -1909 -397
rect -2111 -437 -1909 -431
rect -1843 -397 -1641 -391
rect -1843 -431 -1831 -397
rect -1653 -431 -1641 -397
rect -1843 -437 -1641 -431
rect -1575 -397 -1373 -391
rect -1575 -431 -1563 -397
rect -1385 -431 -1373 -397
rect -1575 -437 -1373 -431
rect -1307 -397 -1105 -391
rect -1307 -431 -1295 -397
rect -1117 -431 -1105 -397
rect -1307 -437 -1105 -431
rect -1039 -397 -837 -391
rect -1039 -431 -1027 -397
rect -849 -431 -837 -397
rect -1039 -437 -837 -431
rect -771 -397 -569 -391
rect -771 -431 -759 -397
rect -581 -431 -569 -397
rect -771 -437 -569 -431
rect -503 -397 -301 -391
rect -503 -431 -491 -397
rect -313 -431 -301 -397
rect -503 -437 -301 -431
rect -235 -397 -33 -391
rect -235 -431 -223 -397
rect -45 -431 -33 -397
rect -235 -437 -33 -431
rect 33 -397 235 -391
rect 33 -431 45 -397
rect 223 -431 235 -397
rect 33 -437 235 -431
rect 301 -397 503 -391
rect 301 -431 313 -397
rect 491 -431 503 -397
rect 301 -437 503 -431
rect 569 -397 771 -391
rect 569 -431 581 -397
rect 759 -431 771 -397
rect 569 -437 771 -431
rect 837 -397 1039 -391
rect 837 -431 849 -397
rect 1027 -431 1039 -397
rect 837 -437 1039 -431
rect 1105 -397 1307 -391
rect 1105 -431 1117 -397
rect 1295 -431 1307 -397
rect 1105 -437 1307 -431
rect 1373 -397 1575 -391
rect 1373 -431 1385 -397
rect 1563 -431 1575 -397
rect 1373 -437 1575 -431
rect 1641 -397 1843 -391
rect 1641 -431 1653 -397
rect 1831 -431 1843 -397
rect 1641 -437 1843 -431
rect 1909 -397 2111 -391
rect 1909 -431 1921 -397
rect 2099 -431 2111 -397
rect 1909 -437 2111 -431
rect 2177 -397 2379 -391
rect 2177 -431 2189 -397
rect 2367 -431 2379 -397
rect 2177 -437 2379 -431
rect 2445 -397 2647 -391
rect 2445 -431 2457 -397
rect 2635 -431 2647 -397
rect 2445 -437 2647 -431
rect 2713 -397 2915 -391
rect 2713 -431 2725 -397
rect 2903 -431 2915 -397
rect 2713 -437 2915 -431
rect 2981 -397 3183 -391
rect 2981 -431 2993 -397
rect 3171 -431 3183 -397
rect 2981 -437 3183 -431
rect 3249 -397 3451 -391
rect 3249 -431 3261 -397
rect 3439 -431 3451 -397
rect 3249 -437 3451 -431
rect 3517 -397 3719 -391
rect 3517 -431 3529 -397
rect 3707 -431 3719 -397
rect 3517 -437 3719 -431
rect 3785 -397 3987 -391
rect 3785 -431 3797 -397
rect 3975 -431 3987 -397
rect 3785 -437 3987 -431
rect 4053 -397 4255 -391
rect 4053 -431 4065 -397
rect 4243 -431 4255 -397
rect 4053 -437 4255 -431
rect 4321 -397 4523 -391
rect 4321 -431 4333 -397
rect 4511 -431 4523 -397
rect 4321 -437 4523 -431
rect 4589 -397 4791 -391
rect 4589 -431 4601 -397
rect 4779 -431 4791 -397
rect 4589 -437 4791 -431
rect 4857 -397 5059 -391
rect 4857 -431 4869 -397
rect 5047 -431 5059 -397
rect 4857 -437 5059 -431
rect 5125 -397 5327 -391
rect 5125 -431 5137 -397
rect 5315 -431 5327 -397
rect 5125 -437 5327 -431
rect 5393 -397 5595 -391
rect 5393 -431 5405 -397
rect 5583 -431 5595 -397
rect 5393 -437 5595 -431
rect 5661 -397 5863 -391
rect 5661 -431 5673 -397
rect 5851 -431 5863 -397
rect 5661 -437 5863 -431
rect 5929 -397 6131 -391
rect 5929 -431 5941 -397
rect 6119 -431 6131 -397
rect 5929 -437 6131 -431
rect 6197 -397 6399 -391
rect 6197 -431 6209 -397
rect 6387 -431 6399 -397
rect 6197 -437 6399 -431
rect 6465 -397 6667 -391
rect 6465 -431 6477 -397
rect 6655 -431 6667 -397
rect 6465 -437 6667 -431
rect 6733 -397 6935 -391
rect 6733 -431 6745 -397
rect 6923 -431 6935 -397
rect 6733 -437 6935 -431
rect 7001 -397 7203 -391
rect 7001 -431 7013 -397
rect 7191 -431 7203 -397
rect 7001 -437 7203 -431
rect 7269 -397 7471 -391
rect 7269 -431 7281 -397
rect 7459 -431 7471 -397
rect 7269 -437 7471 -431
rect 7537 -397 7739 -391
rect 7537 -431 7549 -397
rect 7727 -431 7739 -397
rect 7537 -437 7739 -431
rect 7805 -397 8007 -391
rect 7805 -431 7817 -397
rect 7995 -431 8007 -397
rect 7805 -437 8007 -431
rect 8073 -397 8275 -391
rect 8073 -431 8085 -397
rect 8263 -431 8275 -397
rect 8073 -437 8275 -431
rect 8341 -397 8543 -391
rect 8341 -431 8353 -397
rect 8531 -431 8543 -397
rect 8341 -437 8543 -431
rect 8609 -397 8811 -391
rect 8609 -431 8621 -397
rect 8799 -431 8811 -397
rect 8609 -437 8811 -431
rect 8877 -397 9079 -391
rect 8877 -431 8889 -397
rect 9067 -431 9079 -397
rect 8877 -437 9079 -431
rect 9145 -397 9347 -391
rect 9145 -431 9157 -397
rect 9335 -431 9347 -397
rect 9145 -437 9347 -431
rect 9413 -397 9615 -391
rect 9413 -431 9425 -397
rect 9603 -431 9615 -397
rect 9413 -437 9615 -431
rect 9681 -397 9883 -391
rect 9681 -431 9693 -397
rect 9871 -431 9883 -397
rect 9681 -437 9883 -431
rect 9949 -397 10151 -391
rect 9949 -431 9961 -397
rect 10139 -431 10151 -397
rect 9949 -437 10151 -431
rect 10217 -397 10419 -391
rect 10217 -431 10229 -397
rect 10407 -431 10419 -397
rect 10217 -437 10419 -431
rect 10485 -397 10687 -391
rect 10485 -431 10497 -397
rect 10675 -431 10687 -397
rect 10485 -437 10687 -431
rect 10753 -397 10955 -391
rect 10753 -431 10765 -397
rect 10943 -431 10955 -397
rect 10753 -437 10955 -431
rect 11021 -397 11223 -391
rect 11021 -431 11033 -397
rect 11211 -431 11223 -397
rect 11021 -437 11223 -431
rect 11289 -397 11491 -391
rect 11289 -431 11301 -397
rect 11479 -431 11491 -397
rect 11289 -437 11491 -431
rect 11557 -397 11759 -391
rect 11557 -431 11569 -397
rect 11747 -431 11759 -397
rect 11557 -437 11759 -431
rect 11825 -397 12027 -391
rect 11825 -431 11837 -397
rect 12015 -431 12027 -397
rect 11825 -437 12027 -431
rect 12093 -397 12295 -391
rect 12093 -431 12105 -397
rect 12283 -431 12295 -397
rect 12093 -437 12295 -431
rect 12361 -397 12563 -391
rect 12361 -431 12373 -397
rect 12551 -431 12563 -397
rect 12361 -437 12563 -431
rect 12629 -397 12831 -391
rect 12629 -431 12641 -397
rect 12819 -431 12831 -397
rect 12629 -437 12831 -431
rect 12897 -397 13099 -391
rect 12897 -431 12909 -397
rect 13087 -431 13099 -397
rect 12897 -437 13099 -431
rect 13165 -397 13367 -391
rect 13165 -431 13177 -397
rect 13355 -431 13367 -397
rect 13165 -437 13367 -431
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -13514 -516 13514 516
string parameters w 3.5 l 1.05 m 1 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
