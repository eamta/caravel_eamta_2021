magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect -1044 1639 -844 1652
rect -1044 1618 -819 1639
rect -701 1605 -648 1606
rect -1034 1584 -648 1605
rect -844 1582 -648 1584
rect -855 1577 -648 1582
rect -855 1571 -803 1577
rect -719 1571 -648 1577
rect -718 1570 -648 1571
rect -631 1570 -349 1577
rect -701 1566 -315 1570
rect -701 1563 -349 1566
rect -1034 1419 -1000 1563
rect -718 1553 -349 1563
rect -718 1535 -315 1553
rect -926 1509 -914 1513
rect -718 1509 -279 1535
rect -926 1503 -902 1509
rect -888 1503 -880 1509
rect -926 1491 -908 1503
rect -926 1457 -914 1491
rect -907 1459 -902 1503
rect -892 1469 -880 1503
rect -876 1469 -830 1503
rect -880 1459 -814 1469
rect -908 1457 -814 1459
rect -948 1449 -914 1457
rect -907 1449 -902 1457
rect -948 1431 -886 1449
rect -880 1441 -814 1457
rect -832 1431 -798 1435
rect -914 1426 -874 1431
rect -844 1426 -792 1431
rect -914 1419 -880 1426
rect -1001 1267 -1000 1419
rect -920 1413 -880 1419
rect -838 1413 -792 1426
rect -920 1393 -886 1413
rect -832 1407 -798 1413
rect -836 1334 -786 1372
rect -818 1284 -786 1334
rect -768 1300 -764 1334
rect -718 1330 -631 1509
rect -630 1502 -596 1509
rect -542 1502 -508 1509
rect -454 1506 -420 1509
rect -473 1502 -420 1506
rect -366 1502 -279 1509
rect -630 1330 -597 1502
rect -542 1484 -508 1497
rect -542 1468 -496 1484
rect -473 1474 -423 1502
rect -350 1499 -279 1502
rect 80 1500 108 1553
rect 2440 1549 2475 1583
rect 37 1499 459 1500
rect -488 1468 -423 1474
rect -542 1434 -423 1468
rect -542 1418 -496 1434
rect -488 1428 -423 1434
rect -466 1418 -423 1428
rect -542 1409 -508 1418
rect -505 1409 -496 1418
rect -460 1409 -423 1418
rect -349 1465 -261 1499
rect -166 1465 -20 1499
rect 19 1465 459 1499
rect 2071 1496 2106 1530
rect 1298 1475 1386 1478
rect -542 1387 -483 1409
rect -460 1400 -395 1409
rect -454 1387 -395 1400
rect -563 1341 -395 1387
rect -563 1330 -417 1341
rect -349 1330 -262 1465
rect -154 1435 -120 1465
rect 20 1464 459 1465
rect -166 1431 -78 1435
rect -166 1419 -54 1431
rect 20 1419 34 1464
rect 37 1447 459 1464
rect 466 1447 506 1465
rect 1279 1463 1386 1475
rect -154 1415 -120 1419
rect -66 1415 -54 1419
rect -120 1397 -92 1403
rect -154 1381 -88 1397
rect 37 1376 828 1447
rect 1702 1443 1737 1477
rect 1333 1407 1339 1424
rect 20 1363 828 1376
rect 9 1354 828 1363
rect 928 1379 1350 1407
rect 928 1354 1367 1379
rect -718 1329 -262 1330
rect -801 1269 -786 1284
rect -718 1291 -631 1329
rect -630 1325 -597 1329
rect -563 1303 -554 1329
rect -718 1284 -642 1291
rect -563 1288 -548 1303
rect -718 1273 -707 1284
rect -1034 1261 -1023 1267
rect -1011 1261 -1000 1267
rect -701 1261 -631 1284
rect -1070 1186 -631 1261
rect -563 1261 -548 1276
rect -563 1231 -505 1261
rect -475 1231 -466 1329
rect -423 1288 -417 1329
rect -349 1261 -262 1329
rect -128 1261 -120 1353
rect 9 1341 1367 1354
rect 1373 1341 1401 1345
rect 1433 1341 1441 1348
rect -106 1310 -63 1325
rect -106 1261 -78 1310
rect 6 1295 111 1341
rect 6 1261 107 1295
rect 191 1294 214 1341
rect 219 1328 242 1341
rect 219 1322 277 1328
rect -563 1222 -554 1231
rect -563 1207 -539 1222
rect -457 1207 -417 1213
rect -349 1212 107 1261
rect 175 1212 183 1281
rect 192 1212 221 1285
rect 307 1277 315 1281
rect 307 1269 321 1277
rect 288 1265 321 1269
rect 335 1265 343 1309
rect 389 1265 423 1341
rect 442 1265 476 1341
rect 651 1318 692 1341
rect 760 1318 792 1341
rect 964 1337 999 1341
rect 595 1304 902 1318
rect 595 1299 911 1304
rect 584 1286 911 1299
rect 930 1286 945 1318
rect 964 1286 998 1337
rect 1117 1288 1196 1303
rect 584 1284 1197 1286
rect 584 1275 650 1284
rect 595 1273 629 1275
rect 595 1269 660 1273
rect 672 1269 692 1284
rect 714 1269 748 1273
rect 758 1269 1197 1284
rect -1070 1179 -642 1186
rect -638 1179 -631 1186
rect -1070 1106 -631 1179
rect -565 1176 -554 1207
rect -349 1178 111 1212
rect 127 1201 221 1212
rect 138 1189 168 1201
rect 175 1189 221 1201
rect 127 1178 221 1189
rect -523 1159 -512 1176
rect -488 1160 -461 1166
rect -507 1159 -416 1160
rect -349 1159 107 1178
rect -630 1106 -597 1145
rect -523 1141 107 1159
rect -538 1129 107 1141
rect 173 1168 221 1178
rect 226 1231 321 1265
rect 322 1231 480 1265
rect 226 1168 260 1231
rect 275 1168 294 1231
rect 307 1183 315 1231
rect 306 1168 321 1183
rect 173 1129 260 1168
rect 263 1134 321 1168
rect -542 1125 107 1129
rect -542 1120 -433 1125
rect -542 1106 -478 1120
rect -466 1110 -433 1120
rect -1070 1088 -478 1106
rect -460 1092 -433 1110
rect -349 1104 107 1125
rect -379 1095 107 1104
rect 146 1113 260 1129
rect 275 1113 321 1134
rect 146 1097 221 1113
rect 146 1095 214 1097
rect 226 1095 260 1113
rect 274 1101 321 1113
rect 275 1097 294 1101
rect 306 1097 309 1101
rect -1070 1072 -531 1088
rect -1070 1058 -631 1072
rect -630 1058 -596 1072
rect -565 1058 -531 1072
rect -512 1058 -478 1088
rect -454 1088 -435 1092
rect -379 1091 141 1095
rect -454 1058 -444 1088
rect -388 1058 141 1091
rect -1070 1041 141 1058
rect -915 957 -914 1041
rect -906 961 -902 1041
rect -881 1018 -847 1041
rect -718 1038 -672 1041
rect -665 1038 141 1041
rect -718 1035 141 1038
rect -730 1024 141 1035
rect -730 1020 -655 1024
rect -881 1010 -848 1018
rect -881 852 -847 1010
rect -730 977 -642 1020
rect -599 977 -596 1024
rect -730 973 -596 977
rect -730 961 -584 973
rect -565 961 -531 1024
rect -718 957 -684 961
rect -672 954 -642 961
rect -630 957 -611 961
rect -599 957 -596 961
rect -752 923 -733 927
rect -746 911 -727 923
rect -767 908 -727 911
rect -969 818 -847 852
rect -779 893 -727 908
rect -779 863 -721 893
rect -779 858 -727 863
rect -718 858 -699 951
rect -672 935 -649 954
rect -679 923 -645 927
rect -687 920 -633 923
rect -658 911 -639 920
rect -679 908 -639 911
rect -679 893 -633 908
rect -630 899 -611 951
rect -691 885 -633 893
rect -691 863 -631 885
rect -779 851 -733 858
rect -679 851 -631 863
rect -565 852 -554 961
rect -779 848 -622 851
rect -881 771 -847 818
rect -767 817 -622 848
rect -767 773 -733 817
rect -911 737 -847 771
rect -789 755 -733 773
rect -679 755 -645 817
rect -565 775 -554 786
rect -789 753 -767 755
rect -770 737 -743 743
rect -673 739 -645 755
rect -633 753 -621 773
rect -565 771 -563 775
rect -546 771 -531 957
rect -585 753 -531 771
rect -639 737 -611 753
rect -585 737 -517 753
rect -512 749 -478 1024
rect -454 957 -444 1024
rect -370 1017 141 1024
rect -370 1014 107 1017
rect 126 1014 141 1017
rect 173 1015 260 1095
rect 335 1082 343 1231
rect 389 1201 423 1231
rect 344 1163 368 1197
rect 382 1169 423 1201
rect 372 1163 423 1169
rect 344 1133 423 1163
rect 442 1201 476 1231
rect 442 1133 484 1201
rect 344 1129 434 1133
rect 344 1095 368 1129
rect 372 1123 423 1129
rect 389 1108 423 1123
rect 442 1108 468 1133
rect 389 1086 476 1108
rect 334 1074 343 1082
rect 371 1074 476 1086
rect 372 1070 510 1074
rect 265 1020 294 1054
rect -432 1004 -420 1014
rect -370 1007 126 1014
rect -432 1002 -414 1004
rect -352 1002 126 1007
rect -436 973 -414 1002
rect -366 991 126 1002
rect -398 980 126 991
rect -398 976 -386 980
rect -404 975 -386 976
rect -432 961 -414 973
rect -408 964 -378 975
rect -366 973 126 980
rect -352 964 126 973
rect -404 961 -364 964
rect -432 899 -420 961
rect -408 935 -364 961
rect -344 952 126 964
rect 173 1004 281 1015
rect 340 1004 476 1070
rect 173 952 260 1004
rect 279 973 313 986
rect 328 973 476 1004
rect 263 961 476 973
rect 494 961 510 1070
rect 522 1020 536 1256
rect 550 1241 576 1265
rect 561 1232 576 1241
rect 595 1259 672 1269
rect 702 1259 1197 1269
rect 595 1257 665 1259
rect 595 1256 660 1257
rect 561 1228 590 1232
rect 544 1203 590 1228
rect 595 1216 663 1256
rect 672 1216 678 1227
rect 595 1203 678 1216
rect 544 1163 678 1203
rect 680 1163 684 1228
rect 544 1140 684 1163
rect 542 1060 684 1140
rect 708 1135 712 1256
rect 698 1123 702 1134
rect 703 1123 712 1135
rect 714 1232 748 1259
rect 758 1232 1197 1259
rect 714 1166 1197 1232
rect 714 1123 748 1166
rect 542 1044 590 1060
rect 542 1035 576 1044
rect 595 1035 663 1060
rect 675 1048 684 1060
rect 675 1044 678 1048
rect 542 1001 668 1035
rect 703 1020 748 1123
rect 263 957 494 961
rect 263 952 298 957
rect 302 953 494 957
rect 302 952 506 953
rect -344 935 506 952
rect -404 923 -386 935
rect -404 908 -392 923
rect -410 893 -392 908
rect -410 863 -352 893
rect -410 848 -395 863
rect -344 858 -332 935
rect -316 893 -276 935
rect -271 934 -238 935
rect -271 918 -242 934
rect -230 918 -205 935
rect -271 893 -264 918
rect -322 863 -264 893
rect -316 858 -304 863
rect -279 848 -264 863
rect -196 863 -162 935
rect -196 852 -185 863
rect -366 749 -308 755
rect -512 737 -483 749
rect -881 594 -843 737
rect -789 722 -743 737
rect -795 717 -743 722
rect -823 628 -817 694
rect -795 628 -789 717
rect -773 631 -743 717
rect -735 696 -677 702
rect -739 662 -696 696
rect -651 662 -642 737
rect -639 717 -607 737
rect -639 705 -611 717
rect -735 656 -677 662
rect -565 656 -483 737
rect -366 715 -354 749
rect -366 709 -308 715
rect -773 628 -749 631
rect -823 615 -789 628
rect -761 624 -755 628
rect -823 594 -755 615
rect -639 594 -593 628
rect -565 594 -517 656
rect -512 613 -483 656
rect -177 632 -162 863
rect -143 700 -109 935
rect -29 923 2 935
rect 47 927 506 935
rect 47 918 105 927
rect 127 918 506 927
rect 47 861 93 918
rect 47 849 79 861
rect -25 811 89 836
rect 3 783 61 808
rect 3 768 15 783
rect 3 762 61 768
rect 64 756 65 768
rect 173 762 207 918
rect 106 752 107 756
rect 173 755 184 762
rect 192 755 207 762
rect 173 725 207 755
rect 173 714 184 725
rect -143 666 -108 700
rect 23 689 75 700
rect 95 689 147 700
rect 34 677 64 689
rect 106 677 136 689
rect 192 685 207 725
rect 226 753 260 918
rect 263 907 294 918
rect 306 907 329 918
rect 340 914 374 918
rect 340 907 363 914
rect 328 905 363 907
rect 394 906 412 918
rect 418 917 506 918
rect 416 906 506 917
rect 328 902 368 905
rect 394 902 406 906
rect 416 902 494 906
rect 340 898 363 902
rect 418 899 476 902
rect 542 899 576 1001
rect 584 967 668 1001
rect 709 967 748 1020
rect 595 953 663 967
rect 714 955 748 967
rect 755 1161 1197 1166
rect 1297 1254 1466 1341
rect 1475 1328 1483 1338
rect 1475 1322 1537 1328
rect 1475 1288 1491 1322
rect 1475 1282 1537 1288
rect 1475 1278 1483 1282
rect 1297 1245 1473 1254
rect 755 1107 1212 1161
rect 1297 1129 1466 1245
rect 755 955 1197 1107
rect 1240 1008 1266 1107
rect 1280 973 1466 1129
rect 1479 1032 1537 1038
rect 1479 998 1491 1032
rect 1479 992 1537 998
rect 706 953 1197 955
rect 595 909 672 953
rect 702 909 1197 953
rect 1252 939 1466 973
rect 1280 927 1466 939
rect 595 905 660 909
rect 714 908 1197 909
rect 714 905 744 908
rect 595 899 629 905
rect 737 899 744 905
rect 753 899 1197 908
rect 418 880 1197 899
rect 442 865 1197 880
rect 364 851 434 855
rect 542 852 576 865
rect 310 821 434 851
rect 469 831 576 852
rect 310 817 337 821
rect 357 817 434 821
rect 377 805 434 817
rect 339 753 480 785
rect 542 753 576 831
rect 595 806 629 865
rect 775 859 1197 865
rect 1297 860 1466 927
rect 1668 915 1683 1424
rect 1702 983 1736 1443
rect 1848 1375 1906 1381
rect 1848 1341 1860 1375
rect 1848 1335 1906 1341
rect 1848 1085 1906 1091
rect 1848 1051 1860 1085
rect 2037 1058 2052 1477
rect 2071 1126 2105 1496
rect 2217 1428 2275 1434
rect 2217 1394 2229 1428
rect 2217 1388 2275 1394
rect 2217 1228 2275 1234
rect 2217 1194 2229 1228
rect 2217 1188 2275 1194
rect 2071 1092 2106 1126
rect 2406 1111 2421 1530
rect 2440 1179 2474 1549
rect 2586 1481 2644 1487
rect 2586 1447 2598 1481
rect 2586 1441 2644 1447
rect 2586 1281 2644 1287
rect 2586 1247 2598 1281
rect 2586 1241 2644 1247
rect 2440 1145 2475 1179
rect 2775 1145 2790 1583
rect 2809 1145 2837 1636
rect 2809 1111 2824 1145
rect 1848 1045 1906 1051
rect 1702 949 1737 983
rect 713 853 1218 859
rect 639 852 1218 853
rect 639 840 1197 852
rect 1201 851 1218 852
rect 639 819 722 840
rect 595 797 756 806
rect 775 797 1197 840
rect 1235 825 1252 851
rect 1210 817 1215 825
rect 595 776 1197 797
rect 595 772 871 776
rect 888 772 945 776
rect 226 742 310 753
rect 339 751 507 753
rect 226 725 299 742
rect 226 719 322 725
rect 339 719 514 751
rect 561 738 576 753
rect 655 738 689 747
rect 743 738 777 747
rect 831 736 871 772
rect 942 747 945 763
rect 954 738 979 767
rect 846 730 1085 736
rect 871 725 1085 730
rect 23 666 75 677
rect 95 666 147 677
rect -881 569 -743 594
rect -651 579 -517 594
rect -651 569 -531 579
rect 6 577 128 630
rect -881 560 -790 569
rect -604 560 -552 569
rect -823 541 -817 560
rect -877 315 -789 322
rect -905 287 -817 294
rect -823 94 -817 287
rect -795 107 -789 287
<< pwell >>
rect -1083 329 6 356
rect -469 6 6 329
<< metal1 >>
rect -517 1612 -220 1658
rect -32 1612 23 1659
rect 1462 1393 1471 1427
rect 99 1278 100 1349
rect -1059 1197 -1049 1249
rect -997 1197 -987 1249
rect -1084 811 -170 858
rect -98 852 1467 858
rect -98 818 322 852
rect 561 818 906 852
rect 1370 818 1467 852
rect -98 811 1467 818
rect -762 454 -752 506
rect -700 454 -690 506
rect -37 391 -27 443
rect 25 425 35 443
rect 25 392 64 425
rect 25 391 63 392
rect -1029 337 -1019 389
rect -967 337 -957 389
rect -551 356 -477 387
rect -469 13 5 58
rect 1103 52 1496 58
rect 1103 18 1115 52
rect 1484 18 1496 52
rect 1103 12 1496 18
<< via1 >>
rect -1049 1197 -997 1249
rect -752 454 -700 506
rect -27 391 25 443
rect -1019 337 -967 389
<< metal2 >>
rect -1040 1553 1423 1587
rect -1040 1259 -1006 1553
rect -1049 1249 -997 1259
rect -1049 1187 -997 1197
rect -1040 399 -1006 1187
rect -768 506 -700 516
rect -768 464 -752 506
rect -255 498 -221 968
rect -700 464 -221 498
rect -752 444 -700 454
rect -17 453 17 1314
rect 1389 1295 1423 1553
rect -27 443 25 453
rect -1040 389 -967 399
rect -1040 345 -1019 389
rect -27 381 25 391
rect -1019 327 -967 337
rect 31 182 32 216
use xor_lede  xor_lede_0
timestamp 1624053917
transform 1 0 -864 0 -1 1689
box -220 -2000 4428 1165
use and_lede  and_lede_0
timestamp 1624053917
transform 1 0 -1017 0 1 494
box -67 -2000 2214 1147
use ffd  ffd_0
timestamp 1624053917
transform 1 0 -1403 0 1 -1111
box 1310 1103 2980 2788
<< labels >>
rlabel metal2 1389 1295 1423 1587 1 Dn
rlabel space 1246 1393 1466 1427 1 Dnb
rlabel metal2 -700 464 -221 498 1 CE
rlabel metal1 -480 356 -477 387 1 Sout
rlabel metal1 1470 1393 1471 1427 1 Dnb
rlabel metal2 31 182 32 216 1 CLR
rlabel metal1 99 1278 100 1349 1 CLK
<< end >>
