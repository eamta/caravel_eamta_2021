magic
tech sky130A
magscale 1 2
timestamp 1616030774
<< nwell >>
rect -1784 -5513 34024 3239
<< pmos >>
rect 11495 740 11635 2140
rect 11693 740 11833 2140
rect 11891 740 12031 2140
rect 12089 740 12229 2140
rect 12287 740 12427 2140
rect 12485 740 12625 2140
rect 12683 740 12823 2140
rect 12881 740 13021 2140
rect 13079 740 13219 2140
rect 13277 740 13417 2140
rect 13475 740 13615 2140
rect 13673 740 13813 2140
rect 13871 740 14011 2140
rect 14069 740 14209 2140
rect 14267 740 14407 2140
rect 14465 740 14605 2140
rect 14663 740 14803 2140
rect 14861 740 15001 2140
rect 15059 740 15199 2140
rect 15257 740 15397 2140
rect 15455 740 15595 2140
rect 15653 740 15793 2140
rect 15851 740 15991 2140
rect 16049 740 16189 2140
rect 16247 740 16387 2140
rect 16445 740 16585 2140
rect 16643 740 16783 2140
rect 16841 740 16981 2140
rect 17039 740 17179 2140
rect 17237 740 17377 2140
rect 17435 740 17575 2140
rect 17633 740 17773 2140
rect 17831 740 17971 2140
rect 18029 740 18169 2140
rect 18227 740 18367 2140
rect 18425 740 18565 2140
rect 18623 740 18763 2140
rect 18821 740 18961 2140
rect 19019 740 19159 2140
rect 19217 740 19357 2140
rect 19415 740 19555 2140
rect 19613 740 19753 2140
rect 11495 -896 11635 504
rect 11693 -896 11833 504
rect 11891 -896 12031 504
rect 12089 -896 12229 504
rect 12287 -896 12427 504
rect 12485 -896 12625 504
rect 12683 -896 12823 504
rect 12881 -896 13021 504
rect 13079 -896 13219 504
rect 13277 -896 13417 504
rect 13475 -896 13615 504
rect 13673 -896 13813 504
rect 13871 -896 14011 504
rect 14069 -896 14209 504
rect 14267 -896 14407 504
rect 14465 -896 14605 504
rect 14663 -896 14803 504
rect 14861 -896 15001 504
rect 15059 -896 15199 504
rect 15257 -896 15397 504
rect 15455 -896 15595 504
rect 15653 -896 15793 504
rect 15851 -896 15991 504
rect 16049 -896 16189 504
rect 16247 -896 16387 504
rect 16445 -896 16585 504
rect 16643 -896 16783 504
rect 16841 -896 16981 504
rect 17039 -896 17179 504
rect 17237 -896 17377 504
rect 17435 -896 17575 504
rect 17633 -896 17773 504
rect 17831 -896 17971 504
rect 18029 -896 18169 504
rect 18227 -896 18367 504
rect 18425 -896 18565 504
rect 18623 -896 18763 504
rect 18821 -896 18961 504
rect 19019 -896 19159 504
rect 19217 -896 19357 504
rect 19415 -896 19555 504
rect 19613 -896 19753 504
rect 11495 -2532 11635 -1132
rect 11693 -2532 11833 -1132
rect 11891 -2532 12031 -1132
rect 12089 -2532 12229 -1132
rect 12287 -2532 12427 -1132
rect 12485 -2532 12625 -1132
rect 12683 -2532 12823 -1132
rect 12881 -2532 13021 -1132
rect 13079 -2532 13219 -1132
rect 13277 -2532 13417 -1132
rect 13475 -2532 13615 -1132
rect 13673 -2532 13813 -1132
rect 13871 -2532 14011 -1132
rect 14069 -2532 14209 -1132
rect 14267 -2532 14407 -1132
rect 14465 -2532 14605 -1132
rect 14663 -2532 14803 -1132
rect 14861 -2532 15001 -1132
rect 15059 -2532 15199 -1132
rect 15257 -2532 15397 -1132
rect 15455 -2532 15595 -1132
rect 15653 -2532 15793 -1132
rect 15851 -2532 15991 -1132
rect 16049 -2532 16189 -1132
rect 16247 -2532 16387 -1132
rect 16445 -2532 16585 -1132
rect 16643 -2532 16783 -1132
rect 16841 -2532 16981 -1132
rect 17039 -2532 17179 -1132
rect 17237 -2532 17377 -1132
rect 17435 -2532 17575 -1132
rect 17633 -2532 17773 -1132
rect 17831 -2532 17971 -1132
rect 18029 -2532 18169 -1132
rect 18227 -2532 18367 -1132
rect 18425 -2532 18565 -1132
rect 18623 -2532 18763 -1132
rect 18821 -2532 18961 -1132
rect 19019 -2532 19159 -1132
rect 19217 -2532 19357 -1132
rect 19415 -2532 19555 -1132
rect 19613 -2532 19753 -1132
rect 11495 -4168 11635 -2768
rect 11693 -4168 11833 -2768
rect 11891 -4168 12031 -2768
rect 12089 -4168 12229 -2768
rect 12287 -4168 12427 -2768
rect 12485 -4168 12625 -2768
rect 12683 -4168 12823 -2768
rect 12881 -4168 13021 -2768
rect 13079 -4168 13219 -2768
rect 13277 -4168 13417 -2768
rect 13475 -4168 13615 -2768
rect 13673 -4168 13813 -2768
rect 13871 -4168 14011 -2768
rect 14069 -4168 14209 -2768
rect 14267 -4168 14407 -2768
rect 14465 -4168 14605 -2768
rect 14663 -4168 14803 -2768
rect 14861 -4168 15001 -2768
rect 15059 -4168 15199 -2768
rect 15257 -4168 15397 -2768
rect 15455 -4168 15595 -2768
rect 15653 -4168 15793 -2768
rect 15851 -4168 15991 -2768
rect 16049 -4168 16189 -2768
rect 16247 -4168 16387 -2768
rect 16445 -4168 16585 -2768
rect 16643 -4168 16783 -2768
rect 16841 -4168 16981 -2768
rect 17039 -4168 17179 -2768
rect 17237 -4168 17377 -2768
rect 17435 -4168 17575 -2768
rect 17633 -4168 17773 -2768
rect 17831 -4168 17971 -2768
rect 18029 -4168 18169 -2768
rect 18227 -4168 18367 -2768
rect 18425 -4168 18565 -2768
rect 18623 -4168 18763 -2768
rect 18821 -4168 18961 -2768
rect 19019 -4168 19159 -2768
rect 19217 -4168 19357 -2768
rect 19415 -4168 19555 -2768
rect 19613 -4168 19753 -2768
rect 23345 740 23485 2140
rect 23543 740 23683 2140
rect 23741 740 23881 2140
rect 23939 740 24079 2140
rect 24137 740 24277 2140
rect 24335 740 24475 2140
rect 24533 740 24673 2140
rect 24731 740 24871 2140
rect 24929 740 25069 2140
rect 25127 740 25267 2140
rect 25325 740 25465 2140
rect 25523 740 25663 2140
rect 25721 740 25861 2140
rect 25919 740 26059 2140
rect 26117 740 26257 2140
rect 26315 740 26455 2140
rect 26513 740 26653 2140
rect 26711 740 26851 2140
rect 26909 740 27049 2140
rect 27107 740 27247 2140
rect 27305 740 27445 2140
rect 27503 740 27643 2140
rect 27701 740 27841 2140
rect 27899 740 28039 2140
rect 28097 740 28237 2140
rect 28295 740 28435 2140
rect 28493 740 28633 2140
rect 28691 740 28831 2140
rect 28889 740 29029 2140
rect 29087 740 29227 2140
rect 29285 740 29425 2140
rect 29483 740 29623 2140
rect 29681 740 29821 2140
rect 29879 740 30019 2140
rect 30077 740 30217 2140
rect 30275 740 30415 2140
rect 30473 740 30613 2140
rect 30671 740 30811 2140
rect 30869 740 31009 2140
rect 31067 740 31207 2140
rect 31265 740 31405 2140
rect 31463 740 31603 2140
rect 23345 -896 23485 504
rect 23543 -896 23683 504
rect 23741 -896 23881 504
rect 23939 -896 24079 504
rect 24137 -896 24277 504
rect 24335 -896 24475 504
rect 24533 -896 24673 504
rect 24731 -896 24871 504
rect 24929 -896 25069 504
rect 25127 -896 25267 504
rect 25325 -896 25465 504
rect 25523 -896 25663 504
rect 25721 -896 25861 504
rect 25919 -896 26059 504
rect 26117 -896 26257 504
rect 26315 -896 26455 504
rect 26513 -896 26653 504
rect 26711 -896 26851 504
rect 26909 -896 27049 504
rect 27107 -896 27247 504
rect 27305 -896 27445 504
rect 27503 -896 27643 504
rect 27701 -896 27841 504
rect 27899 -896 28039 504
rect 28097 -896 28237 504
rect 28295 -896 28435 504
rect 28493 -896 28633 504
rect 28691 -896 28831 504
rect 28889 -896 29029 504
rect 29087 -896 29227 504
rect 29285 -896 29425 504
rect 29483 -896 29623 504
rect 29681 -896 29821 504
rect 29879 -896 30019 504
rect 30077 -896 30217 504
rect 30275 -896 30415 504
rect 30473 -896 30613 504
rect 30671 -896 30811 504
rect 30869 -896 31009 504
rect 31067 -896 31207 504
rect 31265 -896 31405 504
rect 31463 -896 31603 504
rect 23345 -2532 23485 -1132
rect 23543 -2532 23683 -1132
rect 23741 -2532 23881 -1132
rect 23939 -2532 24079 -1132
rect 24137 -2532 24277 -1132
rect 24335 -2532 24475 -1132
rect 24533 -2532 24673 -1132
rect 24731 -2532 24871 -1132
rect 24929 -2532 25069 -1132
rect 25127 -2532 25267 -1132
rect 25325 -2532 25465 -1132
rect 25523 -2532 25663 -1132
rect 25721 -2532 25861 -1132
rect 25919 -2532 26059 -1132
rect 26117 -2532 26257 -1132
rect 26315 -2532 26455 -1132
rect 26513 -2532 26653 -1132
rect 26711 -2532 26851 -1132
rect 26909 -2532 27049 -1132
rect 27107 -2532 27247 -1132
rect 27305 -2532 27445 -1132
rect 27503 -2532 27643 -1132
rect 27701 -2532 27841 -1132
rect 27899 -2532 28039 -1132
rect 28097 -2532 28237 -1132
rect 28295 -2532 28435 -1132
rect 28493 -2532 28633 -1132
rect 28691 -2532 28831 -1132
rect 28889 -2532 29029 -1132
rect 29087 -2532 29227 -1132
rect 29285 -2532 29425 -1132
rect 29483 -2532 29623 -1132
rect 29681 -2532 29821 -1132
rect 29879 -2532 30019 -1132
rect 30077 -2532 30217 -1132
rect 30275 -2532 30415 -1132
rect 30473 -2532 30613 -1132
rect 30671 -2532 30811 -1132
rect 30869 -2532 31009 -1132
rect 31067 -2532 31207 -1132
rect 31265 -2532 31405 -1132
rect 31463 -2532 31603 -1132
rect 23345 -4168 23485 -2768
rect 23543 -4168 23683 -2768
rect 23741 -4168 23881 -2768
rect 23939 -4168 24079 -2768
rect 24137 -4168 24277 -2768
rect 24335 -4168 24475 -2768
rect 24533 -4168 24673 -2768
rect 24731 -4168 24871 -2768
rect 24929 -4168 25069 -2768
rect 25127 -4168 25267 -2768
rect 25325 -4168 25465 -2768
rect 25523 -4168 25663 -2768
rect 25721 -4168 25861 -2768
rect 25919 -4168 26059 -2768
rect 26117 -4168 26257 -2768
rect 26315 -4168 26455 -2768
rect 26513 -4168 26653 -2768
rect 26711 -4168 26851 -2768
rect 26909 -4168 27049 -2768
rect 27107 -4168 27247 -2768
rect 27305 -4168 27445 -2768
rect 27503 -4168 27643 -2768
rect 27701 -4168 27841 -2768
rect 27899 -4168 28039 -2768
rect 28097 -4168 28237 -2768
rect 28295 -4168 28435 -2768
rect 28493 -4168 28633 -2768
rect 28691 -4168 28831 -2768
rect 28889 -4168 29029 -2768
rect 29087 -4168 29227 -2768
rect 29285 -4168 29425 -2768
rect 29483 -4168 29623 -2768
rect 29681 -4168 29821 -2768
rect 29879 -4168 30019 -2768
rect 30077 -4168 30217 -2768
rect 30275 -4168 30415 -2768
rect 30473 -4168 30613 -2768
rect 30671 -4168 30811 -2768
rect 30869 -4168 31009 -2768
rect 31067 -4168 31207 -2768
rect 31265 -4168 31405 -2768
rect 31463 -4168 31603 -2768
<< pdiff >>
rect 11437 2128 11495 2140
rect 11437 752 11449 2128
rect 11483 752 11495 2128
rect 11437 740 11495 752
rect 11635 2128 11693 2140
rect 11635 752 11647 2128
rect 11681 752 11693 2128
rect 11635 740 11693 752
rect 11833 2128 11891 2140
rect 11833 752 11845 2128
rect 11879 752 11891 2128
rect 11833 740 11891 752
rect 12031 2128 12089 2140
rect 12031 752 12043 2128
rect 12077 752 12089 2128
rect 12031 740 12089 752
rect 12229 2128 12287 2140
rect 12229 752 12241 2128
rect 12275 752 12287 2128
rect 12229 740 12287 752
rect 12427 2128 12485 2140
rect 12427 752 12439 2128
rect 12473 752 12485 2128
rect 12427 740 12485 752
rect 12625 2128 12683 2140
rect 12625 752 12637 2128
rect 12671 752 12683 2128
rect 12625 740 12683 752
rect 12823 2128 12881 2140
rect 12823 752 12835 2128
rect 12869 752 12881 2128
rect 12823 740 12881 752
rect 13021 2128 13079 2140
rect 13021 752 13033 2128
rect 13067 752 13079 2128
rect 13021 740 13079 752
rect 13219 2128 13277 2140
rect 13219 752 13231 2128
rect 13265 752 13277 2128
rect 13219 740 13277 752
rect 13417 2128 13475 2140
rect 13417 752 13429 2128
rect 13463 752 13475 2128
rect 13417 740 13475 752
rect 13615 2128 13673 2140
rect 13615 752 13627 2128
rect 13661 752 13673 2128
rect 13615 740 13673 752
rect 13813 2128 13871 2140
rect 13813 752 13825 2128
rect 13859 752 13871 2128
rect 13813 740 13871 752
rect 14011 2128 14069 2140
rect 14011 752 14023 2128
rect 14057 752 14069 2128
rect 14011 740 14069 752
rect 14209 2128 14267 2140
rect 14209 752 14221 2128
rect 14255 752 14267 2128
rect 14209 740 14267 752
rect 14407 2128 14465 2140
rect 14407 752 14419 2128
rect 14453 752 14465 2128
rect 14407 740 14465 752
rect 14605 2128 14663 2140
rect 14605 752 14617 2128
rect 14651 752 14663 2128
rect 14605 740 14663 752
rect 14803 2128 14861 2140
rect 14803 752 14815 2128
rect 14849 752 14861 2128
rect 14803 740 14861 752
rect 15001 2128 15059 2140
rect 15001 752 15013 2128
rect 15047 752 15059 2128
rect 15001 740 15059 752
rect 15199 2128 15257 2140
rect 15199 752 15211 2128
rect 15245 752 15257 2128
rect 15199 740 15257 752
rect 15397 2128 15455 2140
rect 15397 752 15409 2128
rect 15443 752 15455 2128
rect 15397 740 15455 752
rect 15595 2128 15653 2140
rect 15595 752 15607 2128
rect 15641 752 15653 2128
rect 15595 740 15653 752
rect 15793 2128 15851 2140
rect 15793 752 15805 2128
rect 15839 752 15851 2128
rect 15793 740 15851 752
rect 15991 2128 16049 2140
rect 15991 752 16003 2128
rect 16037 752 16049 2128
rect 15991 740 16049 752
rect 16189 2128 16247 2140
rect 16189 752 16201 2128
rect 16235 752 16247 2128
rect 16189 740 16247 752
rect 16387 2128 16445 2140
rect 16387 752 16399 2128
rect 16433 752 16445 2128
rect 16387 740 16445 752
rect 16585 2128 16643 2140
rect 16585 752 16597 2128
rect 16631 752 16643 2128
rect 16585 740 16643 752
rect 16783 2128 16841 2140
rect 16783 752 16795 2128
rect 16829 752 16841 2128
rect 16783 740 16841 752
rect 16981 2128 17039 2140
rect 16981 752 16993 2128
rect 17027 752 17039 2128
rect 16981 740 17039 752
rect 17179 2128 17237 2140
rect 17179 752 17191 2128
rect 17225 752 17237 2128
rect 17179 740 17237 752
rect 17377 2128 17435 2140
rect 17377 752 17389 2128
rect 17423 752 17435 2128
rect 17377 740 17435 752
rect 17575 2128 17633 2140
rect 17575 752 17587 2128
rect 17621 752 17633 2128
rect 17575 740 17633 752
rect 17773 2128 17831 2140
rect 17773 752 17785 2128
rect 17819 752 17831 2128
rect 17773 740 17831 752
rect 17971 2128 18029 2140
rect 17971 752 17983 2128
rect 18017 752 18029 2128
rect 17971 740 18029 752
rect 18169 2128 18227 2140
rect 18169 752 18181 2128
rect 18215 752 18227 2128
rect 18169 740 18227 752
rect 18367 2128 18425 2140
rect 18367 752 18379 2128
rect 18413 752 18425 2128
rect 18367 740 18425 752
rect 18565 2128 18623 2140
rect 18565 752 18577 2128
rect 18611 752 18623 2128
rect 18565 740 18623 752
rect 18763 2128 18821 2140
rect 18763 752 18775 2128
rect 18809 752 18821 2128
rect 18763 740 18821 752
rect 18961 2128 19019 2140
rect 18961 752 18973 2128
rect 19007 752 19019 2128
rect 18961 740 19019 752
rect 19159 2128 19217 2140
rect 19159 752 19171 2128
rect 19205 752 19217 2128
rect 19159 740 19217 752
rect 19357 2128 19415 2140
rect 19357 752 19369 2128
rect 19403 752 19415 2128
rect 19357 740 19415 752
rect 19555 2128 19613 2140
rect 19555 752 19567 2128
rect 19601 752 19613 2128
rect 19555 740 19613 752
rect 19753 2128 19811 2140
rect 19753 752 19765 2128
rect 19799 752 19811 2128
rect 19753 740 19811 752
rect 11437 492 11495 504
rect 11437 -884 11449 492
rect 11483 -884 11495 492
rect 11437 -896 11495 -884
rect 11635 492 11693 504
rect 11635 -884 11647 492
rect 11681 -884 11693 492
rect 11635 -896 11693 -884
rect 11833 492 11891 504
rect 11833 -884 11845 492
rect 11879 -884 11891 492
rect 11833 -896 11891 -884
rect 12031 492 12089 504
rect 12031 -884 12043 492
rect 12077 -884 12089 492
rect 12031 -896 12089 -884
rect 12229 492 12287 504
rect 12229 -884 12241 492
rect 12275 -884 12287 492
rect 12229 -896 12287 -884
rect 12427 492 12485 504
rect 12427 -884 12439 492
rect 12473 -884 12485 492
rect 12427 -896 12485 -884
rect 12625 492 12683 504
rect 12625 -884 12637 492
rect 12671 -884 12683 492
rect 12625 -896 12683 -884
rect 12823 492 12881 504
rect 12823 -884 12835 492
rect 12869 -884 12881 492
rect 12823 -896 12881 -884
rect 13021 492 13079 504
rect 13021 -884 13033 492
rect 13067 -884 13079 492
rect 13021 -896 13079 -884
rect 13219 492 13277 504
rect 13219 -884 13231 492
rect 13265 -884 13277 492
rect 13219 -896 13277 -884
rect 13417 492 13475 504
rect 13417 -884 13429 492
rect 13463 -884 13475 492
rect 13417 -896 13475 -884
rect 13615 492 13673 504
rect 13615 -884 13627 492
rect 13661 -884 13673 492
rect 13615 -896 13673 -884
rect 13813 492 13871 504
rect 13813 -884 13825 492
rect 13859 -884 13871 492
rect 13813 -896 13871 -884
rect 14011 492 14069 504
rect 14011 -884 14023 492
rect 14057 -884 14069 492
rect 14011 -896 14069 -884
rect 14209 492 14267 504
rect 14209 -884 14221 492
rect 14255 -884 14267 492
rect 14209 -896 14267 -884
rect 14407 492 14465 504
rect 14407 -884 14419 492
rect 14453 -884 14465 492
rect 14407 -896 14465 -884
rect 14605 492 14663 504
rect 14605 -884 14617 492
rect 14651 -884 14663 492
rect 14605 -896 14663 -884
rect 14803 492 14861 504
rect 14803 -884 14815 492
rect 14849 -884 14861 492
rect 14803 -896 14861 -884
rect 15001 492 15059 504
rect 15001 -884 15013 492
rect 15047 -884 15059 492
rect 15001 -896 15059 -884
rect 15199 492 15257 504
rect 15199 -884 15211 492
rect 15245 -884 15257 492
rect 15199 -896 15257 -884
rect 15397 492 15455 504
rect 15397 -884 15409 492
rect 15443 -884 15455 492
rect 15397 -896 15455 -884
rect 15595 492 15653 504
rect 15595 -884 15607 492
rect 15641 -884 15653 492
rect 15595 -896 15653 -884
rect 15793 492 15851 504
rect 15793 -884 15805 492
rect 15839 -884 15851 492
rect 15793 -896 15851 -884
rect 15991 492 16049 504
rect 15991 -884 16003 492
rect 16037 -884 16049 492
rect 15991 -896 16049 -884
rect 16189 492 16247 504
rect 16189 -884 16201 492
rect 16235 -884 16247 492
rect 16189 -896 16247 -884
rect 16387 492 16445 504
rect 16387 -884 16399 492
rect 16433 -884 16445 492
rect 16387 -896 16445 -884
rect 16585 492 16643 504
rect 16585 -884 16597 492
rect 16631 -884 16643 492
rect 16585 -896 16643 -884
rect 16783 492 16841 504
rect 16783 -884 16795 492
rect 16829 -884 16841 492
rect 16783 -896 16841 -884
rect 16981 492 17039 504
rect 16981 -884 16993 492
rect 17027 -884 17039 492
rect 16981 -896 17039 -884
rect 17179 492 17237 504
rect 17179 -884 17191 492
rect 17225 -884 17237 492
rect 17179 -896 17237 -884
rect 17377 492 17435 504
rect 17377 -884 17389 492
rect 17423 -884 17435 492
rect 17377 -896 17435 -884
rect 17575 492 17633 504
rect 17575 -884 17587 492
rect 17621 -884 17633 492
rect 17575 -896 17633 -884
rect 17773 492 17831 504
rect 17773 -884 17785 492
rect 17819 -884 17831 492
rect 17773 -896 17831 -884
rect 17971 492 18029 504
rect 17971 -884 17983 492
rect 18017 -884 18029 492
rect 17971 -896 18029 -884
rect 18169 492 18227 504
rect 18169 -884 18181 492
rect 18215 -884 18227 492
rect 18169 -896 18227 -884
rect 18367 492 18425 504
rect 18367 -884 18379 492
rect 18413 -884 18425 492
rect 18367 -896 18425 -884
rect 18565 492 18623 504
rect 18565 -884 18577 492
rect 18611 -884 18623 492
rect 18565 -896 18623 -884
rect 18763 492 18821 504
rect 18763 -884 18775 492
rect 18809 -884 18821 492
rect 18763 -896 18821 -884
rect 18961 492 19019 504
rect 18961 -884 18973 492
rect 19007 -884 19019 492
rect 18961 -896 19019 -884
rect 19159 492 19217 504
rect 19159 -884 19171 492
rect 19205 -884 19217 492
rect 19159 -896 19217 -884
rect 19357 492 19415 504
rect 19357 -884 19369 492
rect 19403 -884 19415 492
rect 19357 -896 19415 -884
rect 19555 492 19613 504
rect 19555 -884 19567 492
rect 19601 -884 19613 492
rect 19555 -896 19613 -884
rect 19753 492 19811 504
rect 19753 -884 19765 492
rect 19799 -884 19811 492
rect 19753 -896 19811 -884
rect 11437 -1144 11495 -1132
rect 11437 -2520 11449 -1144
rect 11483 -2520 11495 -1144
rect 11437 -2532 11495 -2520
rect 11635 -1144 11693 -1132
rect 11635 -2520 11647 -1144
rect 11681 -2520 11693 -1144
rect 11635 -2532 11693 -2520
rect 11833 -1144 11891 -1132
rect 11833 -2520 11845 -1144
rect 11879 -2520 11891 -1144
rect 11833 -2532 11891 -2520
rect 12031 -1144 12089 -1132
rect 12031 -2520 12043 -1144
rect 12077 -2520 12089 -1144
rect 12031 -2532 12089 -2520
rect 12229 -1144 12287 -1132
rect 12229 -2520 12241 -1144
rect 12275 -2520 12287 -1144
rect 12229 -2532 12287 -2520
rect 12427 -1144 12485 -1132
rect 12427 -2520 12439 -1144
rect 12473 -2520 12485 -1144
rect 12427 -2532 12485 -2520
rect 12625 -1144 12683 -1132
rect 12625 -2520 12637 -1144
rect 12671 -2520 12683 -1144
rect 12625 -2532 12683 -2520
rect 12823 -1144 12881 -1132
rect 12823 -2520 12835 -1144
rect 12869 -2520 12881 -1144
rect 12823 -2532 12881 -2520
rect 13021 -1144 13079 -1132
rect 13021 -2520 13033 -1144
rect 13067 -2520 13079 -1144
rect 13021 -2532 13079 -2520
rect 13219 -1144 13277 -1132
rect 13219 -2520 13231 -1144
rect 13265 -2520 13277 -1144
rect 13219 -2532 13277 -2520
rect 13417 -1144 13475 -1132
rect 13417 -2520 13429 -1144
rect 13463 -2520 13475 -1144
rect 13417 -2532 13475 -2520
rect 13615 -1144 13673 -1132
rect 13615 -2520 13627 -1144
rect 13661 -2520 13673 -1144
rect 13615 -2532 13673 -2520
rect 13813 -1144 13871 -1132
rect 13813 -2520 13825 -1144
rect 13859 -2520 13871 -1144
rect 13813 -2532 13871 -2520
rect 14011 -1144 14069 -1132
rect 14011 -2520 14023 -1144
rect 14057 -2520 14069 -1144
rect 14011 -2532 14069 -2520
rect 14209 -1144 14267 -1132
rect 14209 -2520 14221 -1144
rect 14255 -2520 14267 -1144
rect 14209 -2532 14267 -2520
rect 14407 -1144 14465 -1132
rect 14407 -2520 14419 -1144
rect 14453 -2520 14465 -1144
rect 14407 -2532 14465 -2520
rect 14605 -1144 14663 -1132
rect 14605 -2520 14617 -1144
rect 14651 -2520 14663 -1144
rect 14605 -2532 14663 -2520
rect 14803 -1144 14861 -1132
rect 14803 -2520 14815 -1144
rect 14849 -2520 14861 -1144
rect 14803 -2532 14861 -2520
rect 15001 -1144 15059 -1132
rect 15001 -2520 15013 -1144
rect 15047 -2520 15059 -1144
rect 15001 -2532 15059 -2520
rect 15199 -1144 15257 -1132
rect 15199 -2520 15211 -1144
rect 15245 -2520 15257 -1144
rect 15199 -2532 15257 -2520
rect 15397 -1144 15455 -1132
rect 15397 -2520 15409 -1144
rect 15443 -2520 15455 -1144
rect 15397 -2532 15455 -2520
rect 15595 -1144 15653 -1132
rect 15595 -2520 15607 -1144
rect 15641 -2520 15653 -1144
rect 15595 -2532 15653 -2520
rect 15793 -1144 15851 -1132
rect 15793 -2520 15805 -1144
rect 15839 -2520 15851 -1144
rect 15793 -2532 15851 -2520
rect 15991 -1144 16049 -1132
rect 15991 -2520 16003 -1144
rect 16037 -2520 16049 -1144
rect 15991 -2532 16049 -2520
rect 16189 -1144 16247 -1132
rect 16189 -2520 16201 -1144
rect 16235 -2520 16247 -1144
rect 16189 -2532 16247 -2520
rect 16387 -1144 16445 -1132
rect 16387 -2520 16399 -1144
rect 16433 -2520 16445 -1144
rect 16387 -2532 16445 -2520
rect 16585 -1144 16643 -1132
rect 16585 -2520 16597 -1144
rect 16631 -2520 16643 -1144
rect 16585 -2532 16643 -2520
rect 16783 -1144 16841 -1132
rect 16783 -2520 16795 -1144
rect 16829 -2520 16841 -1144
rect 16783 -2532 16841 -2520
rect 16981 -1144 17039 -1132
rect 16981 -2520 16993 -1144
rect 17027 -2520 17039 -1144
rect 16981 -2532 17039 -2520
rect 17179 -1144 17237 -1132
rect 17179 -2520 17191 -1144
rect 17225 -2520 17237 -1144
rect 17179 -2532 17237 -2520
rect 17377 -1144 17435 -1132
rect 17377 -2520 17389 -1144
rect 17423 -2520 17435 -1144
rect 17377 -2532 17435 -2520
rect 17575 -1144 17633 -1132
rect 17575 -2520 17587 -1144
rect 17621 -2520 17633 -1144
rect 17575 -2532 17633 -2520
rect 17773 -1144 17831 -1132
rect 17773 -2520 17785 -1144
rect 17819 -2520 17831 -1144
rect 17773 -2532 17831 -2520
rect 17971 -1144 18029 -1132
rect 17971 -2520 17983 -1144
rect 18017 -2520 18029 -1144
rect 17971 -2532 18029 -2520
rect 18169 -1144 18227 -1132
rect 18169 -2520 18181 -1144
rect 18215 -2520 18227 -1144
rect 18169 -2532 18227 -2520
rect 18367 -1144 18425 -1132
rect 18367 -2520 18379 -1144
rect 18413 -2520 18425 -1144
rect 18367 -2532 18425 -2520
rect 18565 -1144 18623 -1132
rect 18565 -2520 18577 -1144
rect 18611 -2520 18623 -1144
rect 18565 -2532 18623 -2520
rect 18763 -1144 18821 -1132
rect 18763 -2520 18775 -1144
rect 18809 -2520 18821 -1144
rect 18763 -2532 18821 -2520
rect 18961 -1144 19019 -1132
rect 18961 -2520 18973 -1144
rect 19007 -2520 19019 -1144
rect 18961 -2532 19019 -2520
rect 19159 -1144 19217 -1132
rect 19159 -2520 19171 -1144
rect 19205 -2520 19217 -1144
rect 19159 -2532 19217 -2520
rect 19357 -1144 19415 -1132
rect 19357 -2520 19369 -1144
rect 19403 -2520 19415 -1144
rect 19357 -2532 19415 -2520
rect 19555 -1144 19613 -1132
rect 19555 -2520 19567 -1144
rect 19601 -2520 19613 -1144
rect 19555 -2532 19613 -2520
rect 19753 -1144 19811 -1132
rect 19753 -2520 19765 -1144
rect 19799 -2520 19811 -1144
rect 19753 -2532 19811 -2520
rect 11437 -2780 11495 -2768
rect 11437 -4156 11449 -2780
rect 11483 -4156 11495 -2780
rect 11437 -4168 11495 -4156
rect 11635 -2780 11693 -2768
rect 11635 -4156 11647 -2780
rect 11681 -4156 11693 -2780
rect 11635 -4168 11693 -4156
rect 11833 -2780 11891 -2768
rect 11833 -4156 11845 -2780
rect 11879 -4156 11891 -2780
rect 11833 -4168 11891 -4156
rect 12031 -2780 12089 -2768
rect 12031 -4156 12043 -2780
rect 12077 -4156 12089 -2780
rect 12031 -4168 12089 -4156
rect 12229 -2780 12287 -2768
rect 12229 -4156 12241 -2780
rect 12275 -4156 12287 -2780
rect 12229 -4168 12287 -4156
rect 12427 -2780 12485 -2768
rect 12427 -4156 12439 -2780
rect 12473 -4156 12485 -2780
rect 12427 -4168 12485 -4156
rect 12625 -2780 12683 -2768
rect 12625 -4156 12637 -2780
rect 12671 -4156 12683 -2780
rect 12625 -4168 12683 -4156
rect 12823 -2780 12881 -2768
rect 12823 -4156 12835 -2780
rect 12869 -4156 12881 -2780
rect 12823 -4168 12881 -4156
rect 13021 -2780 13079 -2768
rect 13021 -4156 13033 -2780
rect 13067 -4156 13079 -2780
rect 13021 -4168 13079 -4156
rect 13219 -2780 13277 -2768
rect 13219 -4156 13231 -2780
rect 13265 -4156 13277 -2780
rect 13219 -4168 13277 -4156
rect 13417 -2780 13475 -2768
rect 13417 -4156 13429 -2780
rect 13463 -4156 13475 -2780
rect 13417 -4168 13475 -4156
rect 13615 -2780 13673 -2768
rect 13615 -4156 13627 -2780
rect 13661 -4156 13673 -2780
rect 13615 -4168 13673 -4156
rect 13813 -2780 13871 -2768
rect 13813 -4156 13825 -2780
rect 13859 -4156 13871 -2780
rect 13813 -4168 13871 -4156
rect 14011 -2780 14069 -2768
rect 14011 -4156 14023 -2780
rect 14057 -4156 14069 -2780
rect 14011 -4168 14069 -4156
rect 14209 -2780 14267 -2768
rect 14209 -4156 14221 -2780
rect 14255 -4156 14267 -2780
rect 14209 -4168 14267 -4156
rect 14407 -2780 14465 -2768
rect 14407 -4156 14419 -2780
rect 14453 -4156 14465 -2780
rect 14407 -4168 14465 -4156
rect 14605 -2780 14663 -2768
rect 14605 -4156 14617 -2780
rect 14651 -4156 14663 -2780
rect 14605 -4168 14663 -4156
rect 14803 -2780 14861 -2768
rect 14803 -4156 14815 -2780
rect 14849 -4156 14861 -2780
rect 14803 -4168 14861 -4156
rect 15001 -2780 15059 -2768
rect 15001 -4156 15013 -2780
rect 15047 -4156 15059 -2780
rect 15001 -4168 15059 -4156
rect 15199 -2780 15257 -2768
rect 15199 -4156 15211 -2780
rect 15245 -4156 15257 -2780
rect 15199 -4168 15257 -4156
rect 15397 -2780 15455 -2768
rect 15397 -4156 15409 -2780
rect 15443 -4156 15455 -2780
rect 15397 -4168 15455 -4156
rect 15595 -2780 15653 -2768
rect 15595 -4156 15607 -2780
rect 15641 -4156 15653 -2780
rect 15595 -4168 15653 -4156
rect 15793 -2780 15851 -2768
rect 15793 -4156 15805 -2780
rect 15839 -4156 15851 -2780
rect 15793 -4168 15851 -4156
rect 15991 -2780 16049 -2768
rect 15991 -4156 16003 -2780
rect 16037 -4156 16049 -2780
rect 15991 -4168 16049 -4156
rect 16189 -2780 16247 -2768
rect 16189 -4156 16201 -2780
rect 16235 -4156 16247 -2780
rect 16189 -4168 16247 -4156
rect 16387 -2780 16445 -2768
rect 16387 -4156 16399 -2780
rect 16433 -4156 16445 -2780
rect 16387 -4168 16445 -4156
rect 16585 -2780 16643 -2768
rect 16585 -4156 16597 -2780
rect 16631 -4156 16643 -2780
rect 16585 -4168 16643 -4156
rect 16783 -2780 16841 -2768
rect 16783 -4156 16795 -2780
rect 16829 -4156 16841 -2780
rect 16783 -4168 16841 -4156
rect 16981 -2780 17039 -2768
rect 16981 -4156 16993 -2780
rect 17027 -4156 17039 -2780
rect 16981 -4168 17039 -4156
rect 17179 -2780 17237 -2768
rect 17179 -4156 17191 -2780
rect 17225 -4156 17237 -2780
rect 17179 -4168 17237 -4156
rect 17377 -2780 17435 -2768
rect 17377 -4156 17389 -2780
rect 17423 -4156 17435 -2780
rect 17377 -4168 17435 -4156
rect 17575 -2780 17633 -2768
rect 17575 -4156 17587 -2780
rect 17621 -4156 17633 -2780
rect 17575 -4168 17633 -4156
rect 17773 -2780 17831 -2768
rect 17773 -4156 17785 -2780
rect 17819 -4156 17831 -2780
rect 17773 -4168 17831 -4156
rect 17971 -2780 18029 -2768
rect 17971 -4156 17983 -2780
rect 18017 -4156 18029 -2780
rect 17971 -4168 18029 -4156
rect 18169 -2780 18227 -2768
rect 18169 -4156 18181 -2780
rect 18215 -4156 18227 -2780
rect 18169 -4168 18227 -4156
rect 18367 -2780 18425 -2768
rect 18367 -4156 18379 -2780
rect 18413 -4156 18425 -2780
rect 18367 -4168 18425 -4156
rect 18565 -2780 18623 -2768
rect 18565 -4156 18577 -2780
rect 18611 -4156 18623 -2780
rect 18565 -4168 18623 -4156
rect 18763 -2780 18821 -2768
rect 18763 -4156 18775 -2780
rect 18809 -4156 18821 -2780
rect 18763 -4168 18821 -4156
rect 18961 -2780 19019 -2768
rect 18961 -4156 18973 -2780
rect 19007 -4156 19019 -2780
rect 18961 -4168 19019 -4156
rect 19159 -2780 19217 -2768
rect 19159 -4156 19171 -2780
rect 19205 -4156 19217 -2780
rect 19159 -4168 19217 -4156
rect 19357 -2780 19415 -2768
rect 19357 -4156 19369 -2780
rect 19403 -4156 19415 -2780
rect 19357 -4168 19415 -4156
rect 19555 -2780 19613 -2768
rect 19555 -4156 19567 -2780
rect 19601 -4156 19613 -2780
rect 19555 -4168 19613 -4156
rect 19753 -2780 19811 -2768
rect 19753 -4156 19765 -2780
rect 19799 -4156 19811 -2780
rect 19753 -4168 19811 -4156
rect 23287 2128 23345 2140
rect 23287 752 23299 2128
rect 23333 752 23345 2128
rect 23287 740 23345 752
rect 23485 2128 23543 2140
rect 23485 752 23497 2128
rect 23531 752 23543 2128
rect 23485 740 23543 752
rect 23683 2128 23741 2140
rect 23683 752 23695 2128
rect 23729 752 23741 2128
rect 23683 740 23741 752
rect 23881 2128 23939 2140
rect 23881 752 23893 2128
rect 23927 752 23939 2128
rect 23881 740 23939 752
rect 24079 2128 24137 2140
rect 24079 752 24091 2128
rect 24125 752 24137 2128
rect 24079 740 24137 752
rect 24277 2128 24335 2140
rect 24277 752 24289 2128
rect 24323 752 24335 2128
rect 24277 740 24335 752
rect 24475 2128 24533 2140
rect 24475 752 24487 2128
rect 24521 752 24533 2128
rect 24475 740 24533 752
rect 24673 2128 24731 2140
rect 24673 752 24685 2128
rect 24719 752 24731 2128
rect 24673 740 24731 752
rect 24871 2128 24929 2140
rect 24871 752 24883 2128
rect 24917 752 24929 2128
rect 24871 740 24929 752
rect 25069 2128 25127 2140
rect 25069 752 25081 2128
rect 25115 752 25127 2128
rect 25069 740 25127 752
rect 25267 2128 25325 2140
rect 25267 752 25279 2128
rect 25313 752 25325 2128
rect 25267 740 25325 752
rect 25465 2128 25523 2140
rect 25465 752 25477 2128
rect 25511 752 25523 2128
rect 25465 740 25523 752
rect 25663 2128 25721 2140
rect 25663 752 25675 2128
rect 25709 752 25721 2128
rect 25663 740 25721 752
rect 25861 2128 25919 2140
rect 25861 752 25873 2128
rect 25907 752 25919 2128
rect 25861 740 25919 752
rect 26059 2128 26117 2140
rect 26059 752 26071 2128
rect 26105 752 26117 2128
rect 26059 740 26117 752
rect 26257 2128 26315 2140
rect 26257 752 26269 2128
rect 26303 752 26315 2128
rect 26257 740 26315 752
rect 26455 2128 26513 2140
rect 26455 752 26467 2128
rect 26501 752 26513 2128
rect 26455 740 26513 752
rect 26653 2128 26711 2140
rect 26653 752 26665 2128
rect 26699 752 26711 2128
rect 26653 740 26711 752
rect 26851 2128 26909 2140
rect 26851 752 26863 2128
rect 26897 752 26909 2128
rect 26851 740 26909 752
rect 27049 2128 27107 2140
rect 27049 752 27061 2128
rect 27095 752 27107 2128
rect 27049 740 27107 752
rect 27247 2128 27305 2140
rect 27247 752 27259 2128
rect 27293 752 27305 2128
rect 27247 740 27305 752
rect 27445 2128 27503 2140
rect 27445 752 27457 2128
rect 27491 752 27503 2128
rect 27445 740 27503 752
rect 27643 2128 27701 2140
rect 27643 752 27655 2128
rect 27689 752 27701 2128
rect 27643 740 27701 752
rect 27841 2128 27899 2140
rect 27841 752 27853 2128
rect 27887 752 27899 2128
rect 27841 740 27899 752
rect 28039 2128 28097 2140
rect 28039 752 28051 2128
rect 28085 752 28097 2128
rect 28039 740 28097 752
rect 28237 2128 28295 2140
rect 28237 752 28249 2128
rect 28283 752 28295 2128
rect 28237 740 28295 752
rect 28435 2128 28493 2140
rect 28435 752 28447 2128
rect 28481 752 28493 2128
rect 28435 740 28493 752
rect 28633 2128 28691 2140
rect 28633 752 28645 2128
rect 28679 752 28691 2128
rect 28633 740 28691 752
rect 28831 2128 28889 2140
rect 28831 752 28843 2128
rect 28877 752 28889 2128
rect 28831 740 28889 752
rect 29029 2128 29087 2140
rect 29029 752 29041 2128
rect 29075 752 29087 2128
rect 29029 740 29087 752
rect 29227 2128 29285 2140
rect 29227 752 29239 2128
rect 29273 752 29285 2128
rect 29227 740 29285 752
rect 29425 2128 29483 2140
rect 29425 752 29437 2128
rect 29471 752 29483 2128
rect 29425 740 29483 752
rect 29623 2128 29681 2140
rect 29623 752 29635 2128
rect 29669 752 29681 2128
rect 29623 740 29681 752
rect 29821 2128 29879 2140
rect 29821 752 29833 2128
rect 29867 752 29879 2128
rect 29821 740 29879 752
rect 30019 2128 30077 2140
rect 30019 752 30031 2128
rect 30065 752 30077 2128
rect 30019 740 30077 752
rect 30217 2128 30275 2140
rect 30217 752 30229 2128
rect 30263 752 30275 2128
rect 30217 740 30275 752
rect 30415 2128 30473 2140
rect 30415 752 30427 2128
rect 30461 752 30473 2128
rect 30415 740 30473 752
rect 30613 2128 30671 2140
rect 30613 752 30625 2128
rect 30659 752 30671 2128
rect 30613 740 30671 752
rect 30811 2128 30869 2140
rect 30811 752 30823 2128
rect 30857 752 30869 2128
rect 30811 740 30869 752
rect 31009 2128 31067 2140
rect 31009 752 31021 2128
rect 31055 752 31067 2128
rect 31009 740 31067 752
rect 31207 2128 31265 2140
rect 31207 752 31219 2128
rect 31253 752 31265 2128
rect 31207 740 31265 752
rect 31405 2128 31463 2140
rect 31405 752 31417 2128
rect 31451 752 31463 2128
rect 31405 740 31463 752
rect 31603 2128 31661 2140
rect 31603 752 31615 2128
rect 31649 752 31661 2128
rect 31603 740 31661 752
rect 23287 492 23345 504
rect 23287 -884 23299 492
rect 23333 -884 23345 492
rect 23287 -896 23345 -884
rect 23485 492 23543 504
rect 23485 -884 23497 492
rect 23531 -884 23543 492
rect 23485 -896 23543 -884
rect 23683 492 23741 504
rect 23683 -884 23695 492
rect 23729 -884 23741 492
rect 23683 -896 23741 -884
rect 23881 492 23939 504
rect 23881 -884 23893 492
rect 23927 -884 23939 492
rect 23881 -896 23939 -884
rect 24079 492 24137 504
rect 24079 -884 24091 492
rect 24125 -884 24137 492
rect 24079 -896 24137 -884
rect 24277 492 24335 504
rect 24277 -884 24289 492
rect 24323 -884 24335 492
rect 24277 -896 24335 -884
rect 24475 492 24533 504
rect 24475 -884 24487 492
rect 24521 -884 24533 492
rect 24475 -896 24533 -884
rect 24673 492 24731 504
rect 24673 -884 24685 492
rect 24719 -884 24731 492
rect 24673 -896 24731 -884
rect 24871 492 24929 504
rect 24871 -884 24883 492
rect 24917 -884 24929 492
rect 24871 -896 24929 -884
rect 25069 492 25127 504
rect 25069 -884 25081 492
rect 25115 -884 25127 492
rect 25069 -896 25127 -884
rect 25267 492 25325 504
rect 25267 -884 25279 492
rect 25313 -884 25325 492
rect 25267 -896 25325 -884
rect 25465 492 25523 504
rect 25465 -884 25477 492
rect 25511 -884 25523 492
rect 25465 -896 25523 -884
rect 25663 492 25721 504
rect 25663 -884 25675 492
rect 25709 -884 25721 492
rect 25663 -896 25721 -884
rect 25861 492 25919 504
rect 25861 -884 25873 492
rect 25907 -884 25919 492
rect 25861 -896 25919 -884
rect 26059 492 26117 504
rect 26059 -884 26071 492
rect 26105 -884 26117 492
rect 26059 -896 26117 -884
rect 26257 492 26315 504
rect 26257 -884 26269 492
rect 26303 -884 26315 492
rect 26257 -896 26315 -884
rect 26455 492 26513 504
rect 26455 -884 26467 492
rect 26501 -884 26513 492
rect 26455 -896 26513 -884
rect 26653 492 26711 504
rect 26653 -884 26665 492
rect 26699 -884 26711 492
rect 26653 -896 26711 -884
rect 26851 492 26909 504
rect 26851 -884 26863 492
rect 26897 -884 26909 492
rect 26851 -896 26909 -884
rect 27049 492 27107 504
rect 27049 -884 27061 492
rect 27095 -884 27107 492
rect 27049 -896 27107 -884
rect 27247 492 27305 504
rect 27247 -884 27259 492
rect 27293 -884 27305 492
rect 27247 -896 27305 -884
rect 27445 492 27503 504
rect 27445 -884 27457 492
rect 27491 -884 27503 492
rect 27445 -896 27503 -884
rect 27643 492 27701 504
rect 27643 -884 27655 492
rect 27689 -884 27701 492
rect 27643 -896 27701 -884
rect 27841 492 27899 504
rect 27841 -884 27853 492
rect 27887 -884 27899 492
rect 27841 -896 27899 -884
rect 28039 492 28097 504
rect 28039 -884 28051 492
rect 28085 -884 28097 492
rect 28039 -896 28097 -884
rect 28237 492 28295 504
rect 28237 -884 28249 492
rect 28283 -884 28295 492
rect 28237 -896 28295 -884
rect 28435 492 28493 504
rect 28435 -884 28447 492
rect 28481 -884 28493 492
rect 28435 -896 28493 -884
rect 28633 492 28691 504
rect 28633 -884 28645 492
rect 28679 -884 28691 492
rect 28633 -896 28691 -884
rect 28831 492 28889 504
rect 28831 -884 28843 492
rect 28877 -884 28889 492
rect 28831 -896 28889 -884
rect 29029 492 29087 504
rect 29029 -884 29041 492
rect 29075 -884 29087 492
rect 29029 -896 29087 -884
rect 29227 492 29285 504
rect 29227 -884 29239 492
rect 29273 -884 29285 492
rect 29227 -896 29285 -884
rect 29425 492 29483 504
rect 29425 -884 29437 492
rect 29471 -884 29483 492
rect 29425 -896 29483 -884
rect 29623 492 29681 504
rect 29623 -884 29635 492
rect 29669 -884 29681 492
rect 29623 -896 29681 -884
rect 29821 492 29879 504
rect 29821 -884 29833 492
rect 29867 -884 29879 492
rect 29821 -896 29879 -884
rect 30019 492 30077 504
rect 30019 -884 30031 492
rect 30065 -884 30077 492
rect 30019 -896 30077 -884
rect 30217 492 30275 504
rect 30217 -884 30229 492
rect 30263 -884 30275 492
rect 30217 -896 30275 -884
rect 30415 492 30473 504
rect 30415 -884 30427 492
rect 30461 -884 30473 492
rect 30415 -896 30473 -884
rect 30613 492 30671 504
rect 30613 -884 30625 492
rect 30659 -884 30671 492
rect 30613 -896 30671 -884
rect 30811 492 30869 504
rect 30811 -884 30823 492
rect 30857 -884 30869 492
rect 30811 -896 30869 -884
rect 31009 492 31067 504
rect 31009 -884 31021 492
rect 31055 -884 31067 492
rect 31009 -896 31067 -884
rect 31207 492 31265 504
rect 31207 -884 31219 492
rect 31253 -884 31265 492
rect 31207 -896 31265 -884
rect 31405 492 31463 504
rect 31405 -884 31417 492
rect 31451 -884 31463 492
rect 31405 -896 31463 -884
rect 31603 492 31661 504
rect 31603 -884 31615 492
rect 31649 -884 31661 492
rect 31603 -896 31661 -884
rect 23287 -1144 23345 -1132
rect 23287 -2520 23299 -1144
rect 23333 -2520 23345 -1144
rect 23287 -2532 23345 -2520
rect 23485 -1144 23543 -1132
rect 23485 -2520 23497 -1144
rect 23531 -2520 23543 -1144
rect 23485 -2532 23543 -2520
rect 23683 -1144 23741 -1132
rect 23683 -2520 23695 -1144
rect 23729 -2520 23741 -1144
rect 23683 -2532 23741 -2520
rect 23881 -1144 23939 -1132
rect 23881 -2520 23893 -1144
rect 23927 -2520 23939 -1144
rect 23881 -2532 23939 -2520
rect 24079 -1144 24137 -1132
rect 24079 -2520 24091 -1144
rect 24125 -2520 24137 -1144
rect 24079 -2532 24137 -2520
rect 24277 -1144 24335 -1132
rect 24277 -2520 24289 -1144
rect 24323 -2520 24335 -1144
rect 24277 -2532 24335 -2520
rect 24475 -1144 24533 -1132
rect 24475 -2520 24487 -1144
rect 24521 -2520 24533 -1144
rect 24475 -2532 24533 -2520
rect 24673 -1144 24731 -1132
rect 24673 -2520 24685 -1144
rect 24719 -2520 24731 -1144
rect 24673 -2532 24731 -2520
rect 24871 -1144 24929 -1132
rect 24871 -2520 24883 -1144
rect 24917 -2520 24929 -1144
rect 24871 -2532 24929 -2520
rect 25069 -1144 25127 -1132
rect 25069 -2520 25081 -1144
rect 25115 -2520 25127 -1144
rect 25069 -2532 25127 -2520
rect 25267 -1144 25325 -1132
rect 25267 -2520 25279 -1144
rect 25313 -2520 25325 -1144
rect 25267 -2532 25325 -2520
rect 25465 -1144 25523 -1132
rect 25465 -2520 25477 -1144
rect 25511 -2520 25523 -1144
rect 25465 -2532 25523 -2520
rect 25663 -1144 25721 -1132
rect 25663 -2520 25675 -1144
rect 25709 -2520 25721 -1144
rect 25663 -2532 25721 -2520
rect 25861 -1144 25919 -1132
rect 25861 -2520 25873 -1144
rect 25907 -2520 25919 -1144
rect 25861 -2532 25919 -2520
rect 26059 -1144 26117 -1132
rect 26059 -2520 26071 -1144
rect 26105 -2520 26117 -1144
rect 26059 -2532 26117 -2520
rect 26257 -1144 26315 -1132
rect 26257 -2520 26269 -1144
rect 26303 -2520 26315 -1144
rect 26257 -2532 26315 -2520
rect 26455 -1144 26513 -1132
rect 26455 -2520 26467 -1144
rect 26501 -2520 26513 -1144
rect 26455 -2532 26513 -2520
rect 26653 -1144 26711 -1132
rect 26653 -2520 26665 -1144
rect 26699 -2520 26711 -1144
rect 26653 -2532 26711 -2520
rect 26851 -1144 26909 -1132
rect 26851 -2520 26863 -1144
rect 26897 -2520 26909 -1144
rect 26851 -2532 26909 -2520
rect 27049 -1144 27107 -1132
rect 27049 -2520 27061 -1144
rect 27095 -2520 27107 -1144
rect 27049 -2532 27107 -2520
rect 27247 -1144 27305 -1132
rect 27247 -2520 27259 -1144
rect 27293 -2520 27305 -1144
rect 27247 -2532 27305 -2520
rect 27445 -1144 27503 -1132
rect 27445 -2520 27457 -1144
rect 27491 -2520 27503 -1144
rect 27445 -2532 27503 -2520
rect 27643 -1144 27701 -1132
rect 27643 -2520 27655 -1144
rect 27689 -2520 27701 -1144
rect 27643 -2532 27701 -2520
rect 27841 -1144 27899 -1132
rect 27841 -2520 27853 -1144
rect 27887 -2520 27899 -1144
rect 27841 -2532 27899 -2520
rect 28039 -1144 28097 -1132
rect 28039 -2520 28051 -1144
rect 28085 -2520 28097 -1144
rect 28039 -2532 28097 -2520
rect 28237 -1144 28295 -1132
rect 28237 -2520 28249 -1144
rect 28283 -2520 28295 -1144
rect 28237 -2532 28295 -2520
rect 28435 -1144 28493 -1132
rect 28435 -2520 28447 -1144
rect 28481 -2520 28493 -1144
rect 28435 -2532 28493 -2520
rect 28633 -1144 28691 -1132
rect 28633 -2520 28645 -1144
rect 28679 -2520 28691 -1144
rect 28633 -2532 28691 -2520
rect 28831 -1144 28889 -1132
rect 28831 -2520 28843 -1144
rect 28877 -2520 28889 -1144
rect 28831 -2532 28889 -2520
rect 29029 -1144 29087 -1132
rect 29029 -2520 29041 -1144
rect 29075 -2520 29087 -1144
rect 29029 -2532 29087 -2520
rect 29227 -1144 29285 -1132
rect 29227 -2520 29239 -1144
rect 29273 -2520 29285 -1144
rect 29227 -2532 29285 -2520
rect 29425 -1144 29483 -1132
rect 29425 -2520 29437 -1144
rect 29471 -2520 29483 -1144
rect 29425 -2532 29483 -2520
rect 29623 -1144 29681 -1132
rect 29623 -2520 29635 -1144
rect 29669 -2520 29681 -1144
rect 29623 -2532 29681 -2520
rect 29821 -1144 29879 -1132
rect 29821 -2520 29833 -1144
rect 29867 -2520 29879 -1144
rect 29821 -2532 29879 -2520
rect 30019 -1144 30077 -1132
rect 30019 -2520 30031 -1144
rect 30065 -2520 30077 -1144
rect 30019 -2532 30077 -2520
rect 30217 -1144 30275 -1132
rect 30217 -2520 30229 -1144
rect 30263 -2520 30275 -1144
rect 30217 -2532 30275 -2520
rect 30415 -1144 30473 -1132
rect 30415 -2520 30427 -1144
rect 30461 -2520 30473 -1144
rect 30415 -2532 30473 -2520
rect 30613 -1144 30671 -1132
rect 30613 -2520 30625 -1144
rect 30659 -2520 30671 -1144
rect 30613 -2532 30671 -2520
rect 30811 -1144 30869 -1132
rect 30811 -2520 30823 -1144
rect 30857 -2520 30869 -1144
rect 30811 -2532 30869 -2520
rect 31009 -1144 31067 -1132
rect 31009 -2520 31021 -1144
rect 31055 -2520 31067 -1144
rect 31009 -2532 31067 -2520
rect 31207 -1144 31265 -1132
rect 31207 -2520 31219 -1144
rect 31253 -2520 31265 -1144
rect 31207 -2532 31265 -2520
rect 31405 -1144 31463 -1132
rect 31405 -2520 31417 -1144
rect 31451 -2520 31463 -1144
rect 31405 -2532 31463 -2520
rect 31603 -1144 31661 -1132
rect 31603 -2520 31615 -1144
rect 31649 -2520 31661 -1144
rect 31603 -2532 31661 -2520
rect 23287 -2780 23345 -2768
rect 23287 -4156 23299 -2780
rect 23333 -4156 23345 -2780
rect 23287 -4168 23345 -4156
rect 23485 -2780 23543 -2768
rect 23485 -4156 23497 -2780
rect 23531 -4156 23543 -2780
rect 23485 -4168 23543 -4156
rect 23683 -2780 23741 -2768
rect 23683 -4156 23695 -2780
rect 23729 -4156 23741 -2780
rect 23683 -4168 23741 -4156
rect 23881 -2780 23939 -2768
rect 23881 -4156 23893 -2780
rect 23927 -4156 23939 -2780
rect 23881 -4168 23939 -4156
rect 24079 -2780 24137 -2768
rect 24079 -4156 24091 -2780
rect 24125 -4156 24137 -2780
rect 24079 -4168 24137 -4156
rect 24277 -2780 24335 -2768
rect 24277 -4156 24289 -2780
rect 24323 -4156 24335 -2780
rect 24277 -4168 24335 -4156
rect 24475 -2780 24533 -2768
rect 24475 -4156 24487 -2780
rect 24521 -4156 24533 -2780
rect 24475 -4168 24533 -4156
rect 24673 -2780 24731 -2768
rect 24673 -4156 24685 -2780
rect 24719 -4156 24731 -2780
rect 24673 -4168 24731 -4156
rect 24871 -2780 24929 -2768
rect 24871 -4156 24883 -2780
rect 24917 -4156 24929 -2780
rect 24871 -4168 24929 -4156
rect 25069 -2780 25127 -2768
rect 25069 -4156 25081 -2780
rect 25115 -4156 25127 -2780
rect 25069 -4168 25127 -4156
rect 25267 -2780 25325 -2768
rect 25267 -4156 25279 -2780
rect 25313 -4156 25325 -2780
rect 25267 -4168 25325 -4156
rect 25465 -2780 25523 -2768
rect 25465 -4156 25477 -2780
rect 25511 -4156 25523 -2780
rect 25465 -4168 25523 -4156
rect 25663 -2780 25721 -2768
rect 25663 -4156 25675 -2780
rect 25709 -4156 25721 -2780
rect 25663 -4168 25721 -4156
rect 25861 -2780 25919 -2768
rect 25861 -4156 25873 -2780
rect 25907 -4156 25919 -2780
rect 25861 -4168 25919 -4156
rect 26059 -2780 26117 -2768
rect 26059 -4156 26071 -2780
rect 26105 -4156 26117 -2780
rect 26059 -4168 26117 -4156
rect 26257 -2780 26315 -2768
rect 26257 -4156 26269 -2780
rect 26303 -4156 26315 -2780
rect 26257 -4168 26315 -4156
rect 26455 -2780 26513 -2768
rect 26455 -4156 26467 -2780
rect 26501 -4156 26513 -2780
rect 26455 -4168 26513 -4156
rect 26653 -2780 26711 -2768
rect 26653 -4156 26665 -2780
rect 26699 -4156 26711 -2780
rect 26653 -4168 26711 -4156
rect 26851 -2780 26909 -2768
rect 26851 -4156 26863 -2780
rect 26897 -4156 26909 -2780
rect 26851 -4168 26909 -4156
rect 27049 -2780 27107 -2768
rect 27049 -4156 27061 -2780
rect 27095 -4156 27107 -2780
rect 27049 -4168 27107 -4156
rect 27247 -2780 27305 -2768
rect 27247 -4156 27259 -2780
rect 27293 -4156 27305 -2780
rect 27247 -4168 27305 -4156
rect 27445 -2780 27503 -2768
rect 27445 -4156 27457 -2780
rect 27491 -4156 27503 -2780
rect 27445 -4168 27503 -4156
rect 27643 -2780 27701 -2768
rect 27643 -4156 27655 -2780
rect 27689 -4156 27701 -2780
rect 27643 -4168 27701 -4156
rect 27841 -2780 27899 -2768
rect 27841 -4156 27853 -2780
rect 27887 -4156 27899 -2780
rect 27841 -4168 27899 -4156
rect 28039 -2780 28097 -2768
rect 28039 -4156 28051 -2780
rect 28085 -4156 28097 -2780
rect 28039 -4168 28097 -4156
rect 28237 -2780 28295 -2768
rect 28237 -4156 28249 -2780
rect 28283 -4156 28295 -2780
rect 28237 -4168 28295 -4156
rect 28435 -2780 28493 -2768
rect 28435 -4156 28447 -2780
rect 28481 -4156 28493 -2780
rect 28435 -4168 28493 -4156
rect 28633 -2780 28691 -2768
rect 28633 -4156 28645 -2780
rect 28679 -4156 28691 -2780
rect 28633 -4168 28691 -4156
rect 28831 -2780 28889 -2768
rect 28831 -4156 28843 -2780
rect 28877 -4156 28889 -2780
rect 28831 -4168 28889 -4156
rect 29029 -2780 29087 -2768
rect 29029 -4156 29041 -2780
rect 29075 -4156 29087 -2780
rect 29029 -4168 29087 -4156
rect 29227 -2780 29285 -2768
rect 29227 -4156 29239 -2780
rect 29273 -4156 29285 -2780
rect 29227 -4168 29285 -4156
rect 29425 -2780 29483 -2768
rect 29425 -4156 29437 -2780
rect 29471 -4156 29483 -2780
rect 29425 -4168 29483 -4156
rect 29623 -2780 29681 -2768
rect 29623 -4156 29635 -2780
rect 29669 -4156 29681 -2780
rect 29623 -4168 29681 -4156
rect 29821 -2780 29879 -2768
rect 29821 -4156 29833 -2780
rect 29867 -4156 29879 -2780
rect 29821 -4168 29879 -4156
rect 30019 -2780 30077 -2768
rect 30019 -4156 30031 -2780
rect 30065 -4156 30077 -2780
rect 30019 -4168 30077 -4156
rect 30217 -2780 30275 -2768
rect 30217 -4156 30229 -2780
rect 30263 -4156 30275 -2780
rect 30217 -4168 30275 -4156
rect 30415 -2780 30473 -2768
rect 30415 -4156 30427 -2780
rect 30461 -4156 30473 -2780
rect 30415 -4168 30473 -4156
rect 30613 -2780 30671 -2768
rect 30613 -4156 30625 -2780
rect 30659 -4156 30671 -2780
rect 30613 -4168 30671 -4156
rect 30811 -2780 30869 -2768
rect 30811 -4156 30823 -2780
rect 30857 -4156 30869 -2780
rect 30811 -4168 30869 -4156
rect 31009 -2780 31067 -2768
rect 31009 -4156 31021 -2780
rect 31055 -4156 31067 -2780
rect 31009 -4168 31067 -4156
rect 31207 -2780 31265 -2768
rect 31207 -4156 31219 -2780
rect 31253 -4156 31265 -2780
rect 31207 -4168 31265 -4156
rect 31405 -2780 31463 -2768
rect 31405 -4156 31417 -2780
rect 31451 -4156 31463 -2780
rect 31405 -4168 31463 -4156
rect 31603 -2780 31661 -2768
rect 31603 -4156 31615 -2780
rect 31649 -4156 31661 -2780
rect 31603 -4168 31661 -4156
<< pdiffc >>
rect 11449 752 11483 2128
rect 11647 752 11681 2128
rect 11845 752 11879 2128
rect 12043 752 12077 2128
rect 12241 752 12275 2128
rect 12439 752 12473 2128
rect 12637 752 12671 2128
rect 12835 752 12869 2128
rect 13033 752 13067 2128
rect 13231 752 13265 2128
rect 13429 752 13463 2128
rect 13627 752 13661 2128
rect 13825 752 13859 2128
rect 14023 752 14057 2128
rect 14221 752 14255 2128
rect 14419 752 14453 2128
rect 14617 752 14651 2128
rect 14815 752 14849 2128
rect 15013 752 15047 2128
rect 15211 752 15245 2128
rect 15409 752 15443 2128
rect 15607 752 15641 2128
rect 15805 752 15839 2128
rect 16003 752 16037 2128
rect 16201 752 16235 2128
rect 16399 752 16433 2128
rect 16597 752 16631 2128
rect 16795 752 16829 2128
rect 16993 752 17027 2128
rect 17191 752 17225 2128
rect 17389 752 17423 2128
rect 17587 752 17621 2128
rect 17785 752 17819 2128
rect 17983 752 18017 2128
rect 18181 752 18215 2128
rect 18379 752 18413 2128
rect 18577 752 18611 2128
rect 18775 752 18809 2128
rect 18973 752 19007 2128
rect 19171 752 19205 2128
rect 19369 752 19403 2128
rect 19567 752 19601 2128
rect 19765 752 19799 2128
rect 11449 -884 11483 492
rect 11647 -884 11681 492
rect 11845 -884 11879 492
rect 12043 -884 12077 492
rect 12241 -884 12275 492
rect 12439 -884 12473 492
rect 12637 -884 12671 492
rect 12835 -884 12869 492
rect 13033 -884 13067 492
rect 13231 -884 13265 492
rect 13429 -884 13463 492
rect 13627 -884 13661 492
rect 13825 -884 13859 492
rect 14023 -884 14057 492
rect 14221 -884 14255 492
rect 14419 -884 14453 492
rect 14617 -884 14651 492
rect 14815 -884 14849 492
rect 15013 -884 15047 492
rect 15211 -884 15245 492
rect 15409 -884 15443 492
rect 15607 -884 15641 492
rect 15805 -884 15839 492
rect 16003 -884 16037 492
rect 16201 -884 16235 492
rect 16399 -884 16433 492
rect 16597 -884 16631 492
rect 16795 -884 16829 492
rect 16993 -884 17027 492
rect 17191 -884 17225 492
rect 17389 -884 17423 492
rect 17587 -884 17621 492
rect 17785 -884 17819 492
rect 17983 -884 18017 492
rect 18181 -884 18215 492
rect 18379 -884 18413 492
rect 18577 -884 18611 492
rect 18775 -884 18809 492
rect 18973 -884 19007 492
rect 19171 -884 19205 492
rect 19369 -884 19403 492
rect 19567 -884 19601 492
rect 19765 -884 19799 492
rect 11449 -2520 11483 -1144
rect 11647 -2520 11681 -1144
rect 11845 -2520 11879 -1144
rect 12043 -2520 12077 -1144
rect 12241 -2520 12275 -1144
rect 12439 -2520 12473 -1144
rect 12637 -2520 12671 -1144
rect 12835 -2520 12869 -1144
rect 13033 -2520 13067 -1144
rect 13231 -2520 13265 -1144
rect 13429 -2520 13463 -1144
rect 13627 -2520 13661 -1144
rect 13825 -2520 13859 -1144
rect 14023 -2520 14057 -1144
rect 14221 -2520 14255 -1144
rect 14419 -2520 14453 -1144
rect 14617 -2520 14651 -1144
rect 14815 -2520 14849 -1144
rect 15013 -2520 15047 -1144
rect 15211 -2520 15245 -1144
rect 15409 -2520 15443 -1144
rect 15607 -2520 15641 -1144
rect 15805 -2520 15839 -1144
rect 16003 -2520 16037 -1144
rect 16201 -2520 16235 -1144
rect 16399 -2520 16433 -1144
rect 16597 -2520 16631 -1144
rect 16795 -2520 16829 -1144
rect 16993 -2520 17027 -1144
rect 17191 -2520 17225 -1144
rect 17389 -2520 17423 -1144
rect 17587 -2520 17621 -1144
rect 17785 -2520 17819 -1144
rect 17983 -2520 18017 -1144
rect 18181 -2520 18215 -1144
rect 18379 -2520 18413 -1144
rect 18577 -2520 18611 -1144
rect 18775 -2520 18809 -1144
rect 18973 -2520 19007 -1144
rect 19171 -2520 19205 -1144
rect 19369 -2520 19403 -1144
rect 19567 -2520 19601 -1144
rect 19765 -2520 19799 -1144
rect 11449 -4156 11483 -2780
rect 11647 -4156 11681 -2780
rect 11845 -4156 11879 -2780
rect 12043 -4156 12077 -2780
rect 12241 -4156 12275 -2780
rect 12439 -4156 12473 -2780
rect 12637 -4156 12671 -2780
rect 12835 -4156 12869 -2780
rect 13033 -4156 13067 -2780
rect 13231 -4156 13265 -2780
rect 13429 -4156 13463 -2780
rect 13627 -4156 13661 -2780
rect 13825 -4156 13859 -2780
rect 14023 -4156 14057 -2780
rect 14221 -4156 14255 -2780
rect 14419 -4156 14453 -2780
rect 14617 -4156 14651 -2780
rect 14815 -4156 14849 -2780
rect 15013 -4156 15047 -2780
rect 15211 -4156 15245 -2780
rect 15409 -4156 15443 -2780
rect 15607 -4156 15641 -2780
rect 15805 -4156 15839 -2780
rect 16003 -4156 16037 -2780
rect 16201 -4156 16235 -2780
rect 16399 -4156 16433 -2780
rect 16597 -4156 16631 -2780
rect 16795 -4156 16829 -2780
rect 16993 -4156 17027 -2780
rect 17191 -4156 17225 -2780
rect 17389 -4156 17423 -2780
rect 17587 -4156 17621 -2780
rect 17785 -4156 17819 -2780
rect 17983 -4156 18017 -2780
rect 18181 -4156 18215 -2780
rect 18379 -4156 18413 -2780
rect 18577 -4156 18611 -2780
rect 18775 -4156 18809 -2780
rect 18973 -4156 19007 -2780
rect 19171 -4156 19205 -2780
rect 19369 -4156 19403 -2780
rect 19567 -4156 19601 -2780
rect 19765 -4156 19799 -2780
rect 23299 752 23333 2128
rect 23497 752 23531 2128
rect 23695 752 23729 2128
rect 23893 752 23927 2128
rect 24091 752 24125 2128
rect 24289 752 24323 2128
rect 24487 752 24521 2128
rect 24685 752 24719 2128
rect 24883 752 24917 2128
rect 25081 752 25115 2128
rect 25279 752 25313 2128
rect 25477 752 25511 2128
rect 25675 752 25709 2128
rect 25873 752 25907 2128
rect 26071 752 26105 2128
rect 26269 752 26303 2128
rect 26467 752 26501 2128
rect 26665 752 26699 2128
rect 26863 752 26897 2128
rect 27061 752 27095 2128
rect 27259 752 27293 2128
rect 27457 752 27491 2128
rect 27655 752 27689 2128
rect 27853 752 27887 2128
rect 28051 752 28085 2128
rect 28249 752 28283 2128
rect 28447 752 28481 2128
rect 28645 752 28679 2128
rect 28843 752 28877 2128
rect 29041 752 29075 2128
rect 29239 752 29273 2128
rect 29437 752 29471 2128
rect 29635 752 29669 2128
rect 29833 752 29867 2128
rect 30031 752 30065 2128
rect 30229 752 30263 2128
rect 30427 752 30461 2128
rect 30625 752 30659 2128
rect 30823 752 30857 2128
rect 31021 752 31055 2128
rect 31219 752 31253 2128
rect 31417 752 31451 2128
rect 31615 752 31649 2128
rect 23299 -884 23333 492
rect 23497 -884 23531 492
rect 23695 -884 23729 492
rect 23893 -884 23927 492
rect 24091 -884 24125 492
rect 24289 -884 24323 492
rect 24487 -884 24521 492
rect 24685 -884 24719 492
rect 24883 -884 24917 492
rect 25081 -884 25115 492
rect 25279 -884 25313 492
rect 25477 -884 25511 492
rect 25675 -884 25709 492
rect 25873 -884 25907 492
rect 26071 -884 26105 492
rect 26269 -884 26303 492
rect 26467 -884 26501 492
rect 26665 -884 26699 492
rect 26863 -884 26897 492
rect 27061 -884 27095 492
rect 27259 -884 27293 492
rect 27457 -884 27491 492
rect 27655 -884 27689 492
rect 27853 -884 27887 492
rect 28051 -884 28085 492
rect 28249 -884 28283 492
rect 28447 -884 28481 492
rect 28645 -884 28679 492
rect 28843 -884 28877 492
rect 29041 -884 29075 492
rect 29239 -884 29273 492
rect 29437 -884 29471 492
rect 29635 -884 29669 492
rect 29833 -884 29867 492
rect 30031 -884 30065 492
rect 30229 -884 30263 492
rect 30427 -884 30461 492
rect 30625 -884 30659 492
rect 30823 -884 30857 492
rect 31021 -884 31055 492
rect 31219 -884 31253 492
rect 31417 -884 31451 492
rect 31615 -884 31649 492
rect 23299 -2520 23333 -1144
rect 23497 -2520 23531 -1144
rect 23695 -2520 23729 -1144
rect 23893 -2520 23927 -1144
rect 24091 -2520 24125 -1144
rect 24289 -2520 24323 -1144
rect 24487 -2520 24521 -1144
rect 24685 -2520 24719 -1144
rect 24883 -2520 24917 -1144
rect 25081 -2520 25115 -1144
rect 25279 -2520 25313 -1144
rect 25477 -2520 25511 -1144
rect 25675 -2520 25709 -1144
rect 25873 -2520 25907 -1144
rect 26071 -2520 26105 -1144
rect 26269 -2520 26303 -1144
rect 26467 -2520 26501 -1144
rect 26665 -2520 26699 -1144
rect 26863 -2520 26897 -1144
rect 27061 -2520 27095 -1144
rect 27259 -2520 27293 -1144
rect 27457 -2520 27491 -1144
rect 27655 -2520 27689 -1144
rect 27853 -2520 27887 -1144
rect 28051 -2520 28085 -1144
rect 28249 -2520 28283 -1144
rect 28447 -2520 28481 -1144
rect 28645 -2520 28679 -1144
rect 28843 -2520 28877 -1144
rect 29041 -2520 29075 -1144
rect 29239 -2520 29273 -1144
rect 29437 -2520 29471 -1144
rect 29635 -2520 29669 -1144
rect 29833 -2520 29867 -1144
rect 30031 -2520 30065 -1144
rect 30229 -2520 30263 -1144
rect 30427 -2520 30461 -1144
rect 30625 -2520 30659 -1144
rect 30823 -2520 30857 -1144
rect 31021 -2520 31055 -1144
rect 31219 -2520 31253 -1144
rect 31417 -2520 31451 -1144
rect 31615 -2520 31649 -1144
rect 23299 -4156 23333 -2780
rect 23497 -4156 23531 -2780
rect 23695 -4156 23729 -2780
rect 23893 -4156 23927 -2780
rect 24091 -4156 24125 -2780
rect 24289 -4156 24323 -2780
rect 24487 -4156 24521 -2780
rect 24685 -4156 24719 -2780
rect 24883 -4156 24917 -2780
rect 25081 -4156 25115 -2780
rect 25279 -4156 25313 -2780
rect 25477 -4156 25511 -2780
rect 25675 -4156 25709 -2780
rect 25873 -4156 25907 -2780
rect 26071 -4156 26105 -2780
rect 26269 -4156 26303 -2780
rect 26467 -4156 26501 -2780
rect 26665 -4156 26699 -2780
rect 26863 -4156 26897 -2780
rect 27061 -4156 27095 -2780
rect 27259 -4156 27293 -2780
rect 27457 -4156 27491 -2780
rect 27655 -4156 27689 -2780
rect 27853 -4156 27887 -2780
rect 28051 -4156 28085 -2780
rect 28249 -4156 28283 -2780
rect 28447 -4156 28481 -2780
rect 28645 -4156 28679 -2780
rect 28843 -4156 28877 -2780
rect 29041 -4156 29075 -2780
rect 29239 -4156 29273 -2780
rect 29437 -4156 29471 -2780
rect 29635 -4156 29669 -2780
rect 29833 -4156 29867 -2780
rect 30031 -4156 30065 -2780
rect 30229 -4156 30263 -2780
rect 30427 -4156 30461 -2780
rect 30625 -4156 30659 -2780
rect 30823 -4156 30857 -2780
rect 31021 -4156 31055 -2780
rect 31219 -4156 31253 -2780
rect 31417 -4156 31451 -2780
rect 31615 -4156 31649 -2780
<< nsubdiff >>
rect -848 2237 -752 2271
rect 8337 2237 8433 2271
rect -848 2175 -814 2237
rect -848 -4415 -814 -4353
rect 8399 2175 8433 2237
rect 8399 -4415 8433 -4353
rect -848 -4449 -752 -4415
rect 8337 -4449 8433 -4415
rect 10991 2237 11087 2271
rect 20176 2237 20272 2271
rect 10991 2175 11025 2237
rect 20238 2175 20272 2237
rect 10991 -4415 11025 -4353
rect 20238 -4415 20272 -4353
rect 10991 -4449 11087 -4415
rect 20176 -4449 20272 -4415
rect 22841 2237 22937 2271
rect 32026 2237 32122 2271
rect 22841 2175 22875 2237
rect 32088 2175 32122 2237
rect 22841 -4415 22875 -4353
rect 32088 -4415 32122 -4353
rect 22841 -4449 22937 -4415
rect 32026 -4449 32122 -4415
<< nsubdiffcont >>
rect -752 2237 8337 2271
rect -848 -4353 -814 2175
rect 8399 -4353 8433 2175
rect -752 -4449 8337 -4415
rect 11087 2237 20176 2271
rect 10991 -4353 11025 2175
rect 20238 -4353 20272 2175
rect 11087 -4449 20176 -4415
rect 22937 2237 32026 2271
rect 22841 -4353 22875 2175
rect 32088 -4353 32122 2175
rect 22937 -4449 32026 -4415
<< poly >>
rect 11495 2140 11635 2166
rect 11693 2140 11833 2166
rect 11891 2140 12031 2166
rect 12089 2140 12229 2166
rect 12287 2140 12427 2166
rect 12485 2140 12625 2166
rect 12683 2140 12823 2166
rect 12881 2140 13021 2166
rect 13079 2140 13219 2166
rect 13277 2140 13417 2166
rect 13475 2140 13615 2166
rect 13673 2140 13813 2166
rect 13871 2140 14011 2166
rect 14069 2140 14209 2166
rect 14267 2140 14407 2166
rect 14465 2140 14605 2166
rect 14663 2140 14803 2166
rect 14861 2140 15001 2166
rect 15059 2140 15199 2166
rect 15257 2140 15397 2166
rect 15455 2140 15595 2166
rect 15653 2140 15793 2166
rect 15851 2140 15991 2166
rect 16049 2140 16189 2166
rect 16247 2140 16387 2166
rect 16445 2140 16585 2166
rect 16643 2140 16783 2166
rect 16841 2140 16981 2166
rect 17039 2140 17179 2166
rect 17237 2140 17377 2166
rect 17435 2140 17575 2166
rect 17633 2140 17773 2166
rect 17831 2140 17971 2166
rect 18029 2140 18169 2166
rect 18227 2140 18367 2166
rect 18425 2140 18565 2166
rect 18623 2140 18763 2166
rect 18821 2140 18961 2166
rect 19019 2140 19159 2166
rect 19217 2140 19357 2166
rect 19415 2140 19555 2166
rect 19613 2140 19753 2166
rect 11495 693 11635 740
rect 11495 659 11511 693
rect 11619 659 11635 693
rect 11495 643 11635 659
rect 11693 693 11833 740
rect 11693 659 11709 693
rect 11817 659 11833 693
rect 11693 643 11833 659
rect 11891 693 12031 740
rect 11891 659 11907 693
rect 12015 659 12031 693
rect 11891 643 12031 659
rect 12089 693 12229 740
rect 12089 659 12105 693
rect 12213 659 12229 693
rect 12089 643 12229 659
rect 12287 693 12427 740
rect 12287 659 12303 693
rect 12411 659 12427 693
rect 12287 643 12427 659
rect 12485 693 12625 740
rect 12485 659 12501 693
rect 12609 659 12625 693
rect 12485 643 12625 659
rect 12683 693 12823 740
rect 12683 659 12699 693
rect 12807 659 12823 693
rect 12683 643 12823 659
rect 12881 693 13021 740
rect 12881 659 12897 693
rect 13005 659 13021 693
rect 12881 643 13021 659
rect 13079 693 13219 740
rect 13079 659 13095 693
rect 13203 659 13219 693
rect 13079 643 13219 659
rect 13277 693 13417 740
rect 13277 659 13293 693
rect 13401 659 13417 693
rect 13277 643 13417 659
rect 13475 693 13615 740
rect 13475 659 13491 693
rect 13599 659 13615 693
rect 13475 643 13615 659
rect 13673 693 13813 740
rect 13673 659 13689 693
rect 13797 659 13813 693
rect 13673 643 13813 659
rect 13871 693 14011 740
rect 13871 659 13887 693
rect 13995 659 14011 693
rect 13871 643 14011 659
rect 14069 693 14209 740
rect 14069 659 14085 693
rect 14193 659 14209 693
rect 14069 643 14209 659
rect 14267 693 14407 740
rect 14267 659 14283 693
rect 14391 659 14407 693
rect 14267 643 14407 659
rect 14465 693 14605 740
rect 14465 659 14481 693
rect 14589 659 14605 693
rect 14465 643 14605 659
rect 14663 693 14803 740
rect 14663 659 14679 693
rect 14787 659 14803 693
rect 14663 643 14803 659
rect 14861 693 15001 740
rect 14861 659 14877 693
rect 14985 659 15001 693
rect 14861 643 15001 659
rect 15059 693 15199 740
rect 15059 659 15075 693
rect 15183 659 15199 693
rect 15059 643 15199 659
rect 15257 693 15397 740
rect 15257 659 15273 693
rect 15381 659 15397 693
rect 15257 643 15397 659
rect 15455 693 15595 740
rect 15455 659 15471 693
rect 15579 659 15595 693
rect 15455 643 15595 659
rect 15653 693 15793 740
rect 15653 659 15669 693
rect 15777 659 15793 693
rect 15653 643 15793 659
rect 15851 693 15991 740
rect 15851 659 15867 693
rect 15975 659 15991 693
rect 15851 643 15991 659
rect 16049 693 16189 740
rect 16049 659 16065 693
rect 16173 659 16189 693
rect 16049 643 16189 659
rect 16247 693 16387 740
rect 16247 659 16263 693
rect 16371 659 16387 693
rect 16247 643 16387 659
rect 16445 693 16585 740
rect 16445 659 16461 693
rect 16569 659 16585 693
rect 16445 643 16585 659
rect 16643 693 16783 740
rect 16643 659 16659 693
rect 16767 659 16783 693
rect 16643 643 16783 659
rect 16841 693 16981 740
rect 16841 659 16857 693
rect 16965 659 16981 693
rect 16841 643 16981 659
rect 17039 693 17179 740
rect 17039 659 17055 693
rect 17163 659 17179 693
rect 17039 643 17179 659
rect 17237 693 17377 740
rect 17237 659 17253 693
rect 17361 659 17377 693
rect 17237 643 17377 659
rect 17435 693 17575 740
rect 17435 659 17451 693
rect 17559 659 17575 693
rect 17435 643 17575 659
rect 17633 693 17773 740
rect 17633 659 17649 693
rect 17757 659 17773 693
rect 17633 643 17773 659
rect 17831 693 17971 740
rect 17831 659 17847 693
rect 17955 659 17971 693
rect 17831 643 17971 659
rect 18029 693 18169 740
rect 18029 659 18045 693
rect 18153 659 18169 693
rect 18029 643 18169 659
rect 18227 693 18367 740
rect 18227 659 18243 693
rect 18351 659 18367 693
rect 18227 643 18367 659
rect 18425 693 18565 740
rect 18425 659 18441 693
rect 18549 659 18565 693
rect 18425 643 18565 659
rect 18623 693 18763 740
rect 18623 659 18639 693
rect 18747 659 18763 693
rect 18623 643 18763 659
rect 18821 693 18961 740
rect 18821 659 18837 693
rect 18945 659 18961 693
rect 18821 643 18961 659
rect 19019 693 19159 740
rect 19019 659 19035 693
rect 19143 659 19159 693
rect 19019 643 19159 659
rect 19217 693 19357 740
rect 19217 659 19233 693
rect 19341 659 19357 693
rect 19217 643 19357 659
rect 19415 693 19555 740
rect 19415 659 19431 693
rect 19539 659 19555 693
rect 19415 643 19555 659
rect 19613 693 19753 740
rect 19613 659 19629 693
rect 19737 659 19753 693
rect 19613 643 19753 659
rect 11495 585 11635 601
rect 11495 551 11511 585
rect 11619 551 11635 585
rect 11495 504 11635 551
rect 11693 585 11833 601
rect 11693 551 11709 585
rect 11817 551 11833 585
rect 11693 504 11833 551
rect 11891 585 12031 601
rect 11891 551 11907 585
rect 12015 551 12031 585
rect 11891 504 12031 551
rect 12089 585 12229 601
rect 12089 551 12105 585
rect 12213 551 12229 585
rect 12089 504 12229 551
rect 12287 585 12427 601
rect 12287 551 12303 585
rect 12411 551 12427 585
rect 12287 504 12427 551
rect 12485 585 12625 601
rect 12485 551 12501 585
rect 12609 551 12625 585
rect 12485 504 12625 551
rect 12683 585 12823 601
rect 12683 551 12699 585
rect 12807 551 12823 585
rect 12683 504 12823 551
rect 12881 585 13021 601
rect 12881 551 12897 585
rect 13005 551 13021 585
rect 12881 504 13021 551
rect 13079 585 13219 601
rect 13079 551 13095 585
rect 13203 551 13219 585
rect 13079 504 13219 551
rect 13277 585 13417 601
rect 13277 551 13293 585
rect 13401 551 13417 585
rect 13277 504 13417 551
rect 13475 585 13615 601
rect 13475 551 13491 585
rect 13599 551 13615 585
rect 13475 504 13615 551
rect 13673 585 13813 601
rect 13673 551 13689 585
rect 13797 551 13813 585
rect 13673 504 13813 551
rect 13871 585 14011 601
rect 13871 551 13887 585
rect 13995 551 14011 585
rect 13871 504 14011 551
rect 14069 585 14209 601
rect 14069 551 14085 585
rect 14193 551 14209 585
rect 14069 504 14209 551
rect 14267 585 14407 601
rect 14267 551 14283 585
rect 14391 551 14407 585
rect 14267 504 14407 551
rect 14465 585 14605 601
rect 14465 551 14481 585
rect 14589 551 14605 585
rect 14465 504 14605 551
rect 14663 585 14803 601
rect 14663 551 14679 585
rect 14787 551 14803 585
rect 14663 504 14803 551
rect 14861 585 15001 601
rect 14861 551 14877 585
rect 14985 551 15001 585
rect 14861 504 15001 551
rect 15059 585 15199 601
rect 15059 551 15075 585
rect 15183 551 15199 585
rect 15059 504 15199 551
rect 15257 585 15397 601
rect 15257 551 15273 585
rect 15381 551 15397 585
rect 15257 504 15397 551
rect 15455 585 15595 601
rect 15455 551 15471 585
rect 15579 551 15595 585
rect 15455 504 15595 551
rect 15653 585 15793 601
rect 15653 551 15669 585
rect 15777 551 15793 585
rect 15653 504 15793 551
rect 15851 585 15991 601
rect 15851 551 15867 585
rect 15975 551 15991 585
rect 15851 504 15991 551
rect 16049 585 16189 601
rect 16049 551 16065 585
rect 16173 551 16189 585
rect 16049 504 16189 551
rect 16247 585 16387 601
rect 16247 551 16263 585
rect 16371 551 16387 585
rect 16247 504 16387 551
rect 16445 585 16585 601
rect 16445 551 16461 585
rect 16569 551 16585 585
rect 16445 504 16585 551
rect 16643 585 16783 601
rect 16643 551 16659 585
rect 16767 551 16783 585
rect 16643 504 16783 551
rect 16841 585 16981 601
rect 16841 551 16857 585
rect 16965 551 16981 585
rect 16841 504 16981 551
rect 17039 585 17179 601
rect 17039 551 17055 585
rect 17163 551 17179 585
rect 17039 504 17179 551
rect 17237 585 17377 601
rect 17237 551 17253 585
rect 17361 551 17377 585
rect 17237 504 17377 551
rect 17435 585 17575 601
rect 17435 551 17451 585
rect 17559 551 17575 585
rect 17435 504 17575 551
rect 17633 585 17773 601
rect 17633 551 17649 585
rect 17757 551 17773 585
rect 17633 504 17773 551
rect 17831 585 17971 601
rect 17831 551 17847 585
rect 17955 551 17971 585
rect 17831 504 17971 551
rect 18029 585 18169 601
rect 18029 551 18045 585
rect 18153 551 18169 585
rect 18029 504 18169 551
rect 18227 585 18367 601
rect 18227 551 18243 585
rect 18351 551 18367 585
rect 18227 504 18367 551
rect 18425 585 18565 601
rect 18425 551 18441 585
rect 18549 551 18565 585
rect 18425 504 18565 551
rect 18623 585 18763 601
rect 18623 551 18639 585
rect 18747 551 18763 585
rect 18623 504 18763 551
rect 18821 585 18961 601
rect 18821 551 18837 585
rect 18945 551 18961 585
rect 18821 504 18961 551
rect 19019 585 19159 601
rect 19019 551 19035 585
rect 19143 551 19159 585
rect 19019 504 19159 551
rect 19217 585 19357 601
rect 19217 551 19233 585
rect 19341 551 19357 585
rect 19217 504 19357 551
rect 19415 585 19555 601
rect 19415 551 19431 585
rect 19539 551 19555 585
rect 19415 504 19555 551
rect 19613 585 19753 601
rect 19613 551 19629 585
rect 19737 551 19753 585
rect 19613 504 19753 551
rect 11495 -943 11635 -896
rect 11495 -977 11511 -943
rect 11619 -977 11635 -943
rect 11495 -993 11635 -977
rect 11693 -943 11833 -896
rect 11693 -977 11709 -943
rect 11817 -977 11833 -943
rect 11693 -993 11833 -977
rect 11891 -943 12031 -896
rect 11891 -977 11907 -943
rect 12015 -977 12031 -943
rect 11891 -993 12031 -977
rect 12089 -943 12229 -896
rect 12089 -977 12105 -943
rect 12213 -977 12229 -943
rect 12089 -993 12229 -977
rect 12287 -943 12427 -896
rect 12287 -977 12303 -943
rect 12411 -977 12427 -943
rect 12287 -993 12427 -977
rect 12485 -943 12625 -896
rect 12485 -977 12501 -943
rect 12609 -977 12625 -943
rect 12485 -993 12625 -977
rect 12683 -943 12823 -896
rect 12683 -977 12699 -943
rect 12807 -977 12823 -943
rect 12683 -993 12823 -977
rect 12881 -943 13021 -896
rect 12881 -977 12897 -943
rect 13005 -977 13021 -943
rect 12881 -993 13021 -977
rect 13079 -943 13219 -896
rect 13079 -977 13095 -943
rect 13203 -977 13219 -943
rect 13079 -993 13219 -977
rect 13277 -943 13417 -896
rect 13277 -977 13293 -943
rect 13401 -977 13417 -943
rect 13277 -993 13417 -977
rect 13475 -943 13615 -896
rect 13475 -977 13491 -943
rect 13599 -977 13615 -943
rect 13475 -993 13615 -977
rect 13673 -943 13813 -896
rect 13673 -977 13689 -943
rect 13797 -977 13813 -943
rect 13673 -993 13813 -977
rect 13871 -943 14011 -896
rect 13871 -977 13887 -943
rect 13995 -977 14011 -943
rect 13871 -993 14011 -977
rect 14069 -943 14209 -896
rect 14069 -977 14085 -943
rect 14193 -977 14209 -943
rect 14069 -993 14209 -977
rect 14267 -943 14407 -896
rect 14267 -977 14283 -943
rect 14391 -977 14407 -943
rect 14267 -993 14407 -977
rect 14465 -943 14605 -896
rect 14465 -977 14481 -943
rect 14589 -977 14605 -943
rect 14465 -993 14605 -977
rect 14663 -943 14803 -896
rect 14663 -977 14679 -943
rect 14787 -977 14803 -943
rect 14663 -993 14803 -977
rect 14861 -943 15001 -896
rect 14861 -977 14877 -943
rect 14985 -977 15001 -943
rect 14861 -993 15001 -977
rect 15059 -943 15199 -896
rect 15059 -977 15075 -943
rect 15183 -977 15199 -943
rect 15059 -993 15199 -977
rect 15257 -943 15397 -896
rect 15257 -977 15273 -943
rect 15381 -977 15397 -943
rect 15257 -993 15397 -977
rect 15455 -943 15595 -896
rect 15455 -977 15471 -943
rect 15579 -977 15595 -943
rect 15455 -993 15595 -977
rect 15653 -943 15793 -896
rect 15653 -977 15669 -943
rect 15777 -977 15793 -943
rect 15653 -993 15793 -977
rect 15851 -943 15991 -896
rect 15851 -977 15867 -943
rect 15975 -977 15991 -943
rect 15851 -993 15991 -977
rect 16049 -943 16189 -896
rect 16049 -977 16065 -943
rect 16173 -977 16189 -943
rect 16049 -993 16189 -977
rect 16247 -943 16387 -896
rect 16247 -977 16263 -943
rect 16371 -977 16387 -943
rect 16247 -993 16387 -977
rect 16445 -943 16585 -896
rect 16445 -977 16461 -943
rect 16569 -977 16585 -943
rect 16445 -993 16585 -977
rect 16643 -943 16783 -896
rect 16643 -977 16659 -943
rect 16767 -977 16783 -943
rect 16643 -993 16783 -977
rect 16841 -943 16981 -896
rect 16841 -977 16857 -943
rect 16965 -977 16981 -943
rect 16841 -993 16981 -977
rect 17039 -943 17179 -896
rect 17039 -977 17055 -943
rect 17163 -977 17179 -943
rect 17039 -993 17179 -977
rect 17237 -943 17377 -896
rect 17237 -977 17253 -943
rect 17361 -977 17377 -943
rect 17237 -993 17377 -977
rect 17435 -943 17575 -896
rect 17435 -977 17451 -943
rect 17559 -977 17575 -943
rect 17435 -993 17575 -977
rect 17633 -943 17773 -896
rect 17633 -977 17649 -943
rect 17757 -977 17773 -943
rect 17633 -993 17773 -977
rect 17831 -943 17971 -896
rect 17831 -977 17847 -943
rect 17955 -977 17971 -943
rect 17831 -993 17971 -977
rect 18029 -943 18169 -896
rect 18029 -977 18045 -943
rect 18153 -977 18169 -943
rect 18029 -993 18169 -977
rect 18227 -943 18367 -896
rect 18227 -977 18243 -943
rect 18351 -977 18367 -943
rect 18227 -993 18367 -977
rect 18425 -943 18565 -896
rect 18425 -977 18441 -943
rect 18549 -977 18565 -943
rect 18425 -993 18565 -977
rect 18623 -943 18763 -896
rect 18623 -977 18639 -943
rect 18747 -977 18763 -943
rect 18623 -993 18763 -977
rect 18821 -943 18961 -896
rect 18821 -977 18837 -943
rect 18945 -977 18961 -943
rect 18821 -993 18961 -977
rect 19019 -943 19159 -896
rect 19019 -977 19035 -943
rect 19143 -977 19159 -943
rect 19019 -993 19159 -977
rect 19217 -943 19357 -896
rect 19217 -977 19233 -943
rect 19341 -977 19357 -943
rect 19217 -993 19357 -977
rect 19415 -943 19555 -896
rect 19415 -977 19431 -943
rect 19539 -977 19555 -943
rect 19415 -993 19555 -977
rect 19613 -943 19753 -896
rect 19613 -977 19629 -943
rect 19737 -977 19753 -943
rect 19613 -993 19753 -977
rect 11495 -1051 11635 -1035
rect 11495 -1085 11511 -1051
rect 11619 -1085 11635 -1051
rect 11495 -1132 11635 -1085
rect 11693 -1051 11833 -1035
rect 11693 -1085 11709 -1051
rect 11817 -1085 11833 -1051
rect 11693 -1132 11833 -1085
rect 11891 -1051 12031 -1035
rect 11891 -1085 11907 -1051
rect 12015 -1085 12031 -1051
rect 11891 -1132 12031 -1085
rect 12089 -1051 12229 -1035
rect 12089 -1085 12105 -1051
rect 12213 -1085 12229 -1051
rect 12089 -1132 12229 -1085
rect 12287 -1051 12427 -1035
rect 12287 -1085 12303 -1051
rect 12411 -1085 12427 -1051
rect 12287 -1132 12427 -1085
rect 12485 -1051 12625 -1035
rect 12485 -1085 12501 -1051
rect 12609 -1085 12625 -1051
rect 12485 -1132 12625 -1085
rect 12683 -1051 12823 -1035
rect 12683 -1085 12699 -1051
rect 12807 -1085 12823 -1051
rect 12683 -1132 12823 -1085
rect 12881 -1051 13021 -1035
rect 12881 -1085 12897 -1051
rect 13005 -1085 13021 -1051
rect 12881 -1132 13021 -1085
rect 13079 -1051 13219 -1035
rect 13079 -1085 13095 -1051
rect 13203 -1085 13219 -1051
rect 13079 -1132 13219 -1085
rect 13277 -1051 13417 -1035
rect 13277 -1085 13293 -1051
rect 13401 -1085 13417 -1051
rect 13277 -1132 13417 -1085
rect 13475 -1051 13615 -1035
rect 13475 -1085 13491 -1051
rect 13599 -1085 13615 -1051
rect 13475 -1132 13615 -1085
rect 13673 -1051 13813 -1035
rect 13673 -1085 13689 -1051
rect 13797 -1085 13813 -1051
rect 13673 -1132 13813 -1085
rect 13871 -1051 14011 -1035
rect 13871 -1085 13887 -1051
rect 13995 -1085 14011 -1051
rect 13871 -1132 14011 -1085
rect 14069 -1051 14209 -1035
rect 14069 -1085 14085 -1051
rect 14193 -1085 14209 -1051
rect 14069 -1132 14209 -1085
rect 14267 -1051 14407 -1035
rect 14267 -1085 14283 -1051
rect 14391 -1085 14407 -1051
rect 14267 -1132 14407 -1085
rect 14465 -1051 14605 -1035
rect 14465 -1085 14481 -1051
rect 14589 -1085 14605 -1051
rect 14465 -1132 14605 -1085
rect 14663 -1051 14803 -1035
rect 14663 -1085 14679 -1051
rect 14787 -1085 14803 -1051
rect 14663 -1132 14803 -1085
rect 14861 -1051 15001 -1035
rect 14861 -1085 14877 -1051
rect 14985 -1085 15001 -1051
rect 14861 -1132 15001 -1085
rect 15059 -1051 15199 -1035
rect 15059 -1085 15075 -1051
rect 15183 -1085 15199 -1051
rect 15059 -1132 15199 -1085
rect 15257 -1051 15397 -1035
rect 15257 -1085 15273 -1051
rect 15381 -1085 15397 -1051
rect 15257 -1132 15397 -1085
rect 15455 -1051 15595 -1035
rect 15455 -1085 15471 -1051
rect 15579 -1085 15595 -1051
rect 15455 -1132 15595 -1085
rect 15653 -1051 15793 -1035
rect 15653 -1085 15669 -1051
rect 15777 -1085 15793 -1051
rect 15653 -1132 15793 -1085
rect 15851 -1051 15991 -1035
rect 15851 -1085 15867 -1051
rect 15975 -1085 15991 -1051
rect 15851 -1132 15991 -1085
rect 16049 -1051 16189 -1035
rect 16049 -1085 16065 -1051
rect 16173 -1085 16189 -1051
rect 16049 -1132 16189 -1085
rect 16247 -1051 16387 -1035
rect 16247 -1085 16263 -1051
rect 16371 -1085 16387 -1051
rect 16247 -1132 16387 -1085
rect 16445 -1051 16585 -1035
rect 16445 -1085 16461 -1051
rect 16569 -1085 16585 -1051
rect 16445 -1132 16585 -1085
rect 16643 -1051 16783 -1035
rect 16643 -1085 16659 -1051
rect 16767 -1085 16783 -1051
rect 16643 -1132 16783 -1085
rect 16841 -1051 16981 -1035
rect 16841 -1085 16857 -1051
rect 16965 -1085 16981 -1051
rect 16841 -1132 16981 -1085
rect 17039 -1051 17179 -1035
rect 17039 -1085 17055 -1051
rect 17163 -1085 17179 -1051
rect 17039 -1132 17179 -1085
rect 17237 -1051 17377 -1035
rect 17237 -1085 17253 -1051
rect 17361 -1085 17377 -1051
rect 17237 -1132 17377 -1085
rect 17435 -1051 17575 -1035
rect 17435 -1085 17451 -1051
rect 17559 -1085 17575 -1051
rect 17435 -1132 17575 -1085
rect 17633 -1051 17773 -1035
rect 17633 -1085 17649 -1051
rect 17757 -1085 17773 -1051
rect 17633 -1132 17773 -1085
rect 17831 -1051 17971 -1035
rect 17831 -1085 17847 -1051
rect 17955 -1085 17971 -1051
rect 17831 -1132 17971 -1085
rect 18029 -1051 18169 -1035
rect 18029 -1085 18045 -1051
rect 18153 -1085 18169 -1051
rect 18029 -1132 18169 -1085
rect 18227 -1051 18367 -1035
rect 18227 -1085 18243 -1051
rect 18351 -1085 18367 -1051
rect 18227 -1132 18367 -1085
rect 18425 -1051 18565 -1035
rect 18425 -1085 18441 -1051
rect 18549 -1085 18565 -1051
rect 18425 -1132 18565 -1085
rect 18623 -1051 18763 -1035
rect 18623 -1085 18639 -1051
rect 18747 -1085 18763 -1051
rect 18623 -1132 18763 -1085
rect 18821 -1051 18961 -1035
rect 18821 -1085 18837 -1051
rect 18945 -1085 18961 -1051
rect 18821 -1132 18961 -1085
rect 19019 -1051 19159 -1035
rect 19019 -1085 19035 -1051
rect 19143 -1085 19159 -1051
rect 19019 -1132 19159 -1085
rect 19217 -1051 19357 -1035
rect 19217 -1085 19233 -1051
rect 19341 -1085 19357 -1051
rect 19217 -1132 19357 -1085
rect 19415 -1051 19555 -1035
rect 19415 -1085 19431 -1051
rect 19539 -1085 19555 -1051
rect 19415 -1132 19555 -1085
rect 19613 -1051 19753 -1035
rect 19613 -1085 19629 -1051
rect 19737 -1085 19753 -1051
rect 19613 -1132 19753 -1085
rect 11495 -2579 11635 -2532
rect 11495 -2613 11511 -2579
rect 11619 -2613 11635 -2579
rect 11495 -2629 11635 -2613
rect 11693 -2579 11833 -2532
rect 11693 -2613 11709 -2579
rect 11817 -2613 11833 -2579
rect 11693 -2629 11833 -2613
rect 11891 -2579 12031 -2532
rect 11891 -2613 11907 -2579
rect 12015 -2613 12031 -2579
rect 11891 -2629 12031 -2613
rect 12089 -2579 12229 -2532
rect 12089 -2613 12105 -2579
rect 12213 -2613 12229 -2579
rect 12089 -2629 12229 -2613
rect 12287 -2579 12427 -2532
rect 12287 -2613 12303 -2579
rect 12411 -2613 12427 -2579
rect 12287 -2629 12427 -2613
rect 12485 -2579 12625 -2532
rect 12485 -2613 12501 -2579
rect 12609 -2613 12625 -2579
rect 12485 -2629 12625 -2613
rect 12683 -2579 12823 -2532
rect 12683 -2613 12699 -2579
rect 12807 -2613 12823 -2579
rect 12683 -2629 12823 -2613
rect 12881 -2579 13021 -2532
rect 12881 -2613 12897 -2579
rect 13005 -2613 13021 -2579
rect 12881 -2629 13021 -2613
rect 13079 -2579 13219 -2532
rect 13079 -2613 13095 -2579
rect 13203 -2613 13219 -2579
rect 13079 -2629 13219 -2613
rect 13277 -2579 13417 -2532
rect 13277 -2613 13293 -2579
rect 13401 -2613 13417 -2579
rect 13277 -2629 13417 -2613
rect 13475 -2579 13615 -2532
rect 13475 -2613 13491 -2579
rect 13599 -2613 13615 -2579
rect 13475 -2629 13615 -2613
rect 13673 -2579 13813 -2532
rect 13673 -2613 13689 -2579
rect 13797 -2613 13813 -2579
rect 13673 -2629 13813 -2613
rect 13871 -2579 14011 -2532
rect 13871 -2613 13887 -2579
rect 13995 -2613 14011 -2579
rect 13871 -2629 14011 -2613
rect 14069 -2579 14209 -2532
rect 14069 -2613 14085 -2579
rect 14193 -2613 14209 -2579
rect 14069 -2629 14209 -2613
rect 14267 -2579 14407 -2532
rect 14267 -2613 14283 -2579
rect 14391 -2613 14407 -2579
rect 14267 -2629 14407 -2613
rect 14465 -2579 14605 -2532
rect 14465 -2613 14481 -2579
rect 14589 -2613 14605 -2579
rect 14465 -2629 14605 -2613
rect 14663 -2579 14803 -2532
rect 14663 -2613 14679 -2579
rect 14787 -2613 14803 -2579
rect 14663 -2629 14803 -2613
rect 14861 -2579 15001 -2532
rect 14861 -2613 14877 -2579
rect 14985 -2613 15001 -2579
rect 14861 -2629 15001 -2613
rect 15059 -2579 15199 -2532
rect 15059 -2613 15075 -2579
rect 15183 -2613 15199 -2579
rect 15059 -2629 15199 -2613
rect 15257 -2579 15397 -2532
rect 15257 -2613 15273 -2579
rect 15381 -2613 15397 -2579
rect 15257 -2629 15397 -2613
rect 15455 -2579 15595 -2532
rect 15455 -2613 15471 -2579
rect 15579 -2613 15595 -2579
rect 15455 -2629 15595 -2613
rect 15653 -2579 15793 -2532
rect 15653 -2613 15669 -2579
rect 15777 -2613 15793 -2579
rect 15653 -2629 15793 -2613
rect 15851 -2579 15991 -2532
rect 15851 -2613 15867 -2579
rect 15975 -2613 15991 -2579
rect 15851 -2629 15991 -2613
rect 16049 -2579 16189 -2532
rect 16049 -2613 16065 -2579
rect 16173 -2613 16189 -2579
rect 16049 -2629 16189 -2613
rect 16247 -2579 16387 -2532
rect 16247 -2613 16263 -2579
rect 16371 -2613 16387 -2579
rect 16247 -2629 16387 -2613
rect 16445 -2579 16585 -2532
rect 16445 -2613 16461 -2579
rect 16569 -2613 16585 -2579
rect 16445 -2629 16585 -2613
rect 16643 -2579 16783 -2532
rect 16643 -2613 16659 -2579
rect 16767 -2613 16783 -2579
rect 16643 -2629 16783 -2613
rect 16841 -2579 16981 -2532
rect 16841 -2613 16857 -2579
rect 16965 -2613 16981 -2579
rect 16841 -2629 16981 -2613
rect 17039 -2579 17179 -2532
rect 17039 -2613 17055 -2579
rect 17163 -2613 17179 -2579
rect 17039 -2629 17179 -2613
rect 17237 -2579 17377 -2532
rect 17237 -2613 17253 -2579
rect 17361 -2613 17377 -2579
rect 17237 -2629 17377 -2613
rect 17435 -2579 17575 -2532
rect 17435 -2613 17451 -2579
rect 17559 -2613 17575 -2579
rect 17435 -2629 17575 -2613
rect 17633 -2579 17773 -2532
rect 17633 -2613 17649 -2579
rect 17757 -2613 17773 -2579
rect 17633 -2629 17773 -2613
rect 17831 -2579 17971 -2532
rect 17831 -2613 17847 -2579
rect 17955 -2613 17971 -2579
rect 17831 -2629 17971 -2613
rect 18029 -2579 18169 -2532
rect 18029 -2613 18045 -2579
rect 18153 -2613 18169 -2579
rect 18029 -2629 18169 -2613
rect 18227 -2579 18367 -2532
rect 18227 -2613 18243 -2579
rect 18351 -2613 18367 -2579
rect 18227 -2629 18367 -2613
rect 18425 -2579 18565 -2532
rect 18425 -2613 18441 -2579
rect 18549 -2613 18565 -2579
rect 18425 -2629 18565 -2613
rect 18623 -2579 18763 -2532
rect 18623 -2613 18639 -2579
rect 18747 -2613 18763 -2579
rect 18623 -2629 18763 -2613
rect 18821 -2579 18961 -2532
rect 18821 -2613 18837 -2579
rect 18945 -2613 18961 -2579
rect 18821 -2629 18961 -2613
rect 19019 -2579 19159 -2532
rect 19019 -2613 19035 -2579
rect 19143 -2613 19159 -2579
rect 19019 -2629 19159 -2613
rect 19217 -2579 19357 -2532
rect 19217 -2613 19233 -2579
rect 19341 -2613 19357 -2579
rect 19217 -2629 19357 -2613
rect 19415 -2579 19555 -2532
rect 19415 -2613 19431 -2579
rect 19539 -2613 19555 -2579
rect 19415 -2629 19555 -2613
rect 19613 -2579 19753 -2532
rect 19613 -2613 19629 -2579
rect 19737 -2613 19753 -2579
rect 19613 -2629 19753 -2613
rect 11495 -2687 11635 -2671
rect 11495 -2721 11511 -2687
rect 11619 -2721 11635 -2687
rect 11495 -2768 11635 -2721
rect 11693 -2687 11833 -2671
rect 11693 -2721 11709 -2687
rect 11817 -2721 11833 -2687
rect 11693 -2768 11833 -2721
rect 11891 -2687 12031 -2671
rect 11891 -2721 11907 -2687
rect 12015 -2721 12031 -2687
rect 11891 -2768 12031 -2721
rect 12089 -2687 12229 -2671
rect 12089 -2721 12105 -2687
rect 12213 -2721 12229 -2687
rect 12089 -2768 12229 -2721
rect 12287 -2687 12427 -2671
rect 12287 -2721 12303 -2687
rect 12411 -2721 12427 -2687
rect 12287 -2768 12427 -2721
rect 12485 -2687 12625 -2671
rect 12485 -2721 12501 -2687
rect 12609 -2721 12625 -2687
rect 12485 -2768 12625 -2721
rect 12683 -2687 12823 -2671
rect 12683 -2721 12699 -2687
rect 12807 -2721 12823 -2687
rect 12683 -2768 12823 -2721
rect 12881 -2687 13021 -2671
rect 12881 -2721 12897 -2687
rect 13005 -2721 13021 -2687
rect 12881 -2768 13021 -2721
rect 13079 -2687 13219 -2671
rect 13079 -2721 13095 -2687
rect 13203 -2721 13219 -2687
rect 13079 -2768 13219 -2721
rect 13277 -2687 13417 -2671
rect 13277 -2721 13293 -2687
rect 13401 -2721 13417 -2687
rect 13277 -2768 13417 -2721
rect 13475 -2687 13615 -2671
rect 13475 -2721 13491 -2687
rect 13599 -2721 13615 -2687
rect 13475 -2768 13615 -2721
rect 13673 -2687 13813 -2671
rect 13673 -2721 13689 -2687
rect 13797 -2721 13813 -2687
rect 13673 -2768 13813 -2721
rect 13871 -2687 14011 -2671
rect 13871 -2721 13887 -2687
rect 13995 -2721 14011 -2687
rect 13871 -2768 14011 -2721
rect 14069 -2687 14209 -2671
rect 14069 -2721 14085 -2687
rect 14193 -2721 14209 -2687
rect 14069 -2768 14209 -2721
rect 14267 -2687 14407 -2671
rect 14267 -2721 14283 -2687
rect 14391 -2721 14407 -2687
rect 14267 -2768 14407 -2721
rect 14465 -2687 14605 -2671
rect 14465 -2721 14481 -2687
rect 14589 -2721 14605 -2687
rect 14465 -2768 14605 -2721
rect 14663 -2687 14803 -2671
rect 14663 -2721 14679 -2687
rect 14787 -2721 14803 -2687
rect 14663 -2768 14803 -2721
rect 14861 -2687 15001 -2671
rect 14861 -2721 14877 -2687
rect 14985 -2721 15001 -2687
rect 14861 -2768 15001 -2721
rect 15059 -2687 15199 -2671
rect 15059 -2721 15075 -2687
rect 15183 -2721 15199 -2687
rect 15059 -2768 15199 -2721
rect 15257 -2687 15397 -2671
rect 15257 -2721 15273 -2687
rect 15381 -2721 15397 -2687
rect 15257 -2768 15397 -2721
rect 15455 -2687 15595 -2671
rect 15455 -2721 15471 -2687
rect 15579 -2721 15595 -2687
rect 15455 -2768 15595 -2721
rect 15653 -2687 15793 -2671
rect 15653 -2721 15669 -2687
rect 15777 -2721 15793 -2687
rect 15653 -2768 15793 -2721
rect 15851 -2687 15991 -2671
rect 15851 -2721 15867 -2687
rect 15975 -2721 15991 -2687
rect 15851 -2768 15991 -2721
rect 16049 -2687 16189 -2671
rect 16049 -2721 16065 -2687
rect 16173 -2721 16189 -2687
rect 16049 -2768 16189 -2721
rect 16247 -2687 16387 -2671
rect 16247 -2721 16263 -2687
rect 16371 -2721 16387 -2687
rect 16247 -2768 16387 -2721
rect 16445 -2687 16585 -2671
rect 16445 -2721 16461 -2687
rect 16569 -2721 16585 -2687
rect 16445 -2768 16585 -2721
rect 16643 -2687 16783 -2671
rect 16643 -2721 16659 -2687
rect 16767 -2721 16783 -2687
rect 16643 -2768 16783 -2721
rect 16841 -2687 16981 -2671
rect 16841 -2721 16857 -2687
rect 16965 -2721 16981 -2687
rect 16841 -2768 16981 -2721
rect 17039 -2687 17179 -2671
rect 17039 -2721 17055 -2687
rect 17163 -2721 17179 -2687
rect 17039 -2768 17179 -2721
rect 17237 -2687 17377 -2671
rect 17237 -2721 17253 -2687
rect 17361 -2721 17377 -2687
rect 17237 -2768 17377 -2721
rect 17435 -2687 17575 -2671
rect 17435 -2721 17451 -2687
rect 17559 -2721 17575 -2687
rect 17435 -2768 17575 -2721
rect 17633 -2687 17773 -2671
rect 17633 -2721 17649 -2687
rect 17757 -2721 17773 -2687
rect 17633 -2768 17773 -2721
rect 17831 -2687 17971 -2671
rect 17831 -2721 17847 -2687
rect 17955 -2721 17971 -2687
rect 17831 -2768 17971 -2721
rect 18029 -2687 18169 -2671
rect 18029 -2721 18045 -2687
rect 18153 -2721 18169 -2687
rect 18029 -2768 18169 -2721
rect 18227 -2687 18367 -2671
rect 18227 -2721 18243 -2687
rect 18351 -2721 18367 -2687
rect 18227 -2768 18367 -2721
rect 18425 -2687 18565 -2671
rect 18425 -2721 18441 -2687
rect 18549 -2721 18565 -2687
rect 18425 -2768 18565 -2721
rect 18623 -2687 18763 -2671
rect 18623 -2721 18639 -2687
rect 18747 -2721 18763 -2687
rect 18623 -2768 18763 -2721
rect 18821 -2687 18961 -2671
rect 18821 -2721 18837 -2687
rect 18945 -2721 18961 -2687
rect 18821 -2768 18961 -2721
rect 19019 -2687 19159 -2671
rect 19019 -2721 19035 -2687
rect 19143 -2721 19159 -2687
rect 19019 -2768 19159 -2721
rect 19217 -2687 19357 -2671
rect 19217 -2721 19233 -2687
rect 19341 -2721 19357 -2687
rect 19217 -2768 19357 -2721
rect 19415 -2687 19555 -2671
rect 19415 -2721 19431 -2687
rect 19539 -2721 19555 -2687
rect 19415 -2768 19555 -2721
rect 19613 -2687 19753 -2671
rect 19613 -2721 19629 -2687
rect 19737 -2721 19753 -2687
rect 19613 -2768 19753 -2721
rect 11495 -4194 11635 -4168
rect 11693 -4194 11833 -4168
rect 11891 -4194 12031 -4168
rect 12089 -4194 12229 -4168
rect 12287 -4194 12427 -4168
rect 12485 -4194 12625 -4168
rect 12683 -4194 12823 -4168
rect 12881 -4194 13021 -4168
rect 13079 -4194 13219 -4168
rect 13277 -4194 13417 -4168
rect 13475 -4194 13615 -4168
rect 13673 -4194 13813 -4168
rect 13871 -4194 14011 -4168
rect 14069 -4194 14209 -4168
rect 14267 -4194 14407 -4168
rect 14465 -4194 14605 -4168
rect 14663 -4194 14803 -4168
rect 14861 -4194 15001 -4168
rect 15059 -4194 15199 -4168
rect 15257 -4194 15397 -4168
rect 15455 -4194 15595 -4168
rect 15653 -4194 15793 -4168
rect 15851 -4194 15991 -4168
rect 16049 -4194 16189 -4168
rect 16247 -4194 16387 -4168
rect 16445 -4194 16585 -4168
rect 16643 -4194 16783 -4168
rect 16841 -4194 16981 -4168
rect 17039 -4194 17179 -4168
rect 17237 -4194 17377 -4168
rect 17435 -4194 17575 -4168
rect 17633 -4194 17773 -4168
rect 17831 -4194 17971 -4168
rect 18029 -4194 18169 -4168
rect 18227 -4194 18367 -4168
rect 18425 -4194 18565 -4168
rect 18623 -4194 18763 -4168
rect 18821 -4194 18961 -4168
rect 19019 -4194 19159 -4168
rect 19217 -4194 19357 -4168
rect 19415 -4194 19555 -4168
rect 19613 -4194 19753 -4168
rect 23345 2140 23485 2166
rect 23543 2140 23683 2166
rect 23741 2140 23881 2166
rect 23939 2140 24079 2166
rect 24137 2140 24277 2166
rect 24335 2140 24475 2166
rect 24533 2140 24673 2166
rect 24731 2140 24871 2166
rect 24929 2140 25069 2166
rect 25127 2140 25267 2166
rect 25325 2140 25465 2166
rect 25523 2140 25663 2166
rect 25721 2140 25861 2166
rect 25919 2140 26059 2166
rect 26117 2140 26257 2166
rect 26315 2140 26455 2166
rect 26513 2140 26653 2166
rect 26711 2140 26851 2166
rect 26909 2140 27049 2166
rect 27107 2140 27247 2166
rect 27305 2140 27445 2166
rect 27503 2140 27643 2166
rect 27701 2140 27841 2166
rect 27899 2140 28039 2166
rect 28097 2140 28237 2166
rect 28295 2140 28435 2166
rect 28493 2140 28633 2166
rect 28691 2140 28831 2166
rect 28889 2140 29029 2166
rect 29087 2140 29227 2166
rect 29285 2140 29425 2166
rect 29483 2140 29623 2166
rect 29681 2140 29821 2166
rect 29879 2140 30019 2166
rect 30077 2140 30217 2166
rect 30275 2140 30415 2166
rect 30473 2140 30613 2166
rect 30671 2140 30811 2166
rect 30869 2140 31009 2166
rect 31067 2140 31207 2166
rect 31265 2140 31405 2166
rect 31463 2140 31603 2166
rect 23345 693 23485 740
rect 23345 659 23361 693
rect 23469 659 23485 693
rect 23345 643 23485 659
rect 23543 693 23683 740
rect 23543 659 23559 693
rect 23667 659 23683 693
rect 23543 643 23683 659
rect 23741 693 23881 740
rect 23741 659 23757 693
rect 23865 659 23881 693
rect 23741 643 23881 659
rect 23939 693 24079 740
rect 23939 659 23955 693
rect 24063 659 24079 693
rect 23939 643 24079 659
rect 24137 693 24277 740
rect 24137 659 24153 693
rect 24261 659 24277 693
rect 24137 643 24277 659
rect 24335 693 24475 740
rect 24335 659 24351 693
rect 24459 659 24475 693
rect 24335 643 24475 659
rect 24533 693 24673 740
rect 24533 659 24549 693
rect 24657 659 24673 693
rect 24533 643 24673 659
rect 24731 693 24871 740
rect 24731 659 24747 693
rect 24855 659 24871 693
rect 24731 643 24871 659
rect 24929 693 25069 740
rect 24929 659 24945 693
rect 25053 659 25069 693
rect 24929 643 25069 659
rect 25127 693 25267 740
rect 25127 659 25143 693
rect 25251 659 25267 693
rect 25127 643 25267 659
rect 25325 693 25465 740
rect 25325 659 25341 693
rect 25449 659 25465 693
rect 25325 643 25465 659
rect 25523 693 25663 740
rect 25523 659 25539 693
rect 25647 659 25663 693
rect 25523 643 25663 659
rect 25721 693 25861 740
rect 25721 659 25737 693
rect 25845 659 25861 693
rect 25721 643 25861 659
rect 25919 693 26059 740
rect 25919 659 25935 693
rect 26043 659 26059 693
rect 25919 643 26059 659
rect 26117 693 26257 740
rect 26117 659 26133 693
rect 26241 659 26257 693
rect 26117 643 26257 659
rect 26315 693 26455 740
rect 26315 659 26331 693
rect 26439 659 26455 693
rect 26315 643 26455 659
rect 26513 693 26653 740
rect 26513 659 26529 693
rect 26637 659 26653 693
rect 26513 643 26653 659
rect 26711 693 26851 740
rect 26711 659 26727 693
rect 26835 659 26851 693
rect 26711 643 26851 659
rect 26909 693 27049 740
rect 26909 659 26925 693
rect 27033 659 27049 693
rect 26909 643 27049 659
rect 27107 693 27247 740
rect 27107 659 27123 693
rect 27231 659 27247 693
rect 27107 643 27247 659
rect 27305 693 27445 740
rect 27305 659 27321 693
rect 27429 659 27445 693
rect 27305 643 27445 659
rect 27503 693 27643 740
rect 27503 659 27519 693
rect 27627 659 27643 693
rect 27503 643 27643 659
rect 27701 693 27841 740
rect 27701 659 27717 693
rect 27825 659 27841 693
rect 27701 643 27841 659
rect 27899 693 28039 740
rect 27899 659 27915 693
rect 28023 659 28039 693
rect 27899 643 28039 659
rect 28097 693 28237 740
rect 28097 659 28113 693
rect 28221 659 28237 693
rect 28097 643 28237 659
rect 28295 693 28435 740
rect 28295 659 28311 693
rect 28419 659 28435 693
rect 28295 643 28435 659
rect 28493 693 28633 740
rect 28493 659 28509 693
rect 28617 659 28633 693
rect 28493 643 28633 659
rect 28691 693 28831 740
rect 28691 659 28707 693
rect 28815 659 28831 693
rect 28691 643 28831 659
rect 28889 693 29029 740
rect 28889 659 28905 693
rect 29013 659 29029 693
rect 28889 643 29029 659
rect 29087 693 29227 740
rect 29087 659 29103 693
rect 29211 659 29227 693
rect 29087 643 29227 659
rect 29285 693 29425 740
rect 29285 659 29301 693
rect 29409 659 29425 693
rect 29285 643 29425 659
rect 29483 693 29623 740
rect 29483 659 29499 693
rect 29607 659 29623 693
rect 29483 643 29623 659
rect 29681 693 29821 740
rect 29681 659 29697 693
rect 29805 659 29821 693
rect 29681 643 29821 659
rect 29879 693 30019 740
rect 29879 659 29895 693
rect 30003 659 30019 693
rect 29879 643 30019 659
rect 30077 693 30217 740
rect 30077 659 30093 693
rect 30201 659 30217 693
rect 30077 643 30217 659
rect 30275 693 30415 740
rect 30275 659 30291 693
rect 30399 659 30415 693
rect 30275 643 30415 659
rect 30473 693 30613 740
rect 30473 659 30489 693
rect 30597 659 30613 693
rect 30473 643 30613 659
rect 30671 693 30811 740
rect 30671 659 30687 693
rect 30795 659 30811 693
rect 30671 643 30811 659
rect 30869 693 31009 740
rect 30869 659 30885 693
rect 30993 659 31009 693
rect 30869 643 31009 659
rect 31067 693 31207 740
rect 31067 659 31083 693
rect 31191 659 31207 693
rect 31067 643 31207 659
rect 31265 693 31405 740
rect 31265 659 31281 693
rect 31389 659 31405 693
rect 31265 643 31405 659
rect 31463 693 31603 740
rect 31463 659 31479 693
rect 31587 659 31603 693
rect 31463 643 31603 659
rect 23345 585 23485 601
rect 23345 551 23361 585
rect 23469 551 23485 585
rect 23345 504 23485 551
rect 23543 585 23683 601
rect 23543 551 23559 585
rect 23667 551 23683 585
rect 23543 504 23683 551
rect 23741 585 23881 601
rect 23741 551 23757 585
rect 23865 551 23881 585
rect 23741 504 23881 551
rect 23939 585 24079 601
rect 23939 551 23955 585
rect 24063 551 24079 585
rect 23939 504 24079 551
rect 24137 585 24277 601
rect 24137 551 24153 585
rect 24261 551 24277 585
rect 24137 504 24277 551
rect 24335 585 24475 601
rect 24335 551 24351 585
rect 24459 551 24475 585
rect 24335 504 24475 551
rect 24533 585 24673 601
rect 24533 551 24549 585
rect 24657 551 24673 585
rect 24533 504 24673 551
rect 24731 585 24871 601
rect 24731 551 24747 585
rect 24855 551 24871 585
rect 24731 504 24871 551
rect 24929 585 25069 601
rect 24929 551 24945 585
rect 25053 551 25069 585
rect 24929 504 25069 551
rect 25127 585 25267 601
rect 25127 551 25143 585
rect 25251 551 25267 585
rect 25127 504 25267 551
rect 25325 585 25465 601
rect 25325 551 25341 585
rect 25449 551 25465 585
rect 25325 504 25465 551
rect 25523 585 25663 601
rect 25523 551 25539 585
rect 25647 551 25663 585
rect 25523 504 25663 551
rect 25721 585 25861 601
rect 25721 551 25737 585
rect 25845 551 25861 585
rect 25721 504 25861 551
rect 25919 585 26059 601
rect 25919 551 25935 585
rect 26043 551 26059 585
rect 25919 504 26059 551
rect 26117 585 26257 601
rect 26117 551 26133 585
rect 26241 551 26257 585
rect 26117 504 26257 551
rect 26315 585 26455 601
rect 26315 551 26331 585
rect 26439 551 26455 585
rect 26315 504 26455 551
rect 26513 585 26653 601
rect 26513 551 26529 585
rect 26637 551 26653 585
rect 26513 504 26653 551
rect 26711 585 26851 601
rect 26711 551 26727 585
rect 26835 551 26851 585
rect 26711 504 26851 551
rect 26909 585 27049 601
rect 26909 551 26925 585
rect 27033 551 27049 585
rect 26909 504 27049 551
rect 27107 585 27247 601
rect 27107 551 27123 585
rect 27231 551 27247 585
rect 27107 504 27247 551
rect 27305 585 27445 601
rect 27305 551 27321 585
rect 27429 551 27445 585
rect 27305 504 27445 551
rect 27503 585 27643 601
rect 27503 551 27519 585
rect 27627 551 27643 585
rect 27503 504 27643 551
rect 27701 585 27841 601
rect 27701 551 27717 585
rect 27825 551 27841 585
rect 27701 504 27841 551
rect 27899 585 28039 601
rect 27899 551 27915 585
rect 28023 551 28039 585
rect 27899 504 28039 551
rect 28097 585 28237 601
rect 28097 551 28113 585
rect 28221 551 28237 585
rect 28097 504 28237 551
rect 28295 585 28435 601
rect 28295 551 28311 585
rect 28419 551 28435 585
rect 28295 504 28435 551
rect 28493 585 28633 601
rect 28493 551 28509 585
rect 28617 551 28633 585
rect 28493 504 28633 551
rect 28691 585 28831 601
rect 28691 551 28707 585
rect 28815 551 28831 585
rect 28691 504 28831 551
rect 28889 585 29029 601
rect 28889 551 28905 585
rect 29013 551 29029 585
rect 28889 504 29029 551
rect 29087 585 29227 601
rect 29087 551 29103 585
rect 29211 551 29227 585
rect 29087 504 29227 551
rect 29285 585 29425 601
rect 29285 551 29301 585
rect 29409 551 29425 585
rect 29285 504 29425 551
rect 29483 585 29623 601
rect 29483 551 29499 585
rect 29607 551 29623 585
rect 29483 504 29623 551
rect 29681 585 29821 601
rect 29681 551 29697 585
rect 29805 551 29821 585
rect 29681 504 29821 551
rect 29879 585 30019 601
rect 29879 551 29895 585
rect 30003 551 30019 585
rect 29879 504 30019 551
rect 30077 585 30217 601
rect 30077 551 30093 585
rect 30201 551 30217 585
rect 30077 504 30217 551
rect 30275 585 30415 601
rect 30275 551 30291 585
rect 30399 551 30415 585
rect 30275 504 30415 551
rect 30473 585 30613 601
rect 30473 551 30489 585
rect 30597 551 30613 585
rect 30473 504 30613 551
rect 30671 585 30811 601
rect 30671 551 30687 585
rect 30795 551 30811 585
rect 30671 504 30811 551
rect 30869 585 31009 601
rect 30869 551 30885 585
rect 30993 551 31009 585
rect 30869 504 31009 551
rect 31067 585 31207 601
rect 31067 551 31083 585
rect 31191 551 31207 585
rect 31067 504 31207 551
rect 31265 585 31405 601
rect 31265 551 31281 585
rect 31389 551 31405 585
rect 31265 504 31405 551
rect 31463 585 31603 601
rect 31463 551 31479 585
rect 31587 551 31603 585
rect 31463 504 31603 551
rect 23345 -943 23485 -896
rect 23345 -977 23361 -943
rect 23469 -977 23485 -943
rect 23345 -993 23485 -977
rect 23543 -943 23683 -896
rect 23543 -977 23559 -943
rect 23667 -977 23683 -943
rect 23543 -993 23683 -977
rect 23741 -943 23881 -896
rect 23741 -977 23757 -943
rect 23865 -977 23881 -943
rect 23741 -993 23881 -977
rect 23939 -943 24079 -896
rect 23939 -977 23955 -943
rect 24063 -977 24079 -943
rect 23939 -993 24079 -977
rect 24137 -943 24277 -896
rect 24137 -977 24153 -943
rect 24261 -977 24277 -943
rect 24137 -993 24277 -977
rect 24335 -943 24475 -896
rect 24335 -977 24351 -943
rect 24459 -977 24475 -943
rect 24335 -993 24475 -977
rect 24533 -943 24673 -896
rect 24533 -977 24549 -943
rect 24657 -977 24673 -943
rect 24533 -993 24673 -977
rect 24731 -943 24871 -896
rect 24731 -977 24747 -943
rect 24855 -977 24871 -943
rect 24731 -993 24871 -977
rect 24929 -943 25069 -896
rect 24929 -977 24945 -943
rect 25053 -977 25069 -943
rect 24929 -993 25069 -977
rect 25127 -943 25267 -896
rect 25127 -977 25143 -943
rect 25251 -977 25267 -943
rect 25127 -993 25267 -977
rect 25325 -943 25465 -896
rect 25325 -977 25341 -943
rect 25449 -977 25465 -943
rect 25325 -993 25465 -977
rect 25523 -943 25663 -896
rect 25523 -977 25539 -943
rect 25647 -977 25663 -943
rect 25523 -993 25663 -977
rect 25721 -943 25861 -896
rect 25721 -977 25737 -943
rect 25845 -977 25861 -943
rect 25721 -993 25861 -977
rect 25919 -943 26059 -896
rect 25919 -977 25935 -943
rect 26043 -977 26059 -943
rect 25919 -993 26059 -977
rect 26117 -943 26257 -896
rect 26117 -977 26133 -943
rect 26241 -977 26257 -943
rect 26117 -993 26257 -977
rect 26315 -943 26455 -896
rect 26315 -977 26331 -943
rect 26439 -977 26455 -943
rect 26315 -993 26455 -977
rect 26513 -943 26653 -896
rect 26513 -977 26529 -943
rect 26637 -977 26653 -943
rect 26513 -993 26653 -977
rect 26711 -943 26851 -896
rect 26711 -977 26727 -943
rect 26835 -977 26851 -943
rect 26711 -993 26851 -977
rect 26909 -943 27049 -896
rect 26909 -977 26925 -943
rect 27033 -977 27049 -943
rect 26909 -993 27049 -977
rect 27107 -943 27247 -896
rect 27107 -977 27123 -943
rect 27231 -977 27247 -943
rect 27107 -993 27247 -977
rect 27305 -943 27445 -896
rect 27305 -977 27321 -943
rect 27429 -977 27445 -943
rect 27305 -993 27445 -977
rect 27503 -943 27643 -896
rect 27503 -977 27519 -943
rect 27627 -977 27643 -943
rect 27503 -993 27643 -977
rect 27701 -943 27841 -896
rect 27701 -977 27717 -943
rect 27825 -977 27841 -943
rect 27701 -993 27841 -977
rect 27899 -943 28039 -896
rect 27899 -977 27915 -943
rect 28023 -977 28039 -943
rect 27899 -993 28039 -977
rect 28097 -943 28237 -896
rect 28097 -977 28113 -943
rect 28221 -977 28237 -943
rect 28097 -993 28237 -977
rect 28295 -943 28435 -896
rect 28295 -977 28311 -943
rect 28419 -977 28435 -943
rect 28295 -993 28435 -977
rect 28493 -943 28633 -896
rect 28493 -977 28509 -943
rect 28617 -977 28633 -943
rect 28493 -993 28633 -977
rect 28691 -943 28831 -896
rect 28691 -977 28707 -943
rect 28815 -977 28831 -943
rect 28691 -993 28831 -977
rect 28889 -943 29029 -896
rect 28889 -977 28905 -943
rect 29013 -977 29029 -943
rect 28889 -993 29029 -977
rect 29087 -943 29227 -896
rect 29087 -977 29103 -943
rect 29211 -977 29227 -943
rect 29087 -993 29227 -977
rect 29285 -943 29425 -896
rect 29285 -977 29301 -943
rect 29409 -977 29425 -943
rect 29285 -993 29425 -977
rect 29483 -943 29623 -896
rect 29483 -977 29499 -943
rect 29607 -977 29623 -943
rect 29483 -993 29623 -977
rect 29681 -943 29821 -896
rect 29681 -977 29697 -943
rect 29805 -977 29821 -943
rect 29681 -993 29821 -977
rect 29879 -943 30019 -896
rect 29879 -977 29895 -943
rect 30003 -977 30019 -943
rect 29879 -993 30019 -977
rect 30077 -943 30217 -896
rect 30077 -977 30093 -943
rect 30201 -977 30217 -943
rect 30077 -993 30217 -977
rect 30275 -943 30415 -896
rect 30275 -977 30291 -943
rect 30399 -977 30415 -943
rect 30275 -993 30415 -977
rect 30473 -943 30613 -896
rect 30473 -977 30489 -943
rect 30597 -977 30613 -943
rect 30473 -993 30613 -977
rect 30671 -943 30811 -896
rect 30671 -977 30687 -943
rect 30795 -977 30811 -943
rect 30671 -993 30811 -977
rect 30869 -943 31009 -896
rect 30869 -977 30885 -943
rect 30993 -977 31009 -943
rect 30869 -993 31009 -977
rect 31067 -943 31207 -896
rect 31067 -977 31083 -943
rect 31191 -977 31207 -943
rect 31067 -993 31207 -977
rect 31265 -943 31405 -896
rect 31265 -977 31281 -943
rect 31389 -977 31405 -943
rect 31265 -993 31405 -977
rect 31463 -943 31603 -896
rect 31463 -977 31479 -943
rect 31587 -977 31603 -943
rect 31463 -993 31603 -977
rect 23345 -1051 23485 -1035
rect 23345 -1085 23361 -1051
rect 23469 -1085 23485 -1051
rect 23345 -1132 23485 -1085
rect 23543 -1051 23683 -1035
rect 23543 -1085 23559 -1051
rect 23667 -1085 23683 -1051
rect 23543 -1132 23683 -1085
rect 23741 -1051 23881 -1035
rect 23741 -1085 23757 -1051
rect 23865 -1085 23881 -1051
rect 23741 -1132 23881 -1085
rect 23939 -1051 24079 -1035
rect 23939 -1085 23955 -1051
rect 24063 -1085 24079 -1051
rect 23939 -1132 24079 -1085
rect 24137 -1051 24277 -1035
rect 24137 -1085 24153 -1051
rect 24261 -1085 24277 -1051
rect 24137 -1132 24277 -1085
rect 24335 -1051 24475 -1035
rect 24335 -1085 24351 -1051
rect 24459 -1085 24475 -1051
rect 24335 -1132 24475 -1085
rect 24533 -1051 24673 -1035
rect 24533 -1085 24549 -1051
rect 24657 -1085 24673 -1051
rect 24533 -1132 24673 -1085
rect 24731 -1051 24871 -1035
rect 24731 -1085 24747 -1051
rect 24855 -1085 24871 -1051
rect 24731 -1132 24871 -1085
rect 24929 -1051 25069 -1035
rect 24929 -1085 24945 -1051
rect 25053 -1085 25069 -1051
rect 24929 -1132 25069 -1085
rect 25127 -1051 25267 -1035
rect 25127 -1085 25143 -1051
rect 25251 -1085 25267 -1051
rect 25127 -1132 25267 -1085
rect 25325 -1051 25465 -1035
rect 25325 -1085 25341 -1051
rect 25449 -1085 25465 -1051
rect 25325 -1132 25465 -1085
rect 25523 -1051 25663 -1035
rect 25523 -1085 25539 -1051
rect 25647 -1085 25663 -1051
rect 25523 -1132 25663 -1085
rect 25721 -1051 25861 -1035
rect 25721 -1085 25737 -1051
rect 25845 -1085 25861 -1051
rect 25721 -1132 25861 -1085
rect 25919 -1051 26059 -1035
rect 25919 -1085 25935 -1051
rect 26043 -1085 26059 -1051
rect 25919 -1132 26059 -1085
rect 26117 -1051 26257 -1035
rect 26117 -1085 26133 -1051
rect 26241 -1085 26257 -1051
rect 26117 -1132 26257 -1085
rect 26315 -1051 26455 -1035
rect 26315 -1085 26331 -1051
rect 26439 -1085 26455 -1051
rect 26315 -1132 26455 -1085
rect 26513 -1051 26653 -1035
rect 26513 -1085 26529 -1051
rect 26637 -1085 26653 -1051
rect 26513 -1132 26653 -1085
rect 26711 -1051 26851 -1035
rect 26711 -1085 26727 -1051
rect 26835 -1085 26851 -1051
rect 26711 -1132 26851 -1085
rect 26909 -1051 27049 -1035
rect 26909 -1085 26925 -1051
rect 27033 -1085 27049 -1051
rect 26909 -1132 27049 -1085
rect 27107 -1051 27247 -1035
rect 27107 -1085 27123 -1051
rect 27231 -1085 27247 -1051
rect 27107 -1132 27247 -1085
rect 27305 -1051 27445 -1035
rect 27305 -1085 27321 -1051
rect 27429 -1085 27445 -1051
rect 27305 -1132 27445 -1085
rect 27503 -1051 27643 -1035
rect 27503 -1085 27519 -1051
rect 27627 -1085 27643 -1051
rect 27503 -1132 27643 -1085
rect 27701 -1051 27841 -1035
rect 27701 -1085 27717 -1051
rect 27825 -1085 27841 -1051
rect 27701 -1132 27841 -1085
rect 27899 -1051 28039 -1035
rect 27899 -1085 27915 -1051
rect 28023 -1085 28039 -1051
rect 27899 -1132 28039 -1085
rect 28097 -1051 28237 -1035
rect 28097 -1085 28113 -1051
rect 28221 -1085 28237 -1051
rect 28097 -1132 28237 -1085
rect 28295 -1051 28435 -1035
rect 28295 -1085 28311 -1051
rect 28419 -1085 28435 -1051
rect 28295 -1132 28435 -1085
rect 28493 -1051 28633 -1035
rect 28493 -1085 28509 -1051
rect 28617 -1085 28633 -1051
rect 28493 -1132 28633 -1085
rect 28691 -1051 28831 -1035
rect 28691 -1085 28707 -1051
rect 28815 -1085 28831 -1051
rect 28691 -1132 28831 -1085
rect 28889 -1051 29029 -1035
rect 28889 -1085 28905 -1051
rect 29013 -1085 29029 -1051
rect 28889 -1132 29029 -1085
rect 29087 -1051 29227 -1035
rect 29087 -1085 29103 -1051
rect 29211 -1085 29227 -1051
rect 29087 -1132 29227 -1085
rect 29285 -1051 29425 -1035
rect 29285 -1085 29301 -1051
rect 29409 -1085 29425 -1051
rect 29285 -1132 29425 -1085
rect 29483 -1051 29623 -1035
rect 29483 -1085 29499 -1051
rect 29607 -1085 29623 -1051
rect 29483 -1132 29623 -1085
rect 29681 -1051 29821 -1035
rect 29681 -1085 29697 -1051
rect 29805 -1085 29821 -1051
rect 29681 -1132 29821 -1085
rect 29879 -1051 30019 -1035
rect 29879 -1085 29895 -1051
rect 30003 -1085 30019 -1051
rect 29879 -1132 30019 -1085
rect 30077 -1051 30217 -1035
rect 30077 -1085 30093 -1051
rect 30201 -1085 30217 -1051
rect 30077 -1132 30217 -1085
rect 30275 -1051 30415 -1035
rect 30275 -1085 30291 -1051
rect 30399 -1085 30415 -1051
rect 30275 -1132 30415 -1085
rect 30473 -1051 30613 -1035
rect 30473 -1085 30489 -1051
rect 30597 -1085 30613 -1051
rect 30473 -1132 30613 -1085
rect 30671 -1051 30811 -1035
rect 30671 -1085 30687 -1051
rect 30795 -1085 30811 -1051
rect 30671 -1132 30811 -1085
rect 30869 -1051 31009 -1035
rect 30869 -1085 30885 -1051
rect 30993 -1085 31009 -1051
rect 30869 -1132 31009 -1085
rect 31067 -1051 31207 -1035
rect 31067 -1085 31083 -1051
rect 31191 -1085 31207 -1051
rect 31067 -1132 31207 -1085
rect 31265 -1051 31405 -1035
rect 31265 -1085 31281 -1051
rect 31389 -1085 31405 -1051
rect 31265 -1132 31405 -1085
rect 31463 -1051 31603 -1035
rect 31463 -1085 31479 -1051
rect 31587 -1085 31603 -1051
rect 31463 -1132 31603 -1085
rect 23345 -2579 23485 -2532
rect 23345 -2613 23361 -2579
rect 23469 -2613 23485 -2579
rect 23345 -2629 23485 -2613
rect 23543 -2579 23683 -2532
rect 23543 -2613 23559 -2579
rect 23667 -2613 23683 -2579
rect 23543 -2629 23683 -2613
rect 23741 -2579 23881 -2532
rect 23741 -2613 23757 -2579
rect 23865 -2613 23881 -2579
rect 23741 -2629 23881 -2613
rect 23939 -2579 24079 -2532
rect 23939 -2613 23955 -2579
rect 24063 -2613 24079 -2579
rect 23939 -2629 24079 -2613
rect 24137 -2579 24277 -2532
rect 24137 -2613 24153 -2579
rect 24261 -2613 24277 -2579
rect 24137 -2629 24277 -2613
rect 24335 -2579 24475 -2532
rect 24335 -2613 24351 -2579
rect 24459 -2613 24475 -2579
rect 24335 -2629 24475 -2613
rect 24533 -2579 24673 -2532
rect 24533 -2613 24549 -2579
rect 24657 -2613 24673 -2579
rect 24533 -2629 24673 -2613
rect 24731 -2579 24871 -2532
rect 24731 -2613 24747 -2579
rect 24855 -2613 24871 -2579
rect 24731 -2629 24871 -2613
rect 24929 -2579 25069 -2532
rect 24929 -2613 24945 -2579
rect 25053 -2613 25069 -2579
rect 24929 -2629 25069 -2613
rect 25127 -2579 25267 -2532
rect 25127 -2613 25143 -2579
rect 25251 -2613 25267 -2579
rect 25127 -2629 25267 -2613
rect 25325 -2579 25465 -2532
rect 25325 -2613 25341 -2579
rect 25449 -2613 25465 -2579
rect 25325 -2629 25465 -2613
rect 25523 -2579 25663 -2532
rect 25523 -2613 25539 -2579
rect 25647 -2613 25663 -2579
rect 25523 -2629 25663 -2613
rect 25721 -2579 25861 -2532
rect 25721 -2613 25737 -2579
rect 25845 -2613 25861 -2579
rect 25721 -2629 25861 -2613
rect 25919 -2579 26059 -2532
rect 25919 -2613 25935 -2579
rect 26043 -2613 26059 -2579
rect 25919 -2629 26059 -2613
rect 26117 -2579 26257 -2532
rect 26117 -2613 26133 -2579
rect 26241 -2613 26257 -2579
rect 26117 -2629 26257 -2613
rect 26315 -2579 26455 -2532
rect 26315 -2613 26331 -2579
rect 26439 -2613 26455 -2579
rect 26315 -2629 26455 -2613
rect 26513 -2579 26653 -2532
rect 26513 -2613 26529 -2579
rect 26637 -2613 26653 -2579
rect 26513 -2629 26653 -2613
rect 26711 -2579 26851 -2532
rect 26711 -2613 26727 -2579
rect 26835 -2613 26851 -2579
rect 26711 -2629 26851 -2613
rect 26909 -2579 27049 -2532
rect 26909 -2613 26925 -2579
rect 27033 -2613 27049 -2579
rect 26909 -2629 27049 -2613
rect 27107 -2579 27247 -2532
rect 27107 -2613 27123 -2579
rect 27231 -2613 27247 -2579
rect 27107 -2629 27247 -2613
rect 27305 -2579 27445 -2532
rect 27305 -2613 27321 -2579
rect 27429 -2613 27445 -2579
rect 27305 -2629 27445 -2613
rect 27503 -2579 27643 -2532
rect 27503 -2613 27519 -2579
rect 27627 -2613 27643 -2579
rect 27503 -2629 27643 -2613
rect 27701 -2579 27841 -2532
rect 27701 -2613 27717 -2579
rect 27825 -2613 27841 -2579
rect 27701 -2629 27841 -2613
rect 27899 -2579 28039 -2532
rect 27899 -2613 27915 -2579
rect 28023 -2613 28039 -2579
rect 27899 -2629 28039 -2613
rect 28097 -2579 28237 -2532
rect 28097 -2613 28113 -2579
rect 28221 -2613 28237 -2579
rect 28097 -2629 28237 -2613
rect 28295 -2579 28435 -2532
rect 28295 -2613 28311 -2579
rect 28419 -2613 28435 -2579
rect 28295 -2629 28435 -2613
rect 28493 -2579 28633 -2532
rect 28493 -2613 28509 -2579
rect 28617 -2613 28633 -2579
rect 28493 -2629 28633 -2613
rect 28691 -2579 28831 -2532
rect 28691 -2613 28707 -2579
rect 28815 -2613 28831 -2579
rect 28691 -2629 28831 -2613
rect 28889 -2579 29029 -2532
rect 28889 -2613 28905 -2579
rect 29013 -2613 29029 -2579
rect 28889 -2629 29029 -2613
rect 29087 -2579 29227 -2532
rect 29087 -2613 29103 -2579
rect 29211 -2613 29227 -2579
rect 29087 -2629 29227 -2613
rect 29285 -2579 29425 -2532
rect 29285 -2613 29301 -2579
rect 29409 -2613 29425 -2579
rect 29285 -2629 29425 -2613
rect 29483 -2579 29623 -2532
rect 29483 -2613 29499 -2579
rect 29607 -2613 29623 -2579
rect 29483 -2629 29623 -2613
rect 29681 -2579 29821 -2532
rect 29681 -2613 29697 -2579
rect 29805 -2613 29821 -2579
rect 29681 -2629 29821 -2613
rect 29879 -2579 30019 -2532
rect 29879 -2613 29895 -2579
rect 30003 -2613 30019 -2579
rect 29879 -2629 30019 -2613
rect 30077 -2579 30217 -2532
rect 30077 -2613 30093 -2579
rect 30201 -2613 30217 -2579
rect 30077 -2629 30217 -2613
rect 30275 -2579 30415 -2532
rect 30275 -2613 30291 -2579
rect 30399 -2613 30415 -2579
rect 30275 -2629 30415 -2613
rect 30473 -2579 30613 -2532
rect 30473 -2613 30489 -2579
rect 30597 -2613 30613 -2579
rect 30473 -2629 30613 -2613
rect 30671 -2579 30811 -2532
rect 30671 -2613 30687 -2579
rect 30795 -2613 30811 -2579
rect 30671 -2629 30811 -2613
rect 30869 -2579 31009 -2532
rect 30869 -2613 30885 -2579
rect 30993 -2613 31009 -2579
rect 30869 -2629 31009 -2613
rect 31067 -2579 31207 -2532
rect 31067 -2613 31083 -2579
rect 31191 -2613 31207 -2579
rect 31067 -2629 31207 -2613
rect 31265 -2579 31405 -2532
rect 31265 -2613 31281 -2579
rect 31389 -2613 31405 -2579
rect 31265 -2629 31405 -2613
rect 31463 -2579 31603 -2532
rect 31463 -2613 31479 -2579
rect 31587 -2613 31603 -2579
rect 31463 -2629 31603 -2613
rect 23345 -2687 23485 -2671
rect 23345 -2721 23361 -2687
rect 23469 -2721 23485 -2687
rect 23345 -2768 23485 -2721
rect 23543 -2687 23683 -2671
rect 23543 -2721 23559 -2687
rect 23667 -2721 23683 -2687
rect 23543 -2768 23683 -2721
rect 23741 -2687 23881 -2671
rect 23741 -2721 23757 -2687
rect 23865 -2721 23881 -2687
rect 23741 -2768 23881 -2721
rect 23939 -2687 24079 -2671
rect 23939 -2721 23955 -2687
rect 24063 -2721 24079 -2687
rect 23939 -2768 24079 -2721
rect 24137 -2687 24277 -2671
rect 24137 -2721 24153 -2687
rect 24261 -2721 24277 -2687
rect 24137 -2768 24277 -2721
rect 24335 -2687 24475 -2671
rect 24335 -2721 24351 -2687
rect 24459 -2721 24475 -2687
rect 24335 -2768 24475 -2721
rect 24533 -2687 24673 -2671
rect 24533 -2721 24549 -2687
rect 24657 -2721 24673 -2687
rect 24533 -2768 24673 -2721
rect 24731 -2687 24871 -2671
rect 24731 -2721 24747 -2687
rect 24855 -2721 24871 -2687
rect 24731 -2768 24871 -2721
rect 24929 -2687 25069 -2671
rect 24929 -2721 24945 -2687
rect 25053 -2721 25069 -2687
rect 24929 -2768 25069 -2721
rect 25127 -2687 25267 -2671
rect 25127 -2721 25143 -2687
rect 25251 -2721 25267 -2687
rect 25127 -2768 25267 -2721
rect 25325 -2687 25465 -2671
rect 25325 -2721 25341 -2687
rect 25449 -2721 25465 -2687
rect 25325 -2768 25465 -2721
rect 25523 -2687 25663 -2671
rect 25523 -2721 25539 -2687
rect 25647 -2721 25663 -2687
rect 25523 -2768 25663 -2721
rect 25721 -2687 25861 -2671
rect 25721 -2721 25737 -2687
rect 25845 -2721 25861 -2687
rect 25721 -2768 25861 -2721
rect 25919 -2687 26059 -2671
rect 25919 -2721 25935 -2687
rect 26043 -2721 26059 -2687
rect 25919 -2768 26059 -2721
rect 26117 -2687 26257 -2671
rect 26117 -2721 26133 -2687
rect 26241 -2721 26257 -2687
rect 26117 -2768 26257 -2721
rect 26315 -2687 26455 -2671
rect 26315 -2721 26331 -2687
rect 26439 -2721 26455 -2687
rect 26315 -2768 26455 -2721
rect 26513 -2687 26653 -2671
rect 26513 -2721 26529 -2687
rect 26637 -2721 26653 -2687
rect 26513 -2768 26653 -2721
rect 26711 -2687 26851 -2671
rect 26711 -2721 26727 -2687
rect 26835 -2721 26851 -2687
rect 26711 -2768 26851 -2721
rect 26909 -2687 27049 -2671
rect 26909 -2721 26925 -2687
rect 27033 -2721 27049 -2687
rect 26909 -2768 27049 -2721
rect 27107 -2687 27247 -2671
rect 27107 -2721 27123 -2687
rect 27231 -2721 27247 -2687
rect 27107 -2768 27247 -2721
rect 27305 -2687 27445 -2671
rect 27305 -2721 27321 -2687
rect 27429 -2721 27445 -2687
rect 27305 -2768 27445 -2721
rect 27503 -2687 27643 -2671
rect 27503 -2721 27519 -2687
rect 27627 -2721 27643 -2687
rect 27503 -2768 27643 -2721
rect 27701 -2687 27841 -2671
rect 27701 -2721 27717 -2687
rect 27825 -2721 27841 -2687
rect 27701 -2768 27841 -2721
rect 27899 -2687 28039 -2671
rect 27899 -2721 27915 -2687
rect 28023 -2721 28039 -2687
rect 27899 -2768 28039 -2721
rect 28097 -2687 28237 -2671
rect 28097 -2721 28113 -2687
rect 28221 -2721 28237 -2687
rect 28097 -2768 28237 -2721
rect 28295 -2687 28435 -2671
rect 28295 -2721 28311 -2687
rect 28419 -2721 28435 -2687
rect 28295 -2768 28435 -2721
rect 28493 -2687 28633 -2671
rect 28493 -2721 28509 -2687
rect 28617 -2721 28633 -2687
rect 28493 -2768 28633 -2721
rect 28691 -2687 28831 -2671
rect 28691 -2721 28707 -2687
rect 28815 -2721 28831 -2687
rect 28691 -2768 28831 -2721
rect 28889 -2687 29029 -2671
rect 28889 -2721 28905 -2687
rect 29013 -2721 29029 -2687
rect 28889 -2768 29029 -2721
rect 29087 -2687 29227 -2671
rect 29087 -2721 29103 -2687
rect 29211 -2721 29227 -2687
rect 29087 -2768 29227 -2721
rect 29285 -2687 29425 -2671
rect 29285 -2721 29301 -2687
rect 29409 -2721 29425 -2687
rect 29285 -2768 29425 -2721
rect 29483 -2687 29623 -2671
rect 29483 -2721 29499 -2687
rect 29607 -2721 29623 -2687
rect 29483 -2768 29623 -2721
rect 29681 -2687 29821 -2671
rect 29681 -2721 29697 -2687
rect 29805 -2721 29821 -2687
rect 29681 -2768 29821 -2721
rect 29879 -2687 30019 -2671
rect 29879 -2721 29895 -2687
rect 30003 -2721 30019 -2687
rect 29879 -2768 30019 -2721
rect 30077 -2687 30217 -2671
rect 30077 -2721 30093 -2687
rect 30201 -2721 30217 -2687
rect 30077 -2768 30217 -2721
rect 30275 -2687 30415 -2671
rect 30275 -2721 30291 -2687
rect 30399 -2721 30415 -2687
rect 30275 -2768 30415 -2721
rect 30473 -2687 30613 -2671
rect 30473 -2721 30489 -2687
rect 30597 -2721 30613 -2687
rect 30473 -2768 30613 -2721
rect 30671 -2687 30811 -2671
rect 30671 -2721 30687 -2687
rect 30795 -2721 30811 -2687
rect 30671 -2768 30811 -2721
rect 30869 -2687 31009 -2671
rect 30869 -2721 30885 -2687
rect 30993 -2721 31009 -2687
rect 30869 -2768 31009 -2721
rect 31067 -2687 31207 -2671
rect 31067 -2721 31083 -2687
rect 31191 -2721 31207 -2687
rect 31067 -2768 31207 -2721
rect 31265 -2687 31405 -2671
rect 31265 -2721 31281 -2687
rect 31389 -2721 31405 -2687
rect 31265 -2768 31405 -2721
rect 31463 -2687 31603 -2671
rect 31463 -2721 31479 -2687
rect 31587 -2721 31603 -2687
rect 31463 -2768 31603 -2721
rect 23345 -4194 23485 -4168
rect 23543 -4194 23683 -4168
rect 23741 -4194 23881 -4168
rect 23939 -4194 24079 -4168
rect 24137 -4194 24277 -4168
rect 24335 -4194 24475 -4168
rect 24533 -4194 24673 -4168
rect 24731 -4194 24871 -4168
rect 24929 -4194 25069 -4168
rect 25127 -4194 25267 -4168
rect 25325 -4194 25465 -4168
rect 25523 -4194 25663 -4168
rect 25721 -4194 25861 -4168
rect 25919 -4194 26059 -4168
rect 26117 -4194 26257 -4168
rect 26315 -4194 26455 -4168
rect 26513 -4194 26653 -4168
rect 26711 -4194 26851 -4168
rect 26909 -4194 27049 -4168
rect 27107 -4194 27247 -4168
rect 27305 -4194 27445 -4168
rect 27503 -4194 27643 -4168
rect 27701 -4194 27841 -4168
rect 27899 -4194 28039 -4168
rect 28097 -4194 28237 -4168
rect 28295 -4194 28435 -4168
rect 28493 -4194 28633 -4168
rect 28691 -4194 28831 -4168
rect 28889 -4194 29029 -4168
rect 29087 -4194 29227 -4168
rect 29285 -4194 29425 -4168
rect 29483 -4194 29623 -4168
rect 29681 -4194 29821 -4168
rect 29879 -4194 30019 -4168
rect 30077 -4194 30217 -4168
rect 30275 -4194 30415 -4168
rect 30473 -4194 30613 -4168
rect 30671 -4194 30811 -4168
rect 30869 -4194 31009 -4168
rect 31067 -4194 31207 -4168
rect 31265 -4194 31405 -4168
rect 31463 -4194 31603 -4168
<< polycont >>
rect 11511 659 11619 693
rect 11709 659 11817 693
rect 11907 659 12015 693
rect 12105 659 12213 693
rect 12303 659 12411 693
rect 12501 659 12609 693
rect 12699 659 12807 693
rect 12897 659 13005 693
rect 13095 659 13203 693
rect 13293 659 13401 693
rect 13491 659 13599 693
rect 13689 659 13797 693
rect 13887 659 13995 693
rect 14085 659 14193 693
rect 14283 659 14391 693
rect 14481 659 14589 693
rect 14679 659 14787 693
rect 14877 659 14985 693
rect 15075 659 15183 693
rect 15273 659 15381 693
rect 15471 659 15579 693
rect 15669 659 15777 693
rect 15867 659 15975 693
rect 16065 659 16173 693
rect 16263 659 16371 693
rect 16461 659 16569 693
rect 16659 659 16767 693
rect 16857 659 16965 693
rect 17055 659 17163 693
rect 17253 659 17361 693
rect 17451 659 17559 693
rect 17649 659 17757 693
rect 17847 659 17955 693
rect 18045 659 18153 693
rect 18243 659 18351 693
rect 18441 659 18549 693
rect 18639 659 18747 693
rect 18837 659 18945 693
rect 19035 659 19143 693
rect 19233 659 19341 693
rect 19431 659 19539 693
rect 19629 659 19737 693
rect 11511 551 11619 585
rect 11709 551 11817 585
rect 11907 551 12015 585
rect 12105 551 12213 585
rect 12303 551 12411 585
rect 12501 551 12609 585
rect 12699 551 12807 585
rect 12897 551 13005 585
rect 13095 551 13203 585
rect 13293 551 13401 585
rect 13491 551 13599 585
rect 13689 551 13797 585
rect 13887 551 13995 585
rect 14085 551 14193 585
rect 14283 551 14391 585
rect 14481 551 14589 585
rect 14679 551 14787 585
rect 14877 551 14985 585
rect 15075 551 15183 585
rect 15273 551 15381 585
rect 15471 551 15579 585
rect 15669 551 15777 585
rect 15867 551 15975 585
rect 16065 551 16173 585
rect 16263 551 16371 585
rect 16461 551 16569 585
rect 16659 551 16767 585
rect 16857 551 16965 585
rect 17055 551 17163 585
rect 17253 551 17361 585
rect 17451 551 17559 585
rect 17649 551 17757 585
rect 17847 551 17955 585
rect 18045 551 18153 585
rect 18243 551 18351 585
rect 18441 551 18549 585
rect 18639 551 18747 585
rect 18837 551 18945 585
rect 19035 551 19143 585
rect 19233 551 19341 585
rect 19431 551 19539 585
rect 19629 551 19737 585
rect 11511 -977 11619 -943
rect 11709 -977 11817 -943
rect 11907 -977 12015 -943
rect 12105 -977 12213 -943
rect 12303 -977 12411 -943
rect 12501 -977 12609 -943
rect 12699 -977 12807 -943
rect 12897 -977 13005 -943
rect 13095 -977 13203 -943
rect 13293 -977 13401 -943
rect 13491 -977 13599 -943
rect 13689 -977 13797 -943
rect 13887 -977 13995 -943
rect 14085 -977 14193 -943
rect 14283 -977 14391 -943
rect 14481 -977 14589 -943
rect 14679 -977 14787 -943
rect 14877 -977 14985 -943
rect 15075 -977 15183 -943
rect 15273 -977 15381 -943
rect 15471 -977 15579 -943
rect 15669 -977 15777 -943
rect 15867 -977 15975 -943
rect 16065 -977 16173 -943
rect 16263 -977 16371 -943
rect 16461 -977 16569 -943
rect 16659 -977 16767 -943
rect 16857 -977 16965 -943
rect 17055 -977 17163 -943
rect 17253 -977 17361 -943
rect 17451 -977 17559 -943
rect 17649 -977 17757 -943
rect 17847 -977 17955 -943
rect 18045 -977 18153 -943
rect 18243 -977 18351 -943
rect 18441 -977 18549 -943
rect 18639 -977 18747 -943
rect 18837 -977 18945 -943
rect 19035 -977 19143 -943
rect 19233 -977 19341 -943
rect 19431 -977 19539 -943
rect 19629 -977 19737 -943
rect 11511 -1085 11619 -1051
rect 11709 -1085 11817 -1051
rect 11907 -1085 12015 -1051
rect 12105 -1085 12213 -1051
rect 12303 -1085 12411 -1051
rect 12501 -1085 12609 -1051
rect 12699 -1085 12807 -1051
rect 12897 -1085 13005 -1051
rect 13095 -1085 13203 -1051
rect 13293 -1085 13401 -1051
rect 13491 -1085 13599 -1051
rect 13689 -1085 13797 -1051
rect 13887 -1085 13995 -1051
rect 14085 -1085 14193 -1051
rect 14283 -1085 14391 -1051
rect 14481 -1085 14589 -1051
rect 14679 -1085 14787 -1051
rect 14877 -1085 14985 -1051
rect 15075 -1085 15183 -1051
rect 15273 -1085 15381 -1051
rect 15471 -1085 15579 -1051
rect 15669 -1085 15777 -1051
rect 15867 -1085 15975 -1051
rect 16065 -1085 16173 -1051
rect 16263 -1085 16371 -1051
rect 16461 -1085 16569 -1051
rect 16659 -1085 16767 -1051
rect 16857 -1085 16965 -1051
rect 17055 -1085 17163 -1051
rect 17253 -1085 17361 -1051
rect 17451 -1085 17559 -1051
rect 17649 -1085 17757 -1051
rect 17847 -1085 17955 -1051
rect 18045 -1085 18153 -1051
rect 18243 -1085 18351 -1051
rect 18441 -1085 18549 -1051
rect 18639 -1085 18747 -1051
rect 18837 -1085 18945 -1051
rect 19035 -1085 19143 -1051
rect 19233 -1085 19341 -1051
rect 19431 -1085 19539 -1051
rect 19629 -1085 19737 -1051
rect 11511 -2613 11619 -2579
rect 11709 -2613 11817 -2579
rect 11907 -2613 12015 -2579
rect 12105 -2613 12213 -2579
rect 12303 -2613 12411 -2579
rect 12501 -2613 12609 -2579
rect 12699 -2613 12807 -2579
rect 12897 -2613 13005 -2579
rect 13095 -2613 13203 -2579
rect 13293 -2613 13401 -2579
rect 13491 -2613 13599 -2579
rect 13689 -2613 13797 -2579
rect 13887 -2613 13995 -2579
rect 14085 -2613 14193 -2579
rect 14283 -2613 14391 -2579
rect 14481 -2613 14589 -2579
rect 14679 -2613 14787 -2579
rect 14877 -2613 14985 -2579
rect 15075 -2613 15183 -2579
rect 15273 -2613 15381 -2579
rect 15471 -2613 15579 -2579
rect 15669 -2613 15777 -2579
rect 15867 -2613 15975 -2579
rect 16065 -2613 16173 -2579
rect 16263 -2613 16371 -2579
rect 16461 -2613 16569 -2579
rect 16659 -2613 16767 -2579
rect 16857 -2613 16965 -2579
rect 17055 -2613 17163 -2579
rect 17253 -2613 17361 -2579
rect 17451 -2613 17559 -2579
rect 17649 -2613 17757 -2579
rect 17847 -2613 17955 -2579
rect 18045 -2613 18153 -2579
rect 18243 -2613 18351 -2579
rect 18441 -2613 18549 -2579
rect 18639 -2613 18747 -2579
rect 18837 -2613 18945 -2579
rect 19035 -2613 19143 -2579
rect 19233 -2613 19341 -2579
rect 19431 -2613 19539 -2579
rect 19629 -2613 19737 -2579
rect 11511 -2721 11619 -2687
rect 11709 -2721 11817 -2687
rect 11907 -2721 12015 -2687
rect 12105 -2721 12213 -2687
rect 12303 -2721 12411 -2687
rect 12501 -2721 12609 -2687
rect 12699 -2721 12807 -2687
rect 12897 -2721 13005 -2687
rect 13095 -2721 13203 -2687
rect 13293 -2721 13401 -2687
rect 13491 -2721 13599 -2687
rect 13689 -2721 13797 -2687
rect 13887 -2721 13995 -2687
rect 14085 -2721 14193 -2687
rect 14283 -2721 14391 -2687
rect 14481 -2721 14589 -2687
rect 14679 -2721 14787 -2687
rect 14877 -2721 14985 -2687
rect 15075 -2721 15183 -2687
rect 15273 -2721 15381 -2687
rect 15471 -2721 15579 -2687
rect 15669 -2721 15777 -2687
rect 15867 -2721 15975 -2687
rect 16065 -2721 16173 -2687
rect 16263 -2721 16371 -2687
rect 16461 -2721 16569 -2687
rect 16659 -2721 16767 -2687
rect 16857 -2721 16965 -2687
rect 17055 -2721 17163 -2687
rect 17253 -2721 17361 -2687
rect 17451 -2721 17559 -2687
rect 17649 -2721 17757 -2687
rect 17847 -2721 17955 -2687
rect 18045 -2721 18153 -2687
rect 18243 -2721 18351 -2687
rect 18441 -2721 18549 -2687
rect 18639 -2721 18747 -2687
rect 18837 -2721 18945 -2687
rect 19035 -2721 19143 -2687
rect 19233 -2721 19341 -2687
rect 19431 -2721 19539 -2687
rect 19629 -2721 19737 -2687
rect 23361 659 23469 693
rect 23559 659 23667 693
rect 23757 659 23865 693
rect 23955 659 24063 693
rect 24153 659 24261 693
rect 24351 659 24459 693
rect 24549 659 24657 693
rect 24747 659 24855 693
rect 24945 659 25053 693
rect 25143 659 25251 693
rect 25341 659 25449 693
rect 25539 659 25647 693
rect 25737 659 25845 693
rect 25935 659 26043 693
rect 26133 659 26241 693
rect 26331 659 26439 693
rect 26529 659 26637 693
rect 26727 659 26835 693
rect 26925 659 27033 693
rect 27123 659 27231 693
rect 27321 659 27429 693
rect 27519 659 27627 693
rect 27717 659 27825 693
rect 27915 659 28023 693
rect 28113 659 28221 693
rect 28311 659 28419 693
rect 28509 659 28617 693
rect 28707 659 28815 693
rect 28905 659 29013 693
rect 29103 659 29211 693
rect 29301 659 29409 693
rect 29499 659 29607 693
rect 29697 659 29805 693
rect 29895 659 30003 693
rect 30093 659 30201 693
rect 30291 659 30399 693
rect 30489 659 30597 693
rect 30687 659 30795 693
rect 30885 659 30993 693
rect 31083 659 31191 693
rect 31281 659 31389 693
rect 31479 659 31587 693
rect 23361 551 23469 585
rect 23559 551 23667 585
rect 23757 551 23865 585
rect 23955 551 24063 585
rect 24153 551 24261 585
rect 24351 551 24459 585
rect 24549 551 24657 585
rect 24747 551 24855 585
rect 24945 551 25053 585
rect 25143 551 25251 585
rect 25341 551 25449 585
rect 25539 551 25647 585
rect 25737 551 25845 585
rect 25935 551 26043 585
rect 26133 551 26241 585
rect 26331 551 26439 585
rect 26529 551 26637 585
rect 26727 551 26835 585
rect 26925 551 27033 585
rect 27123 551 27231 585
rect 27321 551 27429 585
rect 27519 551 27627 585
rect 27717 551 27825 585
rect 27915 551 28023 585
rect 28113 551 28221 585
rect 28311 551 28419 585
rect 28509 551 28617 585
rect 28707 551 28815 585
rect 28905 551 29013 585
rect 29103 551 29211 585
rect 29301 551 29409 585
rect 29499 551 29607 585
rect 29697 551 29805 585
rect 29895 551 30003 585
rect 30093 551 30201 585
rect 30291 551 30399 585
rect 30489 551 30597 585
rect 30687 551 30795 585
rect 30885 551 30993 585
rect 31083 551 31191 585
rect 31281 551 31389 585
rect 31479 551 31587 585
rect 23361 -977 23469 -943
rect 23559 -977 23667 -943
rect 23757 -977 23865 -943
rect 23955 -977 24063 -943
rect 24153 -977 24261 -943
rect 24351 -977 24459 -943
rect 24549 -977 24657 -943
rect 24747 -977 24855 -943
rect 24945 -977 25053 -943
rect 25143 -977 25251 -943
rect 25341 -977 25449 -943
rect 25539 -977 25647 -943
rect 25737 -977 25845 -943
rect 25935 -977 26043 -943
rect 26133 -977 26241 -943
rect 26331 -977 26439 -943
rect 26529 -977 26637 -943
rect 26727 -977 26835 -943
rect 26925 -977 27033 -943
rect 27123 -977 27231 -943
rect 27321 -977 27429 -943
rect 27519 -977 27627 -943
rect 27717 -977 27825 -943
rect 27915 -977 28023 -943
rect 28113 -977 28221 -943
rect 28311 -977 28419 -943
rect 28509 -977 28617 -943
rect 28707 -977 28815 -943
rect 28905 -977 29013 -943
rect 29103 -977 29211 -943
rect 29301 -977 29409 -943
rect 29499 -977 29607 -943
rect 29697 -977 29805 -943
rect 29895 -977 30003 -943
rect 30093 -977 30201 -943
rect 30291 -977 30399 -943
rect 30489 -977 30597 -943
rect 30687 -977 30795 -943
rect 30885 -977 30993 -943
rect 31083 -977 31191 -943
rect 31281 -977 31389 -943
rect 31479 -977 31587 -943
rect 23361 -1085 23469 -1051
rect 23559 -1085 23667 -1051
rect 23757 -1085 23865 -1051
rect 23955 -1085 24063 -1051
rect 24153 -1085 24261 -1051
rect 24351 -1085 24459 -1051
rect 24549 -1085 24657 -1051
rect 24747 -1085 24855 -1051
rect 24945 -1085 25053 -1051
rect 25143 -1085 25251 -1051
rect 25341 -1085 25449 -1051
rect 25539 -1085 25647 -1051
rect 25737 -1085 25845 -1051
rect 25935 -1085 26043 -1051
rect 26133 -1085 26241 -1051
rect 26331 -1085 26439 -1051
rect 26529 -1085 26637 -1051
rect 26727 -1085 26835 -1051
rect 26925 -1085 27033 -1051
rect 27123 -1085 27231 -1051
rect 27321 -1085 27429 -1051
rect 27519 -1085 27627 -1051
rect 27717 -1085 27825 -1051
rect 27915 -1085 28023 -1051
rect 28113 -1085 28221 -1051
rect 28311 -1085 28419 -1051
rect 28509 -1085 28617 -1051
rect 28707 -1085 28815 -1051
rect 28905 -1085 29013 -1051
rect 29103 -1085 29211 -1051
rect 29301 -1085 29409 -1051
rect 29499 -1085 29607 -1051
rect 29697 -1085 29805 -1051
rect 29895 -1085 30003 -1051
rect 30093 -1085 30201 -1051
rect 30291 -1085 30399 -1051
rect 30489 -1085 30597 -1051
rect 30687 -1085 30795 -1051
rect 30885 -1085 30993 -1051
rect 31083 -1085 31191 -1051
rect 31281 -1085 31389 -1051
rect 31479 -1085 31587 -1051
rect 23361 -2613 23469 -2579
rect 23559 -2613 23667 -2579
rect 23757 -2613 23865 -2579
rect 23955 -2613 24063 -2579
rect 24153 -2613 24261 -2579
rect 24351 -2613 24459 -2579
rect 24549 -2613 24657 -2579
rect 24747 -2613 24855 -2579
rect 24945 -2613 25053 -2579
rect 25143 -2613 25251 -2579
rect 25341 -2613 25449 -2579
rect 25539 -2613 25647 -2579
rect 25737 -2613 25845 -2579
rect 25935 -2613 26043 -2579
rect 26133 -2613 26241 -2579
rect 26331 -2613 26439 -2579
rect 26529 -2613 26637 -2579
rect 26727 -2613 26835 -2579
rect 26925 -2613 27033 -2579
rect 27123 -2613 27231 -2579
rect 27321 -2613 27429 -2579
rect 27519 -2613 27627 -2579
rect 27717 -2613 27825 -2579
rect 27915 -2613 28023 -2579
rect 28113 -2613 28221 -2579
rect 28311 -2613 28419 -2579
rect 28509 -2613 28617 -2579
rect 28707 -2613 28815 -2579
rect 28905 -2613 29013 -2579
rect 29103 -2613 29211 -2579
rect 29301 -2613 29409 -2579
rect 29499 -2613 29607 -2579
rect 29697 -2613 29805 -2579
rect 29895 -2613 30003 -2579
rect 30093 -2613 30201 -2579
rect 30291 -2613 30399 -2579
rect 30489 -2613 30597 -2579
rect 30687 -2613 30795 -2579
rect 30885 -2613 30993 -2579
rect 31083 -2613 31191 -2579
rect 31281 -2613 31389 -2579
rect 31479 -2613 31587 -2579
rect 23361 -2721 23469 -2687
rect 23559 -2721 23667 -2687
rect 23757 -2721 23865 -2687
rect 23955 -2721 24063 -2687
rect 24153 -2721 24261 -2687
rect 24351 -2721 24459 -2687
rect 24549 -2721 24657 -2687
rect 24747 -2721 24855 -2687
rect 24945 -2721 25053 -2687
rect 25143 -2721 25251 -2687
rect 25341 -2721 25449 -2687
rect 25539 -2721 25647 -2687
rect 25737 -2721 25845 -2687
rect 25935 -2721 26043 -2687
rect 26133 -2721 26241 -2687
rect 26331 -2721 26439 -2687
rect 26529 -2721 26637 -2687
rect 26727 -2721 26835 -2687
rect 26925 -2721 27033 -2687
rect 27123 -2721 27231 -2687
rect 27321 -2721 27429 -2687
rect 27519 -2721 27627 -2687
rect 27717 -2721 27825 -2687
rect 27915 -2721 28023 -2687
rect 28113 -2721 28221 -2687
rect 28311 -2721 28419 -2687
rect 28509 -2721 28617 -2687
rect 28707 -2721 28815 -2687
rect 28905 -2721 29013 -2687
rect 29103 -2721 29211 -2687
rect 29301 -2721 29409 -2687
rect 29499 -2721 29607 -2687
rect 29697 -2721 29805 -2687
rect 29895 -2721 30003 -2687
rect 30093 -2721 30201 -2687
rect 30291 -2721 30399 -2687
rect 30489 -2721 30597 -2687
rect 30687 -2721 30795 -2687
rect 30885 -2721 30993 -2687
rect 31083 -2721 31191 -2687
rect 31281 -2721 31389 -2687
rect 31479 -2721 31587 -2687
<< locali >>
rect -848 2237 -752 2271
rect 8337 2237 8433 2271
rect -848 2175 -814 2237
rect -848 -4415 -814 -4353
rect 8399 2175 8433 2237
rect 8399 -4415 8433 -4353
rect -848 -4449 -752 -4415
rect 8337 -4449 8433 -4415
rect 10991 2237 11087 2271
rect 20176 2237 20272 2271
rect 10991 2175 11025 2237
rect 20238 2175 20272 2237
rect 11449 2128 11483 2144
rect 11449 736 11483 752
rect 11647 2128 11681 2144
rect 11647 736 11681 752
rect 11845 2128 11879 2144
rect 11845 736 11879 752
rect 12043 2128 12077 2144
rect 12043 736 12077 752
rect 12241 2128 12275 2144
rect 12241 736 12275 752
rect 12439 2128 12473 2144
rect 12439 736 12473 752
rect 12637 2128 12671 2144
rect 12637 736 12671 752
rect 12835 2128 12869 2144
rect 12835 736 12869 752
rect 13033 2128 13067 2144
rect 13033 736 13067 752
rect 13231 2128 13265 2144
rect 13231 736 13265 752
rect 13429 2128 13463 2144
rect 13429 736 13463 752
rect 13627 2128 13661 2144
rect 13627 736 13661 752
rect 13825 2128 13859 2144
rect 13825 736 13859 752
rect 14023 2128 14057 2144
rect 14023 736 14057 752
rect 14221 2128 14255 2144
rect 14221 736 14255 752
rect 14419 2128 14453 2144
rect 14419 736 14453 752
rect 14617 2128 14651 2144
rect 14617 736 14651 752
rect 14815 2128 14849 2144
rect 14815 736 14849 752
rect 15013 2128 15047 2144
rect 15013 736 15047 752
rect 15211 2128 15245 2144
rect 15211 736 15245 752
rect 15409 2128 15443 2144
rect 15409 736 15443 752
rect 15607 2128 15641 2144
rect 15607 736 15641 752
rect 15805 2128 15839 2144
rect 15805 736 15839 752
rect 16003 2128 16037 2144
rect 16003 736 16037 752
rect 16201 2128 16235 2144
rect 16201 736 16235 752
rect 16399 2128 16433 2144
rect 16399 736 16433 752
rect 16597 2128 16631 2144
rect 16597 736 16631 752
rect 16795 2128 16829 2144
rect 16795 736 16829 752
rect 16993 2128 17027 2144
rect 16993 736 17027 752
rect 17191 2128 17225 2144
rect 17191 736 17225 752
rect 17389 2128 17423 2144
rect 17389 736 17423 752
rect 17587 2128 17621 2144
rect 17587 736 17621 752
rect 17785 2128 17819 2144
rect 17785 736 17819 752
rect 17983 2128 18017 2144
rect 17983 736 18017 752
rect 18181 2128 18215 2144
rect 18181 736 18215 752
rect 18379 2128 18413 2144
rect 18379 736 18413 752
rect 18577 2128 18611 2144
rect 18577 736 18611 752
rect 18775 2128 18809 2144
rect 18775 736 18809 752
rect 18973 2128 19007 2144
rect 18973 736 19007 752
rect 19171 2128 19205 2144
rect 19171 736 19205 752
rect 19369 2128 19403 2144
rect 19369 736 19403 752
rect 19567 2128 19601 2144
rect 19567 736 19601 752
rect 19765 2128 19799 2144
rect 19765 736 19799 752
rect 11495 659 11511 693
rect 11619 659 11635 693
rect 11693 659 11709 693
rect 11817 659 11833 693
rect 11891 659 11907 693
rect 12015 659 12031 693
rect 12089 659 12105 693
rect 12213 659 12229 693
rect 12287 659 12303 693
rect 12411 659 12427 693
rect 12485 659 12501 693
rect 12609 659 12625 693
rect 12683 659 12699 693
rect 12807 659 12823 693
rect 12881 659 12897 693
rect 13005 659 13021 693
rect 13079 659 13095 693
rect 13203 659 13219 693
rect 13277 659 13293 693
rect 13401 659 13417 693
rect 13475 659 13491 693
rect 13599 659 13615 693
rect 13673 659 13689 693
rect 13797 659 13813 693
rect 13871 659 13887 693
rect 13995 659 14011 693
rect 14069 659 14085 693
rect 14193 659 14209 693
rect 14267 659 14283 693
rect 14391 659 14407 693
rect 14465 659 14481 693
rect 14589 659 14605 693
rect 14663 659 14679 693
rect 14787 659 14803 693
rect 14861 659 14877 693
rect 14985 659 15001 693
rect 15059 659 15075 693
rect 15183 659 15199 693
rect 15257 659 15273 693
rect 15381 659 15397 693
rect 15455 659 15471 693
rect 15579 659 15595 693
rect 15653 659 15669 693
rect 15777 659 15793 693
rect 15851 659 15867 693
rect 15975 659 15991 693
rect 16049 659 16065 693
rect 16173 659 16189 693
rect 16247 659 16263 693
rect 16371 659 16387 693
rect 16445 659 16461 693
rect 16569 659 16585 693
rect 16643 659 16659 693
rect 16767 659 16783 693
rect 16841 659 16857 693
rect 16965 659 16981 693
rect 17039 659 17055 693
rect 17163 659 17179 693
rect 17237 659 17253 693
rect 17361 659 17377 693
rect 17435 659 17451 693
rect 17559 659 17575 693
rect 17633 659 17649 693
rect 17757 659 17773 693
rect 17831 659 17847 693
rect 17955 659 17971 693
rect 18029 659 18045 693
rect 18153 659 18169 693
rect 18227 659 18243 693
rect 18351 659 18367 693
rect 18425 659 18441 693
rect 18549 659 18565 693
rect 18623 659 18639 693
rect 18747 659 18763 693
rect 18821 659 18837 693
rect 18945 659 18961 693
rect 19019 659 19035 693
rect 19143 659 19159 693
rect 19217 659 19233 693
rect 19341 659 19357 693
rect 19415 659 19431 693
rect 19539 659 19555 693
rect 19613 659 19629 693
rect 19737 659 19753 693
rect 11495 551 11511 585
rect 11619 551 11635 585
rect 11693 551 11709 585
rect 11817 551 11833 585
rect 11891 551 11907 585
rect 12015 551 12031 585
rect 12089 551 12105 585
rect 12213 551 12229 585
rect 12287 551 12303 585
rect 12411 551 12427 585
rect 12485 551 12501 585
rect 12609 551 12625 585
rect 12683 551 12699 585
rect 12807 551 12823 585
rect 12881 551 12897 585
rect 13005 551 13021 585
rect 13079 551 13095 585
rect 13203 551 13219 585
rect 13277 551 13293 585
rect 13401 551 13417 585
rect 13475 551 13491 585
rect 13599 551 13615 585
rect 13673 551 13689 585
rect 13797 551 13813 585
rect 13871 551 13887 585
rect 13995 551 14011 585
rect 14069 551 14085 585
rect 14193 551 14209 585
rect 14267 551 14283 585
rect 14391 551 14407 585
rect 14465 551 14481 585
rect 14589 551 14605 585
rect 14663 551 14679 585
rect 14787 551 14803 585
rect 14861 551 14877 585
rect 14985 551 15001 585
rect 15059 551 15075 585
rect 15183 551 15199 585
rect 15257 551 15273 585
rect 15381 551 15397 585
rect 15455 551 15471 585
rect 15579 551 15595 585
rect 15653 551 15669 585
rect 15777 551 15793 585
rect 15851 551 15867 585
rect 15975 551 15991 585
rect 16049 551 16065 585
rect 16173 551 16189 585
rect 16247 551 16263 585
rect 16371 551 16387 585
rect 16445 551 16461 585
rect 16569 551 16585 585
rect 16643 551 16659 585
rect 16767 551 16783 585
rect 16841 551 16857 585
rect 16965 551 16981 585
rect 17039 551 17055 585
rect 17163 551 17179 585
rect 17237 551 17253 585
rect 17361 551 17377 585
rect 17435 551 17451 585
rect 17559 551 17575 585
rect 17633 551 17649 585
rect 17757 551 17773 585
rect 17831 551 17847 585
rect 17955 551 17971 585
rect 18029 551 18045 585
rect 18153 551 18169 585
rect 18227 551 18243 585
rect 18351 551 18367 585
rect 18425 551 18441 585
rect 18549 551 18565 585
rect 18623 551 18639 585
rect 18747 551 18763 585
rect 18821 551 18837 585
rect 18945 551 18961 585
rect 19019 551 19035 585
rect 19143 551 19159 585
rect 19217 551 19233 585
rect 19341 551 19357 585
rect 19415 551 19431 585
rect 19539 551 19555 585
rect 19613 551 19629 585
rect 19737 551 19753 585
rect 11449 492 11483 508
rect 11449 -900 11483 -884
rect 11647 492 11681 508
rect 11647 -900 11681 -884
rect 11845 492 11879 508
rect 11845 -900 11879 -884
rect 12043 492 12077 508
rect 12043 -900 12077 -884
rect 12241 492 12275 508
rect 12241 -900 12275 -884
rect 12439 492 12473 508
rect 12439 -900 12473 -884
rect 12637 492 12671 508
rect 12637 -900 12671 -884
rect 12835 492 12869 508
rect 12835 -900 12869 -884
rect 13033 492 13067 508
rect 13033 -900 13067 -884
rect 13231 492 13265 508
rect 13231 -900 13265 -884
rect 13429 492 13463 508
rect 13429 -900 13463 -884
rect 13627 492 13661 508
rect 13627 -900 13661 -884
rect 13825 492 13859 508
rect 13825 -900 13859 -884
rect 14023 492 14057 508
rect 14023 -900 14057 -884
rect 14221 492 14255 508
rect 14221 -900 14255 -884
rect 14419 492 14453 508
rect 14419 -900 14453 -884
rect 14617 492 14651 508
rect 14617 -900 14651 -884
rect 14815 492 14849 508
rect 14815 -900 14849 -884
rect 15013 492 15047 508
rect 15013 -900 15047 -884
rect 15211 492 15245 508
rect 15211 -900 15245 -884
rect 15409 492 15443 508
rect 15409 -900 15443 -884
rect 15607 492 15641 508
rect 15607 -900 15641 -884
rect 15805 492 15839 508
rect 15805 -900 15839 -884
rect 16003 492 16037 508
rect 16003 -900 16037 -884
rect 16201 492 16235 508
rect 16201 -900 16235 -884
rect 16399 492 16433 508
rect 16399 -900 16433 -884
rect 16597 492 16631 508
rect 16597 -900 16631 -884
rect 16795 492 16829 508
rect 16795 -900 16829 -884
rect 16993 492 17027 508
rect 16993 -900 17027 -884
rect 17191 492 17225 508
rect 17191 -900 17225 -884
rect 17389 492 17423 508
rect 17389 -900 17423 -884
rect 17587 492 17621 508
rect 17587 -900 17621 -884
rect 17785 492 17819 508
rect 17785 -900 17819 -884
rect 17983 492 18017 508
rect 17983 -900 18017 -884
rect 18181 492 18215 508
rect 18181 -900 18215 -884
rect 18379 492 18413 508
rect 18379 -900 18413 -884
rect 18577 492 18611 508
rect 18577 -900 18611 -884
rect 18775 492 18809 508
rect 18775 -900 18809 -884
rect 18973 492 19007 508
rect 18973 -900 19007 -884
rect 19171 492 19205 508
rect 19171 -900 19205 -884
rect 19369 492 19403 508
rect 19369 -900 19403 -884
rect 19567 492 19601 508
rect 19567 -900 19601 -884
rect 19765 492 19799 508
rect 19765 -900 19799 -884
rect 11495 -977 11511 -943
rect 11619 -977 11635 -943
rect 11693 -977 11709 -943
rect 11817 -977 11833 -943
rect 11891 -977 11907 -943
rect 12015 -977 12031 -943
rect 12089 -977 12105 -943
rect 12213 -977 12229 -943
rect 12287 -977 12303 -943
rect 12411 -977 12427 -943
rect 12485 -977 12501 -943
rect 12609 -977 12625 -943
rect 12683 -977 12699 -943
rect 12807 -977 12823 -943
rect 12881 -977 12897 -943
rect 13005 -977 13021 -943
rect 13079 -977 13095 -943
rect 13203 -977 13219 -943
rect 13277 -977 13293 -943
rect 13401 -977 13417 -943
rect 13475 -977 13491 -943
rect 13599 -977 13615 -943
rect 13673 -977 13689 -943
rect 13797 -977 13813 -943
rect 13871 -977 13887 -943
rect 13995 -977 14011 -943
rect 14069 -977 14085 -943
rect 14193 -977 14209 -943
rect 14267 -977 14283 -943
rect 14391 -977 14407 -943
rect 14465 -977 14481 -943
rect 14589 -977 14605 -943
rect 14663 -977 14679 -943
rect 14787 -977 14803 -943
rect 14861 -977 14877 -943
rect 14985 -977 15001 -943
rect 15059 -977 15075 -943
rect 15183 -977 15199 -943
rect 15257 -977 15273 -943
rect 15381 -977 15397 -943
rect 15455 -977 15471 -943
rect 15579 -977 15595 -943
rect 15653 -977 15669 -943
rect 15777 -977 15793 -943
rect 15851 -977 15867 -943
rect 15975 -977 15991 -943
rect 16049 -977 16065 -943
rect 16173 -977 16189 -943
rect 16247 -977 16263 -943
rect 16371 -977 16387 -943
rect 16445 -977 16461 -943
rect 16569 -977 16585 -943
rect 16643 -977 16659 -943
rect 16767 -977 16783 -943
rect 16841 -977 16857 -943
rect 16965 -977 16981 -943
rect 17039 -977 17055 -943
rect 17163 -977 17179 -943
rect 17237 -977 17253 -943
rect 17361 -977 17377 -943
rect 17435 -977 17451 -943
rect 17559 -977 17575 -943
rect 17633 -977 17649 -943
rect 17757 -977 17773 -943
rect 17831 -977 17847 -943
rect 17955 -977 17971 -943
rect 18029 -977 18045 -943
rect 18153 -977 18169 -943
rect 18227 -977 18243 -943
rect 18351 -977 18367 -943
rect 18425 -977 18441 -943
rect 18549 -977 18565 -943
rect 18623 -977 18639 -943
rect 18747 -977 18763 -943
rect 18821 -977 18837 -943
rect 18945 -977 18961 -943
rect 19019 -977 19035 -943
rect 19143 -977 19159 -943
rect 19217 -977 19233 -943
rect 19341 -977 19357 -943
rect 19415 -977 19431 -943
rect 19539 -977 19555 -943
rect 19613 -977 19629 -943
rect 19737 -977 19753 -943
rect 11495 -1085 11511 -1051
rect 11619 -1085 11635 -1051
rect 11693 -1085 11709 -1051
rect 11817 -1085 11833 -1051
rect 11891 -1085 11907 -1051
rect 12015 -1085 12031 -1051
rect 12089 -1085 12105 -1051
rect 12213 -1085 12229 -1051
rect 12287 -1085 12303 -1051
rect 12411 -1085 12427 -1051
rect 12485 -1085 12501 -1051
rect 12609 -1085 12625 -1051
rect 12683 -1085 12699 -1051
rect 12807 -1085 12823 -1051
rect 12881 -1085 12897 -1051
rect 13005 -1085 13021 -1051
rect 13079 -1085 13095 -1051
rect 13203 -1085 13219 -1051
rect 13277 -1085 13293 -1051
rect 13401 -1085 13417 -1051
rect 13475 -1085 13491 -1051
rect 13599 -1085 13615 -1051
rect 13673 -1085 13689 -1051
rect 13797 -1085 13813 -1051
rect 13871 -1085 13887 -1051
rect 13995 -1085 14011 -1051
rect 14069 -1085 14085 -1051
rect 14193 -1085 14209 -1051
rect 14267 -1085 14283 -1051
rect 14391 -1085 14407 -1051
rect 14465 -1085 14481 -1051
rect 14589 -1085 14605 -1051
rect 14663 -1085 14679 -1051
rect 14787 -1085 14803 -1051
rect 14861 -1085 14877 -1051
rect 14985 -1085 15001 -1051
rect 15059 -1085 15075 -1051
rect 15183 -1085 15199 -1051
rect 15257 -1085 15273 -1051
rect 15381 -1085 15397 -1051
rect 15455 -1085 15471 -1051
rect 15579 -1085 15595 -1051
rect 15653 -1085 15669 -1051
rect 15777 -1085 15793 -1051
rect 15851 -1085 15867 -1051
rect 15975 -1085 15991 -1051
rect 16049 -1085 16065 -1051
rect 16173 -1085 16189 -1051
rect 16247 -1085 16263 -1051
rect 16371 -1085 16387 -1051
rect 16445 -1085 16461 -1051
rect 16569 -1085 16585 -1051
rect 16643 -1085 16659 -1051
rect 16767 -1085 16783 -1051
rect 16841 -1085 16857 -1051
rect 16965 -1085 16981 -1051
rect 17039 -1085 17055 -1051
rect 17163 -1085 17179 -1051
rect 17237 -1085 17253 -1051
rect 17361 -1085 17377 -1051
rect 17435 -1085 17451 -1051
rect 17559 -1085 17575 -1051
rect 17633 -1085 17649 -1051
rect 17757 -1085 17773 -1051
rect 17831 -1085 17847 -1051
rect 17955 -1085 17971 -1051
rect 18029 -1085 18045 -1051
rect 18153 -1085 18169 -1051
rect 18227 -1085 18243 -1051
rect 18351 -1085 18367 -1051
rect 18425 -1085 18441 -1051
rect 18549 -1085 18565 -1051
rect 18623 -1085 18639 -1051
rect 18747 -1085 18763 -1051
rect 18821 -1085 18837 -1051
rect 18945 -1085 18961 -1051
rect 19019 -1085 19035 -1051
rect 19143 -1085 19159 -1051
rect 19217 -1085 19233 -1051
rect 19341 -1085 19357 -1051
rect 19415 -1085 19431 -1051
rect 19539 -1085 19555 -1051
rect 19613 -1085 19629 -1051
rect 19737 -1085 19753 -1051
rect 11449 -1144 11483 -1128
rect 11449 -2536 11483 -2520
rect 11647 -1144 11681 -1128
rect 11647 -2536 11681 -2520
rect 11845 -1144 11879 -1128
rect 11845 -2536 11879 -2520
rect 12043 -1144 12077 -1128
rect 12043 -2536 12077 -2520
rect 12241 -1144 12275 -1128
rect 12241 -2536 12275 -2520
rect 12439 -1144 12473 -1128
rect 12439 -2536 12473 -2520
rect 12637 -1144 12671 -1128
rect 12637 -2536 12671 -2520
rect 12835 -1144 12869 -1128
rect 12835 -2536 12869 -2520
rect 13033 -1144 13067 -1128
rect 13033 -2536 13067 -2520
rect 13231 -1144 13265 -1128
rect 13231 -2536 13265 -2520
rect 13429 -1144 13463 -1128
rect 13429 -2536 13463 -2520
rect 13627 -1144 13661 -1128
rect 13627 -2536 13661 -2520
rect 13825 -1144 13859 -1128
rect 13825 -2536 13859 -2520
rect 14023 -1144 14057 -1128
rect 14023 -2536 14057 -2520
rect 14221 -1144 14255 -1128
rect 14221 -2536 14255 -2520
rect 14419 -1144 14453 -1128
rect 14419 -2536 14453 -2520
rect 14617 -1144 14651 -1128
rect 14617 -2536 14651 -2520
rect 14815 -1144 14849 -1128
rect 14815 -2536 14849 -2520
rect 15013 -1144 15047 -1128
rect 15013 -2536 15047 -2520
rect 15211 -1144 15245 -1128
rect 15211 -2536 15245 -2520
rect 15409 -1144 15443 -1128
rect 15409 -2536 15443 -2520
rect 15607 -1144 15641 -1128
rect 15607 -2536 15641 -2520
rect 15805 -1144 15839 -1128
rect 15805 -2536 15839 -2520
rect 16003 -1144 16037 -1128
rect 16003 -2536 16037 -2520
rect 16201 -1144 16235 -1128
rect 16201 -2536 16235 -2520
rect 16399 -1144 16433 -1128
rect 16399 -2536 16433 -2520
rect 16597 -1144 16631 -1128
rect 16597 -2536 16631 -2520
rect 16795 -1144 16829 -1128
rect 16795 -2536 16829 -2520
rect 16993 -1144 17027 -1128
rect 16993 -2536 17027 -2520
rect 17191 -1144 17225 -1128
rect 17191 -2536 17225 -2520
rect 17389 -1144 17423 -1128
rect 17389 -2536 17423 -2520
rect 17587 -1144 17621 -1128
rect 17587 -2536 17621 -2520
rect 17785 -1144 17819 -1128
rect 17785 -2536 17819 -2520
rect 17983 -1144 18017 -1128
rect 17983 -2536 18017 -2520
rect 18181 -1144 18215 -1128
rect 18181 -2536 18215 -2520
rect 18379 -1144 18413 -1128
rect 18379 -2536 18413 -2520
rect 18577 -1144 18611 -1128
rect 18577 -2536 18611 -2520
rect 18775 -1144 18809 -1128
rect 18775 -2536 18809 -2520
rect 18973 -1144 19007 -1128
rect 18973 -2536 19007 -2520
rect 19171 -1144 19205 -1128
rect 19171 -2536 19205 -2520
rect 19369 -1144 19403 -1128
rect 19369 -2536 19403 -2520
rect 19567 -1144 19601 -1128
rect 19567 -2536 19601 -2520
rect 19765 -1144 19799 -1128
rect 19765 -2536 19799 -2520
rect 11495 -2613 11511 -2579
rect 11619 -2613 11635 -2579
rect 11693 -2613 11709 -2579
rect 11817 -2613 11833 -2579
rect 11891 -2613 11907 -2579
rect 12015 -2613 12031 -2579
rect 12089 -2613 12105 -2579
rect 12213 -2613 12229 -2579
rect 12287 -2613 12303 -2579
rect 12411 -2613 12427 -2579
rect 12485 -2613 12501 -2579
rect 12609 -2613 12625 -2579
rect 12683 -2613 12699 -2579
rect 12807 -2613 12823 -2579
rect 12881 -2613 12897 -2579
rect 13005 -2613 13021 -2579
rect 13079 -2613 13095 -2579
rect 13203 -2613 13219 -2579
rect 13277 -2613 13293 -2579
rect 13401 -2613 13417 -2579
rect 13475 -2613 13491 -2579
rect 13599 -2613 13615 -2579
rect 13673 -2613 13689 -2579
rect 13797 -2613 13813 -2579
rect 13871 -2613 13887 -2579
rect 13995 -2613 14011 -2579
rect 14069 -2613 14085 -2579
rect 14193 -2613 14209 -2579
rect 14267 -2613 14283 -2579
rect 14391 -2613 14407 -2579
rect 14465 -2613 14481 -2579
rect 14589 -2613 14605 -2579
rect 14663 -2613 14679 -2579
rect 14787 -2613 14803 -2579
rect 14861 -2613 14877 -2579
rect 14985 -2613 15001 -2579
rect 15059 -2613 15075 -2579
rect 15183 -2613 15199 -2579
rect 15257 -2613 15273 -2579
rect 15381 -2613 15397 -2579
rect 15455 -2613 15471 -2579
rect 15579 -2613 15595 -2579
rect 15653 -2613 15669 -2579
rect 15777 -2613 15793 -2579
rect 15851 -2613 15867 -2579
rect 15975 -2613 15991 -2579
rect 16049 -2613 16065 -2579
rect 16173 -2613 16189 -2579
rect 16247 -2613 16263 -2579
rect 16371 -2613 16387 -2579
rect 16445 -2613 16461 -2579
rect 16569 -2613 16585 -2579
rect 16643 -2613 16659 -2579
rect 16767 -2613 16783 -2579
rect 16841 -2613 16857 -2579
rect 16965 -2613 16981 -2579
rect 17039 -2613 17055 -2579
rect 17163 -2613 17179 -2579
rect 17237 -2613 17253 -2579
rect 17361 -2613 17377 -2579
rect 17435 -2613 17451 -2579
rect 17559 -2613 17575 -2579
rect 17633 -2613 17649 -2579
rect 17757 -2613 17773 -2579
rect 17831 -2613 17847 -2579
rect 17955 -2613 17971 -2579
rect 18029 -2613 18045 -2579
rect 18153 -2613 18169 -2579
rect 18227 -2613 18243 -2579
rect 18351 -2613 18367 -2579
rect 18425 -2613 18441 -2579
rect 18549 -2613 18565 -2579
rect 18623 -2613 18639 -2579
rect 18747 -2613 18763 -2579
rect 18821 -2613 18837 -2579
rect 18945 -2613 18961 -2579
rect 19019 -2613 19035 -2579
rect 19143 -2613 19159 -2579
rect 19217 -2613 19233 -2579
rect 19341 -2613 19357 -2579
rect 19415 -2613 19431 -2579
rect 19539 -2613 19555 -2579
rect 19613 -2613 19629 -2579
rect 19737 -2613 19753 -2579
rect 11495 -2721 11511 -2687
rect 11619 -2721 11635 -2687
rect 11693 -2721 11709 -2687
rect 11817 -2721 11833 -2687
rect 11891 -2721 11907 -2687
rect 12015 -2721 12031 -2687
rect 12089 -2721 12105 -2687
rect 12213 -2721 12229 -2687
rect 12287 -2721 12303 -2687
rect 12411 -2721 12427 -2687
rect 12485 -2721 12501 -2687
rect 12609 -2721 12625 -2687
rect 12683 -2721 12699 -2687
rect 12807 -2721 12823 -2687
rect 12881 -2721 12897 -2687
rect 13005 -2721 13021 -2687
rect 13079 -2721 13095 -2687
rect 13203 -2721 13219 -2687
rect 13277 -2721 13293 -2687
rect 13401 -2721 13417 -2687
rect 13475 -2721 13491 -2687
rect 13599 -2721 13615 -2687
rect 13673 -2721 13689 -2687
rect 13797 -2721 13813 -2687
rect 13871 -2721 13887 -2687
rect 13995 -2721 14011 -2687
rect 14069 -2721 14085 -2687
rect 14193 -2721 14209 -2687
rect 14267 -2721 14283 -2687
rect 14391 -2721 14407 -2687
rect 14465 -2721 14481 -2687
rect 14589 -2721 14605 -2687
rect 14663 -2721 14679 -2687
rect 14787 -2721 14803 -2687
rect 14861 -2721 14877 -2687
rect 14985 -2721 15001 -2687
rect 15059 -2721 15075 -2687
rect 15183 -2721 15199 -2687
rect 15257 -2721 15273 -2687
rect 15381 -2721 15397 -2687
rect 15455 -2721 15471 -2687
rect 15579 -2721 15595 -2687
rect 15653 -2721 15669 -2687
rect 15777 -2721 15793 -2687
rect 15851 -2721 15867 -2687
rect 15975 -2721 15991 -2687
rect 16049 -2721 16065 -2687
rect 16173 -2721 16189 -2687
rect 16247 -2721 16263 -2687
rect 16371 -2721 16387 -2687
rect 16445 -2721 16461 -2687
rect 16569 -2721 16585 -2687
rect 16643 -2721 16659 -2687
rect 16767 -2721 16783 -2687
rect 16841 -2721 16857 -2687
rect 16965 -2721 16981 -2687
rect 17039 -2721 17055 -2687
rect 17163 -2721 17179 -2687
rect 17237 -2721 17253 -2687
rect 17361 -2721 17377 -2687
rect 17435 -2721 17451 -2687
rect 17559 -2721 17575 -2687
rect 17633 -2721 17649 -2687
rect 17757 -2721 17773 -2687
rect 17831 -2721 17847 -2687
rect 17955 -2721 17971 -2687
rect 18029 -2721 18045 -2687
rect 18153 -2721 18169 -2687
rect 18227 -2721 18243 -2687
rect 18351 -2721 18367 -2687
rect 18425 -2721 18441 -2687
rect 18549 -2721 18565 -2687
rect 18623 -2721 18639 -2687
rect 18747 -2721 18763 -2687
rect 18821 -2721 18837 -2687
rect 18945 -2721 18961 -2687
rect 19019 -2721 19035 -2687
rect 19143 -2721 19159 -2687
rect 19217 -2721 19233 -2687
rect 19341 -2721 19357 -2687
rect 19415 -2721 19431 -2687
rect 19539 -2721 19555 -2687
rect 19613 -2721 19629 -2687
rect 19737 -2721 19753 -2687
rect 11449 -2780 11483 -2764
rect 11449 -4172 11483 -4156
rect 11647 -2780 11681 -2764
rect 11647 -4172 11681 -4156
rect 11845 -2780 11879 -2764
rect 11845 -4172 11879 -4156
rect 12043 -2780 12077 -2764
rect 12043 -4172 12077 -4156
rect 12241 -2780 12275 -2764
rect 12241 -4172 12275 -4156
rect 12439 -2780 12473 -2764
rect 12439 -4172 12473 -4156
rect 12637 -2780 12671 -2764
rect 12637 -4172 12671 -4156
rect 12835 -2780 12869 -2764
rect 12835 -4172 12869 -4156
rect 13033 -2780 13067 -2764
rect 13033 -4172 13067 -4156
rect 13231 -2780 13265 -2764
rect 13231 -4172 13265 -4156
rect 13429 -2780 13463 -2764
rect 13429 -4172 13463 -4156
rect 13627 -2780 13661 -2764
rect 13627 -4172 13661 -4156
rect 13825 -2780 13859 -2764
rect 13825 -4172 13859 -4156
rect 14023 -2780 14057 -2764
rect 14023 -4172 14057 -4156
rect 14221 -2780 14255 -2764
rect 14221 -4172 14255 -4156
rect 14419 -2780 14453 -2764
rect 14419 -4172 14453 -4156
rect 14617 -2780 14651 -2764
rect 14617 -4172 14651 -4156
rect 14815 -2780 14849 -2764
rect 14815 -4172 14849 -4156
rect 15013 -2780 15047 -2764
rect 15013 -4172 15047 -4156
rect 15211 -2780 15245 -2764
rect 15211 -4172 15245 -4156
rect 15409 -2780 15443 -2764
rect 15409 -4172 15443 -4156
rect 15607 -2780 15641 -2764
rect 15607 -4172 15641 -4156
rect 15805 -2780 15839 -2764
rect 15805 -4172 15839 -4156
rect 16003 -2780 16037 -2764
rect 16003 -4172 16037 -4156
rect 16201 -2780 16235 -2764
rect 16201 -4172 16235 -4156
rect 16399 -2780 16433 -2764
rect 16399 -4172 16433 -4156
rect 16597 -2780 16631 -2764
rect 16597 -4172 16631 -4156
rect 16795 -2780 16829 -2764
rect 16795 -4172 16829 -4156
rect 16993 -2780 17027 -2764
rect 16993 -4172 17027 -4156
rect 17191 -2780 17225 -2764
rect 17191 -4172 17225 -4156
rect 17389 -2780 17423 -2764
rect 17389 -4172 17423 -4156
rect 17587 -2780 17621 -2764
rect 17587 -4172 17621 -4156
rect 17785 -2780 17819 -2764
rect 17785 -4172 17819 -4156
rect 17983 -2780 18017 -2764
rect 17983 -4172 18017 -4156
rect 18181 -2780 18215 -2764
rect 18181 -4172 18215 -4156
rect 18379 -2780 18413 -2764
rect 18379 -4172 18413 -4156
rect 18577 -2780 18611 -2764
rect 18577 -4172 18611 -4156
rect 18775 -2780 18809 -2764
rect 18775 -4172 18809 -4156
rect 18973 -2780 19007 -2764
rect 18973 -4172 19007 -4156
rect 19171 -2780 19205 -2764
rect 19171 -4172 19205 -4156
rect 19369 -2780 19403 -2764
rect 19369 -4172 19403 -4156
rect 19567 -2780 19601 -2764
rect 19567 -4172 19601 -4156
rect 19765 -2780 19799 -2764
rect 19765 -4172 19799 -4156
rect 10991 -4415 11025 -4353
rect 20238 -4415 20272 -4353
rect 10991 -4449 11087 -4415
rect 20176 -4449 20272 -4415
rect 22841 2237 22937 2271
rect 32026 2237 32122 2271
rect 22841 2175 22875 2237
rect 32088 2175 32122 2237
rect 23299 2128 23333 2144
rect 23299 736 23333 752
rect 23497 2128 23531 2144
rect 23497 736 23531 752
rect 23695 2128 23729 2144
rect 23695 736 23729 752
rect 23893 2128 23927 2144
rect 23893 736 23927 752
rect 24091 2128 24125 2144
rect 24091 736 24125 752
rect 24289 2128 24323 2144
rect 24289 736 24323 752
rect 24487 2128 24521 2144
rect 24487 736 24521 752
rect 24685 2128 24719 2144
rect 24685 736 24719 752
rect 24883 2128 24917 2144
rect 24883 736 24917 752
rect 25081 2128 25115 2144
rect 25081 736 25115 752
rect 25279 2128 25313 2144
rect 25279 736 25313 752
rect 25477 2128 25511 2144
rect 25477 736 25511 752
rect 25675 2128 25709 2144
rect 25675 736 25709 752
rect 25873 2128 25907 2144
rect 25873 736 25907 752
rect 26071 2128 26105 2144
rect 26071 736 26105 752
rect 26269 2128 26303 2144
rect 26269 736 26303 752
rect 26467 2128 26501 2144
rect 26467 736 26501 752
rect 26665 2128 26699 2144
rect 26665 736 26699 752
rect 26863 2128 26897 2144
rect 26863 736 26897 752
rect 27061 2128 27095 2144
rect 27061 736 27095 752
rect 27259 2128 27293 2144
rect 27259 736 27293 752
rect 27457 2128 27491 2144
rect 27457 736 27491 752
rect 27655 2128 27689 2144
rect 27655 736 27689 752
rect 27853 2128 27887 2144
rect 27853 736 27887 752
rect 28051 2128 28085 2144
rect 28051 736 28085 752
rect 28249 2128 28283 2144
rect 28249 736 28283 752
rect 28447 2128 28481 2144
rect 28447 736 28481 752
rect 28645 2128 28679 2144
rect 28645 736 28679 752
rect 28843 2128 28877 2144
rect 28843 736 28877 752
rect 29041 2128 29075 2144
rect 29041 736 29075 752
rect 29239 2128 29273 2144
rect 29239 736 29273 752
rect 29437 2128 29471 2144
rect 29437 736 29471 752
rect 29635 2128 29669 2144
rect 29635 736 29669 752
rect 29833 2128 29867 2144
rect 29833 736 29867 752
rect 30031 2128 30065 2144
rect 30031 736 30065 752
rect 30229 2128 30263 2144
rect 30229 736 30263 752
rect 30427 2128 30461 2144
rect 30427 736 30461 752
rect 30625 2128 30659 2144
rect 30625 736 30659 752
rect 30823 2128 30857 2144
rect 30823 736 30857 752
rect 31021 2128 31055 2144
rect 31021 736 31055 752
rect 31219 2128 31253 2144
rect 31219 736 31253 752
rect 31417 2128 31451 2144
rect 31417 736 31451 752
rect 31615 2128 31649 2144
rect 31615 736 31649 752
rect 23345 659 23361 693
rect 23469 659 23485 693
rect 23543 659 23559 693
rect 23667 659 23683 693
rect 23741 659 23757 693
rect 23865 659 23881 693
rect 23939 659 23955 693
rect 24063 659 24079 693
rect 24137 659 24153 693
rect 24261 659 24277 693
rect 24335 659 24351 693
rect 24459 659 24475 693
rect 24533 659 24549 693
rect 24657 659 24673 693
rect 24731 659 24747 693
rect 24855 659 24871 693
rect 24929 659 24945 693
rect 25053 659 25069 693
rect 25127 659 25143 693
rect 25251 659 25267 693
rect 25325 659 25341 693
rect 25449 659 25465 693
rect 25523 659 25539 693
rect 25647 659 25663 693
rect 25721 659 25737 693
rect 25845 659 25861 693
rect 25919 659 25935 693
rect 26043 659 26059 693
rect 26117 659 26133 693
rect 26241 659 26257 693
rect 26315 659 26331 693
rect 26439 659 26455 693
rect 26513 659 26529 693
rect 26637 659 26653 693
rect 26711 659 26727 693
rect 26835 659 26851 693
rect 26909 659 26925 693
rect 27033 659 27049 693
rect 27107 659 27123 693
rect 27231 659 27247 693
rect 27305 659 27321 693
rect 27429 659 27445 693
rect 27503 659 27519 693
rect 27627 659 27643 693
rect 27701 659 27717 693
rect 27825 659 27841 693
rect 27899 659 27915 693
rect 28023 659 28039 693
rect 28097 659 28113 693
rect 28221 659 28237 693
rect 28295 659 28311 693
rect 28419 659 28435 693
rect 28493 659 28509 693
rect 28617 659 28633 693
rect 28691 659 28707 693
rect 28815 659 28831 693
rect 28889 659 28905 693
rect 29013 659 29029 693
rect 29087 659 29103 693
rect 29211 659 29227 693
rect 29285 659 29301 693
rect 29409 659 29425 693
rect 29483 659 29499 693
rect 29607 659 29623 693
rect 29681 659 29697 693
rect 29805 659 29821 693
rect 29879 659 29895 693
rect 30003 659 30019 693
rect 30077 659 30093 693
rect 30201 659 30217 693
rect 30275 659 30291 693
rect 30399 659 30415 693
rect 30473 659 30489 693
rect 30597 659 30613 693
rect 30671 659 30687 693
rect 30795 659 30811 693
rect 30869 659 30885 693
rect 30993 659 31009 693
rect 31067 659 31083 693
rect 31191 659 31207 693
rect 31265 659 31281 693
rect 31389 659 31405 693
rect 31463 659 31479 693
rect 31587 659 31603 693
rect 23345 551 23361 585
rect 23469 551 23485 585
rect 23543 551 23559 585
rect 23667 551 23683 585
rect 23741 551 23757 585
rect 23865 551 23881 585
rect 23939 551 23955 585
rect 24063 551 24079 585
rect 24137 551 24153 585
rect 24261 551 24277 585
rect 24335 551 24351 585
rect 24459 551 24475 585
rect 24533 551 24549 585
rect 24657 551 24673 585
rect 24731 551 24747 585
rect 24855 551 24871 585
rect 24929 551 24945 585
rect 25053 551 25069 585
rect 25127 551 25143 585
rect 25251 551 25267 585
rect 25325 551 25341 585
rect 25449 551 25465 585
rect 25523 551 25539 585
rect 25647 551 25663 585
rect 25721 551 25737 585
rect 25845 551 25861 585
rect 25919 551 25935 585
rect 26043 551 26059 585
rect 26117 551 26133 585
rect 26241 551 26257 585
rect 26315 551 26331 585
rect 26439 551 26455 585
rect 26513 551 26529 585
rect 26637 551 26653 585
rect 26711 551 26727 585
rect 26835 551 26851 585
rect 26909 551 26925 585
rect 27033 551 27049 585
rect 27107 551 27123 585
rect 27231 551 27247 585
rect 27305 551 27321 585
rect 27429 551 27445 585
rect 27503 551 27519 585
rect 27627 551 27643 585
rect 27701 551 27717 585
rect 27825 551 27841 585
rect 27899 551 27915 585
rect 28023 551 28039 585
rect 28097 551 28113 585
rect 28221 551 28237 585
rect 28295 551 28311 585
rect 28419 551 28435 585
rect 28493 551 28509 585
rect 28617 551 28633 585
rect 28691 551 28707 585
rect 28815 551 28831 585
rect 28889 551 28905 585
rect 29013 551 29029 585
rect 29087 551 29103 585
rect 29211 551 29227 585
rect 29285 551 29301 585
rect 29409 551 29425 585
rect 29483 551 29499 585
rect 29607 551 29623 585
rect 29681 551 29697 585
rect 29805 551 29821 585
rect 29879 551 29895 585
rect 30003 551 30019 585
rect 30077 551 30093 585
rect 30201 551 30217 585
rect 30275 551 30291 585
rect 30399 551 30415 585
rect 30473 551 30489 585
rect 30597 551 30613 585
rect 30671 551 30687 585
rect 30795 551 30811 585
rect 30869 551 30885 585
rect 30993 551 31009 585
rect 31067 551 31083 585
rect 31191 551 31207 585
rect 31265 551 31281 585
rect 31389 551 31405 585
rect 31463 551 31479 585
rect 31587 551 31603 585
rect 23299 492 23333 508
rect 23299 -900 23333 -884
rect 23497 492 23531 508
rect 23497 -900 23531 -884
rect 23695 492 23729 508
rect 23695 -900 23729 -884
rect 23893 492 23927 508
rect 23893 -900 23927 -884
rect 24091 492 24125 508
rect 24091 -900 24125 -884
rect 24289 492 24323 508
rect 24289 -900 24323 -884
rect 24487 492 24521 508
rect 24487 -900 24521 -884
rect 24685 492 24719 508
rect 24685 -900 24719 -884
rect 24883 492 24917 508
rect 24883 -900 24917 -884
rect 25081 492 25115 508
rect 25081 -900 25115 -884
rect 25279 492 25313 508
rect 25279 -900 25313 -884
rect 25477 492 25511 508
rect 25477 -900 25511 -884
rect 25675 492 25709 508
rect 25675 -900 25709 -884
rect 25873 492 25907 508
rect 25873 -900 25907 -884
rect 26071 492 26105 508
rect 26071 -900 26105 -884
rect 26269 492 26303 508
rect 26269 -900 26303 -884
rect 26467 492 26501 508
rect 26467 -900 26501 -884
rect 26665 492 26699 508
rect 26665 -900 26699 -884
rect 26863 492 26897 508
rect 26863 -900 26897 -884
rect 27061 492 27095 508
rect 27061 -900 27095 -884
rect 27259 492 27293 508
rect 27259 -900 27293 -884
rect 27457 492 27491 508
rect 27457 -900 27491 -884
rect 27655 492 27689 508
rect 27655 -900 27689 -884
rect 27853 492 27887 508
rect 27853 -900 27887 -884
rect 28051 492 28085 508
rect 28051 -900 28085 -884
rect 28249 492 28283 508
rect 28249 -900 28283 -884
rect 28447 492 28481 508
rect 28447 -900 28481 -884
rect 28645 492 28679 508
rect 28645 -900 28679 -884
rect 28843 492 28877 508
rect 28843 -900 28877 -884
rect 29041 492 29075 508
rect 29041 -900 29075 -884
rect 29239 492 29273 508
rect 29239 -900 29273 -884
rect 29437 492 29471 508
rect 29437 -900 29471 -884
rect 29635 492 29669 508
rect 29635 -900 29669 -884
rect 29833 492 29867 508
rect 29833 -900 29867 -884
rect 30031 492 30065 508
rect 30031 -900 30065 -884
rect 30229 492 30263 508
rect 30229 -900 30263 -884
rect 30427 492 30461 508
rect 30427 -900 30461 -884
rect 30625 492 30659 508
rect 30625 -900 30659 -884
rect 30823 492 30857 508
rect 30823 -900 30857 -884
rect 31021 492 31055 508
rect 31021 -900 31055 -884
rect 31219 492 31253 508
rect 31219 -900 31253 -884
rect 31417 492 31451 508
rect 31417 -900 31451 -884
rect 31615 492 31649 508
rect 31615 -900 31649 -884
rect 23345 -977 23361 -943
rect 23469 -977 23485 -943
rect 23543 -977 23559 -943
rect 23667 -977 23683 -943
rect 23741 -977 23757 -943
rect 23865 -977 23881 -943
rect 23939 -977 23955 -943
rect 24063 -977 24079 -943
rect 24137 -977 24153 -943
rect 24261 -977 24277 -943
rect 24335 -977 24351 -943
rect 24459 -977 24475 -943
rect 24533 -977 24549 -943
rect 24657 -977 24673 -943
rect 24731 -977 24747 -943
rect 24855 -977 24871 -943
rect 24929 -977 24945 -943
rect 25053 -977 25069 -943
rect 25127 -977 25143 -943
rect 25251 -977 25267 -943
rect 25325 -977 25341 -943
rect 25449 -977 25465 -943
rect 25523 -977 25539 -943
rect 25647 -977 25663 -943
rect 25721 -977 25737 -943
rect 25845 -977 25861 -943
rect 25919 -977 25935 -943
rect 26043 -977 26059 -943
rect 26117 -977 26133 -943
rect 26241 -977 26257 -943
rect 26315 -977 26331 -943
rect 26439 -977 26455 -943
rect 26513 -977 26529 -943
rect 26637 -977 26653 -943
rect 26711 -977 26727 -943
rect 26835 -977 26851 -943
rect 26909 -977 26925 -943
rect 27033 -977 27049 -943
rect 27107 -977 27123 -943
rect 27231 -977 27247 -943
rect 27305 -977 27321 -943
rect 27429 -977 27445 -943
rect 27503 -977 27519 -943
rect 27627 -977 27643 -943
rect 27701 -977 27717 -943
rect 27825 -977 27841 -943
rect 27899 -977 27915 -943
rect 28023 -977 28039 -943
rect 28097 -977 28113 -943
rect 28221 -977 28237 -943
rect 28295 -977 28311 -943
rect 28419 -977 28435 -943
rect 28493 -977 28509 -943
rect 28617 -977 28633 -943
rect 28691 -977 28707 -943
rect 28815 -977 28831 -943
rect 28889 -977 28905 -943
rect 29013 -977 29029 -943
rect 29087 -977 29103 -943
rect 29211 -977 29227 -943
rect 29285 -977 29301 -943
rect 29409 -977 29425 -943
rect 29483 -977 29499 -943
rect 29607 -977 29623 -943
rect 29681 -977 29697 -943
rect 29805 -977 29821 -943
rect 29879 -977 29895 -943
rect 30003 -977 30019 -943
rect 30077 -977 30093 -943
rect 30201 -977 30217 -943
rect 30275 -977 30291 -943
rect 30399 -977 30415 -943
rect 30473 -977 30489 -943
rect 30597 -977 30613 -943
rect 30671 -977 30687 -943
rect 30795 -977 30811 -943
rect 30869 -977 30885 -943
rect 30993 -977 31009 -943
rect 31067 -977 31083 -943
rect 31191 -977 31207 -943
rect 31265 -977 31281 -943
rect 31389 -977 31405 -943
rect 31463 -977 31479 -943
rect 31587 -977 31603 -943
rect 23345 -1085 23361 -1051
rect 23469 -1085 23485 -1051
rect 23543 -1085 23559 -1051
rect 23667 -1085 23683 -1051
rect 23741 -1085 23757 -1051
rect 23865 -1085 23881 -1051
rect 23939 -1085 23955 -1051
rect 24063 -1085 24079 -1051
rect 24137 -1085 24153 -1051
rect 24261 -1085 24277 -1051
rect 24335 -1085 24351 -1051
rect 24459 -1085 24475 -1051
rect 24533 -1085 24549 -1051
rect 24657 -1085 24673 -1051
rect 24731 -1085 24747 -1051
rect 24855 -1085 24871 -1051
rect 24929 -1085 24945 -1051
rect 25053 -1085 25069 -1051
rect 25127 -1085 25143 -1051
rect 25251 -1085 25267 -1051
rect 25325 -1085 25341 -1051
rect 25449 -1085 25465 -1051
rect 25523 -1085 25539 -1051
rect 25647 -1085 25663 -1051
rect 25721 -1085 25737 -1051
rect 25845 -1085 25861 -1051
rect 25919 -1085 25935 -1051
rect 26043 -1085 26059 -1051
rect 26117 -1085 26133 -1051
rect 26241 -1085 26257 -1051
rect 26315 -1085 26331 -1051
rect 26439 -1085 26455 -1051
rect 26513 -1085 26529 -1051
rect 26637 -1085 26653 -1051
rect 26711 -1085 26727 -1051
rect 26835 -1085 26851 -1051
rect 26909 -1085 26925 -1051
rect 27033 -1085 27049 -1051
rect 27107 -1085 27123 -1051
rect 27231 -1085 27247 -1051
rect 27305 -1085 27321 -1051
rect 27429 -1085 27445 -1051
rect 27503 -1085 27519 -1051
rect 27627 -1085 27643 -1051
rect 27701 -1085 27717 -1051
rect 27825 -1085 27841 -1051
rect 27899 -1085 27915 -1051
rect 28023 -1085 28039 -1051
rect 28097 -1085 28113 -1051
rect 28221 -1085 28237 -1051
rect 28295 -1085 28311 -1051
rect 28419 -1085 28435 -1051
rect 28493 -1085 28509 -1051
rect 28617 -1085 28633 -1051
rect 28691 -1085 28707 -1051
rect 28815 -1085 28831 -1051
rect 28889 -1085 28905 -1051
rect 29013 -1085 29029 -1051
rect 29087 -1085 29103 -1051
rect 29211 -1085 29227 -1051
rect 29285 -1085 29301 -1051
rect 29409 -1085 29425 -1051
rect 29483 -1085 29499 -1051
rect 29607 -1085 29623 -1051
rect 29681 -1085 29697 -1051
rect 29805 -1085 29821 -1051
rect 29879 -1085 29895 -1051
rect 30003 -1085 30019 -1051
rect 30077 -1085 30093 -1051
rect 30201 -1085 30217 -1051
rect 30275 -1085 30291 -1051
rect 30399 -1085 30415 -1051
rect 30473 -1085 30489 -1051
rect 30597 -1085 30613 -1051
rect 30671 -1085 30687 -1051
rect 30795 -1085 30811 -1051
rect 30869 -1085 30885 -1051
rect 30993 -1085 31009 -1051
rect 31067 -1085 31083 -1051
rect 31191 -1085 31207 -1051
rect 31265 -1085 31281 -1051
rect 31389 -1085 31405 -1051
rect 31463 -1085 31479 -1051
rect 31587 -1085 31603 -1051
rect 23299 -1144 23333 -1128
rect 23299 -2536 23333 -2520
rect 23497 -1144 23531 -1128
rect 23497 -2536 23531 -2520
rect 23695 -1144 23729 -1128
rect 23695 -2536 23729 -2520
rect 23893 -1144 23927 -1128
rect 23893 -2536 23927 -2520
rect 24091 -1144 24125 -1128
rect 24091 -2536 24125 -2520
rect 24289 -1144 24323 -1128
rect 24289 -2536 24323 -2520
rect 24487 -1144 24521 -1128
rect 24487 -2536 24521 -2520
rect 24685 -1144 24719 -1128
rect 24685 -2536 24719 -2520
rect 24883 -1144 24917 -1128
rect 24883 -2536 24917 -2520
rect 25081 -1144 25115 -1128
rect 25081 -2536 25115 -2520
rect 25279 -1144 25313 -1128
rect 25279 -2536 25313 -2520
rect 25477 -1144 25511 -1128
rect 25477 -2536 25511 -2520
rect 25675 -1144 25709 -1128
rect 25675 -2536 25709 -2520
rect 25873 -1144 25907 -1128
rect 25873 -2536 25907 -2520
rect 26071 -1144 26105 -1128
rect 26071 -2536 26105 -2520
rect 26269 -1144 26303 -1128
rect 26269 -2536 26303 -2520
rect 26467 -1144 26501 -1128
rect 26467 -2536 26501 -2520
rect 26665 -1144 26699 -1128
rect 26665 -2536 26699 -2520
rect 26863 -1144 26897 -1128
rect 26863 -2536 26897 -2520
rect 27061 -1144 27095 -1128
rect 27061 -2536 27095 -2520
rect 27259 -1144 27293 -1128
rect 27259 -2536 27293 -2520
rect 27457 -1144 27491 -1128
rect 27457 -2536 27491 -2520
rect 27655 -1144 27689 -1128
rect 27655 -2536 27689 -2520
rect 27853 -1144 27887 -1128
rect 27853 -2536 27887 -2520
rect 28051 -1144 28085 -1128
rect 28051 -2536 28085 -2520
rect 28249 -1144 28283 -1128
rect 28249 -2536 28283 -2520
rect 28447 -1144 28481 -1128
rect 28447 -2536 28481 -2520
rect 28645 -1144 28679 -1128
rect 28645 -2536 28679 -2520
rect 28843 -1144 28877 -1128
rect 28843 -2536 28877 -2520
rect 29041 -1144 29075 -1128
rect 29041 -2536 29075 -2520
rect 29239 -1144 29273 -1128
rect 29239 -2536 29273 -2520
rect 29437 -1144 29471 -1128
rect 29437 -2536 29471 -2520
rect 29635 -1144 29669 -1128
rect 29635 -2536 29669 -2520
rect 29833 -1144 29867 -1128
rect 29833 -2536 29867 -2520
rect 30031 -1144 30065 -1128
rect 30031 -2536 30065 -2520
rect 30229 -1144 30263 -1128
rect 30229 -2536 30263 -2520
rect 30427 -1144 30461 -1128
rect 30427 -2536 30461 -2520
rect 30625 -1144 30659 -1128
rect 30625 -2536 30659 -2520
rect 30823 -1144 30857 -1128
rect 30823 -2536 30857 -2520
rect 31021 -1144 31055 -1128
rect 31021 -2536 31055 -2520
rect 31219 -1144 31253 -1128
rect 31219 -2536 31253 -2520
rect 31417 -1144 31451 -1128
rect 31417 -2536 31451 -2520
rect 31615 -1144 31649 -1128
rect 31615 -2536 31649 -2520
rect 23345 -2613 23361 -2579
rect 23469 -2613 23485 -2579
rect 23543 -2613 23559 -2579
rect 23667 -2613 23683 -2579
rect 23741 -2613 23757 -2579
rect 23865 -2613 23881 -2579
rect 23939 -2613 23955 -2579
rect 24063 -2613 24079 -2579
rect 24137 -2613 24153 -2579
rect 24261 -2613 24277 -2579
rect 24335 -2613 24351 -2579
rect 24459 -2613 24475 -2579
rect 24533 -2613 24549 -2579
rect 24657 -2613 24673 -2579
rect 24731 -2613 24747 -2579
rect 24855 -2613 24871 -2579
rect 24929 -2613 24945 -2579
rect 25053 -2613 25069 -2579
rect 25127 -2613 25143 -2579
rect 25251 -2613 25267 -2579
rect 25325 -2613 25341 -2579
rect 25449 -2613 25465 -2579
rect 25523 -2613 25539 -2579
rect 25647 -2613 25663 -2579
rect 25721 -2613 25737 -2579
rect 25845 -2613 25861 -2579
rect 25919 -2613 25935 -2579
rect 26043 -2613 26059 -2579
rect 26117 -2613 26133 -2579
rect 26241 -2613 26257 -2579
rect 26315 -2613 26331 -2579
rect 26439 -2613 26455 -2579
rect 26513 -2613 26529 -2579
rect 26637 -2613 26653 -2579
rect 26711 -2613 26727 -2579
rect 26835 -2613 26851 -2579
rect 26909 -2613 26925 -2579
rect 27033 -2613 27049 -2579
rect 27107 -2613 27123 -2579
rect 27231 -2613 27247 -2579
rect 27305 -2613 27321 -2579
rect 27429 -2613 27445 -2579
rect 27503 -2613 27519 -2579
rect 27627 -2613 27643 -2579
rect 27701 -2613 27717 -2579
rect 27825 -2613 27841 -2579
rect 27899 -2613 27915 -2579
rect 28023 -2613 28039 -2579
rect 28097 -2613 28113 -2579
rect 28221 -2613 28237 -2579
rect 28295 -2613 28311 -2579
rect 28419 -2613 28435 -2579
rect 28493 -2613 28509 -2579
rect 28617 -2613 28633 -2579
rect 28691 -2613 28707 -2579
rect 28815 -2613 28831 -2579
rect 28889 -2613 28905 -2579
rect 29013 -2613 29029 -2579
rect 29087 -2613 29103 -2579
rect 29211 -2613 29227 -2579
rect 29285 -2613 29301 -2579
rect 29409 -2613 29425 -2579
rect 29483 -2613 29499 -2579
rect 29607 -2613 29623 -2579
rect 29681 -2613 29697 -2579
rect 29805 -2613 29821 -2579
rect 29879 -2613 29895 -2579
rect 30003 -2613 30019 -2579
rect 30077 -2613 30093 -2579
rect 30201 -2613 30217 -2579
rect 30275 -2613 30291 -2579
rect 30399 -2613 30415 -2579
rect 30473 -2613 30489 -2579
rect 30597 -2613 30613 -2579
rect 30671 -2613 30687 -2579
rect 30795 -2613 30811 -2579
rect 30869 -2613 30885 -2579
rect 30993 -2613 31009 -2579
rect 31067 -2613 31083 -2579
rect 31191 -2613 31207 -2579
rect 31265 -2613 31281 -2579
rect 31389 -2613 31405 -2579
rect 31463 -2613 31479 -2579
rect 31587 -2613 31603 -2579
rect 23345 -2721 23361 -2687
rect 23469 -2721 23485 -2687
rect 23543 -2721 23559 -2687
rect 23667 -2721 23683 -2687
rect 23741 -2721 23757 -2687
rect 23865 -2721 23881 -2687
rect 23939 -2721 23955 -2687
rect 24063 -2721 24079 -2687
rect 24137 -2721 24153 -2687
rect 24261 -2721 24277 -2687
rect 24335 -2721 24351 -2687
rect 24459 -2721 24475 -2687
rect 24533 -2721 24549 -2687
rect 24657 -2721 24673 -2687
rect 24731 -2721 24747 -2687
rect 24855 -2721 24871 -2687
rect 24929 -2721 24945 -2687
rect 25053 -2721 25069 -2687
rect 25127 -2721 25143 -2687
rect 25251 -2721 25267 -2687
rect 25325 -2721 25341 -2687
rect 25449 -2721 25465 -2687
rect 25523 -2721 25539 -2687
rect 25647 -2721 25663 -2687
rect 25721 -2721 25737 -2687
rect 25845 -2721 25861 -2687
rect 25919 -2721 25935 -2687
rect 26043 -2721 26059 -2687
rect 26117 -2721 26133 -2687
rect 26241 -2721 26257 -2687
rect 26315 -2721 26331 -2687
rect 26439 -2721 26455 -2687
rect 26513 -2721 26529 -2687
rect 26637 -2721 26653 -2687
rect 26711 -2721 26727 -2687
rect 26835 -2721 26851 -2687
rect 26909 -2721 26925 -2687
rect 27033 -2721 27049 -2687
rect 27107 -2721 27123 -2687
rect 27231 -2721 27247 -2687
rect 27305 -2721 27321 -2687
rect 27429 -2721 27445 -2687
rect 27503 -2721 27519 -2687
rect 27627 -2721 27643 -2687
rect 27701 -2721 27717 -2687
rect 27825 -2721 27841 -2687
rect 27899 -2721 27915 -2687
rect 28023 -2721 28039 -2687
rect 28097 -2721 28113 -2687
rect 28221 -2721 28237 -2687
rect 28295 -2721 28311 -2687
rect 28419 -2721 28435 -2687
rect 28493 -2721 28509 -2687
rect 28617 -2721 28633 -2687
rect 28691 -2721 28707 -2687
rect 28815 -2721 28831 -2687
rect 28889 -2721 28905 -2687
rect 29013 -2721 29029 -2687
rect 29087 -2721 29103 -2687
rect 29211 -2721 29227 -2687
rect 29285 -2721 29301 -2687
rect 29409 -2721 29425 -2687
rect 29483 -2721 29499 -2687
rect 29607 -2721 29623 -2687
rect 29681 -2721 29697 -2687
rect 29805 -2721 29821 -2687
rect 29879 -2721 29895 -2687
rect 30003 -2721 30019 -2687
rect 30077 -2721 30093 -2687
rect 30201 -2721 30217 -2687
rect 30275 -2721 30291 -2687
rect 30399 -2721 30415 -2687
rect 30473 -2721 30489 -2687
rect 30597 -2721 30613 -2687
rect 30671 -2721 30687 -2687
rect 30795 -2721 30811 -2687
rect 30869 -2721 30885 -2687
rect 30993 -2721 31009 -2687
rect 31067 -2721 31083 -2687
rect 31191 -2721 31207 -2687
rect 31265 -2721 31281 -2687
rect 31389 -2721 31405 -2687
rect 31463 -2721 31479 -2687
rect 31587 -2721 31603 -2687
rect 23299 -2780 23333 -2764
rect 23299 -4172 23333 -4156
rect 23497 -2780 23531 -2764
rect 23497 -4172 23531 -4156
rect 23695 -2780 23729 -2764
rect 23695 -4172 23729 -4156
rect 23893 -2780 23927 -2764
rect 23893 -4172 23927 -4156
rect 24091 -2780 24125 -2764
rect 24091 -4172 24125 -4156
rect 24289 -2780 24323 -2764
rect 24289 -4172 24323 -4156
rect 24487 -2780 24521 -2764
rect 24487 -4172 24521 -4156
rect 24685 -2780 24719 -2764
rect 24685 -4172 24719 -4156
rect 24883 -2780 24917 -2764
rect 24883 -4172 24917 -4156
rect 25081 -2780 25115 -2764
rect 25081 -4172 25115 -4156
rect 25279 -2780 25313 -2764
rect 25279 -4172 25313 -4156
rect 25477 -2780 25511 -2764
rect 25477 -4172 25511 -4156
rect 25675 -2780 25709 -2764
rect 25675 -4172 25709 -4156
rect 25873 -2780 25907 -2764
rect 25873 -4172 25907 -4156
rect 26071 -2780 26105 -2764
rect 26071 -4172 26105 -4156
rect 26269 -2780 26303 -2764
rect 26269 -4172 26303 -4156
rect 26467 -2780 26501 -2764
rect 26467 -4172 26501 -4156
rect 26665 -2780 26699 -2764
rect 26665 -4172 26699 -4156
rect 26863 -2780 26897 -2764
rect 26863 -4172 26897 -4156
rect 27061 -2780 27095 -2764
rect 27061 -4172 27095 -4156
rect 27259 -2780 27293 -2764
rect 27259 -4172 27293 -4156
rect 27457 -2780 27491 -2764
rect 27457 -4172 27491 -4156
rect 27655 -2780 27689 -2764
rect 27655 -4172 27689 -4156
rect 27853 -2780 27887 -2764
rect 27853 -4172 27887 -4156
rect 28051 -2780 28085 -2764
rect 28051 -4172 28085 -4156
rect 28249 -2780 28283 -2764
rect 28249 -4172 28283 -4156
rect 28447 -2780 28481 -2764
rect 28447 -4172 28481 -4156
rect 28645 -2780 28679 -2764
rect 28645 -4172 28679 -4156
rect 28843 -2780 28877 -2764
rect 28843 -4172 28877 -4156
rect 29041 -2780 29075 -2764
rect 29041 -4172 29075 -4156
rect 29239 -2780 29273 -2764
rect 29239 -4172 29273 -4156
rect 29437 -2780 29471 -2764
rect 29437 -4172 29471 -4156
rect 29635 -2780 29669 -2764
rect 29635 -4172 29669 -4156
rect 29833 -2780 29867 -2764
rect 29833 -4172 29867 -4156
rect 30031 -2780 30065 -2764
rect 30031 -4172 30065 -4156
rect 30229 -2780 30263 -2764
rect 30229 -4172 30263 -4156
rect 30427 -2780 30461 -2764
rect 30427 -4172 30461 -4156
rect 30625 -2780 30659 -2764
rect 30625 -4172 30659 -4156
rect 30823 -2780 30857 -2764
rect 30823 -4172 30857 -4156
rect 31021 -2780 31055 -2764
rect 31021 -4172 31055 -4156
rect 31219 -2780 31253 -2764
rect 31219 -4172 31253 -4156
rect 31417 -2780 31451 -2764
rect 31417 -4172 31451 -4156
rect 31615 -2780 31649 -2764
rect 31615 -4172 31649 -4156
rect 22841 -4415 22875 -4353
rect 32088 -4415 32122 -4353
rect 22841 -4449 22937 -4415
rect 32026 -4449 32122 -4415
<< viali >>
rect 11449 752 11483 2128
rect 11647 752 11681 2128
rect 11845 752 11879 2128
rect 12043 752 12077 2128
rect 12241 752 12275 2128
rect 12439 752 12473 2128
rect 12637 752 12671 2128
rect 12835 752 12869 2128
rect 13033 752 13067 2128
rect 13231 752 13265 2128
rect 13429 752 13463 2128
rect 13627 752 13661 2128
rect 13825 752 13859 2128
rect 14023 752 14057 2128
rect 14221 752 14255 2128
rect 14419 752 14453 2128
rect 14617 752 14651 2128
rect 14815 752 14849 2128
rect 15013 752 15047 2128
rect 15211 752 15245 2128
rect 15409 752 15443 2128
rect 15607 752 15641 2128
rect 15805 752 15839 2128
rect 16003 752 16037 2128
rect 16201 752 16235 2128
rect 16399 752 16433 2128
rect 16597 752 16631 2128
rect 16795 752 16829 2128
rect 16993 752 17027 2128
rect 17191 752 17225 2128
rect 17389 752 17423 2128
rect 17587 752 17621 2128
rect 17785 752 17819 2128
rect 17983 752 18017 2128
rect 18181 752 18215 2128
rect 18379 752 18413 2128
rect 18577 752 18611 2128
rect 18775 752 18809 2128
rect 18973 752 19007 2128
rect 19171 752 19205 2128
rect 19369 752 19403 2128
rect 19567 752 19601 2128
rect 19765 752 19799 2128
rect 11511 659 11619 693
rect 11709 659 11817 693
rect 11907 659 12015 693
rect 12105 659 12213 693
rect 12303 659 12411 693
rect 12501 659 12609 693
rect 12699 659 12807 693
rect 12897 659 13005 693
rect 13095 659 13203 693
rect 13293 659 13401 693
rect 13491 659 13599 693
rect 13689 659 13797 693
rect 13887 659 13995 693
rect 14085 659 14193 693
rect 14283 659 14391 693
rect 14481 659 14589 693
rect 14679 659 14787 693
rect 14877 659 14985 693
rect 15075 659 15183 693
rect 15273 659 15381 693
rect 15471 659 15579 693
rect 15669 659 15777 693
rect 15867 659 15975 693
rect 16065 659 16173 693
rect 16263 659 16371 693
rect 16461 659 16569 693
rect 16659 659 16767 693
rect 16857 659 16965 693
rect 17055 659 17163 693
rect 17253 659 17361 693
rect 17451 659 17559 693
rect 17649 659 17757 693
rect 17847 659 17955 693
rect 18045 659 18153 693
rect 18243 659 18351 693
rect 18441 659 18549 693
rect 18639 659 18747 693
rect 18837 659 18945 693
rect 19035 659 19143 693
rect 19233 659 19341 693
rect 19431 659 19539 693
rect 19629 659 19737 693
rect 11511 551 11619 585
rect 11709 551 11817 585
rect 11907 551 12015 585
rect 12105 551 12213 585
rect 12303 551 12411 585
rect 12501 551 12609 585
rect 12699 551 12807 585
rect 12897 551 13005 585
rect 13095 551 13203 585
rect 13293 551 13401 585
rect 13491 551 13599 585
rect 13689 551 13797 585
rect 13887 551 13995 585
rect 14085 551 14193 585
rect 14283 551 14391 585
rect 14481 551 14589 585
rect 14679 551 14787 585
rect 14877 551 14985 585
rect 15075 551 15183 585
rect 15273 551 15381 585
rect 15471 551 15579 585
rect 15669 551 15777 585
rect 15867 551 15975 585
rect 16065 551 16173 585
rect 16263 551 16371 585
rect 16461 551 16569 585
rect 16659 551 16767 585
rect 16857 551 16965 585
rect 17055 551 17163 585
rect 17253 551 17361 585
rect 17451 551 17559 585
rect 17649 551 17757 585
rect 17847 551 17955 585
rect 18045 551 18153 585
rect 18243 551 18351 585
rect 18441 551 18549 585
rect 18639 551 18747 585
rect 18837 551 18945 585
rect 19035 551 19143 585
rect 19233 551 19341 585
rect 19431 551 19539 585
rect 19629 551 19737 585
rect 11449 -884 11483 492
rect 11647 -884 11681 492
rect 11845 -884 11879 492
rect 12043 -884 12077 492
rect 12241 -884 12275 492
rect 12439 -884 12473 492
rect 12637 -884 12671 492
rect 12835 -884 12869 492
rect 13033 -884 13067 492
rect 13231 -884 13265 492
rect 13429 -884 13463 492
rect 13627 -884 13661 492
rect 13825 -884 13859 492
rect 14023 -884 14057 492
rect 14221 -884 14255 492
rect 14419 -884 14453 492
rect 14617 -884 14651 492
rect 14815 -884 14849 492
rect 15013 -884 15047 492
rect 15211 -884 15245 492
rect 15409 -884 15443 492
rect 15607 -884 15641 492
rect 15805 -884 15839 492
rect 16003 -884 16037 492
rect 16201 -884 16235 492
rect 16399 -884 16433 492
rect 16597 -884 16631 492
rect 16795 -884 16829 492
rect 16993 -884 17027 492
rect 17191 -884 17225 492
rect 17389 -884 17423 492
rect 17587 -884 17621 492
rect 17785 -884 17819 492
rect 17983 -884 18017 492
rect 18181 -884 18215 492
rect 18379 -884 18413 492
rect 18577 -884 18611 492
rect 18775 -884 18809 492
rect 18973 -884 19007 492
rect 19171 -884 19205 492
rect 19369 -884 19403 492
rect 19567 -884 19601 492
rect 19765 -884 19799 492
rect 11511 -977 11619 -943
rect 11709 -977 11817 -943
rect 11907 -977 12015 -943
rect 12105 -977 12213 -943
rect 12303 -977 12411 -943
rect 12501 -977 12609 -943
rect 12699 -977 12807 -943
rect 12897 -977 13005 -943
rect 13095 -977 13203 -943
rect 13293 -977 13401 -943
rect 13491 -977 13599 -943
rect 13689 -977 13797 -943
rect 13887 -977 13995 -943
rect 14085 -977 14193 -943
rect 14283 -977 14391 -943
rect 14481 -977 14589 -943
rect 14679 -977 14787 -943
rect 14877 -977 14985 -943
rect 15075 -977 15183 -943
rect 15273 -977 15381 -943
rect 15471 -977 15579 -943
rect 15669 -977 15777 -943
rect 15867 -977 15975 -943
rect 16065 -977 16173 -943
rect 16263 -977 16371 -943
rect 16461 -977 16569 -943
rect 16659 -977 16767 -943
rect 16857 -977 16965 -943
rect 17055 -977 17163 -943
rect 17253 -977 17361 -943
rect 17451 -977 17559 -943
rect 17649 -977 17757 -943
rect 17847 -977 17955 -943
rect 18045 -977 18153 -943
rect 18243 -977 18351 -943
rect 18441 -977 18549 -943
rect 18639 -977 18747 -943
rect 18837 -977 18945 -943
rect 19035 -977 19143 -943
rect 19233 -977 19341 -943
rect 19431 -977 19539 -943
rect 19629 -977 19737 -943
rect 11511 -1085 11619 -1051
rect 11709 -1085 11817 -1051
rect 11907 -1085 12015 -1051
rect 12105 -1085 12213 -1051
rect 12303 -1085 12411 -1051
rect 12501 -1085 12609 -1051
rect 12699 -1085 12807 -1051
rect 12897 -1085 13005 -1051
rect 13095 -1085 13203 -1051
rect 13293 -1085 13401 -1051
rect 13491 -1085 13599 -1051
rect 13689 -1085 13797 -1051
rect 13887 -1085 13995 -1051
rect 14085 -1085 14193 -1051
rect 14283 -1085 14391 -1051
rect 14481 -1085 14589 -1051
rect 14679 -1085 14787 -1051
rect 14877 -1085 14985 -1051
rect 15075 -1085 15183 -1051
rect 15273 -1085 15381 -1051
rect 15471 -1085 15579 -1051
rect 15669 -1085 15777 -1051
rect 15867 -1085 15975 -1051
rect 16065 -1085 16173 -1051
rect 16263 -1085 16371 -1051
rect 16461 -1085 16569 -1051
rect 16659 -1085 16767 -1051
rect 16857 -1085 16965 -1051
rect 17055 -1085 17163 -1051
rect 17253 -1085 17361 -1051
rect 17451 -1085 17559 -1051
rect 17649 -1085 17757 -1051
rect 17847 -1085 17955 -1051
rect 18045 -1085 18153 -1051
rect 18243 -1085 18351 -1051
rect 18441 -1085 18549 -1051
rect 18639 -1085 18747 -1051
rect 18837 -1085 18945 -1051
rect 19035 -1085 19143 -1051
rect 19233 -1085 19341 -1051
rect 19431 -1085 19539 -1051
rect 19629 -1085 19737 -1051
rect 11449 -2520 11483 -1144
rect 11647 -2520 11681 -1144
rect 11845 -2520 11879 -1144
rect 12043 -2520 12077 -1144
rect 12241 -2520 12275 -1144
rect 12439 -2520 12473 -1144
rect 12637 -2520 12671 -1144
rect 12835 -2520 12869 -1144
rect 13033 -2520 13067 -1144
rect 13231 -2520 13265 -1144
rect 13429 -2520 13463 -1144
rect 13627 -2520 13661 -1144
rect 13825 -2520 13859 -1144
rect 14023 -2520 14057 -1144
rect 14221 -2520 14255 -1144
rect 14419 -2520 14453 -1144
rect 14617 -2520 14651 -1144
rect 14815 -2520 14849 -1144
rect 15013 -2520 15047 -1144
rect 15211 -2520 15245 -1144
rect 15409 -2520 15443 -1144
rect 15607 -2520 15641 -1144
rect 15805 -2520 15839 -1144
rect 16003 -2520 16037 -1144
rect 16201 -2520 16235 -1144
rect 16399 -2520 16433 -1144
rect 16597 -2520 16631 -1144
rect 16795 -2520 16829 -1144
rect 16993 -2520 17027 -1144
rect 17191 -2520 17225 -1144
rect 17389 -2520 17423 -1144
rect 17587 -2520 17621 -1144
rect 17785 -2520 17819 -1144
rect 17983 -2520 18017 -1144
rect 18181 -2520 18215 -1144
rect 18379 -2520 18413 -1144
rect 18577 -2520 18611 -1144
rect 18775 -2520 18809 -1144
rect 18973 -2520 19007 -1144
rect 19171 -2520 19205 -1144
rect 19369 -2520 19403 -1144
rect 19567 -2520 19601 -1144
rect 19765 -2520 19799 -1144
rect 11511 -2613 11619 -2579
rect 11709 -2613 11817 -2579
rect 11907 -2613 12015 -2579
rect 12105 -2613 12213 -2579
rect 12303 -2613 12411 -2579
rect 12501 -2613 12609 -2579
rect 12699 -2613 12807 -2579
rect 12897 -2613 13005 -2579
rect 13095 -2613 13203 -2579
rect 13293 -2613 13401 -2579
rect 13491 -2613 13599 -2579
rect 13689 -2613 13797 -2579
rect 13887 -2613 13995 -2579
rect 14085 -2613 14193 -2579
rect 14283 -2613 14391 -2579
rect 14481 -2613 14589 -2579
rect 14679 -2613 14787 -2579
rect 14877 -2613 14985 -2579
rect 15075 -2613 15183 -2579
rect 15273 -2613 15381 -2579
rect 15471 -2613 15579 -2579
rect 15669 -2613 15777 -2579
rect 15867 -2613 15975 -2579
rect 16065 -2613 16173 -2579
rect 16263 -2613 16371 -2579
rect 16461 -2613 16569 -2579
rect 16659 -2613 16767 -2579
rect 16857 -2613 16965 -2579
rect 17055 -2613 17163 -2579
rect 17253 -2613 17361 -2579
rect 17451 -2613 17559 -2579
rect 17649 -2613 17757 -2579
rect 17847 -2613 17955 -2579
rect 18045 -2613 18153 -2579
rect 18243 -2613 18351 -2579
rect 18441 -2613 18549 -2579
rect 18639 -2613 18747 -2579
rect 18837 -2613 18945 -2579
rect 19035 -2613 19143 -2579
rect 19233 -2613 19341 -2579
rect 19431 -2613 19539 -2579
rect 19629 -2613 19737 -2579
rect 11511 -2721 11619 -2687
rect 11709 -2721 11817 -2687
rect 11907 -2721 12015 -2687
rect 12105 -2721 12213 -2687
rect 12303 -2721 12411 -2687
rect 12501 -2721 12609 -2687
rect 12699 -2721 12807 -2687
rect 12897 -2721 13005 -2687
rect 13095 -2721 13203 -2687
rect 13293 -2721 13401 -2687
rect 13491 -2721 13599 -2687
rect 13689 -2721 13797 -2687
rect 13887 -2721 13995 -2687
rect 14085 -2721 14193 -2687
rect 14283 -2721 14391 -2687
rect 14481 -2721 14589 -2687
rect 14679 -2721 14787 -2687
rect 14877 -2721 14985 -2687
rect 15075 -2721 15183 -2687
rect 15273 -2721 15381 -2687
rect 15471 -2721 15579 -2687
rect 15669 -2721 15777 -2687
rect 15867 -2721 15975 -2687
rect 16065 -2721 16173 -2687
rect 16263 -2721 16371 -2687
rect 16461 -2721 16569 -2687
rect 16659 -2721 16767 -2687
rect 16857 -2721 16965 -2687
rect 17055 -2721 17163 -2687
rect 17253 -2721 17361 -2687
rect 17451 -2721 17559 -2687
rect 17649 -2721 17757 -2687
rect 17847 -2721 17955 -2687
rect 18045 -2721 18153 -2687
rect 18243 -2721 18351 -2687
rect 18441 -2721 18549 -2687
rect 18639 -2721 18747 -2687
rect 18837 -2721 18945 -2687
rect 19035 -2721 19143 -2687
rect 19233 -2721 19341 -2687
rect 19431 -2721 19539 -2687
rect 19629 -2721 19737 -2687
rect 11449 -4156 11483 -2780
rect 11647 -4156 11681 -2780
rect 11845 -4156 11879 -2780
rect 12043 -4156 12077 -2780
rect 12241 -4156 12275 -2780
rect 12439 -4156 12473 -2780
rect 12637 -4156 12671 -2780
rect 12835 -4156 12869 -2780
rect 13033 -4156 13067 -2780
rect 13231 -4156 13265 -2780
rect 13429 -4156 13463 -2780
rect 13627 -4156 13661 -2780
rect 13825 -4156 13859 -2780
rect 14023 -4156 14057 -2780
rect 14221 -4156 14255 -2780
rect 14419 -4156 14453 -2780
rect 14617 -4156 14651 -2780
rect 14815 -4156 14849 -2780
rect 15013 -4156 15047 -2780
rect 15211 -4156 15245 -2780
rect 15409 -4156 15443 -2780
rect 15607 -4156 15641 -2780
rect 15805 -4156 15839 -2780
rect 16003 -4156 16037 -2780
rect 16201 -4156 16235 -2780
rect 16399 -4156 16433 -2780
rect 16597 -4156 16631 -2780
rect 16795 -4156 16829 -2780
rect 16993 -4156 17027 -2780
rect 17191 -4156 17225 -2780
rect 17389 -4156 17423 -2780
rect 17587 -4156 17621 -2780
rect 17785 -4156 17819 -2780
rect 17983 -4156 18017 -2780
rect 18181 -4156 18215 -2780
rect 18379 -4156 18413 -2780
rect 18577 -4156 18611 -2780
rect 18775 -4156 18809 -2780
rect 18973 -4156 19007 -2780
rect 19171 -4156 19205 -2780
rect 19369 -4156 19403 -2780
rect 19567 -4156 19601 -2780
rect 19765 -4156 19799 -2780
rect 23299 752 23333 2128
rect 23497 752 23531 2128
rect 23695 752 23729 2128
rect 23893 752 23927 2128
rect 24091 752 24125 2128
rect 24289 752 24323 2128
rect 24487 752 24521 2128
rect 24685 752 24719 2128
rect 24883 752 24917 2128
rect 25081 752 25115 2128
rect 25279 752 25313 2128
rect 25477 752 25511 2128
rect 25675 752 25709 2128
rect 25873 752 25907 2128
rect 26071 752 26105 2128
rect 26269 752 26303 2128
rect 26467 752 26501 2128
rect 26665 752 26699 2128
rect 26863 752 26897 2128
rect 27061 752 27095 2128
rect 27259 752 27293 2128
rect 27457 752 27491 2128
rect 27655 752 27689 2128
rect 27853 752 27887 2128
rect 28051 752 28085 2128
rect 28249 752 28283 2128
rect 28447 752 28481 2128
rect 28645 752 28679 2128
rect 28843 752 28877 2128
rect 29041 752 29075 2128
rect 29239 752 29273 2128
rect 29437 752 29471 2128
rect 29635 752 29669 2128
rect 29833 752 29867 2128
rect 30031 752 30065 2128
rect 30229 752 30263 2128
rect 30427 752 30461 2128
rect 30625 752 30659 2128
rect 30823 752 30857 2128
rect 31021 752 31055 2128
rect 31219 752 31253 2128
rect 31417 752 31451 2128
rect 31615 752 31649 2128
rect 23361 659 23469 693
rect 23559 659 23667 693
rect 23757 659 23865 693
rect 23955 659 24063 693
rect 24153 659 24261 693
rect 24351 659 24459 693
rect 24549 659 24657 693
rect 24747 659 24855 693
rect 24945 659 25053 693
rect 25143 659 25251 693
rect 25341 659 25449 693
rect 25539 659 25647 693
rect 25737 659 25845 693
rect 25935 659 26043 693
rect 26133 659 26241 693
rect 26331 659 26439 693
rect 26529 659 26637 693
rect 26727 659 26835 693
rect 26925 659 27033 693
rect 27123 659 27231 693
rect 27321 659 27429 693
rect 27519 659 27627 693
rect 27717 659 27825 693
rect 27915 659 28023 693
rect 28113 659 28221 693
rect 28311 659 28419 693
rect 28509 659 28617 693
rect 28707 659 28815 693
rect 28905 659 29013 693
rect 29103 659 29211 693
rect 29301 659 29409 693
rect 29499 659 29607 693
rect 29697 659 29805 693
rect 29895 659 30003 693
rect 30093 659 30201 693
rect 30291 659 30399 693
rect 30489 659 30597 693
rect 30687 659 30795 693
rect 30885 659 30993 693
rect 31083 659 31191 693
rect 31281 659 31389 693
rect 31479 659 31587 693
rect 23361 551 23469 585
rect 23559 551 23667 585
rect 23757 551 23865 585
rect 23955 551 24063 585
rect 24153 551 24261 585
rect 24351 551 24459 585
rect 24549 551 24657 585
rect 24747 551 24855 585
rect 24945 551 25053 585
rect 25143 551 25251 585
rect 25341 551 25449 585
rect 25539 551 25647 585
rect 25737 551 25845 585
rect 25935 551 26043 585
rect 26133 551 26241 585
rect 26331 551 26439 585
rect 26529 551 26637 585
rect 26727 551 26835 585
rect 26925 551 27033 585
rect 27123 551 27231 585
rect 27321 551 27429 585
rect 27519 551 27627 585
rect 27717 551 27825 585
rect 27915 551 28023 585
rect 28113 551 28221 585
rect 28311 551 28419 585
rect 28509 551 28617 585
rect 28707 551 28815 585
rect 28905 551 29013 585
rect 29103 551 29211 585
rect 29301 551 29409 585
rect 29499 551 29607 585
rect 29697 551 29805 585
rect 29895 551 30003 585
rect 30093 551 30201 585
rect 30291 551 30399 585
rect 30489 551 30597 585
rect 30687 551 30795 585
rect 30885 551 30993 585
rect 31083 551 31191 585
rect 31281 551 31389 585
rect 31479 551 31587 585
rect 23299 -884 23333 492
rect 23497 -884 23531 492
rect 23695 -884 23729 492
rect 23893 -884 23927 492
rect 24091 -884 24125 492
rect 24289 -884 24323 492
rect 24487 -884 24521 492
rect 24685 -884 24719 492
rect 24883 -884 24917 492
rect 25081 -884 25115 492
rect 25279 -884 25313 492
rect 25477 -884 25511 492
rect 25675 -884 25709 492
rect 25873 -884 25907 492
rect 26071 -884 26105 492
rect 26269 -884 26303 492
rect 26467 -884 26501 492
rect 26665 -884 26699 492
rect 26863 -884 26897 492
rect 27061 -884 27095 492
rect 27259 -884 27293 492
rect 27457 -884 27491 492
rect 27655 -884 27689 492
rect 27853 -884 27887 492
rect 28051 -884 28085 492
rect 28249 -884 28283 492
rect 28447 -884 28481 492
rect 28645 -884 28679 492
rect 28843 -884 28877 492
rect 29041 -884 29075 492
rect 29239 -884 29273 492
rect 29437 -884 29471 492
rect 29635 -884 29669 492
rect 29833 -884 29867 492
rect 30031 -884 30065 492
rect 30229 -884 30263 492
rect 30427 -884 30461 492
rect 30625 -884 30659 492
rect 30823 -884 30857 492
rect 31021 -884 31055 492
rect 31219 -884 31253 492
rect 31417 -884 31451 492
rect 31615 -884 31649 492
rect 23361 -977 23469 -943
rect 23559 -977 23667 -943
rect 23757 -977 23865 -943
rect 23955 -977 24063 -943
rect 24153 -977 24261 -943
rect 24351 -977 24459 -943
rect 24549 -977 24657 -943
rect 24747 -977 24855 -943
rect 24945 -977 25053 -943
rect 25143 -977 25251 -943
rect 25341 -977 25449 -943
rect 25539 -977 25647 -943
rect 25737 -977 25845 -943
rect 25935 -977 26043 -943
rect 26133 -977 26241 -943
rect 26331 -977 26439 -943
rect 26529 -977 26637 -943
rect 26727 -977 26835 -943
rect 26925 -977 27033 -943
rect 27123 -977 27231 -943
rect 27321 -977 27429 -943
rect 27519 -977 27627 -943
rect 27717 -977 27825 -943
rect 27915 -977 28023 -943
rect 28113 -977 28221 -943
rect 28311 -977 28419 -943
rect 28509 -977 28617 -943
rect 28707 -977 28815 -943
rect 28905 -977 29013 -943
rect 29103 -977 29211 -943
rect 29301 -977 29409 -943
rect 29499 -977 29607 -943
rect 29697 -977 29805 -943
rect 29895 -977 30003 -943
rect 30093 -977 30201 -943
rect 30291 -977 30399 -943
rect 30489 -977 30597 -943
rect 30687 -977 30795 -943
rect 30885 -977 30993 -943
rect 31083 -977 31191 -943
rect 31281 -977 31389 -943
rect 31479 -977 31587 -943
rect 23361 -1085 23469 -1051
rect 23559 -1085 23667 -1051
rect 23757 -1085 23865 -1051
rect 23955 -1085 24063 -1051
rect 24153 -1085 24261 -1051
rect 24351 -1085 24459 -1051
rect 24549 -1085 24657 -1051
rect 24747 -1085 24855 -1051
rect 24945 -1085 25053 -1051
rect 25143 -1085 25251 -1051
rect 25341 -1085 25449 -1051
rect 25539 -1085 25647 -1051
rect 25737 -1085 25845 -1051
rect 25935 -1085 26043 -1051
rect 26133 -1085 26241 -1051
rect 26331 -1085 26439 -1051
rect 26529 -1085 26637 -1051
rect 26727 -1085 26835 -1051
rect 26925 -1085 27033 -1051
rect 27123 -1085 27231 -1051
rect 27321 -1085 27429 -1051
rect 27519 -1085 27627 -1051
rect 27717 -1085 27825 -1051
rect 27915 -1085 28023 -1051
rect 28113 -1085 28221 -1051
rect 28311 -1085 28419 -1051
rect 28509 -1085 28617 -1051
rect 28707 -1085 28815 -1051
rect 28905 -1085 29013 -1051
rect 29103 -1085 29211 -1051
rect 29301 -1085 29409 -1051
rect 29499 -1085 29607 -1051
rect 29697 -1085 29805 -1051
rect 29895 -1085 30003 -1051
rect 30093 -1085 30201 -1051
rect 30291 -1085 30399 -1051
rect 30489 -1085 30597 -1051
rect 30687 -1085 30795 -1051
rect 30885 -1085 30993 -1051
rect 31083 -1085 31191 -1051
rect 31281 -1085 31389 -1051
rect 31479 -1085 31587 -1051
rect 23299 -2520 23333 -1144
rect 23497 -2520 23531 -1144
rect 23695 -2520 23729 -1144
rect 23893 -2520 23927 -1144
rect 24091 -2520 24125 -1144
rect 24289 -2520 24323 -1144
rect 24487 -2520 24521 -1144
rect 24685 -2520 24719 -1144
rect 24883 -2520 24917 -1144
rect 25081 -2520 25115 -1144
rect 25279 -2520 25313 -1144
rect 25477 -2520 25511 -1144
rect 25675 -2520 25709 -1144
rect 25873 -2520 25907 -1144
rect 26071 -2520 26105 -1144
rect 26269 -2520 26303 -1144
rect 26467 -2520 26501 -1144
rect 26665 -2520 26699 -1144
rect 26863 -2520 26897 -1144
rect 27061 -2520 27095 -1144
rect 27259 -2520 27293 -1144
rect 27457 -2520 27491 -1144
rect 27655 -2520 27689 -1144
rect 27853 -2520 27887 -1144
rect 28051 -2520 28085 -1144
rect 28249 -2520 28283 -1144
rect 28447 -2520 28481 -1144
rect 28645 -2520 28679 -1144
rect 28843 -2520 28877 -1144
rect 29041 -2520 29075 -1144
rect 29239 -2520 29273 -1144
rect 29437 -2520 29471 -1144
rect 29635 -2520 29669 -1144
rect 29833 -2520 29867 -1144
rect 30031 -2520 30065 -1144
rect 30229 -2520 30263 -1144
rect 30427 -2520 30461 -1144
rect 30625 -2520 30659 -1144
rect 30823 -2520 30857 -1144
rect 31021 -2520 31055 -1144
rect 31219 -2520 31253 -1144
rect 31417 -2520 31451 -1144
rect 31615 -2520 31649 -1144
rect 23361 -2613 23469 -2579
rect 23559 -2613 23667 -2579
rect 23757 -2613 23865 -2579
rect 23955 -2613 24063 -2579
rect 24153 -2613 24261 -2579
rect 24351 -2613 24459 -2579
rect 24549 -2613 24657 -2579
rect 24747 -2613 24855 -2579
rect 24945 -2613 25053 -2579
rect 25143 -2613 25251 -2579
rect 25341 -2613 25449 -2579
rect 25539 -2613 25647 -2579
rect 25737 -2613 25845 -2579
rect 25935 -2613 26043 -2579
rect 26133 -2613 26241 -2579
rect 26331 -2613 26439 -2579
rect 26529 -2613 26637 -2579
rect 26727 -2613 26835 -2579
rect 26925 -2613 27033 -2579
rect 27123 -2613 27231 -2579
rect 27321 -2613 27429 -2579
rect 27519 -2613 27627 -2579
rect 27717 -2613 27825 -2579
rect 27915 -2613 28023 -2579
rect 28113 -2613 28221 -2579
rect 28311 -2613 28419 -2579
rect 28509 -2613 28617 -2579
rect 28707 -2613 28815 -2579
rect 28905 -2613 29013 -2579
rect 29103 -2613 29211 -2579
rect 29301 -2613 29409 -2579
rect 29499 -2613 29607 -2579
rect 29697 -2613 29805 -2579
rect 29895 -2613 30003 -2579
rect 30093 -2613 30201 -2579
rect 30291 -2613 30399 -2579
rect 30489 -2613 30597 -2579
rect 30687 -2613 30795 -2579
rect 30885 -2613 30993 -2579
rect 31083 -2613 31191 -2579
rect 31281 -2613 31389 -2579
rect 31479 -2613 31587 -2579
rect 23361 -2721 23469 -2687
rect 23559 -2721 23667 -2687
rect 23757 -2721 23865 -2687
rect 23955 -2721 24063 -2687
rect 24153 -2721 24261 -2687
rect 24351 -2721 24459 -2687
rect 24549 -2721 24657 -2687
rect 24747 -2721 24855 -2687
rect 24945 -2721 25053 -2687
rect 25143 -2721 25251 -2687
rect 25341 -2721 25449 -2687
rect 25539 -2721 25647 -2687
rect 25737 -2721 25845 -2687
rect 25935 -2721 26043 -2687
rect 26133 -2721 26241 -2687
rect 26331 -2721 26439 -2687
rect 26529 -2721 26637 -2687
rect 26727 -2721 26835 -2687
rect 26925 -2721 27033 -2687
rect 27123 -2721 27231 -2687
rect 27321 -2721 27429 -2687
rect 27519 -2721 27627 -2687
rect 27717 -2721 27825 -2687
rect 27915 -2721 28023 -2687
rect 28113 -2721 28221 -2687
rect 28311 -2721 28419 -2687
rect 28509 -2721 28617 -2687
rect 28707 -2721 28815 -2687
rect 28905 -2721 29013 -2687
rect 29103 -2721 29211 -2687
rect 29301 -2721 29409 -2687
rect 29499 -2721 29607 -2687
rect 29697 -2721 29805 -2687
rect 29895 -2721 30003 -2687
rect 30093 -2721 30201 -2687
rect 30291 -2721 30399 -2687
rect 30489 -2721 30597 -2687
rect 30687 -2721 30795 -2687
rect 30885 -2721 30993 -2687
rect 31083 -2721 31191 -2687
rect 31281 -2721 31389 -2687
rect 31479 -2721 31587 -2687
rect 23299 -4156 23333 -2780
rect 23497 -4156 23531 -2780
rect 23695 -4156 23729 -2780
rect 23893 -4156 23927 -2780
rect 24091 -4156 24125 -2780
rect 24289 -4156 24323 -2780
rect 24487 -4156 24521 -2780
rect 24685 -4156 24719 -2780
rect 24883 -4156 24917 -2780
rect 25081 -4156 25115 -2780
rect 25279 -4156 25313 -2780
rect 25477 -4156 25511 -2780
rect 25675 -4156 25709 -2780
rect 25873 -4156 25907 -2780
rect 26071 -4156 26105 -2780
rect 26269 -4156 26303 -2780
rect 26467 -4156 26501 -2780
rect 26665 -4156 26699 -2780
rect 26863 -4156 26897 -2780
rect 27061 -4156 27095 -2780
rect 27259 -4156 27293 -2780
rect 27457 -4156 27491 -2780
rect 27655 -4156 27689 -2780
rect 27853 -4156 27887 -2780
rect 28051 -4156 28085 -2780
rect 28249 -4156 28283 -2780
rect 28447 -4156 28481 -2780
rect 28645 -4156 28679 -2780
rect 28843 -4156 28877 -2780
rect 29041 -4156 29075 -2780
rect 29239 -4156 29273 -2780
rect 29437 -4156 29471 -2780
rect 29635 -4156 29669 -2780
rect 29833 -4156 29867 -2780
rect 30031 -4156 30065 -2780
rect 30229 -4156 30263 -2780
rect 30427 -4156 30461 -2780
rect 30625 -4156 30659 -2780
rect 30823 -4156 30857 -2780
rect 31021 -4156 31055 -2780
rect 31219 -4156 31253 -2780
rect 31417 -4156 31451 -2780
rect 31615 -4156 31649 -2780
<< metal1 >>
rect -396 2128 -350 2327
rect 0 2128 46 2327
rect 396 2128 442 2327
rect 792 2128 838 2327
rect 1188 2128 1234 2327
rect 1584 2128 1630 2327
rect 1980 2128 2026 2327
rect 2376 2128 2422 2327
rect 2772 2128 2818 2327
rect 3168 2128 3214 2327
rect 3564 2128 3610 2327
rect 3960 2128 4006 2327
rect 4356 2128 4402 2327
rect 4752 2128 4798 2327
rect 5148 2128 5194 2327
rect 5544 2128 5590 2327
rect 5940 2128 5986 2327
rect 6336 2128 6382 2327
rect 6732 2128 6778 2327
rect 7128 2128 7174 2327
rect 7524 2128 7570 2327
rect 7920 2129 7966 2327
rect -409 752 -399 2128
rect -347 752 -337 2128
rect -211 752 -201 2128
rect -149 752 -139 2128
rect -13 752 -3 2128
rect 49 752 59 2128
rect 185 752 195 2128
rect 247 752 257 2128
rect 383 752 393 2128
rect 445 752 455 2128
rect 581 752 591 2128
rect 643 752 653 2128
rect 779 752 789 2128
rect 841 752 851 2128
rect 977 752 987 2128
rect 1039 752 1049 2128
rect 1175 752 1185 2128
rect 1237 752 1247 2128
rect 1373 752 1383 2128
rect 1435 752 1445 2128
rect 1571 752 1581 2128
rect 1633 752 1643 2128
rect 1769 752 1779 2128
rect 1831 752 1841 2128
rect 1967 752 1977 2128
rect 2029 752 2039 2128
rect 2165 752 2175 2128
rect 2227 752 2237 2128
rect 2363 752 2373 2128
rect 2425 752 2435 2128
rect 2561 752 2571 2128
rect 2623 752 2633 2128
rect 2759 752 2769 2128
rect 2821 752 2831 2128
rect 2957 752 2967 2128
rect 3019 752 3029 2128
rect 3155 752 3165 2128
rect 3217 752 3227 2128
rect 3353 752 3363 2128
rect 3415 752 3425 2128
rect 3551 752 3561 2128
rect 3613 752 3623 2128
rect 3749 752 3759 2128
rect 3811 752 3821 2128
rect 3947 752 3957 2128
rect 4009 752 4019 2128
rect 4145 752 4155 2128
rect 4207 752 4217 2128
rect 4343 752 4353 2128
rect 4405 752 4415 2128
rect 4541 752 4551 2128
rect 4603 752 4613 2128
rect 4739 752 4749 2128
rect 4801 752 4811 2128
rect 4937 752 4947 2128
rect 4999 752 5009 2128
rect 5135 752 5145 2128
rect 5197 752 5207 2128
rect 5333 752 5343 2128
rect 5395 752 5405 2128
rect 5531 752 5541 2128
rect 5593 752 5603 2128
rect 5729 752 5739 2128
rect 5791 752 5801 2128
rect 5927 752 5937 2128
rect 5989 752 5999 2128
rect 6125 752 6135 2128
rect 6187 752 6197 2128
rect 6323 752 6333 2128
rect 6385 752 6395 2128
rect 6521 752 6531 2128
rect 6583 752 6593 2128
rect 6719 752 6729 2128
rect 6781 752 6791 2128
rect 6917 752 6927 2128
rect 6979 752 6989 2128
rect 7115 752 7125 2128
rect 7177 752 7187 2128
rect 7313 752 7323 2128
rect 7375 752 7385 2128
rect 7511 752 7521 2128
rect 7573 752 7583 2128
rect 7709 752 7719 2128
rect 7771 752 7781 2128
rect 7907 753 7917 2129
rect 7969 753 7979 2129
rect -637 545 8207 699
rect -637 -743 -483 545
rect -637 -877 -627 -743
rect -493 -877 -483 -743
rect -637 -937 -483 -877
rect -409 -884 -399 492
rect -347 -884 -337 492
rect -211 -884 -201 492
rect -149 -884 -139 492
rect -13 -884 -3 492
rect 49 -884 59 492
rect 185 -884 195 492
rect 247 -884 257 492
rect 383 -884 393 492
rect 445 -884 455 492
rect 581 -884 591 492
rect 643 -884 653 492
rect 779 -884 789 492
rect 841 -884 851 492
rect 977 -884 987 492
rect 1039 -884 1049 492
rect 1175 -884 1185 492
rect 1237 -884 1247 492
rect 1373 -884 1383 492
rect 1435 -884 1445 492
rect 1571 -884 1581 492
rect 1633 -884 1643 492
rect 1769 -884 1779 492
rect 1831 -884 1841 492
rect 1967 -884 1977 492
rect 2029 -884 2039 492
rect 2165 -884 2175 492
rect 2227 -884 2237 492
rect 2363 -884 2373 492
rect 2425 -884 2435 492
rect 2561 -884 2571 492
rect 2623 -884 2633 492
rect 2759 -884 2769 492
rect 2821 -884 2831 492
rect 2957 -884 2967 492
rect 3019 -884 3029 492
rect 3155 -884 3165 492
rect 3217 -884 3227 492
rect 3353 -884 3363 492
rect 3415 -884 3425 492
rect 3551 -884 3561 492
rect 3613 -884 3623 492
rect 3749 -884 3759 492
rect 3811 -884 3821 492
rect 3947 -884 3957 492
rect 4009 -884 4019 492
rect 4145 -884 4155 492
rect 4207 -884 4217 492
rect 4343 -884 4353 492
rect 4405 -884 4415 492
rect 4541 -884 4551 492
rect 4603 -884 4613 492
rect 4739 -884 4749 492
rect 4801 -884 4811 492
rect 4937 -884 4947 492
rect 4999 -884 5009 492
rect 5135 -884 5145 492
rect 5197 -884 5207 492
rect 5333 -884 5343 492
rect 5395 -884 5405 492
rect 5531 -884 5541 492
rect 5593 -884 5603 492
rect 5729 -884 5739 492
rect 5791 -884 5801 492
rect 5927 -884 5937 492
rect 5989 -884 5999 492
rect 6125 -884 6135 492
rect 6187 -884 6197 492
rect 6323 -884 6333 492
rect 6385 -884 6395 492
rect 6521 -884 6531 492
rect 6583 -884 6593 492
rect 6719 -884 6729 492
rect 6781 -884 6791 492
rect 6917 -884 6927 492
rect 6979 -884 6989 492
rect 7115 -884 7125 492
rect 7177 -884 7187 492
rect 7313 -884 7323 492
rect 7375 -884 7385 492
rect 7511 -884 7521 492
rect 7573 -884 7583 492
rect 7709 -884 7719 492
rect 7771 -884 7781 492
rect 7907 -883 7917 493
rect 7969 -883 7979 493
rect 8053 -743 8207 545
rect 8053 -877 8063 -743
rect 8197 -877 8207 -743
rect 8053 -937 8207 -877
rect -637 -947 8207 -937
rect -637 -1081 -627 -947
rect -493 -1081 8063 -947
rect 8197 -1081 8207 -947
rect -637 -1091 8207 -1081
rect -637 -1151 -483 -1091
rect -637 -1285 -627 -1151
rect -493 -1285 -483 -1151
rect -637 -2573 -483 -1285
rect -409 -2520 -399 -1144
rect -347 -2520 -337 -1144
rect -211 -2520 -201 -1144
rect -149 -2520 -139 -1144
rect -13 -2520 -3 -1144
rect 49 -2520 59 -1144
rect 185 -2520 195 -1144
rect 247 -2520 257 -1144
rect 383 -2520 393 -1144
rect 445 -2520 455 -1144
rect 581 -2520 591 -1144
rect 643 -2520 653 -1144
rect 779 -2520 789 -1144
rect 841 -2520 851 -1144
rect 977 -2520 987 -1144
rect 1039 -2520 1049 -1144
rect 1175 -2520 1185 -1144
rect 1237 -2520 1247 -1144
rect 1373 -2520 1383 -1144
rect 1435 -2520 1445 -1144
rect 1571 -2520 1581 -1144
rect 1633 -2520 1643 -1144
rect 1769 -2520 1779 -1144
rect 1831 -2520 1841 -1144
rect 1967 -2520 1977 -1144
rect 2029 -2520 2039 -1144
rect 2165 -2520 2175 -1144
rect 2227 -2520 2237 -1144
rect 2363 -2520 2373 -1144
rect 2425 -2520 2435 -1144
rect 2561 -2520 2571 -1144
rect 2623 -2520 2633 -1144
rect 2759 -2520 2769 -1144
rect 2821 -2520 2831 -1144
rect 2957 -2520 2967 -1144
rect 3019 -2520 3029 -1144
rect 3155 -2520 3165 -1144
rect 3217 -2520 3227 -1144
rect 3353 -2520 3363 -1144
rect 3415 -2520 3425 -1144
rect 3551 -2520 3561 -1144
rect 3613 -2520 3623 -1144
rect 3749 -2520 3759 -1144
rect 3811 -2520 3821 -1144
rect 3947 -2520 3957 -1144
rect 4009 -2520 4019 -1144
rect 4145 -2520 4155 -1144
rect 4207 -2520 4217 -1144
rect 4343 -2520 4353 -1144
rect 4405 -2520 4415 -1144
rect 4541 -2520 4551 -1144
rect 4603 -2520 4613 -1144
rect 4739 -2520 4749 -1144
rect 4801 -2520 4811 -1144
rect 4937 -2520 4947 -1144
rect 4999 -2520 5009 -1144
rect 5135 -2520 5145 -1144
rect 5197 -2520 5207 -1144
rect 5333 -2520 5343 -1144
rect 5395 -2520 5405 -1144
rect 5531 -2520 5541 -1144
rect 5593 -2520 5603 -1144
rect 5729 -2520 5739 -1144
rect 5791 -2520 5801 -1144
rect 5927 -2520 5937 -1144
rect 5989 -2520 5999 -1144
rect 6125 -2520 6135 -1144
rect 6187 -2520 6197 -1144
rect 6323 -2520 6333 -1144
rect 6385 -2520 6395 -1144
rect 6521 -2520 6531 -1144
rect 6583 -2520 6593 -1144
rect 6719 -2520 6729 -1144
rect 6781 -2520 6791 -1144
rect 6917 -2520 6927 -1144
rect 6979 -2520 6989 -1144
rect 7115 -2520 7125 -1144
rect 7177 -2520 7187 -1144
rect 7313 -2520 7323 -1144
rect 7375 -2520 7385 -1144
rect 7511 -2520 7521 -1144
rect 7573 -2520 7583 -1144
rect 7709 -2520 7719 -1144
rect 7771 -2520 7781 -1144
rect 7907 -2519 7917 -1143
rect 7969 -2519 7979 -1143
rect 8053 -1151 8207 -1091
rect 8053 -1285 8063 -1151
rect 8197 -1285 8207 -1151
rect 8053 -2573 8207 -1285
rect -637 -2727 8207 -2573
rect -409 -4156 -399 -2780
rect -347 -4156 -337 -2780
rect -211 -4156 -201 -2780
rect -149 -4156 -139 -2780
rect -13 -4156 -3 -2780
rect 49 -4156 59 -2780
rect 185 -4156 195 -2780
rect 247 -4156 257 -2780
rect 383 -4156 393 -2780
rect 445 -4156 455 -2780
rect 581 -4156 591 -2780
rect 643 -4156 653 -2780
rect 779 -4156 789 -2780
rect 841 -4156 851 -2780
rect 977 -4156 987 -2780
rect 1039 -4156 1049 -2780
rect 1175 -4156 1185 -2780
rect 1237 -4156 1247 -2780
rect 1373 -4156 1383 -2780
rect 1435 -4156 1445 -2780
rect 1571 -4156 1581 -2780
rect 1633 -4156 1643 -2780
rect 1769 -4156 1779 -2780
rect 1831 -4156 1841 -2780
rect 1967 -4156 1977 -2780
rect 2029 -4156 2039 -2780
rect 2165 -4156 2175 -2780
rect 2227 -4156 2237 -2780
rect 2363 -4156 2373 -2780
rect 2425 -4156 2435 -2780
rect 2561 -4156 2571 -2780
rect 2623 -4156 2633 -2780
rect 2759 -4156 2769 -2780
rect 2821 -4156 2831 -2780
rect 2957 -4156 2967 -2780
rect 3019 -4156 3029 -2780
rect 3155 -4156 3165 -2780
rect 3217 -4156 3227 -2780
rect 3353 -4156 3363 -2780
rect 3415 -4156 3425 -2780
rect 3551 -4156 3561 -2780
rect 3613 -4156 3623 -2780
rect 3749 -4156 3759 -2780
rect 3811 -4156 3821 -2780
rect 3947 -4156 3957 -2780
rect 4009 -4156 4019 -2780
rect 4145 -4156 4155 -2780
rect 4207 -4156 4217 -2780
rect 4343 -4156 4353 -2780
rect 4405 -4156 4415 -2780
rect 4541 -4156 4551 -2780
rect 4603 -4156 4613 -2780
rect 4739 -4156 4749 -2780
rect 4801 -4156 4811 -2780
rect 4937 -4156 4947 -2780
rect 4999 -4156 5009 -2780
rect 5135 -4156 5145 -2780
rect 5197 -4156 5207 -2780
rect 5333 -4156 5343 -2780
rect 5395 -4156 5405 -2780
rect 5531 -4156 5541 -2780
rect 5593 -4156 5603 -2780
rect 5729 -4156 5739 -2780
rect 5791 -4156 5801 -2780
rect 5927 -4156 5937 -2780
rect 5989 -4156 5999 -2780
rect 6125 -4156 6135 -2780
rect 6187 -4156 6197 -2780
rect 6323 -4156 6333 -2780
rect 6385 -4156 6395 -2780
rect 6521 -4156 6531 -2780
rect 6583 -4156 6593 -2780
rect 6719 -4156 6729 -2780
rect 6781 -4156 6791 -2780
rect 6917 -4156 6927 -2780
rect 6979 -4156 6989 -2780
rect 7115 -4156 7125 -2780
rect 7177 -4156 7187 -2780
rect 7313 -4156 7323 -2780
rect 7375 -4156 7385 -2780
rect 7511 -4156 7521 -2780
rect 7573 -4156 7583 -2780
rect 7709 -4156 7719 -2780
rect 7771 -4156 7781 -2780
rect 7907 -4155 7917 -2779
rect 7969 -4155 7979 -2779
rect -396 -4562 -350 -4156
rect 0 -4562 46 -4156
rect 396 -4562 442 -4156
rect 792 -4562 838 -4156
rect 1188 -4562 1234 -4156
rect 1584 -4562 1630 -4156
rect 1980 -4562 2026 -4156
rect 2376 -4562 2422 -4156
rect 2772 -4562 2818 -4156
rect 3168 -4562 3214 -4156
rect 3564 -4562 3610 -4156
rect 3960 -4562 4006 -4156
rect 4356 -4562 4402 -4156
rect 4752 -4562 4798 -4156
rect 5148 -4562 5194 -4156
rect 5544 -4562 5590 -4156
rect 5940 -4562 5986 -4156
rect 6336 -4562 6382 -4156
rect 6732 -4562 6778 -4156
rect 7128 -4562 7174 -4156
rect 7524 -4562 7570 -4156
rect 7920 -4562 7966 -4156
rect 9137 -4562 10357 2327
rect 11443 2128 11489 2327
rect 11641 2128 11687 2140
rect 11839 2128 11885 2327
rect 12037 2128 12083 2140
rect 12235 2128 12281 2327
rect 12433 2128 12479 2140
rect 12631 2128 12677 2327
rect 12829 2128 12875 2140
rect 13027 2128 13073 2327
rect 13225 2128 13271 2140
rect 13423 2128 13469 2327
rect 13621 2128 13667 2140
rect 13819 2128 13865 2327
rect 14017 2128 14063 2140
rect 14215 2128 14261 2327
rect 14413 2128 14459 2140
rect 14611 2128 14657 2327
rect 14809 2128 14855 2140
rect 15007 2128 15053 2327
rect 15205 2128 15251 2140
rect 15403 2128 15449 2327
rect 15601 2128 15647 2140
rect 15799 2128 15845 2327
rect 15997 2128 16043 2140
rect 16195 2128 16241 2327
rect 16393 2128 16439 2140
rect 16591 2128 16637 2327
rect 16789 2128 16835 2140
rect 16987 2128 17033 2327
rect 17185 2128 17231 2140
rect 17383 2128 17429 2327
rect 17581 2128 17627 2140
rect 17779 2128 17825 2327
rect 17977 2128 18023 2140
rect 18175 2128 18221 2327
rect 18373 2128 18419 2140
rect 18571 2128 18617 2327
rect 18769 2128 18815 2140
rect 18967 2128 19013 2327
rect 19165 2128 19211 2140
rect 19363 2128 19409 2327
rect 19561 2128 19607 2140
rect 19759 2129 19805 2327
rect 11430 752 11440 2128
rect 11492 752 11502 2128
rect 11628 752 11638 2128
rect 11690 752 11700 2128
rect 11826 752 11836 2128
rect 11888 752 11898 2128
rect 12024 752 12034 2128
rect 12086 752 12096 2128
rect 12222 752 12232 2128
rect 12284 752 12294 2128
rect 12420 752 12430 2128
rect 12482 752 12492 2128
rect 12618 752 12628 2128
rect 12680 752 12690 2128
rect 12816 752 12826 2128
rect 12878 752 12888 2128
rect 13014 752 13024 2128
rect 13076 752 13086 2128
rect 13212 752 13222 2128
rect 13274 752 13284 2128
rect 13410 752 13420 2128
rect 13472 752 13482 2128
rect 13608 752 13618 2128
rect 13670 752 13680 2128
rect 13806 752 13816 2128
rect 13868 752 13878 2128
rect 14004 752 14014 2128
rect 14066 752 14076 2128
rect 14202 752 14212 2128
rect 14264 752 14274 2128
rect 14400 752 14410 2128
rect 14462 752 14472 2128
rect 14598 752 14608 2128
rect 14660 752 14670 2128
rect 14796 752 14806 2128
rect 14858 752 14868 2128
rect 14994 752 15004 2128
rect 15056 752 15066 2128
rect 15192 752 15202 2128
rect 15254 752 15264 2128
rect 15390 752 15400 2128
rect 15452 752 15462 2128
rect 15588 752 15598 2128
rect 15650 752 15660 2128
rect 15786 752 15796 2128
rect 15848 752 15858 2128
rect 15984 752 15994 2128
rect 16046 752 16056 2128
rect 16182 752 16192 2128
rect 16244 752 16254 2128
rect 16380 752 16390 2128
rect 16442 752 16452 2128
rect 16578 752 16588 2128
rect 16640 752 16650 2128
rect 16776 752 16786 2128
rect 16838 752 16848 2128
rect 16974 752 16984 2128
rect 17036 752 17046 2128
rect 17172 752 17182 2128
rect 17234 752 17244 2128
rect 17370 752 17380 2128
rect 17432 752 17442 2128
rect 17568 752 17578 2128
rect 17630 752 17640 2128
rect 17766 752 17776 2128
rect 17828 752 17838 2128
rect 17964 752 17974 2128
rect 18026 752 18036 2128
rect 18162 752 18172 2128
rect 18224 752 18234 2128
rect 18360 752 18370 2128
rect 18422 752 18432 2128
rect 18558 752 18568 2128
rect 18620 752 18630 2128
rect 18756 752 18766 2128
rect 18818 752 18828 2128
rect 18954 752 18964 2128
rect 19016 752 19026 2128
rect 19152 752 19162 2128
rect 19214 752 19224 2128
rect 19350 752 19360 2128
rect 19412 752 19422 2128
rect 19548 752 19558 2128
rect 19610 752 19620 2128
rect 19746 753 19756 2129
rect 19808 753 19818 2129
rect 19759 752 19765 753
rect 19799 752 19805 753
rect 11443 740 11489 752
rect 11641 740 11687 752
rect 11839 740 11885 752
rect 12037 740 12083 752
rect 12235 740 12281 752
rect 12433 740 12479 752
rect 12631 740 12677 752
rect 12829 740 12875 752
rect 13027 740 13073 752
rect 13225 740 13271 752
rect 13423 740 13469 752
rect 13621 740 13667 752
rect 13819 740 13865 752
rect 14017 740 14063 752
rect 14215 740 14261 752
rect 14413 740 14459 752
rect 14611 740 14657 752
rect 14809 740 14855 752
rect 15007 740 15053 752
rect 15205 740 15251 752
rect 15403 740 15449 752
rect 15601 740 15647 752
rect 15799 740 15845 752
rect 15997 740 16043 752
rect 16195 740 16241 752
rect 16393 740 16439 752
rect 16591 740 16637 752
rect 16789 740 16835 752
rect 16987 740 17033 752
rect 17185 740 17231 752
rect 17383 740 17429 752
rect 17581 740 17627 752
rect 17779 740 17825 752
rect 17977 740 18023 752
rect 18175 740 18221 752
rect 18373 740 18419 752
rect 18571 740 18617 752
rect 18769 740 18815 752
rect 18967 740 19013 752
rect 19165 740 19211 752
rect 19363 740 19409 752
rect 19561 740 19607 752
rect 19759 740 19805 752
rect 11202 693 20046 699
rect 11202 659 11511 693
rect 11619 659 11709 693
rect 11817 659 11907 693
rect 12015 659 12105 693
rect 12213 659 12303 693
rect 12411 659 12501 693
rect 12609 659 12699 693
rect 12807 659 12897 693
rect 13005 659 13095 693
rect 13203 659 13293 693
rect 13401 659 13491 693
rect 13599 659 13689 693
rect 13797 659 13887 693
rect 13995 659 14085 693
rect 14193 659 14283 693
rect 14391 659 14481 693
rect 14589 659 14679 693
rect 14787 659 14877 693
rect 14985 659 15075 693
rect 15183 659 15273 693
rect 15381 659 15471 693
rect 15579 659 15669 693
rect 15777 659 15867 693
rect 15975 659 16065 693
rect 16173 659 16263 693
rect 16371 659 16461 693
rect 16569 659 16659 693
rect 16767 659 16857 693
rect 16965 659 17055 693
rect 17163 659 17253 693
rect 17361 659 17451 693
rect 17559 659 17649 693
rect 17757 659 17847 693
rect 17955 659 18045 693
rect 18153 659 18243 693
rect 18351 659 18441 693
rect 18549 659 18639 693
rect 18747 659 18837 693
rect 18945 659 19035 693
rect 19143 659 19233 693
rect 19341 659 19431 693
rect 19539 659 19629 693
rect 19737 659 20046 693
rect 11202 585 20046 659
rect 11202 551 11511 585
rect 11619 551 11709 585
rect 11817 551 11907 585
rect 12015 551 12105 585
rect 12213 551 12303 585
rect 12411 551 12501 585
rect 12609 551 12699 585
rect 12807 551 12897 585
rect 13005 551 13095 585
rect 13203 551 13293 585
rect 13401 551 13491 585
rect 13599 551 13689 585
rect 13797 551 13887 585
rect 13995 551 14085 585
rect 14193 551 14283 585
rect 14391 551 14481 585
rect 14589 551 14679 585
rect 14787 551 14877 585
rect 14985 551 15075 585
rect 15183 551 15273 585
rect 15381 551 15471 585
rect 15579 551 15669 585
rect 15777 551 15867 585
rect 15975 551 16065 585
rect 16173 551 16263 585
rect 16371 551 16461 585
rect 16569 551 16659 585
rect 16767 551 16857 585
rect 16965 551 17055 585
rect 17163 551 17253 585
rect 17361 551 17451 585
rect 17559 551 17649 585
rect 17757 551 17847 585
rect 17955 551 18045 585
rect 18153 551 18243 585
rect 18351 551 18441 585
rect 18549 551 18639 585
rect 18747 551 18837 585
rect 18945 551 19035 585
rect 19143 551 19233 585
rect 19341 551 19431 585
rect 19539 551 19629 585
rect 19737 551 20046 585
rect 11202 545 20046 551
rect 11202 -743 11356 545
rect 11443 492 11489 504
rect 11641 492 11687 504
rect 11839 492 11885 504
rect 12037 492 12083 504
rect 12235 492 12281 504
rect 12433 492 12479 504
rect 12631 492 12677 504
rect 12829 492 12875 504
rect 13027 492 13073 504
rect 13225 492 13271 504
rect 13423 492 13469 504
rect 13621 492 13667 504
rect 13819 492 13865 504
rect 14017 492 14063 504
rect 14215 492 14261 504
rect 14413 492 14459 504
rect 14611 492 14657 504
rect 14809 492 14855 504
rect 15007 492 15053 504
rect 15205 492 15251 504
rect 15403 492 15449 504
rect 15601 492 15647 504
rect 15799 492 15845 504
rect 15997 492 16043 504
rect 16195 492 16241 504
rect 16393 492 16439 504
rect 16591 492 16637 504
rect 16789 492 16835 504
rect 16987 492 17033 504
rect 17185 492 17231 504
rect 17383 492 17429 504
rect 17581 492 17627 504
rect 17779 492 17825 504
rect 17977 492 18023 504
rect 18175 492 18221 504
rect 18373 492 18419 504
rect 18571 492 18617 504
rect 18769 492 18815 504
rect 18967 492 19013 504
rect 19165 492 19211 504
rect 19363 492 19409 504
rect 19561 492 19607 504
rect 19759 493 19805 504
rect 11202 -877 11212 -743
rect 11346 -877 11356 -743
rect 11202 -937 11356 -877
rect 11430 -884 11440 492
rect 11492 -884 11502 492
rect 11628 -884 11638 492
rect 11690 -884 11700 492
rect 11826 -884 11836 492
rect 11888 -884 11898 492
rect 12024 -884 12034 492
rect 12086 -884 12096 492
rect 12222 -884 12232 492
rect 12284 -884 12294 492
rect 12420 -884 12430 492
rect 12482 -884 12492 492
rect 12618 -884 12628 492
rect 12680 -884 12690 492
rect 12816 -884 12826 492
rect 12878 -884 12888 492
rect 13014 -884 13024 492
rect 13076 -884 13086 492
rect 13212 -884 13222 492
rect 13274 -884 13284 492
rect 13410 -884 13420 492
rect 13472 -884 13482 492
rect 13608 -884 13618 492
rect 13670 -884 13680 492
rect 13806 -884 13816 492
rect 13868 -884 13878 492
rect 14004 -884 14014 492
rect 14066 -884 14076 492
rect 14202 -884 14212 492
rect 14264 -884 14274 492
rect 14400 -884 14410 492
rect 14462 -884 14472 492
rect 14598 -884 14608 492
rect 14660 -884 14670 492
rect 14796 -884 14806 492
rect 14858 -884 14868 492
rect 14994 -884 15004 492
rect 15056 -884 15066 492
rect 15192 -884 15202 492
rect 15254 -884 15264 492
rect 15390 -884 15400 492
rect 15452 -884 15462 492
rect 15588 -884 15598 492
rect 15650 -884 15660 492
rect 15786 -884 15796 492
rect 15848 -884 15858 492
rect 15984 -884 15994 492
rect 16046 -884 16056 492
rect 16182 -884 16192 492
rect 16244 -884 16254 492
rect 16380 -884 16390 492
rect 16442 -884 16452 492
rect 16578 -884 16588 492
rect 16640 -884 16650 492
rect 16776 -884 16786 492
rect 16838 -884 16848 492
rect 16974 -884 16984 492
rect 17036 -884 17046 492
rect 17172 -884 17182 492
rect 17234 -884 17244 492
rect 17370 -884 17380 492
rect 17432 -884 17442 492
rect 17568 -884 17578 492
rect 17630 -884 17640 492
rect 17766 -884 17776 492
rect 17828 -884 17838 492
rect 17964 -884 17974 492
rect 18026 -884 18036 492
rect 18162 -884 18172 492
rect 18224 -884 18234 492
rect 18360 -884 18370 492
rect 18422 -884 18432 492
rect 18558 -884 18568 492
rect 18620 -884 18630 492
rect 18756 -884 18766 492
rect 18818 -884 18828 492
rect 18954 -884 18964 492
rect 19016 -884 19026 492
rect 19152 -884 19162 492
rect 19214 -884 19224 492
rect 19350 -884 19360 492
rect 19412 -884 19422 492
rect 19548 -884 19558 492
rect 19610 -884 19620 492
rect 19746 -883 19756 493
rect 19808 -883 19818 493
rect 19892 -743 20046 545
rect 19892 -877 19902 -743
rect 20036 -877 20046 -743
rect 19759 -884 19765 -883
rect 19799 -884 19805 -883
rect 11443 -896 11489 -884
rect 11641 -896 11687 -884
rect 11839 -896 11885 -884
rect 12037 -896 12083 -884
rect 12235 -896 12281 -884
rect 12433 -896 12479 -884
rect 12631 -896 12677 -884
rect 12829 -896 12875 -884
rect 13027 -896 13073 -884
rect 13225 -896 13271 -884
rect 13423 -896 13469 -884
rect 13621 -896 13667 -884
rect 13819 -896 13865 -884
rect 14017 -896 14063 -884
rect 14215 -896 14261 -884
rect 14413 -896 14459 -884
rect 14611 -896 14657 -884
rect 14809 -896 14855 -884
rect 15007 -896 15053 -884
rect 15205 -896 15251 -884
rect 15403 -896 15449 -884
rect 15601 -896 15647 -884
rect 15799 -896 15845 -884
rect 15997 -896 16043 -884
rect 16195 -896 16241 -884
rect 16393 -896 16439 -884
rect 16591 -896 16637 -884
rect 16789 -896 16835 -884
rect 16987 -896 17033 -884
rect 17185 -896 17231 -884
rect 17383 -896 17429 -884
rect 17581 -896 17627 -884
rect 17779 -896 17825 -884
rect 17977 -896 18023 -884
rect 18175 -896 18221 -884
rect 18373 -896 18419 -884
rect 18571 -896 18617 -884
rect 18769 -896 18815 -884
rect 18967 -896 19013 -884
rect 19165 -896 19211 -884
rect 19363 -896 19409 -884
rect 19561 -896 19607 -884
rect 19759 -896 19805 -884
rect 19892 -937 20046 -877
rect 11202 -943 20046 -937
rect 11202 -947 11511 -943
rect 11202 -1081 11212 -947
rect 11346 -977 11511 -947
rect 11619 -977 11709 -943
rect 11817 -977 11907 -943
rect 12015 -977 12105 -943
rect 12213 -977 12303 -943
rect 12411 -977 12501 -943
rect 12609 -977 12699 -943
rect 12807 -977 12897 -943
rect 13005 -977 13095 -943
rect 13203 -977 13293 -943
rect 13401 -977 13491 -943
rect 13599 -977 13689 -943
rect 13797 -977 13887 -943
rect 13995 -977 14085 -943
rect 14193 -977 14283 -943
rect 14391 -977 14481 -943
rect 14589 -977 14679 -943
rect 14787 -977 14877 -943
rect 14985 -977 15075 -943
rect 15183 -977 15273 -943
rect 15381 -977 15471 -943
rect 15579 -977 15669 -943
rect 15777 -977 15867 -943
rect 15975 -977 16065 -943
rect 16173 -977 16263 -943
rect 16371 -977 16461 -943
rect 16569 -977 16659 -943
rect 16767 -977 16857 -943
rect 16965 -977 17055 -943
rect 17163 -977 17253 -943
rect 17361 -977 17451 -943
rect 17559 -977 17649 -943
rect 17757 -977 17847 -943
rect 17955 -977 18045 -943
rect 18153 -977 18243 -943
rect 18351 -977 18441 -943
rect 18549 -977 18639 -943
rect 18747 -977 18837 -943
rect 18945 -977 19035 -943
rect 19143 -977 19233 -943
rect 19341 -977 19431 -943
rect 19539 -977 19629 -943
rect 19737 -947 20046 -943
rect 19737 -977 19902 -947
rect 11346 -1051 19902 -977
rect 11346 -1081 11511 -1051
rect 11202 -1085 11511 -1081
rect 11619 -1085 11709 -1051
rect 11817 -1085 11907 -1051
rect 12015 -1085 12105 -1051
rect 12213 -1085 12303 -1051
rect 12411 -1085 12501 -1051
rect 12609 -1085 12699 -1051
rect 12807 -1085 12897 -1051
rect 13005 -1085 13095 -1051
rect 13203 -1085 13293 -1051
rect 13401 -1085 13491 -1051
rect 13599 -1085 13689 -1051
rect 13797 -1085 13887 -1051
rect 13995 -1085 14085 -1051
rect 14193 -1085 14283 -1051
rect 14391 -1085 14481 -1051
rect 14589 -1085 14679 -1051
rect 14787 -1085 14877 -1051
rect 14985 -1085 15075 -1051
rect 15183 -1085 15273 -1051
rect 15381 -1085 15471 -1051
rect 15579 -1085 15669 -1051
rect 15777 -1085 15867 -1051
rect 15975 -1085 16065 -1051
rect 16173 -1085 16263 -1051
rect 16371 -1085 16461 -1051
rect 16569 -1085 16659 -1051
rect 16767 -1085 16857 -1051
rect 16965 -1085 17055 -1051
rect 17163 -1085 17253 -1051
rect 17361 -1085 17451 -1051
rect 17559 -1085 17649 -1051
rect 17757 -1085 17847 -1051
rect 17955 -1085 18045 -1051
rect 18153 -1085 18243 -1051
rect 18351 -1085 18441 -1051
rect 18549 -1085 18639 -1051
rect 18747 -1085 18837 -1051
rect 18945 -1085 19035 -1051
rect 19143 -1085 19233 -1051
rect 19341 -1085 19431 -1051
rect 19539 -1085 19629 -1051
rect 19737 -1081 19902 -1051
rect 20036 -1081 20046 -947
rect 19737 -1085 20046 -1081
rect 11202 -1091 20046 -1085
rect 11202 -1151 11356 -1091
rect 11443 -1144 11489 -1132
rect 11641 -1144 11687 -1132
rect 11839 -1144 11885 -1132
rect 12037 -1144 12083 -1132
rect 12235 -1144 12281 -1132
rect 12433 -1144 12479 -1132
rect 12631 -1144 12677 -1132
rect 12829 -1144 12875 -1132
rect 13027 -1144 13073 -1132
rect 13225 -1144 13271 -1132
rect 13423 -1144 13469 -1132
rect 13621 -1144 13667 -1132
rect 13819 -1144 13865 -1132
rect 14017 -1144 14063 -1132
rect 14215 -1144 14261 -1132
rect 14413 -1144 14459 -1132
rect 14611 -1144 14657 -1132
rect 14809 -1144 14855 -1132
rect 15007 -1144 15053 -1132
rect 15205 -1144 15251 -1132
rect 15403 -1144 15449 -1132
rect 15601 -1144 15647 -1132
rect 15799 -1144 15845 -1132
rect 15997 -1144 16043 -1132
rect 16195 -1144 16241 -1132
rect 16393 -1144 16439 -1132
rect 16591 -1144 16637 -1132
rect 16789 -1144 16835 -1132
rect 16987 -1144 17033 -1132
rect 17185 -1144 17231 -1132
rect 17383 -1144 17429 -1132
rect 17581 -1144 17627 -1132
rect 17779 -1144 17825 -1132
rect 17977 -1144 18023 -1132
rect 18175 -1144 18221 -1132
rect 18373 -1144 18419 -1132
rect 18571 -1144 18617 -1132
rect 18769 -1144 18815 -1132
rect 18967 -1144 19013 -1132
rect 19165 -1144 19211 -1132
rect 19363 -1144 19409 -1132
rect 19561 -1144 19607 -1132
rect 19759 -1143 19805 -1132
rect 11202 -1285 11212 -1151
rect 11346 -1285 11356 -1151
rect 11202 -2573 11356 -1285
rect 11430 -2520 11440 -1144
rect 11492 -2520 11502 -1144
rect 11628 -2520 11638 -1144
rect 11690 -2520 11700 -1144
rect 11826 -2520 11836 -1144
rect 11888 -2520 11898 -1144
rect 12024 -2520 12034 -1144
rect 12086 -2520 12096 -1144
rect 12222 -2520 12232 -1144
rect 12284 -2520 12294 -1144
rect 12420 -2520 12430 -1144
rect 12482 -2520 12492 -1144
rect 12618 -2520 12628 -1144
rect 12680 -2520 12690 -1144
rect 12816 -2520 12826 -1144
rect 12878 -2520 12888 -1144
rect 13014 -2520 13024 -1144
rect 13076 -2520 13086 -1144
rect 13212 -2520 13222 -1144
rect 13274 -2520 13284 -1144
rect 13410 -2520 13420 -1144
rect 13472 -2520 13482 -1144
rect 13608 -2520 13618 -1144
rect 13670 -2520 13680 -1144
rect 13806 -2520 13816 -1144
rect 13868 -2520 13878 -1144
rect 14004 -2520 14014 -1144
rect 14066 -2520 14076 -1144
rect 14202 -2520 14212 -1144
rect 14264 -2520 14274 -1144
rect 14400 -2520 14410 -1144
rect 14462 -2520 14472 -1144
rect 14598 -2520 14608 -1144
rect 14660 -2520 14670 -1144
rect 14796 -2520 14806 -1144
rect 14858 -2520 14868 -1144
rect 14994 -2520 15004 -1144
rect 15056 -2520 15066 -1144
rect 15192 -2520 15202 -1144
rect 15254 -2520 15264 -1144
rect 15390 -2520 15400 -1144
rect 15452 -2520 15462 -1144
rect 15588 -2520 15598 -1144
rect 15650 -2520 15660 -1144
rect 15786 -2520 15796 -1144
rect 15848 -2520 15858 -1144
rect 15984 -2520 15994 -1144
rect 16046 -2520 16056 -1144
rect 16182 -2520 16192 -1144
rect 16244 -2520 16254 -1144
rect 16380 -2520 16390 -1144
rect 16442 -2520 16452 -1144
rect 16578 -2520 16588 -1144
rect 16640 -2520 16650 -1144
rect 16776 -2520 16786 -1144
rect 16838 -2520 16848 -1144
rect 16974 -2520 16984 -1144
rect 17036 -2520 17046 -1144
rect 17172 -2520 17182 -1144
rect 17234 -2520 17244 -1144
rect 17370 -2520 17380 -1144
rect 17432 -2520 17442 -1144
rect 17568 -2520 17578 -1144
rect 17630 -2520 17640 -1144
rect 17766 -2520 17776 -1144
rect 17828 -2520 17838 -1144
rect 17964 -2520 17974 -1144
rect 18026 -2520 18036 -1144
rect 18162 -2520 18172 -1144
rect 18224 -2520 18234 -1144
rect 18360 -2520 18370 -1144
rect 18422 -2520 18432 -1144
rect 18558 -2520 18568 -1144
rect 18620 -2520 18630 -1144
rect 18756 -2520 18766 -1144
rect 18818 -2520 18828 -1144
rect 18954 -2520 18964 -1144
rect 19016 -2520 19026 -1144
rect 19152 -2520 19162 -1144
rect 19214 -2520 19224 -1144
rect 19350 -2520 19360 -1144
rect 19412 -2520 19422 -1144
rect 19548 -2520 19558 -1144
rect 19610 -2520 19620 -1144
rect 19746 -2519 19756 -1143
rect 19808 -2519 19818 -1143
rect 19892 -1151 20046 -1091
rect 19892 -1285 19902 -1151
rect 20036 -1285 20046 -1151
rect 19759 -2520 19765 -2519
rect 19799 -2520 19805 -2519
rect 11443 -2532 11489 -2520
rect 11641 -2532 11687 -2520
rect 11839 -2532 11885 -2520
rect 12037 -2532 12083 -2520
rect 12235 -2532 12281 -2520
rect 12433 -2532 12479 -2520
rect 12631 -2532 12677 -2520
rect 12829 -2532 12875 -2520
rect 13027 -2532 13073 -2520
rect 13225 -2532 13271 -2520
rect 13423 -2532 13469 -2520
rect 13621 -2532 13667 -2520
rect 13819 -2532 13865 -2520
rect 14017 -2532 14063 -2520
rect 14215 -2532 14261 -2520
rect 14413 -2532 14459 -2520
rect 14611 -2532 14657 -2520
rect 14809 -2532 14855 -2520
rect 15007 -2532 15053 -2520
rect 15205 -2532 15251 -2520
rect 15403 -2532 15449 -2520
rect 15601 -2532 15647 -2520
rect 15799 -2532 15845 -2520
rect 15997 -2532 16043 -2520
rect 16195 -2532 16241 -2520
rect 16393 -2532 16439 -2520
rect 16591 -2532 16637 -2520
rect 16789 -2532 16835 -2520
rect 16987 -2532 17033 -2520
rect 17185 -2532 17231 -2520
rect 17383 -2532 17429 -2520
rect 17581 -2532 17627 -2520
rect 17779 -2532 17825 -2520
rect 17977 -2532 18023 -2520
rect 18175 -2532 18221 -2520
rect 18373 -2532 18419 -2520
rect 18571 -2532 18617 -2520
rect 18769 -2532 18815 -2520
rect 18967 -2532 19013 -2520
rect 19165 -2532 19211 -2520
rect 19363 -2532 19409 -2520
rect 19561 -2532 19607 -2520
rect 19759 -2532 19805 -2520
rect 19892 -2573 20046 -1285
rect 11202 -2579 20046 -2573
rect 11202 -2613 11511 -2579
rect 11619 -2613 11709 -2579
rect 11817 -2613 11907 -2579
rect 12015 -2613 12105 -2579
rect 12213 -2613 12303 -2579
rect 12411 -2613 12501 -2579
rect 12609 -2613 12699 -2579
rect 12807 -2613 12897 -2579
rect 13005 -2613 13095 -2579
rect 13203 -2613 13293 -2579
rect 13401 -2613 13491 -2579
rect 13599 -2613 13689 -2579
rect 13797 -2613 13887 -2579
rect 13995 -2613 14085 -2579
rect 14193 -2613 14283 -2579
rect 14391 -2613 14481 -2579
rect 14589 -2613 14679 -2579
rect 14787 -2613 14877 -2579
rect 14985 -2613 15075 -2579
rect 15183 -2613 15273 -2579
rect 15381 -2613 15471 -2579
rect 15579 -2613 15669 -2579
rect 15777 -2613 15867 -2579
rect 15975 -2613 16065 -2579
rect 16173 -2613 16263 -2579
rect 16371 -2613 16461 -2579
rect 16569 -2613 16659 -2579
rect 16767 -2613 16857 -2579
rect 16965 -2613 17055 -2579
rect 17163 -2613 17253 -2579
rect 17361 -2613 17451 -2579
rect 17559 -2613 17649 -2579
rect 17757 -2613 17847 -2579
rect 17955 -2613 18045 -2579
rect 18153 -2613 18243 -2579
rect 18351 -2613 18441 -2579
rect 18549 -2613 18639 -2579
rect 18747 -2613 18837 -2579
rect 18945 -2613 19035 -2579
rect 19143 -2613 19233 -2579
rect 19341 -2613 19431 -2579
rect 19539 -2613 19629 -2579
rect 19737 -2613 20046 -2579
rect 11202 -2687 20046 -2613
rect 11202 -2721 11511 -2687
rect 11619 -2721 11709 -2687
rect 11817 -2721 11907 -2687
rect 12015 -2721 12105 -2687
rect 12213 -2721 12303 -2687
rect 12411 -2721 12501 -2687
rect 12609 -2721 12699 -2687
rect 12807 -2721 12897 -2687
rect 13005 -2721 13095 -2687
rect 13203 -2721 13293 -2687
rect 13401 -2721 13491 -2687
rect 13599 -2721 13689 -2687
rect 13797 -2721 13887 -2687
rect 13995 -2721 14085 -2687
rect 14193 -2721 14283 -2687
rect 14391 -2721 14481 -2687
rect 14589 -2721 14679 -2687
rect 14787 -2721 14877 -2687
rect 14985 -2721 15075 -2687
rect 15183 -2721 15273 -2687
rect 15381 -2721 15471 -2687
rect 15579 -2721 15669 -2687
rect 15777 -2721 15867 -2687
rect 15975 -2721 16065 -2687
rect 16173 -2721 16263 -2687
rect 16371 -2721 16461 -2687
rect 16569 -2721 16659 -2687
rect 16767 -2721 16857 -2687
rect 16965 -2721 17055 -2687
rect 17163 -2721 17253 -2687
rect 17361 -2721 17451 -2687
rect 17559 -2721 17649 -2687
rect 17757 -2721 17847 -2687
rect 17955 -2721 18045 -2687
rect 18153 -2721 18243 -2687
rect 18351 -2721 18441 -2687
rect 18549 -2721 18639 -2687
rect 18747 -2721 18837 -2687
rect 18945 -2721 19035 -2687
rect 19143 -2721 19233 -2687
rect 19341 -2721 19431 -2687
rect 19539 -2721 19629 -2687
rect 19737 -2721 20046 -2687
rect 11202 -2727 20046 -2721
rect 11443 -2780 11489 -2768
rect 11641 -2780 11687 -2768
rect 11839 -2780 11885 -2768
rect 12037 -2780 12083 -2768
rect 12235 -2780 12281 -2768
rect 12433 -2780 12479 -2768
rect 12631 -2780 12677 -2768
rect 12829 -2780 12875 -2768
rect 13027 -2780 13073 -2768
rect 13225 -2780 13271 -2768
rect 13423 -2780 13469 -2768
rect 13621 -2780 13667 -2768
rect 13819 -2780 13865 -2768
rect 14017 -2780 14063 -2768
rect 14215 -2780 14261 -2768
rect 14413 -2780 14459 -2768
rect 14611 -2780 14657 -2768
rect 14809 -2780 14855 -2768
rect 15007 -2780 15053 -2768
rect 15205 -2780 15251 -2768
rect 15403 -2780 15449 -2768
rect 15601 -2780 15647 -2768
rect 15799 -2780 15845 -2768
rect 15997 -2780 16043 -2768
rect 16195 -2780 16241 -2768
rect 16393 -2780 16439 -2768
rect 16591 -2780 16637 -2768
rect 16789 -2780 16835 -2768
rect 16987 -2780 17033 -2768
rect 17185 -2780 17231 -2768
rect 17383 -2780 17429 -2768
rect 17581 -2780 17627 -2768
rect 17779 -2780 17825 -2768
rect 17977 -2780 18023 -2768
rect 18175 -2780 18221 -2768
rect 18373 -2780 18419 -2768
rect 18571 -2780 18617 -2768
rect 18769 -2780 18815 -2768
rect 18967 -2780 19013 -2768
rect 19165 -2780 19211 -2768
rect 19363 -2780 19409 -2768
rect 19561 -2780 19607 -2768
rect 19759 -2779 19805 -2768
rect 11430 -4156 11440 -2780
rect 11492 -4156 11502 -2780
rect 11628 -4156 11638 -2780
rect 11690 -4156 11700 -2780
rect 11826 -4156 11836 -2780
rect 11888 -4156 11898 -2780
rect 12024 -4156 12034 -2780
rect 12086 -4156 12096 -2780
rect 12222 -4156 12232 -2780
rect 12284 -4156 12294 -2780
rect 12420 -4156 12430 -2780
rect 12482 -4156 12492 -2780
rect 12618 -4156 12628 -2780
rect 12680 -4156 12690 -2780
rect 12816 -4156 12826 -2780
rect 12878 -4156 12888 -2780
rect 13014 -4156 13024 -2780
rect 13076 -4156 13086 -2780
rect 13212 -4156 13222 -2780
rect 13274 -4156 13284 -2780
rect 13410 -4156 13420 -2780
rect 13472 -4156 13482 -2780
rect 13608 -4156 13618 -2780
rect 13670 -4156 13680 -2780
rect 13806 -4156 13816 -2780
rect 13868 -4156 13878 -2780
rect 14004 -4156 14014 -2780
rect 14066 -4156 14076 -2780
rect 14202 -4156 14212 -2780
rect 14264 -4156 14274 -2780
rect 14400 -4156 14410 -2780
rect 14462 -4156 14472 -2780
rect 14598 -4156 14608 -2780
rect 14660 -4156 14670 -2780
rect 14796 -4156 14806 -2780
rect 14858 -4156 14868 -2780
rect 14994 -4156 15004 -2780
rect 15056 -4156 15066 -2780
rect 15192 -4156 15202 -2780
rect 15254 -4156 15264 -2780
rect 15390 -4156 15400 -2780
rect 15452 -4156 15462 -2780
rect 15588 -4156 15598 -2780
rect 15650 -4156 15660 -2780
rect 15786 -4156 15796 -2780
rect 15848 -4156 15858 -2780
rect 15984 -4156 15994 -2780
rect 16046 -4156 16056 -2780
rect 16182 -4156 16192 -2780
rect 16244 -4156 16254 -2780
rect 16380 -4156 16390 -2780
rect 16442 -4156 16452 -2780
rect 16578 -4156 16588 -2780
rect 16640 -4156 16650 -2780
rect 16776 -4156 16786 -2780
rect 16838 -4156 16848 -2780
rect 16974 -4156 16984 -2780
rect 17036 -4156 17046 -2780
rect 17172 -4156 17182 -2780
rect 17234 -4156 17244 -2780
rect 17370 -4156 17380 -2780
rect 17432 -4156 17442 -2780
rect 17568 -4156 17578 -2780
rect 17630 -4156 17640 -2780
rect 17766 -4156 17776 -2780
rect 17828 -4156 17838 -2780
rect 17964 -4156 17974 -2780
rect 18026 -4156 18036 -2780
rect 18162 -4156 18172 -2780
rect 18224 -4156 18234 -2780
rect 18360 -4156 18370 -2780
rect 18422 -4156 18432 -2780
rect 18558 -4156 18568 -2780
rect 18620 -4156 18630 -2780
rect 18756 -4156 18766 -2780
rect 18818 -4156 18828 -2780
rect 18954 -4156 18964 -2780
rect 19016 -4156 19026 -2780
rect 19152 -4156 19162 -2780
rect 19214 -4156 19224 -2780
rect 19350 -4156 19360 -2780
rect 19412 -4156 19422 -2780
rect 19548 -4156 19558 -2780
rect 19610 -4156 19620 -2780
rect 19746 -4155 19756 -2779
rect 19808 -4155 19818 -2779
rect 19759 -4156 19765 -4155
rect 19799 -4156 19805 -4155
rect 11443 -4562 11489 -4156
rect 11641 -4168 11687 -4156
rect 11839 -4562 11885 -4156
rect 12037 -4168 12083 -4156
rect 12235 -4562 12281 -4156
rect 12433 -4168 12479 -4156
rect 12631 -4562 12677 -4156
rect 12829 -4168 12875 -4156
rect 13027 -4562 13073 -4156
rect 13225 -4168 13271 -4156
rect 13423 -4562 13469 -4156
rect 13621 -4168 13667 -4156
rect 13819 -4562 13865 -4156
rect 14017 -4168 14063 -4156
rect 14215 -4562 14261 -4156
rect 14413 -4168 14459 -4156
rect 14611 -4562 14657 -4156
rect 14809 -4168 14855 -4156
rect 15007 -4562 15053 -4156
rect 15205 -4168 15251 -4156
rect 15403 -4562 15449 -4156
rect 15601 -4168 15647 -4156
rect 15799 -4562 15845 -4156
rect 15997 -4168 16043 -4156
rect 16195 -4562 16241 -4156
rect 16393 -4168 16439 -4156
rect 16591 -4562 16637 -4156
rect 16789 -4168 16835 -4156
rect 16987 -4562 17033 -4156
rect 17185 -4168 17231 -4156
rect 17383 -4562 17429 -4156
rect 17581 -4168 17627 -4156
rect 17779 -4562 17825 -4156
rect 17977 -4168 18023 -4156
rect 18175 -4562 18221 -4156
rect 18373 -4168 18419 -4156
rect 18571 -4562 18617 -4156
rect 18769 -4168 18815 -4156
rect 18967 -4562 19013 -4156
rect 19165 -4168 19211 -4156
rect 19363 -4562 19409 -4156
rect 19561 -4168 19607 -4156
rect 19759 -4562 19805 -4156
rect 20932 -4562 22152 2327
rect 23293 2128 23339 2327
rect 23491 2128 23537 2140
rect 23689 2128 23735 2327
rect 23887 2128 23933 2140
rect 24085 2128 24131 2327
rect 24283 2128 24329 2140
rect 24481 2128 24527 2327
rect 24679 2128 24725 2140
rect 24877 2128 24923 2327
rect 25075 2128 25121 2140
rect 25273 2128 25319 2327
rect 25471 2128 25517 2140
rect 25669 2128 25715 2327
rect 25867 2128 25913 2140
rect 26065 2128 26111 2327
rect 26263 2128 26309 2140
rect 26461 2128 26507 2327
rect 26659 2128 26705 2140
rect 26857 2128 26903 2327
rect 27055 2128 27101 2140
rect 27253 2128 27299 2327
rect 27451 2128 27497 2140
rect 27649 2128 27695 2327
rect 27847 2128 27893 2140
rect 28045 2128 28091 2327
rect 28243 2128 28289 2140
rect 28441 2128 28487 2327
rect 28639 2128 28685 2140
rect 28837 2128 28883 2327
rect 29035 2128 29081 2140
rect 29233 2128 29279 2327
rect 29431 2128 29477 2140
rect 29629 2128 29675 2327
rect 29827 2128 29873 2140
rect 30025 2128 30071 2327
rect 30223 2128 30269 2140
rect 30421 2128 30467 2327
rect 30619 2128 30665 2140
rect 30817 2128 30863 2327
rect 31015 2128 31061 2140
rect 31213 2128 31259 2327
rect 31411 2128 31457 2140
rect 31609 2129 31655 2327
rect 23280 752 23290 2128
rect 23342 752 23352 2128
rect 23478 752 23488 2128
rect 23540 752 23550 2128
rect 23676 752 23686 2128
rect 23738 752 23748 2128
rect 23874 752 23884 2128
rect 23936 752 23946 2128
rect 24072 752 24082 2128
rect 24134 752 24144 2128
rect 24270 752 24280 2128
rect 24332 752 24342 2128
rect 24468 752 24478 2128
rect 24530 752 24540 2128
rect 24666 752 24676 2128
rect 24728 752 24738 2128
rect 24864 752 24874 2128
rect 24926 752 24936 2128
rect 25062 752 25072 2128
rect 25124 752 25134 2128
rect 25260 752 25270 2128
rect 25322 752 25332 2128
rect 25458 752 25468 2128
rect 25520 752 25530 2128
rect 25656 752 25666 2128
rect 25718 752 25728 2128
rect 25854 752 25864 2128
rect 25916 752 25926 2128
rect 26052 752 26062 2128
rect 26114 752 26124 2128
rect 26250 752 26260 2128
rect 26312 752 26322 2128
rect 26448 752 26458 2128
rect 26510 752 26520 2128
rect 26646 752 26656 2128
rect 26708 752 26718 2128
rect 26844 752 26854 2128
rect 26906 752 26916 2128
rect 27042 752 27052 2128
rect 27104 752 27114 2128
rect 27240 752 27250 2128
rect 27302 752 27312 2128
rect 27438 752 27448 2128
rect 27500 752 27510 2128
rect 27636 752 27646 2128
rect 27698 752 27708 2128
rect 27834 752 27844 2128
rect 27896 752 27906 2128
rect 28032 752 28042 2128
rect 28094 752 28104 2128
rect 28230 752 28240 2128
rect 28292 752 28302 2128
rect 28428 752 28438 2128
rect 28490 752 28500 2128
rect 28626 752 28636 2128
rect 28688 752 28698 2128
rect 28824 752 28834 2128
rect 28886 752 28896 2128
rect 29022 752 29032 2128
rect 29084 752 29094 2128
rect 29220 752 29230 2128
rect 29282 752 29292 2128
rect 29418 752 29428 2128
rect 29480 752 29490 2128
rect 29616 752 29626 2128
rect 29678 752 29688 2128
rect 29814 752 29824 2128
rect 29876 752 29886 2128
rect 30012 752 30022 2128
rect 30074 752 30084 2128
rect 30210 752 30220 2128
rect 30272 752 30282 2128
rect 30408 752 30418 2128
rect 30470 752 30480 2128
rect 30606 752 30616 2128
rect 30668 752 30678 2128
rect 30804 752 30814 2128
rect 30866 752 30876 2128
rect 31002 752 31012 2128
rect 31064 752 31074 2128
rect 31200 752 31210 2128
rect 31262 752 31272 2128
rect 31398 752 31408 2128
rect 31460 752 31470 2128
rect 31596 753 31606 2129
rect 31658 753 31668 2129
rect 31609 752 31615 753
rect 31649 752 31655 753
rect 23293 740 23339 752
rect 23491 740 23537 752
rect 23689 740 23735 752
rect 23887 740 23933 752
rect 24085 740 24131 752
rect 24283 740 24329 752
rect 24481 740 24527 752
rect 24679 740 24725 752
rect 24877 740 24923 752
rect 25075 740 25121 752
rect 25273 740 25319 752
rect 25471 740 25517 752
rect 25669 740 25715 752
rect 25867 740 25913 752
rect 26065 740 26111 752
rect 26263 740 26309 752
rect 26461 740 26507 752
rect 26659 740 26705 752
rect 26857 740 26903 752
rect 27055 740 27101 752
rect 27253 740 27299 752
rect 27451 740 27497 752
rect 27649 740 27695 752
rect 27847 740 27893 752
rect 28045 740 28091 752
rect 28243 740 28289 752
rect 28441 740 28487 752
rect 28639 740 28685 752
rect 28837 740 28883 752
rect 29035 740 29081 752
rect 29233 740 29279 752
rect 29431 740 29477 752
rect 29629 740 29675 752
rect 29827 740 29873 752
rect 30025 740 30071 752
rect 30223 740 30269 752
rect 30421 740 30467 752
rect 30619 740 30665 752
rect 30817 740 30863 752
rect 31015 740 31061 752
rect 31213 740 31259 752
rect 31411 740 31457 752
rect 31609 740 31655 752
rect 23052 693 31896 699
rect 23052 659 23361 693
rect 23469 659 23559 693
rect 23667 659 23757 693
rect 23865 659 23955 693
rect 24063 659 24153 693
rect 24261 659 24351 693
rect 24459 659 24549 693
rect 24657 659 24747 693
rect 24855 659 24945 693
rect 25053 659 25143 693
rect 25251 659 25341 693
rect 25449 659 25539 693
rect 25647 659 25737 693
rect 25845 659 25935 693
rect 26043 659 26133 693
rect 26241 659 26331 693
rect 26439 659 26529 693
rect 26637 659 26727 693
rect 26835 659 26925 693
rect 27033 659 27123 693
rect 27231 659 27321 693
rect 27429 659 27519 693
rect 27627 659 27717 693
rect 27825 659 27915 693
rect 28023 659 28113 693
rect 28221 659 28311 693
rect 28419 659 28509 693
rect 28617 659 28707 693
rect 28815 659 28905 693
rect 29013 659 29103 693
rect 29211 659 29301 693
rect 29409 659 29499 693
rect 29607 659 29697 693
rect 29805 659 29895 693
rect 30003 659 30093 693
rect 30201 659 30291 693
rect 30399 659 30489 693
rect 30597 659 30687 693
rect 30795 659 30885 693
rect 30993 659 31083 693
rect 31191 659 31281 693
rect 31389 659 31479 693
rect 31587 659 31896 693
rect 23052 585 31896 659
rect 23052 551 23361 585
rect 23469 551 23559 585
rect 23667 551 23757 585
rect 23865 551 23955 585
rect 24063 551 24153 585
rect 24261 551 24351 585
rect 24459 551 24549 585
rect 24657 551 24747 585
rect 24855 551 24945 585
rect 25053 551 25143 585
rect 25251 551 25341 585
rect 25449 551 25539 585
rect 25647 551 25737 585
rect 25845 551 25935 585
rect 26043 551 26133 585
rect 26241 551 26331 585
rect 26439 551 26529 585
rect 26637 551 26727 585
rect 26835 551 26925 585
rect 27033 551 27123 585
rect 27231 551 27321 585
rect 27429 551 27519 585
rect 27627 551 27717 585
rect 27825 551 27915 585
rect 28023 551 28113 585
rect 28221 551 28311 585
rect 28419 551 28509 585
rect 28617 551 28707 585
rect 28815 551 28905 585
rect 29013 551 29103 585
rect 29211 551 29301 585
rect 29409 551 29499 585
rect 29607 551 29697 585
rect 29805 551 29895 585
rect 30003 551 30093 585
rect 30201 551 30291 585
rect 30399 551 30489 585
rect 30597 551 30687 585
rect 30795 551 30885 585
rect 30993 551 31083 585
rect 31191 551 31281 585
rect 31389 551 31479 585
rect 31587 551 31896 585
rect 23052 545 31896 551
rect 23052 -743 23206 545
rect 23293 492 23339 504
rect 23491 492 23537 504
rect 23689 492 23735 504
rect 23887 492 23933 504
rect 24085 492 24131 504
rect 24283 492 24329 504
rect 24481 492 24527 504
rect 24679 492 24725 504
rect 24877 492 24923 504
rect 25075 492 25121 504
rect 25273 492 25319 504
rect 25471 492 25517 504
rect 25669 492 25715 504
rect 25867 492 25913 504
rect 26065 492 26111 504
rect 26263 492 26309 504
rect 26461 492 26507 504
rect 26659 492 26705 504
rect 26857 492 26903 504
rect 27055 492 27101 504
rect 27253 492 27299 504
rect 27451 492 27497 504
rect 27649 492 27695 504
rect 27847 492 27893 504
rect 28045 492 28091 504
rect 28243 492 28289 504
rect 28441 492 28487 504
rect 28639 492 28685 504
rect 28837 492 28883 504
rect 29035 492 29081 504
rect 29233 492 29279 504
rect 29431 492 29477 504
rect 29629 492 29675 504
rect 29827 492 29873 504
rect 30025 492 30071 504
rect 30223 492 30269 504
rect 30421 492 30467 504
rect 30619 492 30665 504
rect 30817 492 30863 504
rect 31015 492 31061 504
rect 31213 492 31259 504
rect 31411 492 31457 504
rect 31609 493 31655 504
rect 23052 -877 23062 -743
rect 23196 -877 23206 -743
rect 23052 -937 23206 -877
rect 23280 -884 23290 492
rect 23342 -884 23352 492
rect 23478 -884 23488 492
rect 23540 -884 23550 492
rect 23676 -884 23686 492
rect 23738 -884 23748 492
rect 23874 -884 23884 492
rect 23936 -884 23946 492
rect 24072 -884 24082 492
rect 24134 -884 24144 492
rect 24270 -884 24280 492
rect 24332 -884 24342 492
rect 24468 -884 24478 492
rect 24530 -884 24540 492
rect 24666 -884 24676 492
rect 24728 -884 24738 492
rect 24864 -884 24874 492
rect 24926 -884 24936 492
rect 25062 -884 25072 492
rect 25124 -884 25134 492
rect 25260 -884 25270 492
rect 25322 -884 25332 492
rect 25458 -884 25468 492
rect 25520 -884 25530 492
rect 25656 -884 25666 492
rect 25718 -884 25728 492
rect 25854 -884 25864 492
rect 25916 -884 25926 492
rect 26052 -884 26062 492
rect 26114 -884 26124 492
rect 26250 -884 26260 492
rect 26312 -884 26322 492
rect 26448 -884 26458 492
rect 26510 -884 26520 492
rect 26646 -884 26656 492
rect 26708 -884 26718 492
rect 26844 -884 26854 492
rect 26906 -884 26916 492
rect 27042 -884 27052 492
rect 27104 -884 27114 492
rect 27240 -884 27250 492
rect 27302 -884 27312 492
rect 27438 -884 27448 492
rect 27500 -884 27510 492
rect 27636 -884 27646 492
rect 27698 -884 27708 492
rect 27834 -884 27844 492
rect 27896 -884 27906 492
rect 28032 -884 28042 492
rect 28094 -884 28104 492
rect 28230 -884 28240 492
rect 28292 -884 28302 492
rect 28428 -884 28438 492
rect 28490 -884 28500 492
rect 28626 -884 28636 492
rect 28688 -884 28698 492
rect 28824 -884 28834 492
rect 28886 -884 28896 492
rect 29022 -884 29032 492
rect 29084 -884 29094 492
rect 29220 -884 29230 492
rect 29282 -884 29292 492
rect 29418 -884 29428 492
rect 29480 -884 29490 492
rect 29616 -884 29626 492
rect 29678 -884 29688 492
rect 29814 -884 29824 492
rect 29876 -884 29886 492
rect 30012 -884 30022 492
rect 30074 -884 30084 492
rect 30210 -884 30220 492
rect 30272 -884 30282 492
rect 30408 -884 30418 492
rect 30470 -884 30480 492
rect 30606 -884 30616 492
rect 30668 -884 30678 492
rect 30804 -884 30814 492
rect 30866 -884 30876 492
rect 31002 -884 31012 492
rect 31064 -884 31074 492
rect 31200 -884 31210 492
rect 31262 -884 31272 492
rect 31398 -884 31408 492
rect 31460 -884 31470 492
rect 31596 -883 31606 493
rect 31658 -883 31668 493
rect 31609 -884 31615 -883
rect 31649 -884 31655 -883
rect 23293 -896 23339 -884
rect 23491 -896 23537 -884
rect 23689 -896 23735 -884
rect 23887 -896 23933 -884
rect 24085 -896 24131 -884
rect 24283 -896 24329 -884
rect 24481 -896 24527 -884
rect 24679 -896 24725 -884
rect 24877 -896 24923 -884
rect 25075 -896 25121 -884
rect 25273 -896 25319 -884
rect 25471 -896 25517 -884
rect 25669 -896 25715 -884
rect 25867 -896 25913 -884
rect 26065 -896 26111 -884
rect 26263 -896 26309 -884
rect 26461 -896 26507 -884
rect 26659 -896 26705 -884
rect 26857 -896 26903 -884
rect 27055 -896 27101 -884
rect 27253 -896 27299 -884
rect 27451 -896 27497 -884
rect 27649 -896 27695 -884
rect 27847 -896 27893 -884
rect 28045 -896 28091 -884
rect 28243 -896 28289 -884
rect 28441 -896 28487 -884
rect 28639 -896 28685 -884
rect 28837 -896 28883 -884
rect 29035 -896 29081 -884
rect 29233 -896 29279 -884
rect 29431 -896 29477 -884
rect 29629 -896 29675 -884
rect 29827 -896 29873 -884
rect 30025 -896 30071 -884
rect 30223 -896 30269 -884
rect 30421 -896 30467 -884
rect 30619 -896 30665 -884
rect 30817 -896 30863 -884
rect 31015 -896 31061 -884
rect 31213 -896 31259 -884
rect 31411 -896 31457 -884
rect 31609 -896 31655 -884
rect 31742 -937 31896 545
rect 23052 -943 31896 -937
rect 23052 -947 23361 -943
rect 23052 -1081 23062 -947
rect 23196 -977 23361 -947
rect 23469 -977 23559 -943
rect 23667 -977 23757 -943
rect 23865 -977 23955 -943
rect 24063 -977 24153 -943
rect 24261 -977 24351 -943
rect 24459 -977 24549 -943
rect 24657 -977 24747 -943
rect 24855 -977 24945 -943
rect 25053 -977 25143 -943
rect 25251 -977 25341 -943
rect 25449 -977 25539 -943
rect 25647 -977 25737 -943
rect 25845 -977 25935 -943
rect 26043 -977 26133 -943
rect 26241 -977 26331 -943
rect 26439 -977 26529 -943
rect 26637 -977 26727 -943
rect 26835 -977 26925 -943
rect 27033 -977 27123 -943
rect 27231 -977 27321 -943
rect 27429 -977 27519 -943
rect 27627 -977 27717 -943
rect 27825 -977 27915 -943
rect 28023 -977 28113 -943
rect 28221 -977 28311 -943
rect 28419 -977 28509 -943
rect 28617 -977 28707 -943
rect 28815 -977 28905 -943
rect 29013 -977 29103 -943
rect 29211 -977 29301 -943
rect 29409 -977 29499 -943
rect 29607 -977 29697 -943
rect 29805 -977 29895 -943
rect 30003 -977 30093 -943
rect 30201 -977 30291 -943
rect 30399 -977 30489 -943
rect 30597 -977 30687 -943
rect 30795 -977 30885 -943
rect 30993 -977 31083 -943
rect 31191 -977 31281 -943
rect 31389 -977 31479 -943
rect 31587 -977 31896 -943
rect 23196 -1051 31896 -977
rect 23196 -1081 23361 -1051
rect 23052 -1085 23361 -1081
rect 23469 -1085 23559 -1051
rect 23667 -1085 23757 -1051
rect 23865 -1085 23955 -1051
rect 24063 -1085 24153 -1051
rect 24261 -1085 24351 -1051
rect 24459 -1085 24549 -1051
rect 24657 -1085 24747 -1051
rect 24855 -1085 24945 -1051
rect 25053 -1085 25143 -1051
rect 25251 -1085 25341 -1051
rect 25449 -1085 25539 -1051
rect 25647 -1085 25737 -1051
rect 25845 -1085 25935 -1051
rect 26043 -1085 26133 -1051
rect 26241 -1085 26331 -1051
rect 26439 -1085 26529 -1051
rect 26637 -1085 26727 -1051
rect 26835 -1085 26925 -1051
rect 27033 -1085 27123 -1051
rect 27231 -1085 27321 -1051
rect 27429 -1085 27519 -1051
rect 27627 -1085 27717 -1051
rect 27825 -1085 27915 -1051
rect 28023 -1085 28113 -1051
rect 28221 -1085 28311 -1051
rect 28419 -1085 28509 -1051
rect 28617 -1085 28707 -1051
rect 28815 -1085 28905 -1051
rect 29013 -1085 29103 -1051
rect 29211 -1085 29301 -1051
rect 29409 -1085 29499 -1051
rect 29607 -1085 29697 -1051
rect 29805 -1085 29895 -1051
rect 30003 -1085 30093 -1051
rect 30201 -1085 30291 -1051
rect 30399 -1085 30489 -1051
rect 30597 -1085 30687 -1051
rect 30795 -1085 30885 -1051
rect 30993 -1085 31083 -1051
rect 31191 -1085 31281 -1051
rect 31389 -1085 31479 -1051
rect 31587 -1085 31896 -1051
rect 23052 -1091 31896 -1085
rect 23052 -1151 23206 -1091
rect 23293 -1144 23339 -1132
rect 23491 -1144 23537 -1132
rect 23689 -1144 23735 -1132
rect 23887 -1144 23933 -1132
rect 24085 -1144 24131 -1132
rect 24283 -1144 24329 -1132
rect 24481 -1144 24527 -1132
rect 24679 -1144 24725 -1132
rect 24877 -1144 24923 -1132
rect 25075 -1144 25121 -1132
rect 25273 -1144 25319 -1132
rect 25471 -1144 25517 -1132
rect 25669 -1144 25715 -1132
rect 25867 -1144 25913 -1132
rect 26065 -1144 26111 -1132
rect 26263 -1144 26309 -1132
rect 26461 -1144 26507 -1132
rect 26659 -1144 26705 -1132
rect 26857 -1144 26903 -1132
rect 27055 -1144 27101 -1132
rect 27253 -1144 27299 -1132
rect 27451 -1144 27497 -1132
rect 27649 -1144 27695 -1132
rect 27847 -1144 27893 -1132
rect 28045 -1144 28091 -1132
rect 28243 -1144 28289 -1132
rect 28441 -1144 28487 -1132
rect 28639 -1144 28685 -1132
rect 28837 -1144 28883 -1132
rect 29035 -1144 29081 -1132
rect 29233 -1144 29279 -1132
rect 29431 -1144 29477 -1132
rect 29629 -1144 29675 -1132
rect 29827 -1144 29873 -1132
rect 30025 -1144 30071 -1132
rect 30223 -1144 30269 -1132
rect 30421 -1144 30467 -1132
rect 30619 -1144 30665 -1132
rect 30817 -1144 30863 -1132
rect 31015 -1144 31061 -1132
rect 31213 -1144 31259 -1132
rect 31411 -1144 31457 -1132
rect 31609 -1143 31655 -1132
rect 23052 -1285 23062 -1151
rect 23196 -1285 23206 -1151
rect 23052 -2573 23206 -1285
rect 23280 -2520 23290 -1144
rect 23342 -2520 23352 -1144
rect 23478 -2520 23488 -1144
rect 23540 -2520 23550 -1144
rect 23676 -2520 23686 -1144
rect 23738 -2520 23748 -1144
rect 23874 -2520 23884 -1144
rect 23936 -2520 23946 -1144
rect 24072 -2520 24082 -1144
rect 24134 -2520 24144 -1144
rect 24270 -2520 24280 -1144
rect 24332 -2520 24342 -1144
rect 24468 -2520 24478 -1144
rect 24530 -2520 24540 -1144
rect 24666 -2520 24676 -1144
rect 24728 -2520 24738 -1144
rect 24864 -2520 24874 -1144
rect 24926 -2520 24936 -1144
rect 25062 -2520 25072 -1144
rect 25124 -2520 25134 -1144
rect 25260 -2520 25270 -1144
rect 25322 -2520 25332 -1144
rect 25458 -2520 25468 -1144
rect 25520 -2520 25530 -1144
rect 25656 -2520 25666 -1144
rect 25718 -2520 25728 -1144
rect 25854 -2520 25864 -1144
rect 25916 -2520 25926 -1144
rect 26052 -2520 26062 -1144
rect 26114 -2520 26124 -1144
rect 26250 -2520 26260 -1144
rect 26312 -2520 26322 -1144
rect 26448 -2520 26458 -1144
rect 26510 -2520 26520 -1144
rect 26646 -2520 26656 -1144
rect 26708 -2520 26718 -1144
rect 26844 -2520 26854 -1144
rect 26906 -2520 26916 -1144
rect 27042 -2520 27052 -1144
rect 27104 -2520 27114 -1144
rect 27240 -2520 27250 -1144
rect 27302 -2520 27312 -1144
rect 27438 -2520 27448 -1144
rect 27500 -2520 27510 -1144
rect 27636 -2520 27646 -1144
rect 27698 -2520 27708 -1144
rect 27834 -2520 27844 -1144
rect 27896 -2520 27906 -1144
rect 28032 -2520 28042 -1144
rect 28094 -2520 28104 -1144
rect 28230 -2520 28240 -1144
rect 28292 -2520 28302 -1144
rect 28428 -2520 28438 -1144
rect 28490 -2520 28500 -1144
rect 28626 -2520 28636 -1144
rect 28688 -2520 28698 -1144
rect 28824 -2520 28834 -1144
rect 28886 -2520 28896 -1144
rect 29022 -2520 29032 -1144
rect 29084 -2520 29094 -1144
rect 29220 -2520 29230 -1144
rect 29282 -2520 29292 -1144
rect 29418 -2520 29428 -1144
rect 29480 -2520 29490 -1144
rect 29616 -2520 29626 -1144
rect 29678 -2520 29688 -1144
rect 29814 -2520 29824 -1144
rect 29876 -2520 29886 -1144
rect 30012 -2520 30022 -1144
rect 30074 -2520 30084 -1144
rect 30210 -2520 30220 -1144
rect 30272 -2520 30282 -1144
rect 30408 -2520 30418 -1144
rect 30470 -2520 30480 -1144
rect 30606 -2520 30616 -1144
rect 30668 -2520 30678 -1144
rect 30804 -2520 30814 -1144
rect 30866 -2520 30876 -1144
rect 31002 -2520 31012 -1144
rect 31064 -2520 31074 -1144
rect 31200 -2520 31210 -1144
rect 31262 -2520 31272 -1144
rect 31398 -2520 31408 -1144
rect 31460 -2520 31470 -1144
rect 31596 -2519 31606 -1143
rect 31658 -2519 31668 -1143
rect 31609 -2520 31615 -2519
rect 31649 -2520 31655 -2519
rect 23293 -2532 23339 -2520
rect 23491 -2532 23537 -2520
rect 23689 -2532 23735 -2520
rect 23887 -2532 23933 -2520
rect 24085 -2532 24131 -2520
rect 24283 -2532 24329 -2520
rect 24481 -2532 24527 -2520
rect 24679 -2532 24725 -2520
rect 24877 -2532 24923 -2520
rect 25075 -2532 25121 -2520
rect 25273 -2532 25319 -2520
rect 25471 -2532 25517 -2520
rect 25669 -2532 25715 -2520
rect 25867 -2532 25913 -2520
rect 26065 -2532 26111 -2520
rect 26263 -2532 26309 -2520
rect 26461 -2532 26507 -2520
rect 26659 -2532 26705 -2520
rect 26857 -2532 26903 -2520
rect 27055 -2532 27101 -2520
rect 27253 -2532 27299 -2520
rect 27451 -2532 27497 -2520
rect 27649 -2532 27695 -2520
rect 27847 -2532 27893 -2520
rect 28045 -2532 28091 -2520
rect 28243 -2532 28289 -2520
rect 28441 -2532 28487 -2520
rect 28639 -2532 28685 -2520
rect 28837 -2532 28883 -2520
rect 29035 -2532 29081 -2520
rect 29233 -2532 29279 -2520
rect 29431 -2532 29477 -2520
rect 29629 -2532 29675 -2520
rect 29827 -2532 29873 -2520
rect 30025 -2532 30071 -2520
rect 30223 -2532 30269 -2520
rect 30421 -2532 30467 -2520
rect 30619 -2532 30665 -2520
rect 30817 -2532 30863 -2520
rect 31015 -2532 31061 -2520
rect 31213 -2532 31259 -2520
rect 31411 -2532 31457 -2520
rect 31609 -2532 31655 -2520
rect 31742 -2573 31896 -1091
rect 23052 -2579 31896 -2573
rect 23052 -2613 23361 -2579
rect 23469 -2613 23559 -2579
rect 23667 -2613 23757 -2579
rect 23865 -2613 23955 -2579
rect 24063 -2613 24153 -2579
rect 24261 -2613 24351 -2579
rect 24459 -2613 24549 -2579
rect 24657 -2613 24747 -2579
rect 24855 -2613 24945 -2579
rect 25053 -2613 25143 -2579
rect 25251 -2613 25341 -2579
rect 25449 -2613 25539 -2579
rect 25647 -2613 25737 -2579
rect 25845 -2613 25935 -2579
rect 26043 -2613 26133 -2579
rect 26241 -2613 26331 -2579
rect 26439 -2613 26529 -2579
rect 26637 -2613 26727 -2579
rect 26835 -2613 26925 -2579
rect 27033 -2613 27123 -2579
rect 27231 -2613 27321 -2579
rect 27429 -2613 27519 -2579
rect 27627 -2613 27717 -2579
rect 27825 -2613 27915 -2579
rect 28023 -2613 28113 -2579
rect 28221 -2613 28311 -2579
rect 28419 -2613 28509 -2579
rect 28617 -2613 28707 -2579
rect 28815 -2613 28905 -2579
rect 29013 -2613 29103 -2579
rect 29211 -2613 29301 -2579
rect 29409 -2613 29499 -2579
rect 29607 -2613 29697 -2579
rect 29805 -2613 29895 -2579
rect 30003 -2613 30093 -2579
rect 30201 -2613 30291 -2579
rect 30399 -2613 30489 -2579
rect 30597 -2613 30687 -2579
rect 30795 -2613 30885 -2579
rect 30993 -2613 31083 -2579
rect 31191 -2613 31281 -2579
rect 31389 -2613 31479 -2579
rect 31587 -2613 31896 -2579
rect 23052 -2687 31896 -2613
rect 23052 -2721 23361 -2687
rect 23469 -2721 23559 -2687
rect 23667 -2721 23757 -2687
rect 23865 -2721 23955 -2687
rect 24063 -2721 24153 -2687
rect 24261 -2721 24351 -2687
rect 24459 -2721 24549 -2687
rect 24657 -2721 24747 -2687
rect 24855 -2721 24945 -2687
rect 25053 -2721 25143 -2687
rect 25251 -2721 25341 -2687
rect 25449 -2721 25539 -2687
rect 25647 -2721 25737 -2687
rect 25845 -2721 25935 -2687
rect 26043 -2721 26133 -2687
rect 26241 -2721 26331 -2687
rect 26439 -2721 26529 -2687
rect 26637 -2721 26727 -2687
rect 26835 -2721 26925 -2687
rect 27033 -2721 27123 -2687
rect 27231 -2721 27321 -2687
rect 27429 -2721 27519 -2687
rect 27627 -2721 27717 -2687
rect 27825 -2721 27915 -2687
rect 28023 -2721 28113 -2687
rect 28221 -2721 28311 -2687
rect 28419 -2721 28509 -2687
rect 28617 -2721 28707 -2687
rect 28815 -2721 28905 -2687
rect 29013 -2721 29103 -2687
rect 29211 -2721 29301 -2687
rect 29409 -2721 29499 -2687
rect 29607 -2721 29697 -2687
rect 29805 -2721 29895 -2687
rect 30003 -2721 30093 -2687
rect 30201 -2721 30291 -2687
rect 30399 -2721 30489 -2687
rect 30597 -2721 30687 -2687
rect 30795 -2721 30885 -2687
rect 30993 -2721 31083 -2687
rect 31191 -2721 31281 -2687
rect 31389 -2721 31479 -2687
rect 31587 -2721 31896 -2687
rect 23052 -2727 31896 -2721
rect 23293 -2780 23339 -2768
rect 23491 -2780 23537 -2768
rect 23689 -2780 23735 -2768
rect 23887 -2780 23933 -2768
rect 24085 -2780 24131 -2768
rect 24283 -2780 24329 -2768
rect 24481 -2780 24527 -2768
rect 24679 -2780 24725 -2768
rect 24877 -2780 24923 -2768
rect 25075 -2780 25121 -2768
rect 25273 -2780 25319 -2768
rect 25471 -2780 25517 -2768
rect 25669 -2780 25715 -2768
rect 25867 -2780 25913 -2768
rect 26065 -2780 26111 -2768
rect 26263 -2780 26309 -2768
rect 26461 -2780 26507 -2768
rect 26659 -2780 26705 -2768
rect 26857 -2780 26903 -2768
rect 27055 -2780 27101 -2768
rect 27253 -2780 27299 -2768
rect 27451 -2780 27497 -2768
rect 27649 -2780 27695 -2768
rect 27847 -2780 27893 -2768
rect 28045 -2780 28091 -2768
rect 28243 -2780 28289 -2768
rect 28441 -2780 28487 -2768
rect 28639 -2780 28685 -2768
rect 28837 -2780 28883 -2768
rect 29035 -2780 29081 -2768
rect 29233 -2780 29279 -2768
rect 29431 -2780 29477 -2768
rect 29629 -2780 29675 -2768
rect 29827 -2780 29873 -2768
rect 30025 -2780 30071 -2768
rect 30223 -2780 30269 -2768
rect 30421 -2780 30467 -2768
rect 30619 -2780 30665 -2768
rect 30817 -2780 30863 -2768
rect 31015 -2780 31061 -2768
rect 31213 -2780 31259 -2768
rect 31411 -2780 31457 -2768
rect 31609 -2779 31655 -2768
rect 23280 -4156 23290 -2780
rect 23342 -4156 23352 -2780
rect 23478 -4156 23488 -2780
rect 23540 -4156 23550 -2780
rect 23676 -4156 23686 -2780
rect 23738 -4156 23748 -2780
rect 23874 -4156 23884 -2780
rect 23936 -4156 23946 -2780
rect 24072 -4156 24082 -2780
rect 24134 -4156 24144 -2780
rect 24270 -4156 24280 -2780
rect 24332 -4156 24342 -2780
rect 24468 -4156 24478 -2780
rect 24530 -4156 24540 -2780
rect 24666 -4156 24676 -2780
rect 24728 -4156 24738 -2780
rect 24864 -4156 24874 -2780
rect 24926 -4156 24936 -2780
rect 25062 -4156 25072 -2780
rect 25124 -4156 25134 -2780
rect 25260 -4156 25270 -2780
rect 25322 -4156 25332 -2780
rect 25458 -4156 25468 -2780
rect 25520 -4156 25530 -2780
rect 25656 -4156 25666 -2780
rect 25718 -4156 25728 -2780
rect 25854 -4156 25864 -2780
rect 25916 -4156 25926 -2780
rect 26052 -4156 26062 -2780
rect 26114 -4156 26124 -2780
rect 26250 -4156 26260 -2780
rect 26312 -4156 26322 -2780
rect 26448 -4156 26458 -2780
rect 26510 -4156 26520 -2780
rect 26646 -4156 26656 -2780
rect 26708 -4156 26718 -2780
rect 26844 -4156 26854 -2780
rect 26906 -4156 26916 -2780
rect 27042 -4156 27052 -2780
rect 27104 -4156 27114 -2780
rect 27240 -4156 27250 -2780
rect 27302 -4156 27312 -2780
rect 27438 -4156 27448 -2780
rect 27500 -4156 27510 -2780
rect 27636 -4156 27646 -2780
rect 27698 -4156 27708 -2780
rect 27834 -4156 27844 -2780
rect 27896 -4156 27906 -2780
rect 28032 -4156 28042 -2780
rect 28094 -4156 28104 -2780
rect 28230 -4156 28240 -2780
rect 28292 -4156 28302 -2780
rect 28428 -4156 28438 -2780
rect 28490 -4156 28500 -2780
rect 28626 -4156 28636 -2780
rect 28688 -4156 28698 -2780
rect 28824 -4156 28834 -2780
rect 28886 -4156 28896 -2780
rect 29022 -4156 29032 -2780
rect 29084 -4156 29094 -2780
rect 29220 -4156 29230 -2780
rect 29282 -4156 29292 -2780
rect 29418 -4156 29428 -2780
rect 29480 -4156 29490 -2780
rect 29616 -4156 29626 -2780
rect 29678 -4156 29688 -2780
rect 29814 -4156 29824 -2780
rect 29876 -4156 29886 -2780
rect 30012 -4156 30022 -2780
rect 30074 -4156 30084 -2780
rect 30210 -4156 30220 -2780
rect 30272 -4156 30282 -2780
rect 30408 -4156 30418 -2780
rect 30470 -4156 30480 -2780
rect 30606 -4156 30616 -2780
rect 30668 -4156 30678 -2780
rect 30804 -4156 30814 -2780
rect 30866 -4156 30876 -2780
rect 31002 -4156 31012 -2780
rect 31064 -4156 31074 -2780
rect 31200 -4156 31210 -2780
rect 31262 -4156 31272 -2780
rect 31398 -4156 31408 -2780
rect 31460 -4156 31470 -2780
rect 31596 -4155 31606 -2779
rect 31658 -4155 31668 -2779
rect 31609 -4156 31615 -4155
rect 31649 -4156 31655 -4155
rect 23293 -4562 23339 -4156
rect 23491 -4168 23537 -4156
rect 23689 -4562 23735 -4156
rect 23887 -4168 23933 -4156
rect 24085 -4562 24131 -4156
rect 24283 -4168 24329 -4156
rect 24481 -4562 24527 -4156
rect 24679 -4168 24725 -4156
rect 24877 -4562 24923 -4156
rect 25075 -4168 25121 -4156
rect 25273 -4562 25319 -4156
rect 25471 -4168 25517 -4156
rect 25669 -4562 25715 -4156
rect 25867 -4168 25913 -4156
rect 26065 -4562 26111 -4156
rect 26263 -4168 26309 -4156
rect 26461 -4562 26507 -4156
rect 26659 -4168 26705 -4156
rect 26857 -4562 26903 -4156
rect 27055 -4168 27101 -4156
rect 27253 -4562 27299 -4156
rect 27451 -4168 27497 -4156
rect 27649 -4562 27695 -4156
rect 27847 -4168 27893 -4156
rect 28045 -4562 28091 -4156
rect 28243 -4168 28289 -4156
rect 28441 -4562 28487 -4156
rect 28639 -4168 28685 -4156
rect 28837 -4562 28883 -4156
rect 29035 -4168 29081 -4156
rect 29233 -4562 29279 -4156
rect 29431 -4168 29477 -4156
rect 29629 -4562 29675 -4156
rect 29827 -4168 29873 -4156
rect 30025 -4562 30071 -4156
rect 30223 -4168 30269 -4156
rect 30421 -4562 30467 -4156
rect 30619 -4168 30665 -4156
rect 30817 -4562 30863 -4156
rect 31015 -4168 31061 -4156
rect 31213 -4562 31259 -4156
rect 31411 -4168 31457 -4156
rect 31609 -4562 31655 -4156
rect 32606 -4562 33826 2327
rect -753 -5513 33826 -4562
<< via1 >>
rect -399 752 -347 2128
rect -201 752 -149 2128
rect -3 752 49 2128
rect 195 752 247 2128
rect 393 752 445 2128
rect 591 752 643 2128
rect 789 752 841 2128
rect 987 752 1039 2128
rect 1185 752 1237 2128
rect 1383 752 1435 2128
rect 1581 752 1633 2128
rect 1779 752 1831 2128
rect 1977 752 2029 2128
rect 2175 752 2227 2128
rect 2373 752 2425 2128
rect 2571 752 2623 2128
rect 2769 752 2821 2128
rect 2967 752 3019 2128
rect 3165 752 3217 2128
rect 3363 752 3415 2128
rect 3561 752 3613 2128
rect 3759 752 3811 2128
rect 3957 752 4009 2128
rect 4155 752 4207 2128
rect 4353 752 4405 2128
rect 4551 752 4603 2128
rect 4749 752 4801 2128
rect 4947 752 4999 2128
rect 5145 752 5197 2128
rect 5343 752 5395 2128
rect 5541 752 5593 2128
rect 5739 752 5791 2128
rect 5937 752 5989 2128
rect 6135 752 6187 2128
rect 6333 752 6385 2128
rect 6531 752 6583 2128
rect 6729 752 6781 2128
rect 6927 752 6979 2128
rect 7125 752 7177 2128
rect 7323 752 7375 2128
rect 7521 752 7573 2128
rect 7719 752 7771 2128
rect 7917 753 7969 2129
rect -627 -877 -493 -743
rect -399 -884 -347 492
rect -201 -884 -149 492
rect -3 -884 49 492
rect 195 -884 247 492
rect 393 -884 445 492
rect 591 -884 643 492
rect 789 -884 841 492
rect 987 -884 1039 492
rect 1185 -884 1237 492
rect 1383 -884 1435 492
rect 1581 -884 1633 492
rect 1779 -884 1831 492
rect 1977 -884 2029 492
rect 2175 -884 2227 492
rect 2373 -884 2425 492
rect 2571 -884 2623 492
rect 2769 -884 2821 492
rect 2967 -884 3019 492
rect 3165 -884 3217 492
rect 3363 -884 3415 492
rect 3561 -884 3613 492
rect 3759 -884 3811 492
rect 3957 -884 4009 492
rect 4155 -884 4207 492
rect 4353 -884 4405 492
rect 4551 -884 4603 492
rect 4749 -884 4801 492
rect 4947 -884 4999 492
rect 5145 -884 5197 492
rect 5343 -884 5395 492
rect 5541 -884 5593 492
rect 5739 -884 5791 492
rect 5937 -884 5989 492
rect 6135 -884 6187 492
rect 6333 -884 6385 492
rect 6531 -884 6583 492
rect 6729 -884 6781 492
rect 6927 -884 6979 492
rect 7125 -884 7177 492
rect 7323 -884 7375 492
rect 7521 -884 7573 492
rect 7719 -884 7771 492
rect 7917 -883 7969 493
rect 8063 -877 8197 -743
rect -627 -1081 -493 -947
rect 8063 -1081 8197 -947
rect -627 -1285 -493 -1151
rect -399 -2520 -347 -1144
rect -201 -2520 -149 -1144
rect -3 -2520 49 -1144
rect 195 -2520 247 -1144
rect 393 -2520 445 -1144
rect 591 -2520 643 -1144
rect 789 -2520 841 -1144
rect 987 -2520 1039 -1144
rect 1185 -2520 1237 -1144
rect 1383 -2520 1435 -1144
rect 1581 -2520 1633 -1144
rect 1779 -2520 1831 -1144
rect 1977 -2520 2029 -1144
rect 2175 -2520 2227 -1144
rect 2373 -2520 2425 -1144
rect 2571 -2520 2623 -1144
rect 2769 -2520 2821 -1144
rect 2967 -2520 3019 -1144
rect 3165 -2520 3217 -1144
rect 3363 -2520 3415 -1144
rect 3561 -2520 3613 -1144
rect 3759 -2520 3811 -1144
rect 3957 -2520 4009 -1144
rect 4155 -2520 4207 -1144
rect 4353 -2520 4405 -1144
rect 4551 -2520 4603 -1144
rect 4749 -2520 4801 -1144
rect 4947 -2520 4999 -1144
rect 5145 -2520 5197 -1144
rect 5343 -2520 5395 -1144
rect 5541 -2520 5593 -1144
rect 5739 -2520 5791 -1144
rect 5937 -2520 5989 -1144
rect 6135 -2520 6187 -1144
rect 6333 -2520 6385 -1144
rect 6531 -2520 6583 -1144
rect 6729 -2520 6781 -1144
rect 6927 -2520 6979 -1144
rect 7125 -2520 7177 -1144
rect 7323 -2520 7375 -1144
rect 7521 -2520 7573 -1144
rect 7719 -2520 7771 -1144
rect 7917 -2519 7969 -1143
rect 8063 -1285 8197 -1151
rect -399 -4156 -347 -2780
rect -201 -4156 -149 -2780
rect -3 -4156 49 -2780
rect 195 -4156 247 -2780
rect 393 -4156 445 -2780
rect 591 -4156 643 -2780
rect 789 -4156 841 -2780
rect 987 -4156 1039 -2780
rect 1185 -4156 1237 -2780
rect 1383 -4156 1435 -2780
rect 1581 -4156 1633 -2780
rect 1779 -4156 1831 -2780
rect 1977 -4156 2029 -2780
rect 2175 -4156 2227 -2780
rect 2373 -4156 2425 -2780
rect 2571 -4156 2623 -2780
rect 2769 -4156 2821 -2780
rect 2967 -4156 3019 -2780
rect 3165 -4156 3217 -2780
rect 3363 -4156 3415 -2780
rect 3561 -4156 3613 -2780
rect 3759 -4156 3811 -2780
rect 3957 -4156 4009 -2780
rect 4155 -4156 4207 -2780
rect 4353 -4156 4405 -2780
rect 4551 -4156 4603 -2780
rect 4749 -4156 4801 -2780
rect 4947 -4156 4999 -2780
rect 5145 -4156 5197 -2780
rect 5343 -4156 5395 -2780
rect 5541 -4156 5593 -2780
rect 5739 -4156 5791 -2780
rect 5937 -4156 5989 -2780
rect 6135 -4156 6187 -2780
rect 6333 -4156 6385 -2780
rect 6531 -4156 6583 -2780
rect 6729 -4156 6781 -2780
rect 6927 -4156 6979 -2780
rect 7125 -4156 7177 -2780
rect 7323 -4156 7375 -2780
rect 7521 -4156 7573 -2780
rect 7719 -4156 7771 -2780
rect 7917 -4155 7969 -2779
rect 11440 752 11449 2128
rect 11449 752 11483 2128
rect 11483 752 11492 2128
rect 11638 752 11647 2128
rect 11647 752 11681 2128
rect 11681 752 11690 2128
rect 11836 752 11845 2128
rect 11845 752 11879 2128
rect 11879 752 11888 2128
rect 12034 752 12043 2128
rect 12043 752 12077 2128
rect 12077 752 12086 2128
rect 12232 752 12241 2128
rect 12241 752 12275 2128
rect 12275 752 12284 2128
rect 12430 752 12439 2128
rect 12439 752 12473 2128
rect 12473 752 12482 2128
rect 12628 752 12637 2128
rect 12637 752 12671 2128
rect 12671 752 12680 2128
rect 12826 752 12835 2128
rect 12835 752 12869 2128
rect 12869 752 12878 2128
rect 13024 752 13033 2128
rect 13033 752 13067 2128
rect 13067 752 13076 2128
rect 13222 752 13231 2128
rect 13231 752 13265 2128
rect 13265 752 13274 2128
rect 13420 752 13429 2128
rect 13429 752 13463 2128
rect 13463 752 13472 2128
rect 13618 752 13627 2128
rect 13627 752 13661 2128
rect 13661 752 13670 2128
rect 13816 752 13825 2128
rect 13825 752 13859 2128
rect 13859 752 13868 2128
rect 14014 752 14023 2128
rect 14023 752 14057 2128
rect 14057 752 14066 2128
rect 14212 752 14221 2128
rect 14221 752 14255 2128
rect 14255 752 14264 2128
rect 14410 752 14419 2128
rect 14419 752 14453 2128
rect 14453 752 14462 2128
rect 14608 752 14617 2128
rect 14617 752 14651 2128
rect 14651 752 14660 2128
rect 14806 752 14815 2128
rect 14815 752 14849 2128
rect 14849 752 14858 2128
rect 15004 752 15013 2128
rect 15013 752 15047 2128
rect 15047 752 15056 2128
rect 15202 752 15211 2128
rect 15211 752 15245 2128
rect 15245 752 15254 2128
rect 15400 752 15409 2128
rect 15409 752 15443 2128
rect 15443 752 15452 2128
rect 15598 752 15607 2128
rect 15607 752 15641 2128
rect 15641 752 15650 2128
rect 15796 752 15805 2128
rect 15805 752 15839 2128
rect 15839 752 15848 2128
rect 15994 752 16003 2128
rect 16003 752 16037 2128
rect 16037 752 16046 2128
rect 16192 752 16201 2128
rect 16201 752 16235 2128
rect 16235 752 16244 2128
rect 16390 752 16399 2128
rect 16399 752 16433 2128
rect 16433 752 16442 2128
rect 16588 752 16597 2128
rect 16597 752 16631 2128
rect 16631 752 16640 2128
rect 16786 752 16795 2128
rect 16795 752 16829 2128
rect 16829 752 16838 2128
rect 16984 752 16993 2128
rect 16993 752 17027 2128
rect 17027 752 17036 2128
rect 17182 752 17191 2128
rect 17191 752 17225 2128
rect 17225 752 17234 2128
rect 17380 752 17389 2128
rect 17389 752 17423 2128
rect 17423 752 17432 2128
rect 17578 752 17587 2128
rect 17587 752 17621 2128
rect 17621 752 17630 2128
rect 17776 752 17785 2128
rect 17785 752 17819 2128
rect 17819 752 17828 2128
rect 17974 752 17983 2128
rect 17983 752 18017 2128
rect 18017 752 18026 2128
rect 18172 752 18181 2128
rect 18181 752 18215 2128
rect 18215 752 18224 2128
rect 18370 752 18379 2128
rect 18379 752 18413 2128
rect 18413 752 18422 2128
rect 18568 752 18577 2128
rect 18577 752 18611 2128
rect 18611 752 18620 2128
rect 18766 752 18775 2128
rect 18775 752 18809 2128
rect 18809 752 18818 2128
rect 18964 752 18973 2128
rect 18973 752 19007 2128
rect 19007 752 19016 2128
rect 19162 752 19171 2128
rect 19171 752 19205 2128
rect 19205 752 19214 2128
rect 19360 752 19369 2128
rect 19369 752 19403 2128
rect 19403 752 19412 2128
rect 19558 752 19567 2128
rect 19567 752 19601 2128
rect 19601 752 19610 2128
rect 19756 2128 19808 2129
rect 19756 753 19765 2128
rect 19765 753 19799 2128
rect 19799 753 19808 2128
rect 11212 -877 11346 -743
rect 11440 -884 11449 492
rect 11449 -884 11483 492
rect 11483 -884 11492 492
rect 11638 -884 11647 492
rect 11647 -884 11681 492
rect 11681 -884 11690 492
rect 11836 -884 11845 492
rect 11845 -884 11879 492
rect 11879 -884 11888 492
rect 12034 -884 12043 492
rect 12043 -884 12077 492
rect 12077 -884 12086 492
rect 12232 -884 12241 492
rect 12241 -884 12275 492
rect 12275 -884 12284 492
rect 12430 -884 12439 492
rect 12439 -884 12473 492
rect 12473 -884 12482 492
rect 12628 -884 12637 492
rect 12637 -884 12671 492
rect 12671 -884 12680 492
rect 12826 -884 12835 492
rect 12835 -884 12869 492
rect 12869 -884 12878 492
rect 13024 -884 13033 492
rect 13033 -884 13067 492
rect 13067 -884 13076 492
rect 13222 -884 13231 492
rect 13231 -884 13265 492
rect 13265 -884 13274 492
rect 13420 -884 13429 492
rect 13429 -884 13463 492
rect 13463 -884 13472 492
rect 13618 -884 13627 492
rect 13627 -884 13661 492
rect 13661 -884 13670 492
rect 13816 -884 13825 492
rect 13825 -884 13859 492
rect 13859 -884 13868 492
rect 14014 -884 14023 492
rect 14023 -884 14057 492
rect 14057 -884 14066 492
rect 14212 -884 14221 492
rect 14221 -884 14255 492
rect 14255 -884 14264 492
rect 14410 -884 14419 492
rect 14419 -884 14453 492
rect 14453 -884 14462 492
rect 14608 -884 14617 492
rect 14617 -884 14651 492
rect 14651 -884 14660 492
rect 14806 -884 14815 492
rect 14815 -884 14849 492
rect 14849 -884 14858 492
rect 15004 -884 15013 492
rect 15013 -884 15047 492
rect 15047 -884 15056 492
rect 15202 -884 15211 492
rect 15211 -884 15245 492
rect 15245 -884 15254 492
rect 15400 -884 15409 492
rect 15409 -884 15443 492
rect 15443 -884 15452 492
rect 15598 -884 15607 492
rect 15607 -884 15641 492
rect 15641 -884 15650 492
rect 15796 -884 15805 492
rect 15805 -884 15839 492
rect 15839 -884 15848 492
rect 15994 -884 16003 492
rect 16003 -884 16037 492
rect 16037 -884 16046 492
rect 16192 -884 16201 492
rect 16201 -884 16235 492
rect 16235 -884 16244 492
rect 16390 -884 16399 492
rect 16399 -884 16433 492
rect 16433 -884 16442 492
rect 16588 -884 16597 492
rect 16597 -884 16631 492
rect 16631 -884 16640 492
rect 16786 -884 16795 492
rect 16795 -884 16829 492
rect 16829 -884 16838 492
rect 16984 -884 16993 492
rect 16993 -884 17027 492
rect 17027 -884 17036 492
rect 17182 -884 17191 492
rect 17191 -884 17225 492
rect 17225 -884 17234 492
rect 17380 -884 17389 492
rect 17389 -884 17423 492
rect 17423 -884 17432 492
rect 17578 -884 17587 492
rect 17587 -884 17621 492
rect 17621 -884 17630 492
rect 17776 -884 17785 492
rect 17785 -884 17819 492
rect 17819 -884 17828 492
rect 17974 -884 17983 492
rect 17983 -884 18017 492
rect 18017 -884 18026 492
rect 18172 -884 18181 492
rect 18181 -884 18215 492
rect 18215 -884 18224 492
rect 18370 -884 18379 492
rect 18379 -884 18413 492
rect 18413 -884 18422 492
rect 18568 -884 18577 492
rect 18577 -884 18611 492
rect 18611 -884 18620 492
rect 18766 -884 18775 492
rect 18775 -884 18809 492
rect 18809 -884 18818 492
rect 18964 -884 18973 492
rect 18973 -884 19007 492
rect 19007 -884 19016 492
rect 19162 -884 19171 492
rect 19171 -884 19205 492
rect 19205 -884 19214 492
rect 19360 -884 19369 492
rect 19369 -884 19403 492
rect 19403 -884 19412 492
rect 19558 -884 19567 492
rect 19567 -884 19601 492
rect 19601 -884 19610 492
rect 19756 492 19808 493
rect 19756 -883 19765 492
rect 19765 -883 19799 492
rect 19799 -883 19808 492
rect 19902 -877 20036 -743
rect 11212 -1081 11346 -947
rect 19902 -1081 20036 -947
rect 11212 -1285 11346 -1151
rect 11440 -2520 11449 -1144
rect 11449 -2520 11483 -1144
rect 11483 -2520 11492 -1144
rect 11638 -2520 11647 -1144
rect 11647 -2520 11681 -1144
rect 11681 -2520 11690 -1144
rect 11836 -2520 11845 -1144
rect 11845 -2520 11879 -1144
rect 11879 -2520 11888 -1144
rect 12034 -2520 12043 -1144
rect 12043 -2520 12077 -1144
rect 12077 -2520 12086 -1144
rect 12232 -2520 12241 -1144
rect 12241 -2520 12275 -1144
rect 12275 -2520 12284 -1144
rect 12430 -2520 12439 -1144
rect 12439 -2520 12473 -1144
rect 12473 -2520 12482 -1144
rect 12628 -2520 12637 -1144
rect 12637 -2520 12671 -1144
rect 12671 -2520 12680 -1144
rect 12826 -2520 12835 -1144
rect 12835 -2520 12869 -1144
rect 12869 -2520 12878 -1144
rect 13024 -2520 13033 -1144
rect 13033 -2520 13067 -1144
rect 13067 -2520 13076 -1144
rect 13222 -2520 13231 -1144
rect 13231 -2520 13265 -1144
rect 13265 -2520 13274 -1144
rect 13420 -2520 13429 -1144
rect 13429 -2520 13463 -1144
rect 13463 -2520 13472 -1144
rect 13618 -2520 13627 -1144
rect 13627 -2520 13661 -1144
rect 13661 -2520 13670 -1144
rect 13816 -2520 13825 -1144
rect 13825 -2520 13859 -1144
rect 13859 -2520 13868 -1144
rect 14014 -2520 14023 -1144
rect 14023 -2520 14057 -1144
rect 14057 -2520 14066 -1144
rect 14212 -2520 14221 -1144
rect 14221 -2520 14255 -1144
rect 14255 -2520 14264 -1144
rect 14410 -2520 14419 -1144
rect 14419 -2520 14453 -1144
rect 14453 -2520 14462 -1144
rect 14608 -2520 14617 -1144
rect 14617 -2520 14651 -1144
rect 14651 -2520 14660 -1144
rect 14806 -2520 14815 -1144
rect 14815 -2520 14849 -1144
rect 14849 -2520 14858 -1144
rect 15004 -2520 15013 -1144
rect 15013 -2520 15047 -1144
rect 15047 -2520 15056 -1144
rect 15202 -2520 15211 -1144
rect 15211 -2520 15245 -1144
rect 15245 -2520 15254 -1144
rect 15400 -2520 15409 -1144
rect 15409 -2520 15443 -1144
rect 15443 -2520 15452 -1144
rect 15598 -2520 15607 -1144
rect 15607 -2520 15641 -1144
rect 15641 -2520 15650 -1144
rect 15796 -2520 15805 -1144
rect 15805 -2520 15839 -1144
rect 15839 -2520 15848 -1144
rect 15994 -2520 16003 -1144
rect 16003 -2520 16037 -1144
rect 16037 -2520 16046 -1144
rect 16192 -2520 16201 -1144
rect 16201 -2520 16235 -1144
rect 16235 -2520 16244 -1144
rect 16390 -2520 16399 -1144
rect 16399 -2520 16433 -1144
rect 16433 -2520 16442 -1144
rect 16588 -2520 16597 -1144
rect 16597 -2520 16631 -1144
rect 16631 -2520 16640 -1144
rect 16786 -2520 16795 -1144
rect 16795 -2520 16829 -1144
rect 16829 -2520 16838 -1144
rect 16984 -2520 16993 -1144
rect 16993 -2520 17027 -1144
rect 17027 -2520 17036 -1144
rect 17182 -2520 17191 -1144
rect 17191 -2520 17225 -1144
rect 17225 -2520 17234 -1144
rect 17380 -2520 17389 -1144
rect 17389 -2520 17423 -1144
rect 17423 -2520 17432 -1144
rect 17578 -2520 17587 -1144
rect 17587 -2520 17621 -1144
rect 17621 -2520 17630 -1144
rect 17776 -2520 17785 -1144
rect 17785 -2520 17819 -1144
rect 17819 -2520 17828 -1144
rect 17974 -2520 17983 -1144
rect 17983 -2520 18017 -1144
rect 18017 -2520 18026 -1144
rect 18172 -2520 18181 -1144
rect 18181 -2520 18215 -1144
rect 18215 -2520 18224 -1144
rect 18370 -2520 18379 -1144
rect 18379 -2520 18413 -1144
rect 18413 -2520 18422 -1144
rect 18568 -2520 18577 -1144
rect 18577 -2520 18611 -1144
rect 18611 -2520 18620 -1144
rect 18766 -2520 18775 -1144
rect 18775 -2520 18809 -1144
rect 18809 -2520 18818 -1144
rect 18964 -2520 18973 -1144
rect 18973 -2520 19007 -1144
rect 19007 -2520 19016 -1144
rect 19162 -2520 19171 -1144
rect 19171 -2520 19205 -1144
rect 19205 -2520 19214 -1144
rect 19360 -2520 19369 -1144
rect 19369 -2520 19403 -1144
rect 19403 -2520 19412 -1144
rect 19558 -2520 19567 -1144
rect 19567 -2520 19601 -1144
rect 19601 -2520 19610 -1144
rect 19756 -1144 19808 -1143
rect 19756 -2519 19765 -1144
rect 19765 -2519 19799 -1144
rect 19799 -2519 19808 -1144
rect 19902 -1285 20036 -1151
rect 11440 -4156 11449 -2780
rect 11449 -4156 11483 -2780
rect 11483 -4156 11492 -2780
rect 11638 -4156 11647 -2780
rect 11647 -4156 11681 -2780
rect 11681 -4156 11690 -2780
rect 11836 -4156 11845 -2780
rect 11845 -4156 11879 -2780
rect 11879 -4156 11888 -2780
rect 12034 -4156 12043 -2780
rect 12043 -4156 12077 -2780
rect 12077 -4156 12086 -2780
rect 12232 -4156 12241 -2780
rect 12241 -4156 12275 -2780
rect 12275 -4156 12284 -2780
rect 12430 -4156 12439 -2780
rect 12439 -4156 12473 -2780
rect 12473 -4156 12482 -2780
rect 12628 -4156 12637 -2780
rect 12637 -4156 12671 -2780
rect 12671 -4156 12680 -2780
rect 12826 -4156 12835 -2780
rect 12835 -4156 12869 -2780
rect 12869 -4156 12878 -2780
rect 13024 -4156 13033 -2780
rect 13033 -4156 13067 -2780
rect 13067 -4156 13076 -2780
rect 13222 -4156 13231 -2780
rect 13231 -4156 13265 -2780
rect 13265 -4156 13274 -2780
rect 13420 -4156 13429 -2780
rect 13429 -4156 13463 -2780
rect 13463 -4156 13472 -2780
rect 13618 -4156 13627 -2780
rect 13627 -4156 13661 -2780
rect 13661 -4156 13670 -2780
rect 13816 -4156 13825 -2780
rect 13825 -4156 13859 -2780
rect 13859 -4156 13868 -2780
rect 14014 -4156 14023 -2780
rect 14023 -4156 14057 -2780
rect 14057 -4156 14066 -2780
rect 14212 -4156 14221 -2780
rect 14221 -4156 14255 -2780
rect 14255 -4156 14264 -2780
rect 14410 -4156 14419 -2780
rect 14419 -4156 14453 -2780
rect 14453 -4156 14462 -2780
rect 14608 -4156 14617 -2780
rect 14617 -4156 14651 -2780
rect 14651 -4156 14660 -2780
rect 14806 -4156 14815 -2780
rect 14815 -4156 14849 -2780
rect 14849 -4156 14858 -2780
rect 15004 -4156 15013 -2780
rect 15013 -4156 15047 -2780
rect 15047 -4156 15056 -2780
rect 15202 -4156 15211 -2780
rect 15211 -4156 15245 -2780
rect 15245 -4156 15254 -2780
rect 15400 -4156 15409 -2780
rect 15409 -4156 15443 -2780
rect 15443 -4156 15452 -2780
rect 15598 -4156 15607 -2780
rect 15607 -4156 15641 -2780
rect 15641 -4156 15650 -2780
rect 15796 -4156 15805 -2780
rect 15805 -4156 15839 -2780
rect 15839 -4156 15848 -2780
rect 15994 -4156 16003 -2780
rect 16003 -4156 16037 -2780
rect 16037 -4156 16046 -2780
rect 16192 -4156 16201 -2780
rect 16201 -4156 16235 -2780
rect 16235 -4156 16244 -2780
rect 16390 -4156 16399 -2780
rect 16399 -4156 16433 -2780
rect 16433 -4156 16442 -2780
rect 16588 -4156 16597 -2780
rect 16597 -4156 16631 -2780
rect 16631 -4156 16640 -2780
rect 16786 -4156 16795 -2780
rect 16795 -4156 16829 -2780
rect 16829 -4156 16838 -2780
rect 16984 -4156 16993 -2780
rect 16993 -4156 17027 -2780
rect 17027 -4156 17036 -2780
rect 17182 -4156 17191 -2780
rect 17191 -4156 17225 -2780
rect 17225 -4156 17234 -2780
rect 17380 -4156 17389 -2780
rect 17389 -4156 17423 -2780
rect 17423 -4156 17432 -2780
rect 17578 -4156 17587 -2780
rect 17587 -4156 17621 -2780
rect 17621 -4156 17630 -2780
rect 17776 -4156 17785 -2780
rect 17785 -4156 17819 -2780
rect 17819 -4156 17828 -2780
rect 17974 -4156 17983 -2780
rect 17983 -4156 18017 -2780
rect 18017 -4156 18026 -2780
rect 18172 -4156 18181 -2780
rect 18181 -4156 18215 -2780
rect 18215 -4156 18224 -2780
rect 18370 -4156 18379 -2780
rect 18379 -4156 18413 -2780
rect 18413 -4156 18422 -2780
rect 18568 -4156 18577 -2780
rect 18577 -4156 18611 -2780
rect 18611 -4156 18620 -2780
rect 18766 -4156 18775 -2780
rect 18775 -4156 18809 -2780
rect 18809 -4156 18818 -2780
rect 18964 -4156 18973 -2780
rect 18973 -4156 19007 -2780
rect 19007 -4156 19016 -2780
rect 19162 -4156 19171 -2780
rect 19171 -4156 19205 -2780
rect 19205 -4156 19214 -2780
rect 19360 -4156 19369 -2780
rect 19369 -4156 19403 -2780
rect 19403 -4156 19412 -2780
rect 19558 -4156 19567 -2780
rect 19567 -4156 19601 -2780
rect 19601 -4156 19610 -2780
rect 19756 -2780 19808 -2779
rect 19756 -4155 19765 -2780
rect 19765 -4155 19799 -2780
rect 19799 -4155 19808 -2780
rect 23290 752 23299 2128
rect 23299 752 23333 2128
rect 23333 752 23342 2128
rect 23488 752 23497 2128
rect 23497 752 23531 2128
rect 23531 752 23540 2128
rect 23686 752 23695 2128
rect 23695 752 23729 2128
rect 23729 752 23738 2128
rect 23884 752 23893 2128
rect 23893 752 23927 2128
rect 23927 752 23936 2128
rect 24082 752 24091 2128
rect 24091 752 24125 2128
rect 24125 752 24134 2128
rect 24280 752 24289 2128
rect 24289 752 24323 2128
rect 24323 752 24332 2128
rect 24478 752 24487 2128
rect 24487 752 24521 2128
rect 24521 752 24530 2128
rect 24676 752 24685 2128
rect 24685 752 24719 2128
rect 24719 752 24728 2128
rect 24874 752 24883 2128
rect 24883 752 24917 2128
rect 24917 752 24926 2128
rect 25072 752 25081 2128
rect 25081 752 25115 2128
rect 25115 752 25124 2128
rect 25270 752 25279 2128
rect 25279 752 25313 2128
rect 25313 752 25322 2128
rect 25468 752 25477 2128
rect 25477 752 25511 2128
rect 25511 752 25520 2128
rect 25666 752 25675 2128
rect 25675 752 25709 2128
rect 25709 752 25718 2128
rect 25864 752 25873 2128
rect 25873 752 25907 2128
rect 25907 752 25916 2128
rect 26062 752 26071 2128
rect 26071 752 26105 2128
rect 26105 752 26114 2128
rect 26260 752 26269 2128
rect 26269 752 26303 2128
rect 26303 752 26312 2128
rect 26458 752 26467 2128
rect 26467 752 26501 2128
rect 26501 752 26510 2128
rect 26656 752 26665 2128
rect 26665 752 26699 2128
rect 26699 752 26708 2128
rect 26854 752 26863 2128
rect 26863 752 26897 2128
rect 26897 752 26906 2128
rect 27052 752 27061 2128
rect 27061 752 27095 2128
rect 27095 752 27104 2128
rect 27250 752 27259 2128
rect 27259 752 27293 2128
rect 27293 752 27302 2128
rect 27448 752 27457 2128
rect 27457 752 27491 2128
rect 27491 752 27500 2128
rect 27646 752 27655 2128
rect 27655 752 27689 2128
rect 27689 752 27698 2128
rect 27844 752 27853 2128
rect 27853 752 27887 2128
rect 27887 752 27896 2128
rect 28042 752 28051 2128
rect 28051 752 28085 2128
rect 28085 752 28094 2128
rect 28240 752 28249 2128
rect 28249 752 28283 2128
rect 28283 752 28292 2128
rect 28438 752 28447 2128
rect 28447 752 28481 2128
rect 28481 752 28490 2128
rect 28636 752 28645 2128
rect 28645 752 28679 2128
rect 28679 752 28688 2128
rect 28834 752 28843 2128
rect 28843 752 28877 2128
rect 28877 752 28886 2128
rect 29032 752 29041 2128
rect 29041 752 29075 2128
rect 29075 752 29084 2128
rect 29230 752 29239 2128
rect 29239 752 29273 2128
rect 29273 752 29282 2128
rect 29428 752 29437 2128
rect 29437 752 29471 2128
rect 29471 752 29480 2128
rect 29626 752 29635 2128
rect 29635 752 29669 2128
rect 29669 752 29678 2128
rect 29824 752 29833 2128
rect 29833 752 29867 2128
rect 29867 752 29876 2128
rect 30022 752 30031 2128
rect 30031 752 30065 2128
rect 30065 752 30074 2128
rect 30220 752 30229 2128
rect 30229 752 30263 2128
rect 30263 752 30272 2128
rect 30418 752 30427 2128
rect 30427 752 30461 2128
rect 30461 752 30470 2128
rect 30616 752 30625 2128
rect 30625 752 30659 2128
rect 30659 752 30668 2128
rect 30814 752 30823 2128
rect 30823 752 30857 2128
rect 30857 752 30866 2128
rect 31012 752 31021 2128
rect 31021 752 31055 2128
rect 31055 752 31064 2128
rect 31210 752 31219 2128
rect 31219 752 31253 2128
rect 31253 752 31262 2128
rect 31408 752 31417 2128
rect 31417 752 31451 2128
rect 31451 752 31460 2128
rect 31606 2128 31658 2129
rect 31606 753 31615 2128
rect 31615 753 31649 2128
rect 31649 753 31658 2128
rect 23062 -877 23196 -743
rect 23290 -884 23299 492
rect 23299 -884 23333 492
rect 23333 -884 23342 492
rect 23488 -884 23497 492
rect 23497 -884 23531 492
rect 23531 -884 23540 492
rect 23686 -884 23695 492
rect 23695 -884 23729 492
rect 23729 -884 23738 492
rect 23884 -884 23893 492
rect 23893 -884 23927 492
rect 23927 -884 23936 492
rect 24082 -884 24091 492
rect 24091 -884 24125 492
rect 24125 -884 24134 492
rect 24280 -884 24289 492
rect 24289 -884 24323 492
rect 24323 -884 24332 492
rect 24478 -884 24487 492
rect 24487 -884 24521 492
rect 24521 -884 24530 492
rect 24676 -884 24685 492
rect 24685 -884 24719 492
rect 24719 -884 24728 492
rect 24874 -884 24883 492
rect 24883 -884 24917 492
rect 24917 -884 24926 492
rect 25072 -884 25081 492
rect 25081 -884 25115 492
rect 25115 -884 25124 492
rect 25270 -884 25279 492
rect 25279 -884 25313 492
rect 25313 -884 25322 492
rect 25468 -884 25477 492
rect 25477 -884 25511 492
rect 25511 -884 25520 492
rect 25666 -884 25675 492
rect 25675 -884 25709 492
rect 25709 -884 25718 492
rect 25864 -884 25873 492
rect 25873 -884 25907 492
rect 25907 -884 25916 492
rect 26062 -884 26071 492
rect 26071 -884 26105 492
rect 26105 -884 26114 492
rect 26260 -884 26269 492
rect 26269 -884 26303 492
rect 26303 -884 26312 492
rect 26458 -884 26467 492
rect 26467 -884 26501 492
rect 26501 -884 26510 492
rect 26656 -884 26665 492
rect 26665 -884 26699 492
rect 26699 -884 26708 492
rect 26854 -884 26863 492
rect 26863 -884 26897 492
rect 26897 -884 26906 492
rect 27052 -884 27061 492
rect 27061 -884 27095 492
rect 27095 -884 27104 492
rect 27250 -884 27259 492
rect 27259 -884 27293 492
rect 27293 -884 27302 492
rect 27448 -884 27457 492
rect 27457 -884 27491 492
rect 27491 -884 27500 492
rect 27646 -884 27655 492
rect 27655 -884 27689 492
rect 27689 -884 27698 492
rect 27844 -884 27853 492
rect 27853 -884 27887 492
rect 27887 -884 27896 492
rect 28042 -884 28051 492
rect 28051 -884 28085 492
rect 28085 -884 28094 492
rect 28240 -884 28249 492
rect 28249 -884 28283 492
rect 28283 -884 28292 492
rect 28438 -884 28447 492
rect 28447 -884 28481 492
rect 28481 -884 28490 492
rect 28636 -884 28645 492
rect 28645 -884 28679 492
rect 28679 -884 28688 492
rect 28834 -884 28843 492
rect 28843 -884 28877 492
rect 28877 -884 28886 492
rect 29032 -884 29041 492
rect 29041 -884 29075 492
rect 29075 -884 29084 492
rect 29230 -884 29239 492
rect 29239 -884 29273 492
rect 29273 -884 29282 492
rect 29428 -884 29437 492
rect 29437 -884 29471 492
rect 29471 -884 29480 492
rect 29626 -884 29635 492
rect 29635 -884 29669 492
rect 29669 -884 29678 492
rect 29824 -884 29833 492
rect 29833 -884 29867 492
rect 29867 -884 29876 492
rect 30022 -884 30031 492
rect 30031 -884 30065 492
rect 30065 -884 30074 492
rect 30220 -884 30229 492
rect 30229 -884 30263 492
rect 30263 -884 30272 492
rect 30418 -884 30427 492
rect 30427 -884 30461 492
rect 30461 -884 30470 492
rect 30616 -884 30625 492
rect 30625 -884 30659 492
rect 30659 -884 30668 492
rect 30814 -884 30823 492
rect 30823 -884 30857 492
rect 30857 -884 30866 492
rect 31012 -884 31021 492
rect 31021 -884 31055 492
rect 31055 -884 31064 492
rect 31210 -884 31219 492
rect 31219 -884 31253 492
rect 31253 -884 31262 492
rect 31408 -884 31417 492
rect 31417 -884 31451 492
rect 31451 -884 31460 492
rect 31606 492 31658 493
rect 31606 -883 31615 492
rect 31615 -883 31649 492
rect 31649 -883 31658 492
rect 23062 -1081 23196 -947
rect 23062 -1285 23196 -1151
rect 23290 -2520 23299 -1144
rect 23299 -2520 23333 -1144
rect 23333 -2520 23342 -1144
rect 23488 -2520 23497 -1144
rect 23497 -2520 23531 -1144
rect 23531 -2520 23540 -1144
rect 23686 -2520 23695 -1144
rect 23695 -2520 23729 -1144
rect 23729 -2520 23738 -1144
rect 23884 -2520 23893 -1144
rect 23893 -2520 23927 -1144
rect 23927 -2520 23936 -1144
rect 24082 -2520 24091 -1144
rect 24091 -2520 24125 -1144
rect 24125 -2520 24134 -1144
rect 24280 -2520 24289 -1144
rect 24289 -2520 24323 -1144
rect 24323 -2520 24332 -1144
rect 24478 -2520 24487 -1144
rect 24487 -2520 24521 -1144
rect 24521 -2520 24530 -1144
rect 24676 -2520 24685 -1144
rect 24685 -2520 24719 -1144
rect 24719 -2520 24728 -1144
rect 24874 -2520 24883 -1144
rect 24883 -2520 24917 -1144
rect 24917 -2520 24926 -1144
rect 25072 -2520 25081 -1144
rect 25081 -2520 25115 -1144
rect 25115 -2520 25124 -1144
rect 25270 -2520 25279 -1144
rect 25279 -2520 25313 -1144
rect 25313 -2520 25322 -1144
rect 25468 -2520 25477 -1144
rect 25477 -2520 25511 -1144
rect 25511 -2520 25520 -1144
rect 25666 -2520 25675 -1144
rect 25675 -2520 25709 -1144
rect 25709 -2520 25718 -1144
rect 25864 -2520 25873 -1144
rect 25873 -2520 25907 -1144
rect 25907 -2520 25916 -1144
rect 26062 -2520 26071 -1144
rect 26071 -2520 26105 -1144
rect 26105 -2520 26114 -1144
rect 26260 -2520 26269 -1144
rect 26269 -2520 26303 -1144
rect 26303 -2520 26312 -1144
rect 26458 -2520 26467 -1144
rect 26467 -2520 26501 -1144
rect 26501 -2520 26510 -1144
rect 26656 -2520 26665 -1144
rect 26665 -2520 26699 -1144
rect 26699 -2520 26708 -1144
rect 26854 -2520 26863 -1144
rect 26863 -2520 26897 -1144
rect 26897 -2520 26906 -1144
rect 27052 -2520 27061 -1144
rect 27061 -2520 27095 -1144
rect 27095 -2520 27104 -1144
rect 27250 -2520 27259 -1144
rect 27259 -2520 27293 -1144
rect 27293 -2520 27302 -1144
rect 27448 -2520 27457 -1144
rect 27457 -2520 27491 -1144
rect 27491 -2520 27500 -1144
rect 27646 -2520 27655 -1144
rect 27655 -2520 27689 -1144
rect 27689 -2520 27698 -1144
rect 27844 -2520 27853 -1144
rect 27853 -2520 27887 -1144
rect 27887 -2520 27896 -1144
rect 28042 -2520 28051 -1144
rect 28051 -2520 28085 -1144
rect 28085 -2520 28094 -1144
rect 28240 -2520 28249 -1144
rect 28249 -2520 28283 -1144
rect 28283 -2520 28292 -1144
rect 28438 -2520 28447 -1144
rect 28447 -2520 28481 -1144
rect 28481 -2520 28490 -1144
rect 28636 -2520 28645 -1144
rect 28645 -2520 28679 -1144
rect 28679 -2520 28688 -1144
rect 28834 -2520 28843 -1144
rect 28843 -2520 28877 -1144
rect 28877 -2520 28886 -1144
rect 29032 -2520 29041 -1144
rect 29041 -2520 29075 -1144
rect 29075 -2520 29084 -1144
rect 29230 -2520 29239 -1144
rect 29239 -2520 29273 -1144
rect 29273 -2520 29282 -1144
rect 29428 -2520 29437 -1144
rect 29437 -2520 29471 -1144
rect 29471 -2520 29480 -1144
rect 29626 -2520 29635 -1144
rect 29635 -2520 29669 -1144
rect 29669 -2520 29678 -1144
rect 29824 -2520 29833 -1144
rect 29833 -2520 29867 -1144
rect 29867 -2520 29876 -1144
rect 30022 -2520 30031 -1144
rect 30031 -2520 30065 -1144
rect 30065 -2520 30074 -1144
rect 30220 -2520 30229 -1144
rect 30229 -2520 30263 -1144
rect 30263 -2520 30272 -1144
rect 30418 -2520 30427 -1144
rect 30427 -2520 30461 -1144
rect 30461 -2520 30470 -1144
rect 30616 -2520 30625 -1144
rect 30625 -2520 30659 -1144
rect 30659 -2520 30668 -1144
rect 30814 -2520 30823 -1144
rect 30823 -2520 30857 -1144
rect 30857 -2520 30866 -1144
rect 31012 -2520 31021 -1144
rect 31021 -2520 31055 -1144
rect 31055 -2520 31064 -1144
rect 31210 -2520 31219 -1144
rect 31219 -2520 31253 -1144
rect 31253 -2520 31262 -1144
rect 31408 -2520 31417 -1144
rect 31417 -2520 31451 -1144
rect 31451 -2520 31460 -1144
rect 31606 -1144 31658 -1143
rect 31606 -2519 31615 -1144
rect 31615 -2519 31649 -1144
rect 31649 -2519 31658 -1144
rect 23290 -4156 23299 -2780
rect 23299 -4156 23333 -2780
rect 23333 -4156 23342 -2780
rect 23488 -4156 23497 -2780
rect 23497 -4156 23531 -2780
rect 23531 -4156 23540 -2780
rect 23686 -4156 23695 -2780
rect 23695 -4156 23729 -2780
rect 23729 -4156 23738 -2780
rect 23884 -4156 23893 -2780
rect 23893 -4156 23927 -2780
rect 23927 -4156 23936 -2780
rect 24082 -4156 24091 -2780
rect 24091 -4156 24125 -2780
rect 24125 -4156 24134 -2780
rect 24280 -4156 24289 -2780
rect 24289 -4156 24323 -2780
rect 24323 -4156 24332 -2780
rect 24478 -4156 24487 -2780
rect 24487 -4156 24521 -2780
rect 24521 -4156 24530 -2780
rect 24676 -4156 24685 -2780
rect 24685 -4156 24719 -2780
rect 24719 -4156 24728 -2780
rect 24874 -4156 24883 -2780
rect 24883 -4156 24917 -2780
rect 24917 -4156 24926 -2780
rect 25072 -4156 25081 -2780
rect 25081 -4156 25115 -2780
rect 25115 -4156 25124 -2780
rect 25270 -4156 25279 -2780
rect 25279 -4156 25313 -2780
rect 25313 -4156 25322 -2780
rect 25468 -4156 25477 -2780
rect 25477 -4156 25511 -2780
rect 25511 -4156 25520 -2780
rect 25666 -4156 25675 -2780
rect 25675 -4156 25709 -2780
rect 25709 -4156 25718 -2780
rect 25864 -4156 25873 -2780
rect 25873 -4156 25907 -2780
rect 25907 -4156 25916 -2780
rect 26062 -4156 26071 -2780
rect 26071 -4156 26105 -2780
rect 26105 -4156 26114 -2780
rect 26260 -4156 26269 -2780
rect 26269 -4156 26303 -2780
rect 26303 -4156 26312 -2780
rect 26458 -4156 26467 -2780
rect 26467 -4156 26501 -2780
rect 26501 -4156 26510 -2780
rect 26656 -4156 26665 -2780
rect 26665 -4156 26699 -2780
rect 26699 -4156 26708 -2780
rect 26854 -4156 26863 -2780
rect 26863 -4156 26897 -2780
rect 26897 -4156 26906 -2780
rect 27052 -4156 27061 -2780
rect 27061 -4156 27095 -2780
rect 27095 -4156 27104 -2780
rect 27250 -4156 27259 -2780
rect 27259 -4156 27293 -2780
rect 27293 -4156 27302 -2780
rect 27448 -4156 27457 -2780
rect 27457 -4156 27491 -2780
rect 27491 -4156 27500 -2780
rect 27646 -4156 27655 -2780
rect 27655 -4156 27689 -2780
rect 27689 -4156 27698 -2780
rect 27844 -4156 27853 -2780
rect 27853 -4156 27887 -2780
rect 27887 -4156 27896 -2780
rect 28042 -4156 28051 -2780
rect 28051 -4156 28085 -2780
rect 28085 -4156 28094 -2780
rect 28240 -4156 28249 -2780
rect 28249 -4156 28283 -2780
rect 28283 -4156 28292 -2780
rect 28438 -4156 28447 -2780
rect 28447 -4156 28481 -2780
rect 28481 -4156 28490 -2780
rect 28636 -4156 28645 -2780
rect 28645 -4156 28679 -2780
rect 28679 -4156 28688 -2780
rect 28834 -4156 28843 -2780
rect 28843 -4156 28877 -2780
rect 28877 -4156 28886 -2780
rect 29032 -4156 29041 -2780
rect 29041 -4156 29075 -2780
rect 29075 -4156 29084 -2780
rect 29230 -4156 29239 -2780
rect 29239 -4156 29273 -2780
rect 29273 -4156 29282 -2780
rect 29428 -4156 29437 -2780
rect 29437 -4156 29471 -2780
rect 29471 -4156 29480 -2780
rect 29626 -4156 29635 -2780
rect 29635 -4156 29669 -2780
rect 29669 -4156 29678 -2780
rect 29824 -4156 29833 -2780
rect 29833 -4156 29867 -2780
rect 29867 -4156 29876 -2780
rect 30022 -4156 30031 -2780
rect 30031 -4156 30065 -2780
rect 30065 -4156 30074 -2780
rect 30220 -4156 30229 -2780
rect 30229 -4156 30263 -2780
rect 30263 -4156 30272 -2780
rect 30418 -4156 30427 -2780
rect 30427 -4156 30461 -2780
rect 30461 -4156 30470 -2780
rect 30616 -4156 30625 -2780
rect 30625 -4156 30659 -2780
rect 30659 -4156 30668 -2780
rect 30814 -4156 30823 -2780
rect 30823 -4156 30857 -2780
rect 30857 -4156 30866 -2780
rect 31012 -4156 31021 -2780
rect 31021 -4156 31055 -2780
rect 31055 -4156 31064 -2780
rect 31210 -4156 31219 -2780
rect 31219 -4156 31253 -2780
rect 31253 -4156 31262 -2780
rect 31408 -4156 31417 -2780
rect 31417 -4156 31451 -2780
rect 31451 -4156 31460 -2780
rect 31606 -2780 31658 -2779
rect 31606 -4155 31615 -2780
rect 31615 -4155 31649 -2780
rect 31649 -4155 31658 -2780
<< metal2 >>
rect -399 2128 -347 2134
rect -399 492 -347 752
rect -627 -743 -493 -733
rect -627 -887 -493 -877
rect -627 -947 -493 -937
rect -627 -1091 -493 -1081
rect -627 -1151 -493 -1141
rect -627 -1295 -493 -1285
rect -399 -1144 -347 -884
rect -399 -2780 -347 -2520
rect -399 -4166 -347 -4156
rect -201 2128 -149 2138
rect -201 492 -149 752
rect -201 -1144 -149 -884
rect -201 -2780 -149 -2520
rect -201 -4218 -149 -4156
rect -3 2128 49 2134
rect -3 492 49 752
rect -3 -1144 49 -884
rect -3 -2780 49 -2520
rect -3 -4166 49 -4156
rect 195 2128 247 2138
rect 195 492 247 752
rect 195 -1144 247 -884
rect 195 -2780 247 -2520
rect 195 -4218 247 -4156
rect 393 2128 445 2134
rect 393 492 445 752
rect 393 -1144 445 -884
rect 393 -2780 445 -2520
rect 393 -4166 445 -4156
rect 591 2128 643 2138
rect 591 492 643 752
rect 591 -1144 643 -884
rect 591 -2780 643 -2520
rect 591 -4218 643 -4156
rect 789 2128 841 2134
rect 789 492 841 752
rect 789 -1144 841 -884
rect 789 -2780 841 -2520
rect 789 -4166 841 -4156
rect 987 2128 1039 2138
rect 987 492 1039 752
rect 987 -1144 1039 -884
rect 987 -2780 1039 -2520
rect 987 -4218 1039 -4156
rect 1185 2128 1237 2134
rect 1185 492 1237 752
rect 1185 -1144 1237 -884
rect 1185 -2780 1237 -2520
rect 1185 -4166 1237 -4156
rect 1383 2128 1435 2138
rect 1383 492 1435 752
rect 1383 -1144 1435 -884
rect 1383 -2780 1435 -2520
rect 1383 -4218 1435 -4156
rect 1581 2128 1633 2134
rect 1581 492 1633 752
rect 1581 -1144 1633 -884
rect 1581 -2780 1633 -2520
rect 1581 -4166 1633 -4156
rect 1779 2128 1831 2138
rect 1779 492 1831 752
rect 1779 -1144 1831 -884
rect 1779 -2780 1831 -2520
rect 1779 -4218 1831 -4156
rect 1977 2128 2029 2134
rect 1977 492 2029 752
rect 1977 -1144 2029 -884
rect 1977 -2780 2029 -2520
rect 1977 -4166 2029 -4156
rect 2175 2128 2227 2138
rect 2175 492 2227 752
rect 2175 -1144 2227 -884
rect 2175 -2780 2227 -2520
rect 2175 -4218 2227 -4156
rect 2373 2128 2425 2134
rect 2373 492 2425 752
rect 2373 -1144 2425 -884
rect 2373 -2780 2425 -2520
rect 2373 -4166 2425 -4156
rect 2571 2128 2623 2138
rect 2571 492 2623 752
rect 2571 -1144 2623 -884
rect 2571 -2780 2623 -2520
rect 2571 -4218 2623 -4156
rect 2769 2128 2821 2134
rect 2769 492 2821 752
rect 2769 -1144 2821 -884
rect 2769 -2780 2821 -2520
rect 2769 -4166 2821 -4156
rect 2967 2128 3019 2138
rect 2967 492 3019 752
rect 2967 -1144 3019 -884
rect 2967 -2780 3019 -2520
rect 2967 -4218 3019 -4156
rect 3165 2128 3217 2134
rect 3165 492 3217 752
rect 3165 -1144 3217 -884
rect 3165 -2780 3217 -2520
rect 3165 -4166 3217 -4156
rect 3363 2128 3415 2138
rect 3363 492 3415 752
rect 3363 -1144 3415 -884
rect 3363 -2780 3415 -2520
rect 3363 -4218 3415 -4156
rect 3561 2128 3613 2134
rect 3561 492 3613 752
rect 3561 -1144 3613 -884
rect 3561 -2780 3613 -2520
rect 3561 -4166 3613 -4156
rect 3759 2128 3811 2138
rect 3759 492 3811 752
rect 3759 -1144 3811 -884
rect 3759 -2780 3811 -2520
rect 3759 -4218 3811 -4156
rect 3957 2128 4009 2134
rect 3957 492 4009 752
rect 3957 -1144 4009 -884
rect 3957 -2780 4009 -2520
rect 3957 -4166 4009 -4156
rect 4155 2128 4207 2138
rect 4155 492 4207 752
rect 4155 -1144 4207 -884
rect 4155 -2780 4207 -2520
rect 4155 -4218 4207 -4156
rect 4353 2128 4405 2134
rect 4353 492 4405 752
rect 4353 -1144 4405 -884
rect 4353 -2780 4405 -2520
rect 4353 -4166 4405 -4156
rect 4551 2128 4603 2138
rect 4551 492 4603 752
rect 4551 -1144 4603 -884
rect 4551 -2780 4603 -2520
rect 4551 -4218 4603 -4156
rect 4749 2128 4801 2134
rect 4749 492 4801 752
rect 4749 -1144 4801 -884
rect 4749 -2780 4801 -2520
rect 4749 -4166 4801 -4156
rect 4947 2128 4999 2138
rect 4947 492 4999 752
rect 4947 -1144 4999 -884
rect 4947 -2780 4999 -2520
rect 4947 -4218 4999 -4156
rect 5145 2128 5197 2134
rect 5145 492 5197 752
rect 5145 -1144 5197 -884
rect 5145 -2780 5197 -2520
rect 5145 -4166 5197 -4156
rect 5343 2128 5395 2138
rect 5343 492 5395 752
rect 5343 -1144 5395 -884
rect 5343 -2780 5395 -2520
rect 5343 -4218 5395 -4156
rect 5541 2128 5593 2134
rect 5541 492 5593 752
rect 5541 -1144 5593 -884
rect 5541 -2780 5593 -2520
rect 5541 -4166 5593 -4156
rect 5739 2128 5791 2138
rect 5739 492 5791 752
rect 5739 -1144 5791 -884
rect 5739 -2780 5791 -2520
rect 5739 -4218 5791 -4156
rect 5937 2128 5989 2134
rect 5937 492 5989 752
rect 5937 -1144 5989 -884
rect 5937 -2780 5989 -2520
rect 5937 -4166 5989 -4156
rect 6135 2128 6187 2138
rect 6135 492 6187 752
rect 6135 -1144 6187 -884
rect 6135 -2780 6187 -2520
rect 6135 -4218 6187 -4156
rect 6333 2128 6385 2134
rect 6333 492 6385 752
rect 6333 -1144 6385 -884
rect 6333 -2780 6385 -2520
rect 6333 -4166 6385 -4156
rect 6531 2128 6583 2138
rect 6531 492 6583 752
rect 6531 -1144 6583 -884
rect 6531 -2780 6583 -2520
rect 6531 -4218 6583 -4156
rect 6729 2128 6781 2134
rect 6729 492 6781 752
rect 6729 -1144 6781 -884
rect 6729 -2780 6781 -2520
rect 6729 -4166 6781 -4156
rect 6927 2128 6979 2138
rect 6927 492 6979 752
rect 6927 -1144 6979 -884
rect 6927 -2780 6979 -2520
rect 6927 -4218 6979 -4156
rect 7125 2128 7177 2134
rect 7125 492 7177 752
rect 7125 -1144 7177 -884
rect 7125 -2780 7177 -2520
rect 7125 -4166 7177 -4156
rect 7323 2128 7375 2138
rect 7323 492 7375 752
rect 7323 -1144 7375 -884
rect 7323 -2780 7375 -2520
rect 7323 -4218 7375 -4156
rect 7521 2128 7573 2134
rect 7521 492 7573 752
rect 7521 -1144 7573 -884
rect 7521 -2780 7573 -2520
rect 7521 -4166 7573 -4156
rect 7719 2128 7771 2138
rect 7719 492 7771 752
rect 7719 -1144 7771 -884
rect 7719 -2780 7771 -2520
rect 7719 -4218 7771 -4156
rect 7917 2129 7969 2135
rect 7917 493 7969 753
rect 11440 2128 11492 2134
rect 11440 492 11492 752
rect 7917 -1143 7969 -883
rect 8063 -743 8197 -733
rect 8063 -887 8197 -877
rect 11212 -743 11346 -733
rect 11212 -887 11346 -877
rect 8063 -947 8197 -937
rect 8063 -1091 8197 -1081
rect 11212 -947 11346 -937
rect 11212 -1091 11346 -1081
rect 8063 -1151 8197 -1141
rect 8063 -1295 8197 -1285
rect 11212 -1151 11346 -1141
rect 11212 -1295 11346 -1285
rect 11440 -1144 11492 -884
rect 7917 -2779 7969 -2519
rect 7917 -4165 7969 -4155
rect 11440 -2780 11492 -2520
rect 11440 -4166 11492 -4156
rect 11638 2128 11690 2138
rect 11638 492 11690 752
rect 11638 -1144 11690 -884
rect 11638 -2780 11690 -2520
rect 11638 -4218 11690 -4156
rect 11836 2128 11888 2134
rect 11836 492 11888 752
rect 11836 -1144 11888 -884
rect 11836 -2780 11888 -2520
rect 11836 -4166 11888 -4156
rect 12034 2128 12086 2138
rect 12034 492 12086 752
rect 12034 -1144 12086 -884
rect 12034 -2780 12086 -2520
rect 12034 -4218 12086 -4156
rect 12232 2128 12284 2134
rect 12232 492 12284 752
rect 12232 -1144 12284 -884
rect 12232 -2780 12284 -2520
rect 12232 -4166 12284 -4156
rect 12430 2128 12482 2138
rect 12430 492 12482 752
rect 12430 -1144 12482 -884
rect 12430 -2780 12482 -2520
rect 12430 -4218 12482 -4156
rect 12628 2128 12680 2134
rect 12628 492 12680 752
rect 12628 -1144 12680 -884
rect 12628 -2780 12680 -2520
rect 12628 -4166 12680 -4156
rect 12826 2128 12878 2138
rect 12826 492 12878 752
rect 12826 -1144 12878 -884
rect 12826 -2780 12878 -2520
rect 12826 -4218 12878 -4156
rect 13024 2128 13076 2134
rect 13024 492 13076 752
rect 13024 -1144 13076 -884
rect 13024 -2780 13076 -2520
rect 13024 -4166 13076 -4156
rect 13222 2128 13274 2138
rect 13222 492 13274 752
rect 13222 -1144 13274 -884
rect 13222 -2780 13274 -2520
rect 13222 -4218 13274 -4156
rect 13420 2128 13472 2134
rect 13420 492 13472 752
rect 13420 -1144 13472 -884
rect 13420 -2780 13472 -2520
rect 13420 -4166 13472 -4156
rect 13618 2128 13670 2138
rect 13618 492 13670 752
rect 13618 -1144 13670 -884
rect 13618 -2780 13670 -2520
rect 13618 -4218 13670 -4156
rect 13816 2128 13868 2134
rect 13816 492 13868 752
rect 13816 -1144 13868 -884
rect 13816 -2780 13868 -2520
rect 13816 -4166 13868 -4156
rect 14014 2128 14066 2138
rect 14014 492 14066 752
rect 14014 -1144 14066 -884
rect 14014 -2780 14066 -2520
rect 14014 -4218 14066 -4156
rect 14212 2128 14264 2134
rect 14212 492 14264 752
rect 14212 -1144 14264 -884
rect 14212 -2780 14264 -2520
rect 14212 -4166 14264 -4156
rect 14410 2128 14462 2138
rect 14410 492 14462 752
rect 14410 -1144 14462 -884
rect 14410 -2780 14462 -2520
rect 14410 -4218 14462 -4156
rect 14608 2128 14660 2134
rect 14608 492 14660 752
rect 14608 -1144 14660 -884
rect 14608 -2780 14660 -2520
rect 14608 -4166 14660 -4156
rect 14806 2128 14858 2138
rect 14806 492 14858 752
rect 14806 -1144 14858 -884
rect 14806 -2780 14858 -2520
rect 14806 -4218 14858 -4156
rect 15004 2128 15056 2134
rect 15004 492 15056 752
rect 15004 -1144 15056 -884
rect 15004 -2780 15056 -2520
rect 15004 -4166 15056 -4156
rect 15202 2128 15254 2138
rect 15202 492 15254 752
rect 15202 -1144 15254 -884
rect 15202 -2780 15254 -2520
rect 15202 -4218 15254 -4156
rect 15400 2128 15452 2134
rect 15400 492 15452 752
rect 15400 -1144 15452 -884
rect 15400 -2780 15452 -2520
rect 15400 -4166 15452 -4156
rect 15598 2128 15650 2138
rect 15598 492 15650 752
rect 15598 -1144 15650 -884
rect 15598 -2780 15650 -2520
rect 15598 -4218 15650 -4156
rect 15796 2128 15848 2134
rect 15796 492 15848 752
rect 15796 -1144 15848 -884
rect 15796 -2780 15848 -2520
rect 15796 -4166 15848 -4156
rect 15994 2128 16046 2138
rect 15994 492 16046 752
rect 15994 -1144 16046 -884
rect 15994 -2780 16046 -2520
rect 15994 -4218 16046 -4156
rect 16192 2128 16244 2134
rect 16192 492 16244 752
rect 16192 -1144 16244 -884
rect 16192 -2780 16244 -2520
rect 16192 -4166 16244 -4156
rect 16390 2128 16442 2138
rect 16390 492 16442 752
rect 16390 -1144 16442 -884
rect 16390 -2780 16442 -2520
rect 16390 -4218 16442 -4156
rect 16588 2128 16640 2134
rect 16588 492 16640 752
rect 16588 -1144 16640 -884
rect 16588 -2780 16640 -2520
rect 16588 -4166 16640 -4156
rect 16786 2128 16838 2138
rect 16786 492 16838 752
rect 16786 -1144 16838 -884
rect 16786 -2780 16838 -2520
rect 16786 -4218 16838 -4156
rect 16984 2128 17036 2134
rect 16984 492 17036 752
rect 16984 -1144 17036 -884
rect 16984 -2780 17036 -2520
rect 16984 -4166 17036 -4156
rect 17182 2128 17234 2138
rect 17182 492 17234 752
rect 17182 -1144 17234 -884
rect 17182 -2780 17234 -2520
rect 17182 -4218 17234 -4156
rect 17380 2128 17432 2134
rect 17380 492 17432 752
rect 17380 -1144 17432 -884
rect 17380 -2780 17432 -2520
rect 17380 -4166 17432 -4156
rect 17578 2128 17630 2138
rect 17578 492 17630 752
rect 17578 -1144 17630 -884
rect 17578 -2780 17630 -2520
rect 17578 -4218 17630 -4156
rect 17776 2128 17828 2134
rect 17776 492 17828 752
rect 17776 -1144 17828 -884
rect 17776 -2780 17828 -2520
rect 17776 -4166 17828 -4156
rect 17974 2128 18026 2138
rect 17974 492 18026 752
rect 17974 -1144 18026 -884
rect 17974 -2780 18026 -2520
rect 17974 -4218 18026 -4156
rect 18172 2128 18224 2134
rect 18172 492 18224 752
rect 18172 -1144 18224 -884
rect 18172 -2780 18224 -2520
rect 18172 -4166 18224 -4156
rect 18370 2128 18422 2138
rect 18370 492 18422 752
rect 18370 -1144 18422 -884
rect 18370 -2780 18422 -2520
rect 18370 -4218 18422 -4156
rect 18568 2128 18620 2134
rect 18568 492 18620 752
rect 18568 -1144 18620 -884
rect 18568 -2780 18620 -2520
rect 18568 -4166 18620 -4156
rect 18766 2128 18818 2138
rect 18766 492 18818 752
rect 18766 -1144 18818 -884
rect 18766 -2780 18818 -2520
rect 18766 -4218 18818 -4156
rect 18964 2128 19016 2134
rect 18964 492 19016 752
rect 18964 -1144 19016 -884
rect 18964 -2780 19016 -2520
rect 18964 -4166 19016 -4156
rect 19162 2128 19214 2138
rect 19162 492 19214 752
rect 19162 -1144 19214 -884
rect 19162 -2780 19214 -2520
rect 19162 -4218 19214 -4156
rect 19360 2128 19412 2134
rect 19360 492 19412 752
rect 19360 -1144 19412 -884
rect 19360 -2780 19412 -2520
rect 19360 -4166 19412 -4156
rect 19558 2128 19610 2138
rect 19558 492 19610 752
rect 19558 -1144 19610 -884
rect 19558 -2780 19610 -2520
rect 19558 -4218 19610 -4156
rect 19756 2129 19808 2135
rect 19756 493 19808 753
rect 23290 2128 23342 2134
rect 23290 492 23342 752
rect 19756 -1143 19808 -883
rect 19902 -743 20036 -733
rect 19902 -887 20036 -877
rect 23062 -743 23196 -733
rect 23062 -887 23196 -877
rect 19902 -947 20036 -937
rect 19902 -1091 20036 -1081
rect 23062 -947 23196 -937
rect 23062 -1091 23196 -1081
rect 19902 -1151 20036 -1141
rect 19902 -1295 20036 -1285
rect 23062 -1151 23196 -1141
rect 23062 -1295 23196 -1285
rect 23290 -1144 23342 -884
rect 19756 -2779 19808 -2519
rect 19756 -4165 19808 -4155
rect 23290 -2780 23342 -2520
rect 23290 -4166 23342 -4156
rect 23488 2128 23540 2138
rect 23488 492 23540 752
rect 23488 -1144 23540 -884
rect 23488 -2780 23540 -2520
rect 23488 -4218 23540 -4156
rect 23686 2128 23738 2134
rect 23686 492 23738 752
rect 23686 -1144 23738 -884
rect 23686 -2780 23738 -2520
rect 23686 -4166 23738 -4156
rect 23884 2128 23936 2138
rect 23884 492 23936 752
rect 23884 -1144 23936 -884
rect 23884 -2780 23936 -2520
rect 23884 -4218 23936 -4156
rect 24082 2128 24134 2134
rect 24082 492 24134 752
rect 24082 -1144 24134 -884
rect 24082 -2780 24134 -2520
rect 24082 -4166 24134 -4156
rect 24280 2128 24332 2138
rect 24280 492 24332 752
rect 24280 -1144 24332 -884
rect 24280 -2780 24332 -2520
rect 24280 -4218 24332 -4156
rect 24478 2128 24530 2134
rect 24478 492 24530 752
rect 24478 -1144 24530 -884
rect 24478 -2780 24530 -2520
rect 24478 -4166 24530 -4156
rect 24676 2128 24728 2138
rect 24676 492 24728 752
rect 24676 -1144 24728 -884
rect 24676 -2780 24728 -2520
rect 24676 -4218 24728 -4156
rect 24874 2128 24926 2134
rect 24874 492 24926 752
rect 24874 -1144 24926 -884
rect 24874 -2780 24926 -2520
rect 24874 -4166 24926 -4156
rect 25072 2128 25124 2138
rect 25072 492 25124 752
rect 25072 -1144 25124 -884
rect 25072 -2780 25124 -2520
rect 25072 -4218 25124 -4156
rect 25270 2128 25322 2134
rect 25270 492 25322 752
rect 25270 -1144 25322 -884
rect 25270 -2780 25322 -2520
rect 25270 -4166 25322 -4156
rect 25468 2128 25520 2138
rect 25468 492 25520 752
rect 25468 -1144 25520 -884
rect 25468 -2780 25520 -2520
rect 25468 -4218 25520 -4156
rect 25666 2128 25718 2134
rect 25666 492 25718 752
rect 25666 -1144 25718 -884
rect 25666 -2780 25718 -2520
rect 25666 -4166 25718 -4156
rect 25864 2128 25916 2138
rect 25864 492 25916 752
rect 25864 -1144 25916 -884
rect 25864 -2780 25916 -2520
rect 25864 -4218 25916 -4156
rect 26062 2128 26114 2134
rect 26062 492 26114 752
rect 26062 -1144 26114 -884
rect 26062 -2780 26114 -2520
rect 26062 -4166 26114 -4156
rect 26260 2128 26312 2138
rect 26260 492 26312 752
rect 26260 -1144 26312 -884
rect 26260 -2780 26312 -2520
rect 26260 -4218 26312 -4156
rect 26458 2128 26510 2134
rect 26458 492 26510 752
rect 26458 -1144 26510 -884
rect 26458 -2780 26510 -2520
rect 26458 -4166 26510 -4156
rect 26656 2128 26708 2138
rect 26656 492 26708 752
rect 26656 -1144 26708 -884
rect 26656 -2780 26708 -2520
rect 26656 -4218 26708 -4156
rect 26854 2128 26906 2134
rect 26854 492 26906 752
rect 26854 -1144 26906 -884
rect 26854 -2780 26906 -2520
rect 26854 -4166 26906 -4156
rect 27052 2128 27104 2138
rect 27052 492 27104 752
rect 27052 -1144 27104 -884
rect 27052 -2780 27104 -2520
rect 27052 -4218 27104 -4156
rect 27250 2128 27302 2134
rect 27250 492 27302 752
rect 27250 -1144 27302 -884
rect 27250 -2780 27302 -2520
rect 27250 -4166 27302 -4156
rect 27448 2128 27500 2138
rect 27448 492 27500 752
rect 27448 -1144 27500 -884
rect 27448 -2780 27500 -2520
rect 27448 -4218 27500 -4156
rect 27646 2128 27698 2134
rect 27646 492 27698 752
rect 27646 -1144 27698 -884
rect 27646 -2780 27698 -2520
rect 27646 -4166 27698 -4156
rect 27844 2128 27896 2138
rect 27844 492 27896 752
rect 27844 -1144 27896 -884
rect 27844 -2780 27896 -2520
rect 27844 -4218 27896 -4156
rect 28042 2128 28094 2134
rect 28042 492 28094 752
rect 28042 -1144 28094 -884
rect 28042 -2780 28094 -2520
rect 28042 -4166 28094 -4156
rect 28240 2128 28292 2138
rect 28240 492 28292 752
rect 28240 -1144 28292 -884
rect 28240 -2780 28292 -2520
rect 28240 -4218 28292 -4156
rect 28438 2128 28490 2134
rect 28438 492 28490 752
rect 28438 -1144 28490 -884
rect 28438 -2780 28490 -2520
rect 28438 -4166 28490 -4156
rect 28636 2128 28688 2138
rect 28636 492 28688 752
rect 28636 -1144 28688 -884
rect 28636 -2780 28688 -2520
rect 28636 -4218 28688 -4156
rect 28834 2128 28886 2134
rect 28834 492 28886 752
rect 28834 -1144 28886 -884
rect 28834 -2780 28886 -2520
rect 28834 -4166 28886 -4156
rect 29032 2128 29084 2138
rect 29032 492 29084 752
rect 29032 -1144 29084 -884
rect 29032 -2780 29084 -2520
rect 29032 -4218 29084 -4156
rect 29230 2128 29282 2134
rect 29230 492 29282 752
rect 29230 -1144 29282 -884
rect 29230 -2780 29282 -2520
rect 29230 -4166 29282 -4156
rect 29428 2128 29480 2138
rect 29428 492 29480 752
rect 29428 -1144 29480 -884
rect 29428 -2780 29480 -2520
rect 29428 -4218 29480 -4156
rect 29626 2128 29678 2134
rect 29626 492 29678 752
rect 29626 -1144 29678 -884
rect 29626 -2780 29678 -2520
rect 29626 -4166 29678 -4156
rect 29824 2128 29876 2138
rect 29824 492 29876 752
rect 29824 -1144 29876 -884
rect 29824 -2780 29876 -2520
rect 29824 -4218 29876 -4156
rect 30022 2128 30074 2134
rect 30022 492 30074 752
rect 30022 -1144 30074 -884
rect 30022 -2780 30074 -2520
rect 30022 -4166 30074 -4156
rect 30220 2128 30272 2138
rect 30220 492 30272 752
rect 30220 -1144 30272 -884
rect 30220 -2780 30272 -2520
rect 30220 -4218 30272 -4156
rect 30418 2128 30470 2134
rect 30418 492 30470 752
rect 30418 -1144 30470 -884
rect 30418 -2780 30470 -2520
rect 30418 -4166 30470 -4156
rect 30616 2128 30668 2138
rect 30616 492 30668 752
rect 30616 -1144 30668 -884
rect 30616 -2780 30668 -2520
rect 30616 -4218 30668 -4156
rect 30814 2128 30866 2134
rect 30814 492 30866 752
rect 30814 -1144 30866 -884
rect 30814 -2780 30866 -2520
rect 30814 -4166 30866 -4156
rect 31012 2128 31064 2138
rect 31012 492 31064 752
rect 31012 -1144 31064 -884
rect 31012 -2780 31064 -2520
rect 31012 -4218 31064 -4156
rect 31210 2128 31262 2134
rect 31210 492 31262 752
rect 31210 -1144 31262 -884
rect 31210 -2780 31262 -2520
rect 31210 -4166 31262 -4156
rect 31408 2128 31460 2138
rect 31408 492 31460 752
rect 31408 -1144 31460 -884
rect 31408 -2780 31460 -2520
rect 31408 -4218 31460 -4156
rect 31606 2129 31658 2135
rect 31606 493 31658 753
rect 31606 -1143 31658 -883
rect 31606 -2779 31658 -2519
rect 31606 -4165 31658 -4155
rect -225 -4240 -129 -4218
rect -225 -4296 -203 -4240
rect -147 -4296 -129 -4240
rect -225 -4314 -129 -4296
rect 171 -4240 267 -4218
rect 171 -4296 193 -4240
rect 249 -4296 267 -4240
rect 171 -4314 267 -4296
rect 567 -4240 663 -4218
rect 567 -4296 589 -4240
rect 645 -4296 663 -4240
rect 567 -4314 663 -4296
rect 963 -4240 1059 -4218
rect 963 -4296 985 -4240
rect 1041 -4296 1059 -4240
rect 963 -4314 1059 -4296
rect 1359 -4240 1455 -4218
rect 1359 -4296 1381 -4240
rect 1437 -4296 1455 -4240
rect 1359 -4314 1455 -4296
rect 1755 -4240 1851 -4218
rect 1755 -4296 1777 -4240
rect 1833 -4296 1851 -4240
rect 1755 -4314 1851 -4296
rect 2151 -4240 2247 -4218
rect 2151 -4296 2173 -4240
rect 2229 -4296 2247 -4240
rect 2151 -4314 2247 -4296
rect 2547 -4240 2643 -4218
rect 2547 -4296 2569 -4240
rect 2625 -4296 2643 -4240
rect 2547 -4314 2643 -4296
rect 2943 -4240 3039 -4218
rect 2943 -4296 2965 -4240
rect 3021 -4296 3039 -4240
rect 2943 -4314 3039 -4296
rect 3339 -4240 3435 -4218
rect 3339 -4296 3361 -4240
rect 3417 -4296 3435 -4240
rect 3339 -4314 3435 -4296
rect 3735 -4240 3831 -4218
rect 3735 -4296 3757 -4240
rect 3813 -4296 3831 -4240
rect 3735 -4314 3831 -4296
rect 4131 -4240 4227 -4218
rect 4131 -4296 4153 -4240
rect 4209 -4296 4227 -4240
rect 4131 -4314 4227 -4296
rect 4527 -4240 4623 -4218
rect 4527 -4296 4549 -4240
rect 4605 -4296 4623 -4240
rect 4527 -4314 4623 -4296
rect 4923 -4240 5019 -4218
rect 4923 -4296 4945 -4240
rect 5001 -4296 5019 -4240
rect 4923 -4314 5019 -4296
rect 5319 -4240 5415 -4218
rect 5319 -4296 5341 -4240
rect 5397 -4296 5415 -4240
rect 5319 -4314 5415 -4296
rect 5715 -4240 5811 -4218
rect 5715 -4296 5737 -4240
rect 5793 -4296 5811 -4240
rect 5715 -4314 5811 -4296
rect 6111 -4240 6207 -4218
rect 6111 -4296 6133 -4240
rect 6189 -4296 6207 -4240
rect 6111 -4314 6207 -4296
rect 6507 -4240 6603 -4218
rect 6507 -4296 6529 -4240
rect 6585 -4296 6603 -4240
rect 6507 -4314 6603 -4296
rect 6903 -4240 6999 -4218
rect 6903 -4296 6925 -4240
rect 6981 -4296 6999 -4240
rect 6903 -4314 6999 -4296
rect 7299 -4240 7395 -4218
rect 7299 -4296 7321 -4240
rect 7377 -4296 7395 -4240
rect 7299 -4314 7395 -4296
rect 7695 -4240 7791 -4218
rect 7695 -4296 7717 -4240
rect 7773 -4296 7791 -4240
rect 7695 -4314 7791 -4296
rect 11614 -4240 11710 -4218
rect 11614 -4296 11636 -4240
rect 11692 -4296 11710 -4240
rect 11614 -4314 11710 -4296
rect 12010 -4240 12106 -4218
rect 12010 -4296 12032 -4240
rect 12088 -4296 12106 -4240
rect 12010 -4314 12106 -4296
rect 12406 -4240 12502 -4218
rect 12406 -4296 12428 -4240
rect 12484 -4296 12502 -4240
rect 12406 -4314 12502 -4296
rect 12802 -4240 12898 -4218
rect 12802 -4296 12824 -4240
rect 12880 -4296 12898 -4240
rect 12802 -4314 12898 -4296
rect 13198 -4240 13294 -4218
rect 13198 -4296 13220 -4240
rect 13276 -4296 13294 -4240
rect 13198 -4314 13294 -4296
rect 13594 -4240 13690 -4218
rect 13594 -4296 13616 -4240
rect 13672 -4296 13690 -4240
rect 13594 -4314 13690 -4296
rect 13990 -4240 14086 -4218
rect 13990 -4296 14012 -4240
rect 14068 -4296 14086 -4240
rect 13990 -4314 14086 -4296
rect 14386 -4240 14482 -4218
rect 14386 -4296 14408 -4240
rect 14464 -4296 14482 -4240
rect 14386 -4314 14482 -4296
rect 14782 -4240 14878 -4218
rect 14782 -4296 14804 -4240
rect 14860 -4296 14878 -4240
rect 14782 -4314 14878 -4296
rect 15178 -4240 15274 -4218
rect 15178 -4296 15200 -4240
rect 15256 -4296 15274 -4240
rect 15178 -4314 15274 -4296
rect 15574 -4240 15670 -4218
rect 15574 -4296 15596 -4240
rect 15652 -4296 15670 -4240
rect 15574 -4314 15670 -4296
rect 15970 -4240 16066 -4218
rect 15970 -4296 15992 -4240
rect 16048 -4296 16066 -4240
rect 15970 -4314 16066 -4296
rect 16366 -4240 16462 -4218
rect 16366 -4296 16388 -4240
rect 16444 -4296 16462 -4240
rect 16366 -4314 16462 -4296
rect 16762 -4240 16858 -4218
rect 16762 -4296 16784 -4240
rect 16840 -4296 16858 -4240
rect 16762 -4314 16858 -4296
rect 17158 -4240 17254 -4218
rect 17158 -4296 17180 -4240
rect 17236 -4296 17254 -4240
rect 17158 -4314 17254 -4296
rect 17554 -4240 17650 -4218
rect 17554 -4296 17576 -4240
rect 17632 -4296 17650 -4240
rect 17554 -4314 17650 -4296
rect 17950 -4240 18046 -4218
rect 17950 -4296 17972 -4240
rect 18028 -4296 18046 -4240
rect 17950 -4314 18046 -4296
rect 18346 -4240 18442 -4218
rect 18346 -4296 18368 -4240
rect 18424 -4296 18442 -4240
rect 18346 -4314 18442 -4296
rect 18742 -4240 18838 -4218
rect 18742 -4296 18764 -4240
rect 18820 -4296 18838 -4240
rect 18742 -4314 18838 -4296
rect 19138 -4240 19234 -4218
rect 19138 -4296 19160 -4240
rect 19216 -4296 19234 -4240
rect 19138 -4314 19234 -4296
rect 19534 -4240 19630 -4218
rect 19534 -4296 19556 -4240
rect 19612 -4296 19630 -4240
rect 19534 -4314 19630 -4296
rect 23464 -4240 23560 -4218
rect 23464 -4296 23486 -4240
rect 23542 -4296 23560 -4240
rect 23464 -4314 23560 -4296
rect 23860 -4240 23956 -4218
rect 23860 -4296 23882 -4240
rect 23938 -4296 23956 -4240
rect 23860 -4314 23956 -4296
rect 24256 -4240 24352 -4218
rect 24256 -4296 24278 -4240
rect 24334 -4296 24352 -4240
rect 24256 -4314 24352 -4296
rect 24652 -4240 24748 -4218
rect 24652 -4296 24674 -4240
rect 24730 -4296 24748 -4240
rect 24652 -4314 24748 -4296
rect 25048 -4240 25144 -4218
rect 25048 -4296 25070 -4240
rect 25126 -4296 25144 -4240
rect 25048 -4314 25144 -4296
rect 25444 -4240 25540 -4218
rect 25444 -4296 25466 -4240
rect 25522 -4296 25540 -4240
rect 25444 -4314 25540 -4296
rect 25840 -4240 25936 -4218
rect 25840 -4296 25862 -4240
rect 25918 -4296 25936 -4240
rect 25840 -4314 25936 -4296
rect 26236 -4240 26332 -4218
rect 26236 -4296 26258 -4240
rect 26314 -4296 26332 -4240
rect 26236 -4314 26332 -4296
rect 26632 -4240 26728 -4218
rect 26632 -4296 26654 -4240
rect 26710 -4296 26728 -4240
rect 26632 -4314 26728 -4296
rect 27028 -4240 27124 -4218
rect 27028 -4296 27050 -4240
rect 27106 -4296 27124 -4240
rect 27028 -4314 27124 -4296
rect 27424 -4240 27520 -4218
rect 27424 -4296 27446 -4240
rect 27502 -4296 27520 -4240
rect 27424 -4314 27520 -4296
rect 27820 -4240 27916 -4218
rect 27820 -4296 27842 -4240
rect 27898 -4296 27916 -4240
rect 27820 -4314 27916 -4296
rect 28216 -4240 28312 -4218
rect 28216 -4296 28238 -4240
rect 28294 -4296 28312 -4240
rect 28216 -4314 28312 -4296
rect 28612 -4240 28708 -4218
rect 28612 -4296 28634 -4240
rect 28690 -4296 28708 -4240
rect 28612 -4314 28708 -4296
rect 29008 -4240 29104 -4218
rect 29008 -4296 29030 -4240
rect 29086 -4296 29104 -4240
rect 29008 -4314 29104 -4296
rect 29404 -4240 29500 -4218
rect 29404 -4296 29426 -4240
rect 29482 -4296 29500 -4240
rect 29404 -4314 29500 -4296
rect 29800 -4240 29896 -4218
rect 29800 -4296 29822 -4240
rect 29878 -4296 29896 -4240
rect 29800 -4314 29896 -4296
rect 30196 -4240 30292 -4218
rect 30196 -4296 30218 -4240
rect 30274 -4296 30292 -4240
rect 30196 -4314 30292 -4296
rect 30592 -4240 30688 -4218
rect 30592 -4296 30614 -4240
rect 30670 -4296 30688 -4240
rect 30592 -4314 30688 -4296
rect 30988 -4240 31084 -4218
rect 30988 -4296 31010 -4240
rect 31066 -4296 31084 -4240
rect 30988 -4314 31084 -4296
rect 31384 -4240 31480 -4218
rect 31384 -4296 31406 -4240
rect 31462 -4296 31480 -4240
rect 31384 -4314 31480 -4296
<< via2 >>
rect -627 -877 -493 -743
rect -627 -1081 -493 -947
rect -627 -1285 -493 -1151
rect 8063 -877 8197 -743
rect 11212 -877 11346 -743
rect 8063 -1081 8197 -947
rect 11212 -1081 11346 -947
rect 8063 -1285 8197 -1151
rect 11212 -1285 11346 -1151
rect 19902 -877 20036 -743
rect 23062 -877 23196 -743
rect 19902 -1081 20036 -947
rect 23062 -1081 23196 -947
rect 19902 -1285 20036 -1151
rect 23062 -1285 23196 -1151
rect -203 -4296 -147 -4240
rect 193 -4296 249 -4240
rect 589 -4296 645 -4240
rect 985 -4296 1041 -4240
rect 1381 -4296 1437 -4240
rect 1777 -4296 1833 -4240
rect 2173 -4296 2229 -4240
rect 2569 -4296 2625 -4240
rect 2965 -4296 3021 -4240
rect 3361 -4296 3417 -4240
rect 3757 -4296 3813 -4240
rect 4153 -4296 4209 -4240
rect 4549 -4296 4605 -4240
rect 4945 -4296 5001 -4240
rect 5341 -4296 5397 -4240
rect 5737 -4296 5793 -4240
rect 6133 -4296 6189 -4240
rect 6529 -4296 6585 -4240
rect 6925 -4296 6981 -4240
rect 7321 -4296 7377 -4240
rect 7717 -4296 7773 -4240
rect 11636 -4296 11692 -4240
rect 12032 -4296 12088 -4240
rect 12428 -4296 12484 -4240
rect 12824 -4296 12880 -4240
rect 13220 -4296 13276 -4240
rect 13616 -4296 13672 -4240
rect 14012 -4296 14068 -4240
rect 14408 -4296 14464 -4240
rect 14804 -4296 14860 -4240
rect 15200 -4296 15256 -4240
rect 15596 -4296 15652 -4240
rect 15992 -4296 16048 -4240
rect 16388 -4296 16444 -4240
rect 16784 -4296 16840 -4240
rect 17180 -4296 17236 -4240
rect 17576 -4296 17632 -4240
rect 17972 -4296 18028 -4240
rect 18368 -4296 18424 -4240
rect 18764 -4296 18820 -4240
rect 19160 -4296 19216 -4240
rect 19556 -4296 19612 -4240
rect 23486 -4296 23542 -4240
rect 23882 -4296 23938 -4240
rect 24278 -4296 24334 -4240
rect 24674 -4296 24730 -4240
rect 25070 -4296 25126 -4240
rect 25466 -4296 25522 -4240
rect 25862 -4296 25918 -4240
rect 26258 -4296 26314 -4240
rect 26654 -4296 26710 -4240
rect 27050 -4296 27106 -4240
rect 27446 -4296 27502 -4240
rect 27842 -4296 27898 -4240
rect 28238 -4296 28294 -4240
rect 28634 -4296 28690 -4240
rect 29030 -4296 29086 -4240
rect 29426 -4296 29482 -4240
rect 29822 -4296 29878 -4240
rect 30218 -4296 30274 -4240
rect 30614 -4296 30670 -4240
rect 31010 -4296 31066 -4240
rect 31406 -4296 31462 -4240
<< metal3 >>
rect -637 -743 -483 -738
rect -637 -877 -627 -743
rect -493 -877 -483 -743
rect -637 -882 -483 -877
rect 8053 -743 11356 -738
rect 8053 -877 8063 -743
rect 8197 -877 11212 -743
rect 11346 -877 11356 -743
rect -637 -947 -483 -942
rect -637 -1081 -627 -947
rect -493 -1081 -483 -947
rect -637 -1086 -483 -1081
rect 8053 -947 11356 -877
rect 19892 -743 23206 -738
rect 19892 -877 19902 -743
rect 20036 -877 23062 -743
rect 23196 -877 23206 -743
rect 19892 -882 23206 -877
rect 20036 -942 23062 -882
rect 8053 -1081 8063 -947
rect 8197 -1081 11212 -947
rect 11346 -1081 11356 -947
rect -637 -1151 -483 -1146
rect -637 -1285 -627 -1151
rect -493 -1285 -483 -1151
rect -637 -1290 -483 -1285
rect 8053 -1151 11356 -1081
rect 19892 -947 23206 -942
rect 19892 -1081 19902 -947
rect 20036 -1081 23062 -947
rect 23196 -1081 23206 -947
rect 19892 -1086 23206 -1081
rect 20036 -1146 23062 -1086
rect 8053 -1285 8063 -1151
rect 8197 -1285 11212 -1151
rect 11346 -1285 11356 -1151
rect 8053 -1290 11356 -1285
rect 19892 -1151 23206 -1146
rect 19892 -1285 19902 -1151
rect 20036 -1285 23062 -1151
rect 23196 -1285 23206 -1151
rect 19892 -1290 23206 -1285
rect -225 -4240 7791 -4218
rect -225 -4296 -203 -4240
rect -147 -4296 193 -4240
rect 249 -4296 589 -4240
rect 645 -4296 985 -4240
rect 1041 -4296 1381 -4240
rect 1437 -4296 1777 -4240
rect 1833 -4296 2173 -4240
rect 2229 -4296 2569 -4240
rect 2625 -4296 2965 -4240
rect 3021 -4296 3361 -4240
rect 3417 -4296 3757 -4240
rect 3813 -4296 4153 -4240
rect 4209 -4296 4549 -4240
rect 4605 -4296 4945 -4240
rect 5001 -4296 5341 -4240
rect 5397 -4296 5737 -4240
rect 5793 -4296 6133 -4240
rect 6189 -4296 6529 -4240
rect 6585 -4296 6925 -4240
rect 6981 -4296 7321 -4240
rect 7377 -4296 7717 -4240
rect 7773 -4296 7791 -4240
rect -225 -4314 7791 -4296
rect 11614 -4240 19630 -4218
rect 11614 -4296 11636 -4240
rect 11692 -4296 12032 -4240
rect 12088 -4296 12428 -4240
rect 12484 -4296 12824 -4240
rect 12880 -4296 13220 -4240
rect 13276 -4296 13616 -4240
rect 13672 -4296 14012 -4240
rect 14068 -4296 14408 -4240
rect 14464 -4296 14804 -4240
rect 14860 -4296 15200 -4240
rect 15256 -4296 15596 -4240
rect 15652 -4296 15992 -4240
rect 16048 -4296 16388 -4240
rect 16444 -4296 16784 -4240
rect 16840 -4296 17180 -4240
rect 17236 -4296 17576 -4240
rect 17632 -4296 17972 -4240
rect 18028 -4296 18368 -4240
rect 18424 -4296 18764 -4240
rect 18820 -4296 19160 -4240
rect 19216 -4296 19556 -4240
rect 19612 -4296 19630 -4240
rect 11614 -4314 19630 -4296
rect 23464 -4240 31480 -4218
rect 23464 -4296 23486 -4240
rect 23542 -4296 23882 -4240
rect 23938 -4296 24278 -4240
rect 24334 -4296 24674 -4240
rect 24730 -4296 25070 -4240
rect 25126 -4296 25466 -4240
rect 25522 -4296 25862 -4240
rect 25918 -4296 26258 -4240
rect 26314 -4296 26654 -4240
rect 26710 -4296 27050 -4240
rect 27106 -4296 27446 -4240
rect 27502 -4296 27842 -4240
rect 27898 -4296 28238 -4240
rect 28294 -4296 28634 -4240
rect 28690 -4296 29030 -4240
rect 29086 -4296 29426 -4240
rect 29482 -4296 29822 -4240
rect 29878 -4296 30218 -4240
rect 30274 -4296 30614 -4240
rect 30670 -4296 31010 -4240
rect 31066 -4296 31406 -4240
rect 31462 -4296 31480 -4240
rect 23464 -4314 31480 -4296
use sky130_fd_pr__pfet_01v8_ZYZ5C6  sky130_fd_pr__pfet_01v8_ZYZ5C6_1
timestamp 1615920820
transform -1 0 3785 0 -1 -3432
box -4223 -764 4223 798
use sky130_fd_pr__pfet_01v8_ZYZ5C6  sky130_fd_pr__pfet_01v8_ZYZ5C6_0
timestamp 1615920820
transform 1 0 3785 0 1 1404
box -4223 -764 4223 798
use sky130_fd_pr__pfet_01v8_9JQ4XZ  sky130_fd_pr__pfet_01v8_9JQ4XZ_0
timestamp 1615920820
transform 1 0 3785 0 1 -1014
box -4223 -1618 4223 1618
<< end >>
