magic
tech sky130A
magscale 1 2
timestamp 1616093313
<< nwell >>
rect -203 -890 14571 1187
rect -944 -1621 14571 -890
rect -203 -3703 14571 -1621
rect -162 -3705 14202 -3703
<< pmoslvt >>
rect 143 -2531 223 -1731
rect 281 -2531 361 -1731
rect 419 -2531 499 -1731
rect 557 -2531 637 -1731
rect 695 -2531 775 -1731
rect 833 -2531 913 -1731
rect 971 -2531 1051 -1731
rect 1109 -2531 1189 -1731
rect 1247 -2531 1327 -1731
rect 1385 -2531 1465 -1731
rect 1523 -2531 1603 -1731
rect 1661 -2531 1741 -1731
rect 1799 -2531 1879 -1731
rect 1937 -2531 2017 -1731
rect 2075 -2531 2155 -1731
rect 2213 -2531 2293 -1731
rect 2351 -2531 2431 -1731
rect 2489 -2531 2569 -1731
rect 2627 -2531 2707 -1731
rect 2765 -2531 2845 -1731
rect 2903 -2531 2983 -1731
rect 3041 -2531 3121 -1731
rect 3179 -2531 3259 -1731
rect 3317 -2531 3397 -1731
rect 3455 -2531 3535 -1731
rect 3593 -2531 3673 -1731
rect 3731 -2531 3811 -1731
rect 3869 -2531 3949 -1731
rect 4007 -2531 4087 -1731
rect 4145 -2531 4225 -1731
rect 4283 -2531 4363 -1731
rect 4421 -2531 4501 -1731
rect 4559 -2531 4639 -1731
rect 4697 -2531 4777 -1731
rect 4835 -2531 4915 -1731
rect 4973 -2531 5053 -1731
rect 5111 -2531 5191 -1731
rect 5249 -2531 5329 -1731
rect 5387 -2531 5467 -1731
rect 5525 -2531 5605 -1731
rect 5663 -2531 5743 -1731
rect 5801 -2531 5881 -1731
rect 5939 -2531 6019 -1731
rect 6077 -2531 6157 -1731
rect 6215 -2531 6295 -1731
rect 6353 -2531 6433 -1731
rect 6491 -2531 6571 -1731
rect 6629 -2531 6709 -1731
rect 6767 -2531 6847 -1731
rect 6905 -2531 6985 -1731
rect 7043 -2531 7123 -1731
rect 7181 -2531 7261 -1731
rect 7319 -2531 7399 -1731
rect 7457 -2531 7537 -1731
rect 7595 -2531 7675 -1731
rect 7733 -2531 7813 -1731
rect 7871 -2531 7951 -1731
rect 8009 -2531 8089 -1731
rect 8147 -2531 8227 -1731
rect 8285 -2531 8365 -1731
rect 8423 -2531 8503 -1731
rect 8561 -2531 8641 -1731
rect 8699 -2531 8779 -1731
rect 8837 -2531 8917 -1731
rect 8975 -2531 9055 -1731
rect 9113 -2531 9193 -1731
rect 9251 -2531 9331 -1731
rect 9389 -2531 9469 -1731
rect 9527 -2531 9607 -1731
rect 9665 -2531 9745 -1731
rect 9803 -2531 9883 -1731
rect 9941 -2531 10021 -1731
rect 10079 -2531 10159 -1731
rect 10217 -2531 10297 -1731
rect 10355 -2531 10435 -1731
rect 10493 -2531 10573 -1731
rect 10631 -2531 10711 -1731
rect 10769 -2531 10849 -1731
rect 10907 -2531 10987 -1731
rect 11045 -2531 11125 -1731
rect 11183 -2531 11263 -1731
rect 11321 -2531 11401 -1731
rect 11459 -2531 11539 -1731
rect 11597 -2531 11677 -1731
rect 11735 -2531 11815 -1731
rect 11873 -2531 11953 -1731
rect 12011 -2531 12091 -1731
rect 12149 -2531 12229 -1731
rect 12287 -2531 12367 -1731
rect 12425 -2531 12505 -1731
rect 12563 -2531 12643 -1731
rect 12701 -2531 12781 -1731
rect 12839 -2531 12919 -1731
rect 12977 -2531 13057 -1731
rect 13115 -2531 13195 -1731
rect 13253 -2531 13333 -1731
rect 13391 -2531 13471 -1731
rect 13529 -2531 13609 -1731
rect 13667 -2531 13747 -1731
rect 13805 -2531 13885 -1731
rect 143 -3417 223 -2617
rect 281 -3417 361 -2617
rect 419 -3417 499 -2617
rect 557 -3417 637 -2617
rect 695 -3417 775 -2617
rect 833 -3417 913 -2617
rect 971 -3417 1051 -2617
rect 1109 -3417 1189 -2617
rect 1247 -3417 1327 -2617
rect 1385 -3417 1465 -2617
rect 1523 -3417 1603 -2617
rect 1661 -3417 1741 -2617
rect 1799 -3417 1879 -2617
rect 1937 -3417 2017 -2617
rect 2075 -3417 2155 -2617
rect 2213 -3417 2293 -2617
rect 2351 -3417 2431 -2617
rect 2489 -3417 2569 -2617
rect 2627 -3417 2707 -2617
rect 2765 -3417 2845 -2617
rect 2903 -3417 2983 -2617
rect 3041 -3417 3121 -2617
rect 3179 -3417 3259 -2617
rect 3317 -3417 3397 -2617
rect 3455 -3417 3535 -2617
rect 3593 -3417 3673 -2617
rect 3731 -3417 3811 -2617
rect 3869 -3417 3949 -2617
rect 4007 -3417 4087 -2617
rect 4145 -3417 4225 -2617
rect 4283 -3417 4363 -2617
rect 4421 -3417 4501 -2617
rect 4559 -3417 4639 -2617
rect 4697 -3417 4777 -2617
rect 4835 -3417 4915 -2617
rect 4973 -3417 5053 -2617
rect 5111 -3417 5191 -2617
rect 5249 -3417 5329 -2617
rect 5387 -3417 5467 -2617
rect 5525 -3417 5605 -2617
rect 5663 -3417 5743 -2617
rect 5801 -3417 5881 -2617
rect 5939 -3417 6019 -2617
rect 6077 -3417 6157 -2617
rect 6215 -3417 6295 -2617
rect 6353 -3417 6433 -2617
rect 6491 -3417 6571 -2617
rect 6629 -3417 6709 -2617
rect 6767 -3417 6847 -2617
rect 6905 -3417 6985 -2617
rect 7043 -3417 7123 -2617
rect 7181 -3417 7261 -2617
rect 7319 -3417 7399 -2617
rect 7457 -3417 7537 -2617
rect 7595 -3417 7675 -2617
rect 7733 -3417 7813 -2617
rect 7871 -3417 7951 -2617
rect 8009 -3417 8089 -2617
rect 8147 -3417 8227 -2617
rect 8285 -3417 8365 -2617
rect 8423 -3417 8503 -2617
rect 8561 -3417 8641 -2617
rect 8699 -3417 8779 -2617
rect 8837 -3417 8917 -2617
rect 8975 -3417 9055 -2617
rect 9113 -3417 9193 -2617
rect 9251 -3417 9331 -2617
rect 9389 -3417 9469 -2617
rect 9527 -3417 9607 -2617
rect 9665 -3417 9745 -2617
rect 9803 -3417 9883 -2617
rect 9941 -3417 10021 -2617
rect 10079 -3417 10159 -2617
rect 10217 -3417 10297 -2617
rect 10355 -3417 10435 -2617
rect 10493 -3417 10573 -2617
rect 10631 -3417 10711 -2617
rect 10769 -3417 10849 -2617
rect 10907 -3417 10987 -2617
rect 11045 -3417 11125 -2617
rect 11183 -3417 11263 -2617
rect 11321 -3417 11401 -2617
rect 11459 -3417 11539 -2617
rect 11597 -3417 11677 -2617
rect 11735 -3417 11815 -2617
rect 11873 -3417 11953 -2617
rect 12011 -3417 12091 -2617
rect 12149 -3417 12229 -2617
rect 12287 -3417 12367 -2617
rect 12425 -3417 12505 -2617
rect 12563 -3417 12643 -2617
rect 12701 -3417 12781 -2617
rect 12839 -3417 12919 -2617
rect 12977 -3417 13057 -2617
rect 13115 -3417 13195 -2617
rect 13253 -3417 13333 -2617
rect 13391 -3417 13471 -2617
rect 13529 -3417 13609 -2617
rect 13667 -3417 13747 -2617
rect 13805 -3417 13885 -2617
<< pdiff >>
rect 85 -1743 143 -1731
rect 85 -2519 97 -1743
rect 131 -2519 143 -1743
rect 85 -2531 143 -2519
rect 223 -1743 281 -1731
rect 223 -2519 235 -1743
rect 269 -2519 281 -1743
rect 223 -2531 281 -2519
rect 361 -1743 419 -1731
rect 361 -2519 373 -1743
rect 407 -2519 419 -1743
rect 361 -2531 419 -2519
rect 499 -1743 557 -1731
rect 499 -2519 511 -1743
rect 545 -2519 557 -1743
rect 499 -2531 557 -2519
rect 637 -1743 695 -1731
rect 637 -2519 649 -1743
rect 683 -2519 695 -1743
rect 637 -2531 695 -2519
rect 775 -1743 833 -1731
rect 775 -2519 787 -1743
rect 821 -2519 833 -1743
rect 775 -2531 833 -2519
rect 913 -1743 971 -1731
rect 913 -2519 925 -1743
rect 959 -2519 971 -1743
rect 913 -2531 971 -2519
rect 1051 -1743 1109 -1731
rect 1051 -2519 1063 -1743
rect 1097 -2519 1109 -1743
rect 1051 -2531 1109 -2519
rect 1189 -1743 1247 -1731
rect 1189 -2519 1201 -1743
rect 1235 -2519 1247 -1743
rect 1189 -2531 1247 -2519
rect 1327 -1743 1385 -1731
rect 1327 -2519 1339 -1743
rect 1373 -2519 1385 -1743
rect 1327 -2531 1385 -2519
rect 1465 -1743 1523 -1731
rect 1465 -2519 1477 -1743
rect 1511 -2519 1523 -1743
rect 1465 -2531 1523 -2519
rect 1603 -1743 1661 -1731
rect 1603 -2519 1615 -1743
rect 1649 -2519 1661 -1743
rect 1603 -2531 1661 -2519
rect 1741 -1743 1799 -1731
rect 1741 -2519 1753 -1743
rect 1787 -2519 1799 -1743
rect 1741 -2531 1799 -2519
rect 1879 -1743 1937 -1731
rect 1879 -2519 1891 -1743
rect 1925 -2519 1937 -1743
rect 1879 -2531 1937 -2519
rect 2017 -1743 2075 -1731
rect 2017 -2519 2029 -1743
rect 2063 -2519 2075 -1743
rect 2017 -2531 2075 -2519
rect 2155 -1743 2213 -1731
rect 2155 -2519 2167 -1743
rect 2201 -2519 2213 -1743
rect 2155 -2531 2213 -2519
rect 2293 -1743 2351 -1731
rect 2293 -2519 2305 -1743
rect 2339 -2519 2351 -1743
rect 2293 -2531 2351 -2519
rect 2431 -1743 2489 -1731
rect 2431 -2519 2443 -1743
rect 2477 -2519 2489 -1743
rect 2431 -2531 2489 -2519
rect 2569 -1743 2627 -1731
rect 2569 -2519 2581 -1743
rect 2615 -2519 2627 -1743
rect 2569 -2531 2627 -2519
rect 2707 -1743 2765 -1731
rect 2707 -2519 2719 -1743
rect 2753 -2519 2765 -1743
rect 2707 -2531 2765 -2519
rect 2845 -1743 2903 -1731
rect 2845 -2519 2857 -1743
rect 2891 -2519 2903 -1743
rect 2845 -2531 2903 -2519
rect 2983 -1743 3041 -1731
rect 2983 -2519 2995 -1743
rect 3029 -2519 3041 -1743
rect 2983 -2531 3041 -2519
rect 3121 -1743 3179 -1731
rect 3121 -2519 3133 -1743
rect 3167 -2519 3179 -1743
rect 3121 -2531 3179 -2519
rect 3259 -1743 3317 -1731
rect 3259 -2519 3271 -1743
rect 3305 -2519 3317 -1743
rect 3259 -2531 3317 -2519
rect 3397 -1743 3455 -1731
rect 3397 -2519 3409 -1743
rect 3443 -2519 3455 -1743
rect 3397 -2531 3455 -2519
rect 3535 -1743 3593 -1731
rect 3535 -2519 3547 -1743
rect 3581 -2519 3593 -1743
rect 3535 -2531 3593 -2519
rect 3673 -1743 3731 -1731
rect 3673 -2519 3685 -1743
rect 3719 -2519 3731 -1743
rect 3673 -2531 3731 -2519
rect 3811 -1743 3869 -1731
rect 3811 -2519 3823 -1743
rect 3857 -2519 3869 -1743
rect 3811 -2531 3869 -2519
rect 3949 -1743 4007 -1731
rect 3949 -2519 3961 -1743
rect 3995 -2519 4007 -1743
rect 3949 -2531 4007 -2519
rect 4087 -1743 4145 -1731
rect 4087 -2519 4099 -1743
rect 4133 -2519 4145 -1743
rect 4087 -2531 4145 -2519
rect 4225 -1743 4283 -1731
rect 4225 -2519 4237 -1743
rect 4271 -2519 4283 -1743
rect 4225 -2531 4283 -2519
rect 4363 -1743 4421 -1731
rect 4363 -2519 4375 -1743
rect 4409 -2519 4421 -1743
rect 4363 -2531 4421 -2519
rect 4501 -1743 4559 -1731
rect 4501 -2519 4513 -1743
rect 4547 -2519 4559 -1743
rect 4501 -2531 4559 -2519
rect 4639 -1743 4697 -1731
rect 4639 -2519 4651 -1743
rect 4685 -2519 4697 -1743
rect 4639 -2531 4697 -2519
rect 4777 -1743 4835 -1731
rect 4777 -2519 4789 -1743
rect 4823 -2519 4835 -1743
rect 4777 -2531 4835 -2519
rect 4915 -1743 4973 -1731
rect 4915 -2519 4927 -1743
rect 4961 -2519 4973 -1743
rect 4915 -2531 4973 -2519
rect 5053 -1743 5111 -1731
rect 5053 -2519 5065 -1743
rect 5099 -2519 5111 -1743
rect 5053 -2531 5111 -2519
rect 5191 -1743 5249 -1731
rect 5191 -2519 5203 -1743
rect 5237 -2519 5249 -1743
rect 5191 -2531 5249 -2519
rect 5329 -1743 5387 -1731
rect 5329 -2519 5341 -1743
rect 5375 -2519 5387 -1743
rect 5329 -2531 5387 -2519
rect 5467 -1743 5525 -1731
rect 5467 -2519 5479 -1743
rect 5513 -2519 5525 -1743
rect 5467 -2531 5525 -2519
rect 5605 -1743 5663 -1731
rect 5605 -2519 5617 -1743
rect 5651 -2519 5663 -1743
rect 5605 -2531 5663 -2519
rect 5743 -1743 5801 -1731
rect 5743 -2519 5755 -1743
rect 5789 -2519 5801 -1743
rect 5743 -2531 5801 -2519
rect 5881 -1743 5939 -1731
rect 5881 -2519 5893 -1743
rect 5927 -2519 5939 -1743
rect 5881 -2531 5939 -2519
rect 6019 -1743 6077 -1731
rect 6019 -2519 6031 -1743
rect 6065 -2519 6077 -1743
rect 6019 -2531 6077 -2519
rect 6157 -1743 6215 -1731
rect 6157 -2519 6169 -1743
rect 6203 -2519 6215 -1743
rect 6157 -2531 6215 -2519
rect 6295 -1743 6353 -1731
rect 6295 -2519 6307 -1743
rect 6341 -2519 6353 -1743
rect 6295 -2531 6353 -2519
rect 6433 -1743 6491 -1731
rect 6433 -2519 6445 -1743
rect 6479 -2519 6491 -1743
rect 6433 -2531 6491 -2519
rect 6571 -1743 6629 -1731
rect 6571 -2519 6583 -1743
rect 6617 -2519 6629 -1743
rect 6571 -2531 6629 -2519
rect 6709 -1743 6767 -1731
rect 6709 -2519 6721 -1743
rect 6755 -2519 6767 -1743
rect 6709 -2531 6767 -2519
rect 6847 -1743 6905 -1731
rect 6847 -2519 6859 -1743
rect 6893 -2519 6905 -1743
rect 6847 -2531 6905 -2519
rect 6985 -1743 7043 -1731
rect 6985 -2519 6997 -1743
rect 7031 -2519 7043 -1743
rect 6985 -2531 7043 -2519
rect 7123 -1743 7181 -1731
rect 7123 -2519 7135 -1743
rect 7169 -2519 7181 -1743
rect 7123 -2531 7181 -2519
rect 7261 -1743 7319 -1731
rect 7261 -2519 7273 -1743
rect 7307 -2519 7319 -1743
rect 7261 -2531 7319 -2519
rect 7399 -1743 7457 -1731
rect 7399 -2519 7411 -1743
rect 7445 -2519 7457 -1743
rect 7399 -2531 7457 -2519
rect 7537 -1743 7595 -1731
rect 7537 -2519 7549 -1743
rect 7583 -2519 7595 -1743
rect 7537 -2531 7595 -2519
rect 7675 -1743 7733 -1731
rect 7675 -2519 7687 -1743
rect 7721 -2519 7733 -1743
rect 7675 -2531 7733 -2519
rect 7813 -1743 7871 -1731
rect 7813 -2519 7825 -1743
rect 7859 -2519 7871 -1743
rect 7813 -2531 7871 -2519
rect 7951 -1743 8009 -1731
rect 7951 -2519 7963 -1743
rect 7997 -2519 8009 -1743
rect 7951 -2531 8009 -2519
rect 8089 -1743 8147 -1731
rect 8089 -2519 8101 -1743
rect 8135 -2519 8147 -1743
rect 8089 -2531 8147 -2519
rect 8227 -1743 8285 -1731
rect 8227 -2519 8239 -1743
rect 8273 -2519 8285 -1743
rect 8227 -2531 8285 -2519
rect 8365 -1743 8423 -1731
rect 8365 -2519 8377 -1743
rect 8411 -2519 8423 -1743
rect 8365 -2531 8423 -2519
rect 8503 -1743 8561 -1731
rect 8503 -2519 8515 -1743
rect 8549 -2519 8561 -1743
rect 8503 -2531 8561 -2519
rect 8641 -1743 8699 -1731
rect 8641 -2519 8653 -1743
rect 8687 -2519 8699 -1743
rect 8641 -2531 8699 -2519
rect 8779 -1743 8837 -1731
rect 8779 -2519 8791 -1743
rect 8825 -2519 8837 -1743
rect 8779 -2531 8837 -2519
rect 8917 -1743 8975 -1731
rect 8917 -2519 8929 -1743
rect 8963 -2519 8975 -1743
rect 8917 -2531 8975 -2519
rect 9055 -1743 9113 -1731
rect 9055 -2519 9067 -1743
rect 9101 -2519 9113 -1743
rect 9055 -2531 9113 -2519
rect 9193 -1743 9251 -1731
rect 9193 -2519 9205 -1743
rect 9239 -2519 9251 -1743
rect 9193 -2531 9251 -2519
rect 9331 -1743 9389 -1731
rect 9331 -2519 9343 -1743
rect 9377 -2519 9389 -1743
rect 9331 -2531 9389 -2519
rect 9469 -1743 9527 -1731
rect 9469 -2519 9481 -1743
rect 9515 -2519 9527 -1743
rect 9469 -2531 9527 -2519
rect 9607 -1743 9665 -1731
rect 9607 -2519 9619 -1743
rect 9653 -2519 9665 -1743
rect 9607 -2531 9665 -2519
rect 9745 -1743 9803 -1731
rect 9745 -2519 9757 -1743
rect 9791 -2519 9803 -1743
rect 9745 -2531 9803 -2519
rect 9883 -1743 9941 -1731
rect 9883 -2519 9895 -1743
rect 9929 -2519 9941 -1743
rect 9883 -2531 9941 -2519
rect 10021 -1743 10079 -1731
rect 10021 -2519 10033 -1743
rect 10067 -2519 10079 -1743
rect 10021 -2531 10079 -2519
rect 10159 -1743 10217 -1731
rect 10159 -2519 10171 -1743
rect 10205 -2519 10217 -1743
rect 10159 -2531 10217 -2519
rect 10297 -1743 10355 -1731
rect 10297 -2519 10309 -1743
rect 10343 -2519 10355 -1743
rect 10297 -2531 10355 -2519
rect 10435 -1743 10493 -1731
rect 10435 -2519 10447 -1743
rect 10481 -2519 10493 -1743
rect 10435 -2531 10493 -2519
rect 10573 -1743 10631 -1731
rect 10573 -2519 10585 -1743
rect 10619 -2519 10631 -1743
rect 10573 -2531 10631 -2519
rect 10711 -1743 10769 -1731
rect 10711 -2519 10723 -1743
rect 10757 -2519 10769 -1743
rect 10711 -2531 10769 -2519
rect 10849 -1743 10907 -1731
rect 10849 -2519 10861 -1743
rect 10895 -2519 10907 -1743
rect 10849 -2531 10907 -2519
rect 10987 -1743 11045 -1731
rect 10987 -2519 10999 -1743
rect 11033 -2519 11045 -1743
rect 10987 -2531 11045 -2519
rect 11125 -1743 11183 -1731
rect 11125 -2519 11137 -1743
rect 11171 -2519 11183 -1743
rect 11125 -2531 11183 -2519
rect 11263 -1743 11321 -1731
rect 11263 -2519 11275 -1743
rect 11309 -2519 11321 -1743
rect 11263 -2531 11321 -2519
rect 11401 -1743 11459 -1731
rect 11401 -2519 11413 -1743
rect 11447 -2519 11459 -1743
rect 11401 -2531 11459 -2519
rect 11539 -1743 11597 -1731
rect 11539 -2519 11551 -1743
rect 11585 -2519 11597 -1743
rect 11539 -2531 11597 -2519
rect 11677 -1743 11735 -1731
rect 11677 -2519 11689 -1743
rect 11723 -2519 11735 -1743
rect 11677 -2531 11735 -2519
rect 11815 -1743 11873 -1731
rect 11815 -2519 11827 -1743
rect 11861 -2519 11873 -1743
rect 11815 -2531 11873 -2519
rect 11953 -1743 12011 -1731
rect 11953 -2519 11965 -1743
rect 11999 -2519 12011 -1743
rect 11953 -2531 12011 -2519
rect 12091 -1743 12149 -1731
rect 12091 -2519 12103 -1743
rect 12137 -2519 12149 -1743
rect 12091 -2531 12149 -2519
rect 12229 -1743 12287 -1731
rect 12229 -2519 12241 -1743
rect 12275 -2519 12287 -1743
rect 12229 -2531 12287 -2519
rect 12367 -1743 12425 -1731
rect 12367 -2519 12379 -1743
rect 12413 -2519 12425 -1743
rect 12367 -2531 12425 -2519
rect 12505 -1743 12563 -1731
rect 12505 -2519 12517 -1743
rect 12551 -2519 12563 -1743
rect 12505 -2531 12563 -2519
rect 12643 -1743 12701 -1731
rect 12643 -2519 12655 -1743
rect 12689 -2519 12701 -1743
rect 12643 -2531 12701 -2519
rect 12781 -1743 12839 -1731
rect 12781 -2519 12793 -1743
rect 12827 -2519 12839 -1743
rect 12781 -2531 12839 -2519
rect 12919 -1743 12977 -1731
rect 12919 -2519 12931 -1743
rect 12965 -2519 12977 -1743
rect 12919 -2531 12977 -2519
rect 13057 -1743 13115 -1731
rect 13057 -2519 13069 -1743
rect 13103 -2519 13115 -1743
rect 13057 -2531 13115 -2519
rect 13195 -1743 13253 -1731
rect 13195 -2519 13207 -1743
rect 13241 -2519 13253 -1743
rect 13195 -2531 13253 -2519
rect 13333 -1743 13391 -1731
rect 13333 -2519 13345 -1743
rect 13379 -2519 13391 -1743
rect 13333 -2531 13391 -2519
rect 13471 -1743 13529 -1731
rect 13471 -2519 13483 -1743
rect 13517 -2519 13529 -1743
rect 13471 -2531 13529 -2519
rect 13609 -1743 13667 -1731
rect 13609 -2519 13621 -1743
rect 13655 -2519 13667 -1743
rect 13609 -2531 13667 -2519
rect 13747 -1743 13805 -1731
rect 13747 -2519 13759 -1743
rect 13793 -2519 13805 -1743
rect 13747 -2531 13805 -2519
rect 13885 -1743 13943 -1731
rect 13885 -2519 13897 -1743
rect 13931 -2519 13943 -1743
rect 13885 -2531 13943 -2519
rect 85 -2629 143 -2617
rect 85 -3405 97 -2629
rect 131 -3405 143 -2629
rect 85 -3417 143 -3405
rect 223 -2629 281 -2617
rect 223 -3405 235 -2629
rect 269 -3405 281 -2629
rect 223 -3417 281 -3405
rect 361 -2629 419 -2617
rect 361 -3405 373 -2629
rect 407 -3405 419 -2629
rect 361 -3417 419 -3405
rect 499 -2629 557 -2617
rect 499 -3405 511 -2629
rect 545 -3405 557 -2629
rect 499 -3417 557 -3405
rect 637 -2629 695 -2617
rect 637 -3405 649 -2629
rect 683 -3405 695 -2629
rect 637 -3417 695 -3405
rect 775 -2629 833 -2617
rect 775 -3405 787 -2629
rect 821 -3405 833 -2629
rect 775 -3417 833 -3405
rect 913 -2629 971 -2617
rect 913 -3405 925 -2629
rect 959 -3405 971 -2629
rect 913 -3417 971 -3405
rect 1051 -2629 1109 -2617
rect 1051 -3405 1063 -2629
rect 1097 -3405 1109 -2629
rect 1051 -3417 1109 -3405
rect 1189 -2629 1247 -2617
rect 1189 -3405 1201 -2629
rect 1235 -3405 1247 -2629
rect 1189 -3417 1247 -3405
rect 1327 -2629 1385 -2617
rect 1327 -3405 1339 -2629
rect 1373 -3405 1385 -2629
rect 1327 -3417 1385 -3405
rect 1465 -2629 1523 -2617
rect 1465 -3405 1477 -2629
rect 1511 -3405 1523 -2629
rect 1465 -3417 1523 -3405
rect 1603 -2629 1661 -2617
rect 1603 -3405 1615 -2629
rect 1649 -3405 1661 -2629
rect 1603 -3417 1661 -3405
rect 1741 -2629 1799 -2617
rect 1741 -3405 1753 -2629
rect 1787 -3405 1799 -2629
rect 1741 -3417 1799 -3405
rect 1879 -2629 1937 -2617
rect 1879 -3405 1891 -2629
rect 1925 -3405 1937 -2629
rect 1879 -3417 1937 -3405
rect 2017 -2629 2075 -2617
rect 2017 -3405 2029 -2629
rect 2063 -3405 2075 -2629
rect 2017 -3417 2075 -3405
rect 2155 -2629 2213 -2617
rect 2155 -3405 2167 -2629
rect 2201 -3405 2213 -2629
rect 2155 -3417 2213 -3405
rect 2293 -2629 2351 -2617
rect 2293 -3405 2305 -2629
rect 2339 -3405 2351 -2629
rect 2293 -3417 2351 -3405
rect 2431 -2629 2489 -2617
rect 2431 -3405 2443 -2629
rect 2477 -3405 2489 -2629
rect 2431 -3417 2489 -3405
rect 2569 -2629 2627 -2617
rect 2569 -3405 2581 -2629
rect 2615 -3405 2627 -2629
rect 2569 -3417 2627 -3405
rect 2707 -2629 2765 -2617
rect 2707 -3405 2719 -2629
rect 2753 -3405 2765 -2629
rect 2707 -3417 2765 -3405
rect 2845 -2629 2903 -2617
rect 2845 -3405 2857 -2629
rect 2891 -3405 2903 -2629
rect 2845 -3417 2903 -3405
rect 2983 -2629 3041 -2617
rect 2983 -3405 2995 -2629
rect 3029 -3405 3041 -2629
rect 2983 -3417 3041 -3405
rect 3121 -2629 3179 -2617
rect 3121 -3405 3133 -2629
rect 3167 -3405 3179 -2629
rect 3121 -3417 3179 -3405
rect 3259 -2629 3317 -2617
rect 3259 -3405 3271 -2629
rect 3305 -3405 3317 -2629
rect 3259 -3417 3317 -3405
rect 3397 -2629 3455 -2617
rect 3397 -3405 3409 -2629
rect 3443 -3405 3455 -2629
rect 3397 -3417 3455 -3405
rect 3535 -2629 3593 -2617
rect 3535 -3405 3547 -2629
rect 3581 -3405 3593 -2629
rect 3535 -3417 3593 -3405
rect 3673 -2629 3731 -2617
rect 3673 -3405 3685 -2629
rect 3719 -3405 3731 -2629
rect 3673 -3417 3731 -3405
rect 3811 -2629 3869 -2617
rect 3811 -3405 3823 -2629
rect 3857 -3405 3869 -2629
rect 3811 -3417 3869 -3405
rect 3949 -2629 4007 -2617
rect 3949 -3405 3961 -2629
rect 3995 -3405 4007 -2629
rect 3949 -3417 4007 -3405
rect 4087 -2629 4145 -2617
rect 4087 -3405 4099 -2629
rect 4133 -3405 4145 -2629
rect 4087 -3417 4145 -3405
rect 4225 -2629 4283 -2617
rect 4225 -3405 4237 -2629
rect 4271 -3405 4283 -2629
rect 4225 -3417 4283 -3405
rect 4363 -2629 4421 -2617
rect 4363 -3405 4375 -2629
rect 4409 -3405 4421 -2629
rect 4363 -3417 4421 -3405
rect 4501 -2629 4559 -2617
rect 4501 -3405 4513 -2629
rect 4547 -3405 4559 -2629
rect 4501 -3417 4559 -3405
rect 4639 -2629 4697 -2617
rect 4639 -3405 4651 -2629
rect 4685 -3405 4697 -2629
rect 4639 -3417 4697 -3405
rect 4777 -2629 4835 -2617
rect 4777 -3405 4789 -2629
rect 4823 -3405 4835 -2629
rect 4777 -3417 4835 -3405
rect 4915 -2629 4973 -2617
rect 4915 -3405 4927 -2629
rect 4961 -3405 4973 -2629
rect 4915 -3417 4973 -3405
rect 5053 -2629 5111 -2617
rect 5053 -3405 5065 -2629
rect 5099 -3405 5111 -2629
rect 5053 -3417 5111 -3405
rect 5191 -2629 5249 -2617
rect 5191 -3405 5203 -2629
rect 5237 -3405 5249 -2629
rect 5191 -3417 5249 -3405
rect 5329 -2629 5387 -2617
rect 5329 -3405 5341 -2629
rect 5375 -3405 5387 -2629
rect 5329 -3417 5387 -3405
rect 5467 -2629 5525 -2617
rect 5467 -3405 5479 -2629
rect 5513 -3405 5525 -2629
rect 5467 -3417 5525 -3405
rect 5605 -2629 5663 -2617
rect 5605 -3405 5617 -2629
rect 5651 -3405 5663 -2629
rect 5605 -3417 5663 -3405
rect 5743 -2629 5801 -2617
rect 5743 -3405 5755 -2629
rect 5789 -3405 5801 -2629
rect 5743 -3417 5801 -3405
rect 5881 -2629 5939 -2617
rect 5881 -3405 5893 -2629
rect 5927 -3405 5939 -2629
rect 5881 -3417 5939 -3405
rect 6019 -2629 6077 -2617
rect 6019 -3405 6031 -2629
rect 6065 -3405 6077 -2629
rect 6019 -3417 6077 -3405
rect 6157 -2629 6215 -2617
rect 6157 -3405 6169 -2629
rect 6203 -3405 6215 -2629
rect 6157 -3417 6215 -3405
rect 6295 -2629 6353 -2617
rect 6295 -3405 6307 -2629
rect 6341 -3405 6353 -2629
rect 6295 -3417 6353 -3405
rect 6433 -2629 6491 -2617
rect 6433 -3405 6445 -2629
rect 6479 -3405 6491 -2629
rect 6433 -3417 6491 -3405
rect 6571 -2629 6629 -2617
rect 6571 -3405 6583 -2629
rect 6617 -3405 6629 -2629
rect 6571 -3417 6629 -3405
rect 6709 -2629 6767 -2617
rect 6709 -3405 6721 -2629
rect 6755 -3405 6767 -2629
rect 6709 -3417 6767 -3405
rect 6847 -2629 6905 -2617
rect 6847 -3405 6859 -2629
rect 6893 -3405 6905 -2629
rect 6847 -3417 6905 -3405
rect 6985 -2629 7043 -2617
rect 6985 -3405 6997 -2629
rect 7031 -3405 7043 -2629
rect 6985 -3417 7043 -3405
rect 7123 -2629 7181 -2617
rect 7123 -3405 7135 -2629
rect 7169 -3405 7181 -2629
rect 7123 -3417 7181 -3405
rect 7261 -2629 7319 -2617
rect 7261 -3405 7273 -2629
rect 7307 -3405 7319 -2629
rect 7261 -3417 7319 -3405
rect 7399 -2629 7457 -2617
rect 7399 -3405 7411 -2629
rect 7445 -3405 7457 -2629
rect 7399 -3417 7457 -3405
rect 7537 -2629 7595 -2617
rect 7537 -3405 7549 -2629
rect 7583 -3405 7595 -2629
rect 7537 -3417 7595 -3405
rect 7675 -2629 7733 -2617
rect 7675 -3405 7687 -2629
rect 7721 -3405 7733 -2629
rect 7675 -3417 7733 -3405
rect 7813 -2629 7871 -2617
rect 7813 -3405 7825 -2629
rect 7859 -3405 7871 -2629
rect 7813 -3417 7871 -3405
rect 7951 -2629 8009 -2617
rect 7951 -3405 7963 -2629
rect 7997 -3405 8009 -2629
rect 7951 -3417 8009 -3405
rect 8089 -2629 8147 -2617
rect 8089 -3405 8101 -2629
rect 8135 -3405 8147 -2629
rect 8089 -3417 8147 -3405
rect 8227 -2629 8285 -2617
rect 8227 -3405 8239 -2629
rect 8273 -3405 8285 -2629
rect 8227 -3417 8285 -3405
rect 8365 -2629 8423 -2617
rect 8365 -3405 8377 -2629
rect 8411 -3405 8423 -2629
rect 8365 -3417 8423 -3405
rect 8503 -2629 8561 -2617
rect 8503 -3405 8515 -2629
rect 8549 -3405 8561 -2629
rect 8503 -3417 8561 -3405
rect 8641 -2629 8699 -2617
rect 8641 -3405 8653 -2629
rect 8687 -3405 8699 -2629
rect 8641 -3417 8699 -3405
rect 8779 -2629 8837 -2617
rect 8779 -3405 8791 -2629
rect 8825 -3405 8837 -2629
rect 8779 -3417 8837 -3405
rect 8917 -2629 8975 -2617
rect 8917 -3405 8929 -2629
rect 8963 -3405 8975 -2629
rect 8917 -3417 8975 -3405
rect 9055 -2629 9113 -2617
rect 9055 -3405 9067 -2629
rect 9101 -3405 9113 -2629
rect 9055 -3417 9113 -3405
rect 9193 -2629 9251 -2617
rect 9193 -3405 9205 -2629
rect 9239 -3405 9251 -2629
rect 9193 -3417 9251 -3405
rect 9331 -2629 9389 -2617
rect 9331 -3405 9343 -2629
rect 9377 -3405 9389 -2629
rect 9331 -3417 9389 -3405
rect 9469 -2629 9527 -2617
rect 9469 -3405 9481 -2629
rect 9515 -3405 9527 -2629
rect 9469 -3417 9527 -3405
rect 9607 -2629 9665 -2617
rect 9607 -3405 9619 -2629
rect 9653 -3405 9665 -2629
rect 9607 -3417 9665 -3405
rect 9745 -2629 9803 -2617
rect 9745 -3405 9757 -2629
rect 9791 -3405 9803 -2629
rect 9745 -3417 9803 -3405
rect 9883 -2629 9941 -2617
rect 9883 -3405 9895 -2629
rect 9929 -3405 9941 -2629
rect 9883 -3417 9941 -3405
rect 10021 -2629 10079 -2617
rect 10021 -3405 10033 -2629
rect 10067 -3405 10079 -2629
rect 10021 -3417 10079 -3405
rect 10159 -2629 10217 -2617
rect 10159 -3405 10171 -2629
rect 10205 -3405 10217 -2629
rect 10159 -3417 10217 -3405
rect 10297 -2629 10355 -2617
rect 10297 -3405 10309 -2629
rect 10343 -3405 10355 -2629
rect 10297 -3417 10355 -3405
rect 10435 -2629 10493 -2617
rect 10435 -3405 10447 -2629
rect 10481 -3405 10493 -2629
rect 10435 -3417 10493 -3405
rect 10573 -2629 10631 -2617
rect 10573 -3405 10585 -2629
rect 10619 -3405 10631 -2629
rect 10573 -3417 10631 -3405
rect 10711 -2629 10769 -2617
rect 10711 -3405 10723 -2629
rect 10757 -3405 10769 -2629
rect 10711 -3417 10769 -3405
rect 10849 -2629 10907 -2617
rect 10849 -3405 10861 -2629
rect 10895 -3405 10907 -2629
rect 10849 -3417 10907 -3405
rect 10987 -2629 11045 -2617
rect 10987 -3405 10999 -2629
rect 11033 -3405 11045 -2629
rect 10987 -3417 11045 -3405
rect 11125 -2629 11183 -2617
rect 11125 -3405 11137 -2629
rect 11171 -3405 11183 -2629
rect 11125 -3417 11183 -3405
rect 11263 -2629 11321 -2617
rect 11263 -3405 11275 -2629
rect 11309 -3405 11321 -2629
rect 11263 -3417 11321 -3405
rect 11401 -2629 11459 -2617
rect 11401 -3405 11413 -2629
rect 11447 -3405 11459 -2629
rect 11401 -3417 11459 -3405
rect 11539 -2629 11597 -2617
rect 11539 -3405 11551 -2629
rect 11585 -3405 11597 -2629
rect 11539 -3417 11597 -3405
rect 11677 -2629 11735 -2617
rect 11677 -3405 11689 -2629
rect 11723 -3405 11735 -2629
rect 11677 -3417 11735 -3405
rect 11815 -2629 11873 -2617
rect 11815 -3405 11827 -2629
rect 11861 -3405 11873 -2629
rect 11815 -3417 11873 -3405
rect 11953 -2629 12011 -2617
rect 11953 -3405 11965 -2629
rect 11999 -3405 12011 -2629
rect 11953 -3417 12011 -3405
rect 12091 -2629 12149 -2617
rect 12091 -3405 12103 -2629
rect 12137 -3405 12149 -2629
rect 12091 -3417 12149 -3405
rect 12229 -2629 12287 -2617
rect 12229 -3405 12241 -2629
rect 12275 -3405 12287 -2629
rect 12229 -3417 12287 -3405
rect 12367 -2629 12425 -2617
rect 12367 -3405 12379 -2629
rect 12413 -3405 12425 -2629
rect 12367 -3417 12425 -3405
rect 12505 -2629 12563 -2617
rect 12505 -3405 12517 -2629
rect 12551 -3405 12563 -2629
rect 12505 -3417 12563 -3405
rect 12643 -2629 12701 -2617
rect 12643 -3405 12655 -2629
rect 12689 -3405 12701 -2629
rect 12643 -3417 12701 -3405
rect 12781 -2629 12839 -2617
rect 12781 -3405 12793 -2629
rect 12827 -3405 12839 -2629
rect 12781 -3417 12839 -3405
rect 12919 -2629 12977 -2617
rect 12919 -3405 12931 -2629
rect 12965 -3405 12977 -2629
rect 12919 -3417 12977 -3405
rect 13057 -2629 13115 -2617
rect 13057 -3405 13069 -2629
rect 13103 -3405 13115 -2629
rect 13057 -3417 13115 -3405
rect 13195 -2629 13253 -2617
rect 13195 -3405 13207 -2629
rect 13241 -3405 13253 -2629
rect 13195 -3417 13253 -3405
rect 13333 -2629 13391 -2617
rect 13333 -3405 13345 -2629
rect 13379 -3405 13391 -2629
rect 13333 -3417 13391 -3405
rect 13471 -2629 13529 -2617
rect 13471 -3405 13483 -2629
rect 13517 -3405 13529 -2629
rect 13471 -3417 13529 -3405
rect 13609 -2629 13667 -2617
rect 13609 -3405 13621 -2629
rect 13655 -3405 13667 -2629
rect 13609 -3417 13667 -3405
rect 13747 -2629 13805 -2617
rect 13747 -3405 13759 -2629
rect 13793 -3405 13805 -2629
rect 13747 -3417 13805 -3405
rect 13885 -2629 13943 -2617
rect 13885 -3405 13897 -2629
rect 13931 -3405 13943 -2629
rect 13885 -3417 13943 -3405
<< pdiffc >>
rect 97 -2519 131 -1743
rect 235 -2519 269 -1743
rect 373 -2519 407 -1743
rect 511 -2519 545 -1743
rect 649 -2519 683 -1743
rect 787 -2519 821 -1743
rect 925 -2519 959 -1743
rect 1063 -2519 1097 -1743
rect 1201 -2519 1235 -1743
rect 1339 -2519 1373 -1743
rect 1477 -2519 1511 -1743
rect 1615 -2519 1649 -1743
rect 1753 -2519 1787 -1743
rect 1891 -2519 1925 -1743
rect 2029 -2519 2063 -1743
rect 2167 -2519 2201 -1743
rect 2305 -2519 2339 -1743
rect 2443 -2519 2477 -1743
rect 2581 -2519 2615 -1743
rect 2719 -2519 2753 -1743
rect 2857 -2519 2891 -1743
rect 2995 -2519 3029 -1743
rect 3133 -2519 3167 -1743
rect 3271 -2519 3305 -1743
rect 3409 -2519 3443 -1743
rect 3547 -2519 3581 -1743
rect 3685 -2519 3719 -1743
rect 3823 -2519 3857 -1743
rect 3961 -2519 3995 -1743
rect 4099 -2519 4133 -1743
rect 4237 -2519 4271 -1743
rect 4375 -2519 4409 -1743
rect 4513 -2519 4547 -1743
rect 4651 -2519 4685 -1743
rect 4789 -2519 4823 -1743
rect 4927 -2519 4961 -1743
rect 5065 -2519 5099 -1743
rect 5203 -2519 5237 -1743
rect 5341 -2519 5375 -1743
rect 5479 -2519 5513 -1743
rect 5617 -2519 5651 -1743
rect 5755 -2519 5789 -1743
rect 5893 -2519 5927 -1743
rect 6031 -2519 6065 -1743
rect 6169 -2519 6203 -1743
rect 6307 -2519 6341 -1743
rect 6445 -2519 6479 -1743
rect 6583 -2519 6617 -1743
rect 6721 -2519 6755 -1743
rect 6859 -2519 6893 -1743
rect 6997 -2519 7031 -1743
rect 7135 -2519 7169 -1743
rect 7273 -2519 7307 -1743
rect 7411 -2519 7445 -1743
rect 7549 -2519 7583 -1743
rect 7687 -2519 7721 -1743
rect 7825 -2519 7859 -1743
rect 7963 -2519 7997 -1743
rect 8101 -2519 8135 -1743
rect 8239 -2519 8273 -1743
rect 8377 -2519 8411 -1743
rect 8515 -2519 8549 -1743
rect 8653 -2519 8687 -1743
rect 8791 -2519 8825 -1743
rect 8929 -2519 8963 -1743
rect 9067 -2519 9101 -1743
rect 9205 -2519 9239 -1743
rect 9343 -2519 9377 -1743
rect 9481 -2519 9515 -1743
rect 9619 -2519 9653 -1743
rect 9757 -2519 9791 -1743
rect 9895 -2519 9929 -1743
rect 10033 -2519 10067 -1743
rect 10171 -2519 10205 -1743
rect 10309 -2519 10343 -1743
rect 10447 -2519 10481 -1743
rect 10585 -2519 10619 -1743
rect 10723 -2519 10757 -1743
rect 10861 -2519 10895 -1743
rect 10999 -2519 11033 -1743
rect 11137 -2519 11171 -1743
rect 11275 -2519 11309 -1743
rect 11413 -2519 11447 -1743
rect 11551 -2519 11585 -1743
rect 11689 -2519 11723 -1743
rect 11827 -2519 11861 -1743
rect 11965 -2519 11999 -1743
rect 12103 -2519 12137 -1743
rect 12241 -2519 12275 -1743
rect 12379 -2519 12413 -1743
rect 12517 -2519 12551 -1743
rect 12655 -2519 12689 -1743
rect 12793 -2519 12827 -1743
rect 12931 -2519 12965 -1743
rect 13069 -2519 13103 -1743
rect 13207 -2519 13241 -1743
rect 13345 -2519 13379 -1743
rect 13483 -2519 13517 -1743
rect 13621 -2519 13655 -1743
rect 13759 -2519 13793 -1743
rect 13897 -2519 13931 -1743
rect 97 -3405 131 -2629
rect 235 -3405 269 -2629
rect 373 -3405 407 -2629
rect 511 -3405 545 -2629
rect 649 -3405 683 -2629
rect 787 -3405 821 -2629
rect 925 -3405 959 -2629
rect 1063 -3405 1097 -2629
rect 1201 -3405 1235 -2629
rect 1339 -3405 1373 -2629
rect 1477 -3405 1511 -2629
rect 1615 -3405 1649 -2629
rect 1753 -3405 1787 -2629
rect 1891 -3405 1925 -2629
rect 2029 -3405 2063 -2629
rect 2167 -3405 2201 -2629
rect 2305 -3405 2339 -2629
rect 2443 -3405 2477 -2629
rect 2581 -3405 2615 -2629
rect 2719 -3405 2753 -2629
rect 2857 -3405 2891 -2629
rect 2995 -3405 3029 -2629
rect 3133 -3405 3167 -2629
rect 3271 -3405 3305 -2629
rect 3409 -3405 3443 -2629
rect 3547 -3405 3581 -2629
rect 3685 -3405 3719 -2629
rect 3823 -3405 3857 -2629
rect 3961 -3405 3995 -2629
rect 4099 -3405 4133 -2629
rect 4237 -3405 4271 -2629
rect 4375 -3405 4409 -2629
rect 4513 -3405 4547 -2629
rect 4651 -3405 4685 -2629
rect 4789 -3405 4823 -2629
rect 4927 -3405 4961 -2629
rect 5065 -3405 5099 -2629
rect 5203 -3405 5237 -2629
rect 5341 -3405 5375 -2629
rect 5479 -3405 5513 -2629
rect 5617 -3405 5651 -2629
rect 5755 -3405 5789 -2629
rect 5893 -3405 5927 -2629
rect 6031 -3405 6065 -2629
rect 6169 -3405 6203 -2629
rect 6307 -3405 6341 -2629
rect 6445 -3405 6479 -2629
rect 6583 -3405 6617 -2629
rect 6721 -3405 6755 -2629
rect 6859 -3405 6893 -2629
rect 6997 -3405 7031 -2629
rect 7135 -3405 7169 -2629
rect 7273 -3405 7307 -2629
rect 7411 -3405 7445 -2629
rect 7549 -3405 7583 -2629
rect 7687 -3405 7721 -2629
rect 7825 -3405 7859 -2629
rect 7963 -3405 7997 -2629
rect 8101 -3405 8135 -2629
rect 8239 -3405 8273 -2629
rect 8377 -3405 8411 -2629
rect 8515 -3405 8549 -2629
rect 8653 -3405 8687 -2629
rect 8791 -3405 8825 -2629
rect 8929 -3405 8963 -2629
rect 9067 -3405 9101 -2629
rect 9205 -3405 9239 -2629
rect 9343 -3405 9377 -2629
rect 9481 -3405 9515 -2629
rect 9619 -3405 9653 -2629
rect 9757 -3405 9791 -2629
rect 9895 -3405 9929 -2629
rect 10033 -3405 10067 -2629
rect 10171 -3405 10205 -2629
rect 10309 -3405 10343 -2629
rect 10447 -3405 10481 -2629
rect 10585 -3405 10619 -2629
rect 10723 -3405 10757 -2629
rect 10861 -3405 10895 -2629
rect 10999 -3405 11033 -2629
rect 11137 -3405 11171 -2629
rect 11275 -3405 11309 -2629
rect 11413 -3405 11447 -2629
rect 11551 -3405 11585 -2629
rect 11689 -3405 11723 -2629
rect 11827 -3405 11861 -2629
rect 11965 -3405 11999 -2629
rect 12103 -3405 12137 -2629
rect 12241 -3405 12275 -2629
rect 12379 -3405 12413 -2629
rect 12517 -3405 12551 -2629
rect 12655 -3405 12689 -2629
rect 12793 -3405 12827 -2629
rect 12931 -3405 12965 -2629
rect 13069 -3405 13103 -2629
rect 13207 -3405 13241 -2629
rect 13345 -3405 13379 -2629
rect 13483 -3405 13517 -2629
rect 13621 -3405 13655 -2629
rect 13759 -3405 13793 -2629
rect 13897 -3405 13931 -2629
<< nsubdiff >>
rect -12 1023 84 1057
rect 13943 1023 14039 1057
rect -12 961 22 1023
rect 14005 961 14039 1023
rect -12 -874 22 -812
rect 14005 -874 14039 -812
rect -12 -908 84 -874
rect 13943 -908 14039 -874
rect -900 -1551 -876 -970
rect 14374 -1551 14398 -970
rect -12 -1644 84 -1610
rect 13943 -1644 14039 -1610
rect -12 -1706 22 -1644
rect 14005 -1706 14039 -1644
rect -12 -3541 22 -3479
rect 14005 -3541 14039 -3479
rect -12 -3575 84 -3541
rect 13943 -3575 14039 -3541
<< nsubdiffcont >>
rect 84 1023 13943 1057
rect -12 -812 22 961
rect 14005 -812 14039 961
rect 84 -908 13943 -874
rect -876 -1551 14374 -970
rect 84 -1644 13943 -1610
rect -12 -3479 22 -1706
rect 14005 -3479 14039 -1706
rect 84 -3575 13943 -3541
<< poly >>
rect 143 38 13885 74
rect 143 -1731 223 -1705
rect 281 -1731 361 -1705
rect 419 -1731 499 -1705
rect 557 -1731 637 -1705
rect 695 -1731 775 -1705
rect 833 -1731 913 -1705
rect 971 -1731 1051 -1705
rect 1109 -1731 1189 -1705
rect 1247 -1731 1327 -1705
rect 1385 -1731 1465 -1705
rect 1523 -1731 1603 -1705
rect 1661 -1731 1741 -1705
rect 1799 -1731 1879 -1705
rect 1937 -1731 2017 -1705
rect 2075 -1731 2155 -1705
rect 2213 -1731 2293 -1705
rect 2351 -1731 2431 -1705
rect 2489 -1731 2569 -1705
rect 2627 -1731 2707 -1705
rect 2765 -1731 2845 -1705
rect 2903 -1731 2983 -1705
rect 3041 -1731 3121 -1705
rect 3179 -1731 3259 -1705
rect 3317 -1731 3397 -1705
rect 3455 -1731 3535 -1705
rect 3593 -1731 3673 -1705
rect 3731 -1731 3811 -1705
rect 3869 -1731 3949 -1705
rect 4007 -1731 4087 -1705
rect 4145 -1731 4225 -1705
rect 4283 -1731 4363 -1705
rect 4421 -1731 4501 -1705
rect 4559 -1731 4639 -1705
rect 4697 -1731 4777 -1705
rect 4835 -1731 4915 -1705
rect 4973 -1731 5053 -1705
rect 5111 -1731 5191 -1705
rect 5249 -1731 5329 -1705
rect 5387 -1731 5467 -1705
rect 5525 -1731 5605 -1705
rect 5663 -1731 5743 -1705
rect 5801 -1731 5881 -1705
rect 5939 -1731 6019 -1705
rect 6077 -1731 6157 -1705
rect 6215 -1731 6295 -1705
rect 6353 -1731 6433 -1705
rect 6491 -1731 6571 -1705
rect 6629 -1731 6709 -1705
rect 6767 -1731 6847 -1705
rect 6905 -1731 6985 -1705
rect 7043 -1731 7123 -1705
rect 7181 -1731 7261 -1705
rect 7319 -1731 7399 -1705
rect 7457 -1731 7537 -1705
rect 7595 -1731 7675 -1705
rect 7733 -1731 7813 -1705
rect 7871 -1731 7951 -1705
rect 8009 -1731 8089 -1705
rect 8147 -1731 8227 -1705
rect 8285 -1731 8365 -1705
rect 8423 -1731 8503 -1705
rect 8561 -1731 8641 -1705
rect 8699 -1731 8779 -1705
rect 8837 -1731 8917 -1705
rect 8975 -1731 9055 -1705
rect 9113 -1731 9193 -1705
rect 9251 -1731 9331 -1705
rect 9389 -1731 9469 -1705
rect 9527 -1731 9607 -1705
rect 9665 -1731 9745 -1705
rect 9803 -1731 9883 -1705
rect 9941 -1731 10021 -1705
rect 10079 -1731 10159 -1705
rect 10217 -1731 10297 -1705
rect 10355 -1731 10435 -1705
rect 10493 -1731 10573 -1705
rect 10631 -1731 10711 -1705
rect 10769 -1731 10849 -1705
rect 10907 -1731 10987 -1705
rect 11045 -1731 11125 -1705
rect 11183 -1731 11263 -1705
rect 11321 -1731 11401 -1705
rect 11459 -1731 11539 -1705
rect 11597 -1731 11677 -1705
rect 11735 -1731 11815 -1705
rect 11873 -1731 11953 -1705
rect 12011 -1731 12091 -1705
rect 12149 -1731 12229 -1705
rect 12287 -1731 12367 -1705
rect 12425 -1731 12505 -1705
rect 12563 -1731 12643 -1705
rect 12701 -1731 12781 -1705
rect 12839 -1731 12919 -1705
rect 12977 -1731 13057 -1705
rect 13115 -1731 13195 -1705
rect 13253 -1731 13333 -1705
rect 13391 -1731 13471 -1705
rect 13529 -1731 13609 -1705
rect 13667 -1731 13747 -1705
rect 13805 -1731 13885 -1705
rect 143 -2556 223 -2531
rect 281 -2556 361 -2531
rect 419 -2556 499 -2531
rect 557 -2556 637 -2531
rect 695 -2556 775 -2531
rect 833 -2556 913 -2531
rect 971 -2556 1051 -2531
rect 1109 -2556 1189 -2531
rect 1247 -2556 1327 -2531
rect 1385 -2556 1465 -2531
rect 1523 -2556 1603 -2531
rect 1661 -2556 1741 -2531
rect 1799 -2556 1879 -2531
rect 1937 -2556 2017 -2531
rect 2075 -2556 2155 -2531
rect 2213 -2556 2293 -2531
rect 2351 -2556 2431 -2531
rect 2489 -2556 2569 -2531
rect 2627 -2556 2707 -2531
rect 2765 -2556 2845 -2531
rect 2903 -2556 2983 -2531
rect 3041 -2556 3121 -2531
rect 3179 -2556 3259 -2531
rect 3317 -2556 3397 -2531
rect 3455 -2556 3535 -2531
rect 3593 -2556 3673 -2531
rect 3731 -2556 3811 -2531
rect 3869 -2556 3949 -2531
rect 4007 -2556 4087 -2531
rect 4145 -2556 4225 -2531
rect 4283 -2556 4363 -2531
rect 4421 -2556 4501 -2531
rect 4559 -2556 4639 -2531
rect 4697 -2556 4777 -2531
rect 4835 -2556 4915 -2531
rect 4973 -2556 5053 -2531
rect 5111 -2556 5191 -2531
rect 5249 -2556 5329 -2531
rect 5387 -2556 5467 -2531
rect 5525 -2556 5605 -2531
rect 5663 -2556 5743 -2531
rect 5801 -2556 5881 -2531
rect 5939 -2556 6019 -2531
rect 6077 -2556 6157 -2531
rect 6215 -2556 6295 -2531
rect 6353 -2556 6433 -2531
rect 6491 -2556 6571 -2531
rect 6629 -2556 6709 -2531
rect 6767 -2556 6847 -2531
rect 6905 -2556 6985 -2531
rect 7043 -2556 7123 -2531
rect 7181 -2556 7261 -2531
rect 7319 -2556 7399 -2531
rect 7457 -2556 7537 -2531
rect 7595 -2556 7675 -2531
rect 7733 -2556 7813 -2531
rect 7871 -2556 7951 -2531
rect 8009 -2556 8089 -2531
rect 8147 -2556 8227 -2531
rect 8285 -2556 8365 -2531
rect 8423 -2556 8503 -2531
rect 8561 -2556 8641 -2531
rect 8699 -2556 8779 -2531
rect 8837 -2556 8917 -2531
rect 8975 -2556 9055 -2531
rect 9113 -2556 9193 -2531
rect 9251 -2556 9331 -2531
rect 9389 -2556 9469 -2531
rect 9527 -2556 9607 -2531
rect 9665 -2556 9745 -2531
rect 9803 -2556 9883 -2531
rect 9941 -2556 10021 -2531
rect 10079 -2556 10159 -2531
rect 10217 -2556 10297 -2531
rect 10355 -2556 10435 -2531
rect 10493 -2556 10573 -2531
rect 10631 -2556 10711 -2531
rect 10769 -2556 10849 -2531
rect 10907 -2556 10987 -2531
rect 11045 -2556 11125 -2531
rect 11183 -2556 11263 -2531
rect 11321 -2556 11401 -2531
rect 11459 -2556 11539 -2531
rect 11597 -2556 11677 -2531
rect 11735 -2556 11815 -2531
rect 11873 -2556 11953 -2531
rect 12011 -2556 12091 -2531
rect 12149 -2556 12229 -2531
rect 12287 -2556 12367 -2531
rect 12425 -2556 12505 -2531
rect 12563 -2556 12643 -2531
rect 12701 -2556 12781 -2531
rect 12839 -2556 12919 -2531
rect 12977 -2556 13057 -2531
rect 13115 -2556 13195 -2531
rect 13253 -2556 13333 -2531
rect 13391 -2556 13471 -2531
rect 13529 -2556 13609 -2531
rect 13667 -2556 13747 -2531
rect 13805 -2556 13885 -2531
rect 143 -2592 13885 -2556
rect 143 -2617 223 -2592
rect 281 -2617 361 -2592
rect 419 -2617 499 -2592
rect 557 -2617 637 -2592
rect 695 -2617 775 -2592
rect 833 -2617 913 -2592
rect 971 -2617 1051 -2592
rect 1109 -2617 1189 -2592
rect 1247 -2617 1327 -2592
rect 1385 -2617 1465 -2592
rect 1523 -2617 1603 -2592
rect 1661 -2617 1741 -2592
rect 1799 -2617 1879 -2592
rect 1937 -2617 2017 -2592
rect 2075 -2617 2155 -2592
rect 2213 -2617 2293 -2592
rect 2351 -2617 2431 -2592
rect 2489 -2617 2569 -2592
rect 2627 -2617 2707 -2592
rect 2765 -2617 2845 -2592
rect 2903 -2617 2983 -2592
rect 3041 -2617 3121 -2592
rect 3179 -2617 3259 -2592
rect 3317 -2617 3397 -2592
rect 3455 -2617 3535 -2592
rect 3593 -2617 3673 -2592
rect 3731 -2617 3811 -2592
rect 3869 -2617 3949 -2592
rect 4007 -2617 4087 -2592
rect 4145 -2617 4225 -2592
rect 4283 -2617 4363 -2592
rect 4421 -2617 4501 -2592
rect 4559 -2617 4639 -2592
rect 4697 -2617 4777 -2592
rect 4835 -2617 4915 -2592
rect 4973 -2617 5053 -2592
rect 5111 -2617 5191 -2592
rect 5249 -2617 5329 -2592
rect 5387 -2617 5467 -2592
rect 5525 -2617 5605 -2592
rect 5663 -2617 5743 -2592
rect 5801 -2617 5881 -2592
rect 5939 -2617 6019 -2592
rect 6077 -2617 6157 -2592
rect 6215 -2617 6295 -2592
rect 6353 -2617 6433 -2592
rect 6491 -2617 6571 -2592
rect 6629 -2617 6709 -2592
rect 6767 -2617 6847 -2592
rect 6905 -2617 6985 -2592
rect 7043 -2617 7123 -2592
rect 7181 -2617 7261 -2592
rect 7319 -2617 7399 -2592
rect 7457 -2617 7537 -2592
rect 7595 -2617 7675 -2592
rect 7733 -2617 7813 -2592
rect 7871 -2617 7951 -2592
rect 8009 -2617 8089 -2592
rect 8147 -2617 8227 -2592
rect 8285 -2617 8365 -2592
rect 8423 -2617 8503 -2592
rect 8561 -2617 8641 -2592
rect 8699 -2617 8779 -2592
rect 8837 -2617 8917 -2592
rect 8975 -2617 9055 -2592
rect 9113 -2617 9193 -2592
rect 9251 -2617 9331 -2592
rect 9389 -2617 9469 -2592
rect 9527 -2617 9607 -2592
rect 9665 -2617 9745 -2592
rect 9803 -2617 9883 -2592
rect 9941 -2617 10021 -2592
rect 10079 -2617 10159 -2592
rect 10217 -2617 10297 -2592
rect 10355 -2617 10435 -2592
rect 10493 -2617 10573 -2592
rect 10631 -2617 10711 -2592
rect 10769 -2617 10849 -2592
rect 10907 -2617 10987 -2592
rect 11045 -2617 11125 -2592
rect 11183 -2617 11263 -2592
rect 11321 -2617 11401 -2592
rect 11459 -2617 11539 -2592
rect 11597 -2617 11677 -2592
rect 11735 -2617 11815 -2592
rect 11873 -2617 11953 -2592
rect 12011 -2617 12091 -2592
rect 12149 -2617 12229 -2592
rect 12287 -2617 12367 -2592
rect 12425 -2617 12505 -2592
rect 12563 -2617 12643 -2592
rect 12701 -2617 12781 -2592
rect 12839 -2617 12919 -2592
rect 12977 -2617 13057 -2592
rect 13115 -2617 13195 -2592
rect 13253 -2617 13333 -2592
rect 13391 -2617 13471 -2592
rect 13529 -2617 13609 -2592
rect 13667 -2617 13747 -2592
rect 13805 -2617 13885 -2592
rect 143 -3464 223 -3417
rect 143 -3498 159 -3464
rect 207 -3498 223 -3464
rect 143 -3514 223 -3498
rect 281 -3464 361 -3417
rect 281 -3498 297 -3464
rect 345 -3498 361 -3464
rect 281 -3514 361 -3498
rect 419 -3464 499 -3417
rect 419 -3498 435 -3464
rect 483 -3498 499 -3464
rect 419 -3514 499 -3498
rect 557 -3464 637 -3417
rect 557 -3498 573 -3464
rect 621 -3498 637 -3464
rect 557 -3514 637 -3498
rect 695 -3464 775 -3417
rect 695 -3498 711 -3464
rect 759 -3498 775 -3464
rect 695 -3514 775 -3498
rect 833 -3464 913 -3417
rect 833 -3498 849 -3464
rect 897 -3498 913 -3464
rect 833 -3514 913 -3498
rect 971 -3464 1051 -3417
rect 971 -3498 987 -3464
rect 1035 -3498 1051 -3464
rect 971 -3514 1051 -3498
rect 1109 -3464 1189 -3417
rect 1109 -3498 1125 -3464
rect 1173 -3498 1189 -3464
rect 1109 -3514 1189 -3498
rect 1247 -3464 1327 -3417
rect 1247 -3498 1263 -3464
rect 1311 -3498 1327 -3464
rect 1247 -3514 1327 -3498
rect 1385 -3464 1465 -3417
rect 1385 -3498 1401 -3464
rect 1449 -3498 1465 -3464
rect 1385 -3514 1465 -3498
rect 1523 -3464 1603 -3417
rect 1523 -3498 1539 -3464
rect 1587 -3498 1603 -3464
rect 1523 -3514 1603 -3498
rect 1661 -3464 1741 -3417
rect 1661 -3498 1677 -3464
rect 1725 -3498 1741 -3464
rect 1661 -3514 1741 -3498
rect 1799 -3464 1879 -3417
rect 1799 -3498 1815 -3464
rect 1863 -3498 1879 -3464
rect 1799 -3514 1879 -3498
rect 1937 -3464 2017 -3417
rect 1937 -3498 1953 -3464
rect 2001 -3498 2017 -3464
rect 1937 -3514 2017 -3498
rect 2075 -3464 2155 -3417
rect 2075 -3498 2091 -3464
rect 2139 -3498 2155 -3464
rect 2075 -3514 2155 -3498
rect 2213 -3464 2293 -3417
rect 2213 -3498 2229 -3464
rect 2277 -3498 2293 -3464
rect 2213 -3514 2293 -3498
rect 2351 -3464 2431 -3417
rect 2351 -3498 2367 -3464
rect 2415 -3498 2431 -3464
rect 2351 -3514 2431 -3498
rect 2489 -3464 2569 -3417
rect 2489 -3498 2505 -3464
rect 2553 -3498 2569 -3464
rect 2489 -3514 2569 -3498
rect 2627 -3464 2707 -3417
rect 2627 -3498 2643 -3464
rect 2691 -3498 2707 -3464
rect 2627 -3514 2707 -3498
rect 2765 -3464 2845 -3417
rect 2765 -3498 2781 -3464
rect 2829 -3498 2845 -3464
rect 2765 -3514 2845 -3498
rect 2903 -3464 2983 -3417
rect 2903 -3498 2919 -3464
rect 2967 -3498 2983 -3464
rect 2903 -3514 2983 -3498
rect 3041 -3464 3121 -3417
rect 3041 -3498 3057 -3464
rect 3105 -3498 3121 -3464
rect 3041 -3514 3121 -3498
rect 3179 -3464 3259 -3417
rect 3179 -3498 3195 -3464
rect 3243 -3498 3259 -3464
rect 3179 -3514 3259 -3498
rect 3317 -3464 3397 -3417
rect 3317 -3498 3333 -3464
rect 3381 -3498 3397 -3464
rect 3317 -3514 3397 -3498
rect 3455 -3464 3535 -3417
rect 3455 -3498 3471 -3464
rect 3519 -3498 3535 -3464
rect 3455 -3514 3535 -3498
rect 3593 -3464 3673 -3417
rect 3593 -3498 3609 -3464
rect 3657 -3498 3673 -3464
rect 3593 -3514 3673 -3498
rect 3731 -3464 3811 -3417
rect 3731 -3498 3747 -3464
rect 3795 -3498 3811 -3464
rect 3731 -3514 3811 -3498
rect 3869 -3464 3949 -3417
rect 3869 -3498 3885 -3464
rect 3933 -3498 3949 -3464
rect 3869 -3514 3949 -3498
rect 4007 -3464 4087 -3417
rect 4007 -3498 4023 -3464
rect 4071 -3498 4087 -3464
rect 4007 -3514 4087 -3498
rect 4145 -3464 4225 -3417
rect 4145 -3498 4161 -3464
rect 4209 -3498 4225 -3464
rect 4145 -3514 4225 -3498
rect 4283 -3464 4363 -3417
rect 4283 -3498 4299 -3464
rect 4347 -3498 4363 -3464
rect 4283 -3514 4363 -3498
rect 4421 -3464 4501 -3417
rect 4421 -3498 4437 -3464
rect 4485 -3498 4501 -3464
rect 4421 -3514 4501 -3498
rect 4559 -3464 4639 -3417
rect 4559 -3498 4575 -3464
rect 4623 -3498 4639 -3464
rect 4559 -3514 4639 -3498
rect 4697 -3464 4777 -3417
rect 4697 -3498 4713 -3464
rect 4761 -3498 4777 -3464
rect 4697 -3514 4777 -3498
rect 4835 -3464 4915 -3417
rect 4835 -3498 4851 -3464
rect 4899 -3498 4915 -3464
rect 4835 -3514 4915 -3498
rect 4973 -3464 5053 -3417
rect 4973 -3498 4989 -3464
rect 5037 -3498 5053 -3464
rect 4973 -3514 5053 -3498
rect 5111 -3464 5191 -3417
rect 5111 -3498 5127 -3464
rect 5175 -3498 5191 -3464
rect 5111 -3514 5191 -3498
rect 5249 -3464 5329 -3417
rect 5249 -3498 5265 -3464
rect 5313 -3498 5329 -3464
rect 5249 -3514 5329 -3498
rect 5387 -3464 5467 -3417
rect 5387 -3498 5403 -3464
rect 5451 -3498 5467 -3464
rect 5387 -3514 5467 -3498
rect 5525 -3464 5605 -3417
rect 5525 -3498 5541 -3464
rect 5589 -3498 5605 -3464
rect 5525 -3514 5605 -3498
rect 5663 -3464 5743 -3417
rect 5663 -3498 5679 -3464
rect 5727 -3498 5743 -3464
rect 5663 -3514 5743 -3498
rect 5801 -3464 5881 -3417
rect 5801 -3498 5817 -3464
rect 5865 -3498 5881 -3464
rect 5801 -3514 5881 -3498
rect 5939 -3464 6019 -3417
rect 5939 -3498 5955 -3464
rect 6003 -3498 6019 -3464
rect 5939 -3514 6019 -3498
rect 6077 -3464 6157 -3417
rect 6077 -3498 6093 -3464
rect 6141 -3498 6157 -3464
rect 6077 -3514 6157 -3498
rect 6215 -3464 6295 -3417
rect 6215 -3498 6231 -3464
rect 6279 -3498 6295 -3464
rect 6215 -3514 6295 -3498
rect 6353 -3464 6433 -3417
rect 6353 -3498 6369 -3464
rect 6417 -3498 6433 -3464
rect 6353 -3514 6433 -3498
rect 6491 -3464 6571 -3417
rect 6491 -3498 6507 -3464
rect 6555 -3498 6571 -3464
rect 6491 -3514 6571 -3498
rect 6629 -3464 6709 -3417
rect 6629 -3498 6645 -3464
rect 6693 -3498 6709 -3464
rect 6629 -3514 6709 -3498
rect 6767 -3464 6847 -3417
rect 6767 -3498 6783 -3464
rect 6831 -3498 6847 -3464
rect 6767 -3514 6847 -3498
rect 6905 -3464 6985 -3417
rect 6905 -3498 6921 -3464
rect 6969 -3498 6985 -3464
rect 6905 -3514 6985 -3498
rect 7043 -3464 7123 -3417
rect 7043 -3498 7059 -3464
rect 7107 -3498 7123 -3464
rect 7043 -3514 7123 -3498
rect 7181 -3464 7261 -3417
rect 7181 -3498 7197 -3464
rect 7245 -3498 7261 -3464
rect 7181 -3514 7261 -3498
rect 7319 -3464 7399 -3417
rect 7319 -3498 7335 -3464
rect 7383 -3498 7399 -3464
rect 7319 -3514 7399 -3498
rect 7457 -3464 7537 -3417
rect 7457 -3498 7473 -3464
rect 7521 -3498 7537 -3464
rect 7457 -3514 7537 -3498
rect 7595 -3464 7675 -3417
rect 7595 -3498 7611 -3464
rect 7659 -3498 7675 -3464
rect 7595 -3514 7675 -3498
rect 7733 -3464 7813 -3417
rect 7733 -3498 7749 -3464
rect 7797 -3498 7813 -3464
rect 7733 -3514 7813 -3498
rect 7871 -3464 7951 -3417
rect 7871 -3498 7887 -3464
rect 7935 -3498 7951 -3464
rect 7871 -3514 7951 -3498
rect 8009 -3464 8089 -3417
rect 8009 -3498 8025 -3464
rect 8073 -3498 8089 -3464
rect 8009 -3514 8089 -3498
rect 8147 -3464 8227 -3417
rect 8147 -3498 8163 -3464
rect 8211 -3498 8227 -3464
rect 8147 -3514 8227 -3498
rect 8285 -3464 8365 -3417
rect 8285 -3498 8301 -3464
rect 8349 -3498 8365 -3464
rect 8285 -3514 8365 -3498
rect 8423 -3464 8503 -3417
rect 8423 -3498 8439 -3464
rect 8487 -3498 8503 -3464
rect 8423 -3514 8503 -3498
rect 8561 -3464 8641 -3417
rect 8561 -3498 8577 -3464
rect 8625 -3498 8641 -3464
rect 8561 -3514 8641 -3498
rect 8699 -3464 8779 -3417
rect 8699 -3498 8715 -3464
rect 8763 -3498 8779 -3464
rect 8699 -3514 8779 -3498
rect 8837 -3464 8917 -3417
rect 8837 -3498 8853 -3464
rect 8901 -3498 8917 -3464
rect 8837 -3514 8917 -3498
rect 8975 -3464 9055 -3417
rect 8975 -3498 8991 -3464
rect 9039 -3498 9055 -3464
rect 8975 -3514 9055 -3498
rect 9113 -3464 9193 -3417
rect 9113 -3498 9129 -3464
rect 9177 -3498 9193 -3464
rect 9113 -3514 9193 -3498
rect 9251 -3464 9331 -3417
rect 9251 -3498 9267 -3464
rect 9315 -3498 9331 -3464
rect 9251 -3514 9331 -3498
rect 9389 -3464 9469 -3417
rect 9389 -3498 9405 -3464
rect 9453 -3498 9469 -3464
rect 9389 -3514 9469 -3498
rect 9527 -3464 9607 -3417
rect 9527 -3498 9543 -3464
rect 9591 -3498 9607 -3464
rect 9527 -3514 9607 -3498
rect 9665 -3464 9745 -3417
rect 9665 -3498 9681 -3464
rect 9729 -3498 9745 -3464
rect 9665 -3514 9745 -3498
rect 9803 -3464 9883 -3417
rect 9803 -3498 9819 -3464
rect 9867 -3498 9883 -3464
rect 9803 -3514 9883 -3498
rect 9941 -3464 10021 -3417
rect 9941 -3498 9957 -3464
rect 10005 -3498 10021 -3464
rect 9941 -3514 10021 -3498
rect 10079 -3464 10159 -3417
rect 10079 -3498 10095 -3464
rect 10143 -3498 10159 -3464
rect 10079 -3514 10159 -3498
rect 10217 -3464 10297 -3417
rect 10217 -3498 10233 -3464
rect 10281 -3498 10297 -3464
rect 10217 -3514 10297 -3498
rect 10355 -3464 10435 -3417
rect 10355 -3498 10371 -3464
rect 10419 -3498 10435 -3464
rect 10355 -3514 10435 -3498
rect 10493 -3464 10573 -3417
rect 10493 -3498 10509 -3464
rect 10557 -3498 10573 -3464
rect 10493 -3514 10573 -3498
rect 10631 -3464 10711 -3417
rect 10631 -3498 10647 -3464
rect 10695 -3498 10711 -3464
rect 10631 -3514 10711 -3498
rect 10769 -3464 10849 -3417
rect 10769 -3498 10785 -3464
rect 10833 -3498 10849 -3464
rect 10769 -3514 10849 -3498
rect 10907 -3464 10987 -3417
rect 10907 -3498 10923 -3464
rect 10971 -3498 10987 -3464
rect 10907 -3514 10987 -3498
rect 11045 -3464 11125 -3417
rect 11045 -3498 11061 -3464
rect 11109 -3498 11125 -3464
rect 11045 -3514 11125 -3498
rect 11183 -3464 11263 -3417
rect 11183 -3498 11199 -3464
rect 11247 -3498 11263 -3464
rect 11183 -3514 11263 -3498
rect 11321 -3464 11401 -3417
rect 11321 -3498 11337 -3464
rect 11385 -3498 11401 -3464
rect 11321 -3514 11401 -3498
rect 11459 -3464 11539 -3417
rect 11459 -3498 11475 -3464
rect 11523 -3498 11539 -3464
rect 11459 -3514 11539 -3498
rect 11597 -3464 11677 -3417
rect 11597 -3498 11613 -3464
rect 11661 -3498 11677 -3464
rect 11597 -3514 11677 -3498
rect 11735 -3464 11815 -3417
rect 11735 -3498 11751 -3464
rect 11799 -3498 11815 -3464
rect 11735 -3514 11815 -3498
rect 11873 -3464 11953 -3417
rect 11873 -3498 11889 -3464
rect 11937 -3498 11953 -3464
rect 11873 -3514 11953 -3498
rect 12011 -3464 12091 -3417
rect 12011 -3498 12027 -3464
rect 12075 -3498 12091 -3464
rect 12011 -3514 12091 -3498
rect 12149 -3464 12229 -3417
rect 12149 -3498 12165 -3464
rect 12213 -3498 12229 -3464
rect 12149 -3514 12229 -3498
rect 12287 -3464 12367 -3417
rect 12287 -3498 12303 -3464
rect 12351 -3498 12367 -3464
rect 12287 -3514 12367 -3498
rect 12425 -3464 12505 -3417
rect 12425 -3498 12441 -3464
rect 12489 -3498 12505 -3464
rect 12425 -3514 12505 -3498
rect 12563 -3464 12643 -3417
rect 12563 -3498 12579 -3464
rect 12627 -3498 12643 -3464
rect 12563 -3514 12643 -3498
rect 12701 -3464 12781 -3417
rect 12701 -3498 12717 -3464
rect 12765 -3498 12781 -3464
rect 12701 -3514 12781 -3498
rect 12839 -3464 12919 -3417
rect 12839 -3498 12855 -3464
rect 12903 -3498 12919 -3464
rect 12839 -3514 12919 -3498
rect 12977 -3464 13057 -3417
rect 12977 -3498 12993 -3464
rect 13041 -3498 13057 -3464
rect 12977 -3514 13057 -3498
rect 13115 -3464 13195 -3417
rect 13115 -3498 13131 -3464
rect 13179 -3498 13195 -3464
rect 13115 -3514 13195 -3498
rect 13253 -3464 13333 -3417
rect 13253 -3498 13269 -3464
rect 13317 -3498 13333 -3464
rect 13253 -3514 13333 -3498
rect 13391 -3464 13471 -3417
rect 13391 -3498 13407 -3464
rect 13455 -3498 13471 -3464
rect 13391 -3514 13471 -3498
rect 13529 -3464 13609 -3417
rect 13529 -3498 13545 -3464
rect 13593 -3498 13609 -3464
rect 13529 -3514 13609 -3498
rect 13667 -3464 13747 -3417
rect 13667 -3498 13683 -3464
rect 13731 -3498 13747 -3464
rect 13667 -3514 13747 -3498
rect 13805 -3464 13885 -3417
rect 13805 -3498 13821 -3464
rect 13869 -3498 13885 -3464
rect 13805 -3514 13885 -3498
<< polycont >>
rect 159 -3498 207 -3464
rect 297 -3498 345 -3464
rect 435 -3498 483 -3464
rect 573 -3498 621 -3464
rect 711 -3498 759 -3464
rect 849 -3498 897 -3464
rect 987 -3498 1035 -3464
rect 1125 -3498 1173 -3464
rect 1263 -3498 1311 -3464
rect 1401 -3498 1449 -3464
rect 1539 -3498 1587 -3464
rect 1677 -3498 1725 -3464
rect 1815 -3498 1863 -3464
rect 1953 -3498 2001 -3464
rect 2091 -3498 2139 -3464
rect 2229 -3498 2277 -3464
rect 2367 -3498 2415 -3464
rect 2505 -3498 2553 -3464
rect 2643 -3498 2691 -3464
rect 2781 -3498 2829 -3464
rect 2919 -3498 2967 -3464
rect 3057 -3498 3105 -3464
rect 3195 -3498 3243 -3464
rect 3333 -3498 3381 -3464
rect 3471 -3498 3519 -3464
rect 3609 -3498 3657 -3464
rect 3747 -3498 3795 -3464
rect 3885 -3498 3933 -3464
rect 4023 -3498 4071 -3464
rect 4161 -3498 4209 -3464
rect 4299 -3498 4347 -3464
rect 4437 -3498 4485 -3464
rect 4575 -3498 4623 -3464
rect 4713 -3498 4761 -3464
rect 4851 -3498 4899 -3464
rect 4989 -3498 5037 -3464
rect 5127 -3498 5175 -3464
rect 5265 -3498 5313 -3464
rect 5403 -3498 5451 -3464
rect 5541 -3498 5589 -3464
rect 5679 -3498 5727 -3464
rect 5817 -3498 5865 -3464
rect 5955 -3498 6003 -3464
rect 6093 -3498 6141 -3464
rect 6231 -3498 6279 -3464
rect 6369 -3498 6417 -3464
rect 6507 -3498 6555 -3464
rect 6645 -3498 6693 -3464
rect 6783 -3498 6831 -3464
rect 6921 -3498 6969 -3464
rect 7059 -3498 7107 -3464
rect 7197 -3498 7245 -3464
rect 7335 -3498 7383 -3464
rect 7473 -3498 7521 -3464
rect 7611 -3498 7659 -3464
rect 7749 -3498 7797 -3464
rect 7887 -3498 7935 -3464
rect 8025 -3498 8073 -3464
rect 8163 -3498 8211 -3464
rect 8301 -3498 8349 -3464
rect 8439 -3498 8487 -3464
rect 8577 -3498 8625 -3464
rect 8715 -3498 8763 -3464
rect 8853 -3498 8901 -3464
rect 8991 -3498 9039 -3464
rect 9129 -3498 9177 -3464
rect 9267 -3498 9315 -3464
rect 9405 -3498 9453 -3464
rect 9543 -3498 9591 -3464
rect 9681 -3498 9729 -3464
rect 9819 -3498 9867 -3464
rect 9957 -3498 10005 -3464
rect 10095 -3498 10143 -3464
rect 10233 -3498 10281 -3464
rect 10371 -3498 10419 -3464
rect 10509 -3498 10557 -3464
rect 10647 -3498 10695 -3464
rect 10785 -3498 10833 -3464
rect 10923 -3498 10971 -3464
rect 11061 -3498 11109 -3464
rect 11199 -3498 11247 -3464
rect 11337 -3498 11385 -3464
rect 11475 -3498 11523 -3464
rect 11613 -3498 11661 -3464
rect 11751 -3498 11799 -3464
rect 11889 -3498 11937 -3464
rect 12027 -3498 12075 -3464
rect 12165 -3498 12213 -3464
rect 12303 -3498 12351 -3464
rect 12441 -3498 12489 -3464
rect 12579 -3498 12627 -3464
rect 12717 -3498 12765 -3464
rect 12855 -3498 12903 -3464
rect 12993 -3498 13041 -3464
rect 13131 -3498 13179 -3464
rect 13269 -3498 13317 -3464
rect 13407 -3498 13455 -3464
rect 13545 -3498 13593 -3464
rect 13683 -3498 13731 -3464
rect 13821 -3498 13869 -3464
<< locali >>
rect -12 1023 84 1057
rect 13943 1023 14039 1057
rect -12 961 22 1023
rect -12 -874 22 -812
rect 14005 961 14039 1023
rect 14005 -874 14039 -812
rect -12 -908 84 -874
rect 13943 -908 14039 -874
rect -892 -1551 -876 -970
rect 14374 -1551 14390 -970
rect -12 -1644 84 -1610
rect 13943 -1644 14039 -1610
rect -12 -1706 22 -1644
rect 14005 -1706 14039 -1644
rect 97 -1743 131 -1727
rect 97 -2535 131 -2519
rect 235 -1743 269 -1727
rect 235 -2535 269 -2519
rect 373 -1743 407 -1727
rect 373 -2535 407 -2519
rect 511 -1743 545 -1727
rect 511 -2535 545 -2519
rect 649 -1743 683 -1727
rect 649 -2535 683 -2519
rect 787 -1743 821 -1727
rect 787 -2535 821 -2519
rect 925 -1743 959 -1727
rect 925 -2535 959 -2519
rect 1063 -1743 1097 -1727
rect 1063 -2535 1097 -2519
rect 1201 -1743 1235 -1727
rect 1201 -2535 1235 -2519
rect 1339 -1743 1373 -1727
rect 1339 -2535 1373 -2519
rect 1477 -1743 1511 -1727
rect 1477 -2535 1511 -2519
rect 1615 -1743 1649 -1727
rect 1615 -2535 1649 -2519
rect 1753 -1743 1787 -1727
rect 1753 -2535 1787 -2519
rect 1891 -1743 1925 -1727
rect 1891 -2535 1925 -2519
rect 2029 -1743 2063 -1727
rect 2029 -2535 2063 -2519
rect 2167 -1743 2201 -1727
rect 2167 -2535 2201 -2519
rect 2305 -1743 2339 -1727
rect 2305 -2535 2339 -2519
rect 2443 -1743 2477 -1727
rect 2443 -2535 2477 -2519
rect 2581 -1743 2615 -1727
rect 2581 -2535 2615 -2519
rect 2719 -1743 2753 -1727
rect 2719 -2535 2753 -2519
rect 2857 -1743 2891 -1727
rect 2857 -2535 2891 -2519
rect 2995 -1743 3029 -1727
rect 2995 -2535 3029 -2519
rect 3133 -1743 3167 -1727
rect 3133 -2535 3167 -2519
rect 3271 -1743 3305 -1727
rect 3271 -2535 3305 -2519
rect 3409 -1743 3443 -1727
rect 3409 -2535 3443 -2519
rect 3547 -1743 3581 -1727
rect 3547 -2535 3581 -2519
rect 3685 -1743 3719 -1727
rect 3685 -2535 3719 -2519
rect 3823 -1743 3857 -1727
rect 3823 -2535 3857 -2519
rect 3961 -1743 3995 -1727
rect 3961 -2535 3995 -2519
rect 4099 -1743 4133 -1727
rect 4099 -2535 4133 -2519
rect 4237 -1743 4271 -1727
rect 4237 -2535 4271 -2519
rect 4375 -1743 4409 -1727
rect 4375 -2535 4409 -2519
rect 4513 -1743 4547 -1727
rect 4513 -2535 4547 -2519
rect 4651 -1743 4685 -1727
rect 4651 -2535 4685 -2519
rect 4789 -1743 4823 -1727
rect 4789 -2535 4823 -2519
rect 4927 -1743 4961 -1727
rect 4927 -2535 4961 -2519
rect 5065 -1743 5099 -1727
rect 5065 -2535 5099 -2519
rect 5203 -1743 5237 -1727
rect 5203 -2535 5237 -2519
rect 5341 -1743 5375 -1727
rect 5341 -2535 5375 -2519
rect 5479 -1743 5513 -1727
rect 5479 -2535 5513 -2519
rect 5617 -1743 5651 -1727
rect 5617 -2535 5651 -2519
rect 5755 -1743 5789 -1727
rect 5755 -2535 5789 -2519
rect 5893 -1743 5927 -1727
rect 5893 -2535 5927 -2519
rect 6031 -1743 6065 -1727
rect 6031 -2535 6065 -2519
rect 6169 -1743 6203 -1727
rect 6169 -2535 6203 -2519
rect 6307 -1743 6341 -1727
rect 6307 -2535 6341 -2519
rect 6445 -1743 6479 -1727
rect 6445 -2535 6479 -2519
rect 6583 -1743 6617 -1727
rect 6583 -2535 6617 -2519
rect 6721 -1743 6755 -1727
rect 6721 -2535 6755 -2519
rect 6859 -1743 6893 -1727
rect 6859 -2535 6893 -2519
rect 6997 -1743 7031 -1727
rect 6997 -2535 7031 -2519
rect 7135 -1743 7169 -1727
rect 7135 -2535 7169 -2519
rect 7273 -1743 7307 -1727
rect 7273 -2535 7307 -2519
rect 7411 -1743 7445 -1727
rect 7411 -2535 7445 -2519
rect 7549 -1743 7583 -1727
rect 7549 -2535 7583 -2519
rect 7687 -1743 7721 -1727
rect 7687 -2535 7721 -2519
rect 7825 -1743 7859 -1727
rect 7825 -2535 7859 -2519
rect 7963 -1743 7997 -1727
rect 7963 -2535 7997 -2519
rect 8101 -1743 8135 -1727
rect 8101 -2535 8135 -2519
rect 8239 -1743 8273 -1727
rect 8239 -2535 8273 -2519
rect 8377 -1743 8411 -1727
rect 8377 -2535 8411 -2519
rect 8515 -1743 8549 -1727
rect 8515 -2535 8549 -2519
rect 8653 -1743 8687 -1727
rect 8653 -2535 8687 -2519
rect 8791 -1743 8825 -1727
rect 8791 -2535 8825 -2519
rect 8929 -1743 8963 -1727
rect 8929 -2535 8963 -2519
rect 9067 -1743 9101 -1727
rect 9067 -2535 9101 -2519
rect 9205 -1743 9239 -1727
rect 9205 -2535 9239 -2519
rect 9343 -1743 9377 -1727
rect 9343 -2535 9377 -2519
rect 9481 -1743 9515 -1727
rect 9481 -2535 9515 -2519
rect 9619 -1743 9653 -1727
rect 9619 -2535 9653 -2519
rect 9757 -1743 9791 -1727
rect 9757 -2535 9791 -2519
rect 9895 -1743 9929 -1727
rect 9895 -2535 9929 -2519
rect 10033 -1743 10067 -1727
rect 10033 -2535 10067 -2519
rect 10171 -1743 10205 -1727
rect 10171 -2535 10205 -2519
rect 10309 -1743 10343 -1727
rect 10309 -2535 10343 -2519
rect 10447 -1743 10481 -1727
rect 10447 -2535 10481 -2519
rect 10585 -1743 10619 -1727
rect 10585 -2535 10619 -2519
rect 10723 -1743 10757 -1727
rect 10723 -2535 10757 -2519
rect 10861 -1743 10895 -1727
rect 10861 -2535 10895 -2519
rect 10999 -1743 11033 -1727
rect 10999 -2535 11033 -2519
rect 11137 -1743 11171 -1727
rect 11137 -2535 11171 -2519
rect 11275 -1743 11309 -1727
rect 11275 -2535 11309 -2519
rect 11413 -1743 11447 -1727
rect 11413 -2535 11447 -2519
rect 11551 -1743 11585 -1727
rect 11551 -2535 11585 -2519
rect 11689 -1743 11723 -1727
rect 11689 -2535 11723 -2519
rect 11827 -1743 11861 -1727
rect 11827 -2535 11861 -2519
rect 11965 -1743 11999 -1727
rect 11965 -2535 11999 -2519
rect 12103 -1743 12137 -1727
rect 12103 -2535 12137 -2519
rect 12241 -1743 12275 -1727
rect 12241 -2535 12275 -2519
rect 12379 -1743 12413 -1727
rect 12379 -2535 12413 -2519
rect 12517 -1743 12551 -1727
rect 12517 -2535 12551 -2519
rect 12655 -1743 12689 -1727
rect 12655 -2535 12689 -2519
rect 12793 -1743 12827 -1727
rect 12793 -2535 12827 -2519
rect 12931 -1743 12965 -1727
rect 12931 -2535 12965 -2519
rect 13069 -1743 13103 -1727
rect 13069 -2535 13103 -2519
rect 13207 -1743 13241 -1727
rect 13207 -2535 13241 -2519
rect 13345 -1743 13379 -1727
rect 13345 -2535 13379 -2519
rect 13483 -1743 13517 -1727
rect 13483 -2535 13517 -2519
rect 13621 -1743 13655 -1727
rect 13621 -2535 13655 -2519
rect 13759 -1743 13793 -1727
rect 13759 -2535 13793 -2519
rect 13897 -1743 13931 -1727
rect 13897 -2535 13931 -2519
rect 97 -2629 131 -2613
rect 97 -3421 131 -3405
rect 235 -2629 269 -2613
rect 235 -3421 269 -3405
rect 373 -2629 407 -2613
rect 373 -3421 407 -3405
rect 511 -2629 545 -2613
rect 511 -3421 545 -3405
rect 649 -2629 683 -2613
rect 649 -3421 683 -3405
rect 787 -2629 821 -2613
rect 787 -3421 821 -3405
rect 925 -2629 959 -2613
rect 925 -3421 959 -3405
rect 1063 -2629 1097 -2613
rect 1063 -3421 1097 -3405
rect 1201 -2629 1235 -2613
rect 1201 -3421 1235 -3405
rect 1339 -2629 1373 -2613
rect 1339 -3421 1373 -3405
rect 1477 -2629 1511 -2613
rect 1477 -3421 1511 -3405
rect 1615 -2629 1649 -2613
rect 1615 -3421 1649 -3405
rect 1753 -2629 1787 -2613
rect 1753 -3421 1787 -3405
rect 1891 -2629 1925 -2613
rect 1891 -3421 1925 -3405
rect 2029 -2629 2063 -2613
rect 2029 -3421 2063 -3405
rect 2167 -2629 2201 -2613
rect 2167 -3421 2201 -3405
rect 2305 -2629 2339 -2613
rect 2305 -3421 2339 -3405
rect 2443 -2629 2477 -2613
rect 2443 -3421 2477 -3405
rect 2581 -2629 2615 -2613
rect 2581 -3421 2615 -3405
rect 2719 -2629 2753 -2613
rect 2719 -3421 2753 -3405
rect 2857 -2629 2891 -2613
rect 2857 -3421 2891 -3405
rect 2995 -2629 3029 -2613
rect 2995 -3421 3029 -3405
rect 3133 -2629 3167 -2613
rect 3133 -3421 3167 -3405
rect 3271 -2629 3305 -2613
rect 3271 -3421 3305 -3405
rect 3409 -2629 3443 -2613
rect 3409 -3421 3443 -3405
rect 3547 -2629 3581 -2613
rect 3547 -3421 3581 -3405
rect 3685 -2629 3719 -2613
rect 3685 -3421 3719 -3405
rect 3823 -2629 3857 -2613
rect 3823 -3421 3857 -3405
rect 3961 -2629 3995 -2613
rect 3961 -3421 3995 -3405
rect 4099 -2629 4133 -2613
rect 4099 -3421 4133 -3405
rect 4237 -2629 4271 -2613
rect 4237 -3421 4271 -3405
rect 4375 -2629 4409 -2613
rect 4375 -3421 4409 -3405
rect 4513 -2629 4547 -2613
rect 4513 -3421 4547 -3405
rect 4651 -2629 4685 -2613
rect 4651 -3421 4685 -3405
rect 4789 -2629 4823 -2613
rect 4789 -3421 4823 -3405
rect 4927 -2629 4961 -2613
rect 4927 -3421 4961 -3405
rect 5065 -2629 5099 -2613
rect 5065 -3421 5099 -3405
rect 5203 -2629 5237 -2613
rect 5203 -3421 5237 -3405
rect 5341 -2629 5375 -2613
rect 5341 -3421 5375 -3405
rect 5479 -2629 5513 -2613
rect 5479 -3421 5513 -3405
rect 5617 -2629 5651 -2613
rect 5617 -3421 5651 -3405
rect 5755 -2629 5789 -2613
rect 5755 -3421 5789 -3405
rect 5893 -2629 5927 -2613
rect 5893 -3421 5927 -3405
rect 6031 -2629 6065 -2613
rect 6031 -3421 6065 -3405
rect 6169 -2629 6203 -2613
rect 6169 -3421 6203 -3405
rect 6307 -2629 6341 -2613
rect 6307 -3421 6341 -3405
rect 6445 -2629 6479 -2613
rect 6445 -3421 6479 -3405
rect 6583 -2629 6617 -2613
rect 6583 -3421 6617 -3405
rect 6721 -2629 6755 -2613
rect 6721 -3421 6755 -3405
rect 6859 -2629 6893 -2613
rect 6859 -3421 6893 -3405
rect 6997 -2629 7031 -2613
rect 6997 -3421 7031 -3405
rect 7135 -2629 7169 -2613
rect 7135 -3421 7169 -3405
rect 7273 -2629 7307 -2613
rect 7273 -3421 7307 -3405
rect 7411 -2629 7445 -2613
rect 7411 -3421 7445 -3405
rect 7549 -2629 7583 -2613
rect 7549 -3421 7583 -3405
rect 7687 -2629 7721 -2613
rect 7687 -3421 7721 -3405
rect 7825 -2629 7859 -2613
rect 7825 -3421 7859 -3405
rect 7963 -2629 7997 -2613
rect 7963 -3421 7997 -3405
rect 8101 -2629 8135 -2613
rect 8101 -3421 8135 -3405
rect 8239 -2629 8273 -2613
rect 8239 -3421 8273 -3405
rect 8377 -2629 8411 -2613
rect 8377 -3421 8411 -3405
rect 8515 -2629 8549 -2613
rect 8515 -3421 8549 -3405
rect 8653 -2629 8687 -2613
rect 8653 -3421 8687 -3405
rect 8791 -2629 8825 -2613
rect 8791 -3421 8825 -3405
rect 8929 -2629 8963 -2613
rect 8929 -3421 8963 -3405
rect 9067 -2629 9101 -2613
rect 9067 -3421 9101 -3405
rect 9205 -2629 9239 -2613
rect 9205 -3421 9239 -3405
rect 9343 -2629 9377 -2613
rect 9343 -3421 9377 -3405
rect 9481 -2629 9515 -2613
rect 9481 -3421 9515 -3405
rect 9619 -2629 9653 -2613
rect 9619 -3421 9653 -3405
rect 9757 -2629 9791 -2613
rect 9757 -3421 9791 -3405
rect 9895 -2629 9929 -2613
rect 9895 -3421 9929 -3405
rect 10033 -2629 10067 -2613
rect 10033 -3421 10067 -3405
rect 10171 -2629 10205 -2613
rect 10171 -3421 10205 -3405
rect 10309 -2629 10343 -2613
rect 10309 -3421 10343 -3405
rect 10447 -2629 10481 -2613
rect 10447 -3421 10481 -3405
rect 10585 -2629 10619 -2613
rect 10585 -3421 10619 -3405
rect 10723 -2629 10757 -2613
rect 10723 -3421 10757 -3405
rect 10861 -2629 10895 -2613
rect 10861 -3421 10895 -3405
rect 10999 -2629 11033 -2613
rect 10999 -3421 11033 -3405
rect 11137 -2629 11171 -2613
rect 11137 -3421 11171 -3405
rect 11275 -2629 11309 -2613
rect 11275 -3421 11309 -3405
rect 11413 -2629 11447 -2613
rect 11413 -3421 11447 -3405
rect 11551 -2629 11585 -2613
rect 11551 -3421 11585 -3405
rect 11689 -2629 11723 -2613
rect 11689 -3421 11723 -3405
rect 11827 -2629 11861 -2613
rect 11827 -3421 11861 -3405
rect 11965 -2629 11999 -2613
rect 11965 -3421 11999 -3405
rect 12103 -2629 12137 -2613
rect 12103 -3421 12137 -3405
rect 12241 -2629 12275 -2613
rect 12241 -3421 12275 -3405
rect 12379 -2629 12413 -2613
rect 12379 -3421 12413 -3405
rect 12517 -2629 12551 -2613
rect 12517 -3421 12551 -3405
rect 12655 -2629 12689 -2613
rect 12655 -3421 12689 -3405
rect 12793 -2629 12827 -2613
rect 12793 -3421 12827 -3405
rect 12931 -2629 12965 -2613
rect 12931 -3421 12965 -3405
rect 13069 -2629 13103 -2613
rect 13069 -3421 13103 -3405
rect 13207 -2629 13241 -2613
rect 13207 -3421 13241 -3405
rect 13345 -2629 13379 -2613
rect 13345 -3421 13379 -3405
rect 13483 -2629 13517 -2613
rect 13483 -3421 13517 -3405
rect 13621 -2629 13655 -2613
rect 13621 -3421 13655 -3405
rect 13759 -2629 13793 -2613
rect 13759 -3421 13793 -3405
rect 13897 -2629 13931 -2613
rect 13897 -3421 13931 -3405
rect -12 -3541 22 -3479
rect 143 -3498 159 -3464
rect 207 -3498 223 -3464
rect 281 -3498 297 -3464
rect 345 -3498 361 -3464
rect 419 -3498 435 -3464
rect 483 -3498 499 -3464
rect 557 -3498 573 -3464
rect 621 -3498 637 -3464
rect 695 -3498 711 -3464
rect 759 -3498 775 -3464
rect 833 -3498 849 -3464
rect 897 -3498 913 -3464
rect 971 -3498 987 -3464
rect 1035 -3498 1051 -3464
rect 1109 -3498 1125 -3464
rect 1173 -3498 1189 -3464
rect 1247 -3498 1263 -3464
rect 1311 -3498 1327 -3464
rect 1385 -3498 1401 -3464
rect 1449 -3498 1465 -3464
rect 1523 -3498 1539 -3464
rect 1587 -3498 1603 -3464
rect 1661 -3498 1677 -3464
rect 1725 -3498 1741 -3464
rect 1799 -3498 1815 -3464
rect 1863 -3498 1879 -3464
rect 1937 -3498 1953 -3464
rect 2001 -3498 2017 -3464
rect 2075 -3498 2091 -3464
rect 2139 -3498 2155 -3464
rect 2213 -3498 2229 -3464
rect 2277 -3498 2293 -3464
rect 2351 -3498 2367 -3464
rect 2415 -3498 2431 -3464
rect 2489 -3498 2505 -3464
rect 2553 -3498 2569 -3464
rect 2627 -3498 2643 -3464
rect 2691 -3498 2707 -3464
rect 2765 -3498 2781 -3464
rect 2829 -3498 2845 -3464
rect 2903 -3498 2919 -3464
rect 2967 -3498 2983 -3464
rect 3041 -3498 3057 -3464
rect 3105 -3498 3121 -3464
rect 3179 -3498 3195 -3464
rect 3243 -3498 3259 -3464
rect 3317 -3498 3333 -3464
rect 3381 -3498 3397 -3464
rect 3455 -3498 3471 -3464
rect 3519 -3498 3535 -3464
rect 3593 -3498 3609 -3464
rect 3657 -3498 3673 -3464
rect 3731 -3498 3747 -3464
rect 3795 -3498 3811 -3464
rect 3869 -3498 3885 -3464
rect 3933 -3498 3949 -3464
rect 4007 -3498 4023 -3464
rect 4071 -3498 4087 -3464
rect 4145 -3498 4161 -3464
rect 4209 -3498 4225 -3464
rect 4283 -3498 4299 -3464
rect 4347 -3498 4363 -3464
rect 4421 -3498 4437 -3464
rect 4485 -3498 4501 -3464
rect 4559 -3498 4575 -3464
rect 4623 -3498 4639 -3464
rect 4697 -3498 4713 -3464
rect 4761 -3498 4777 -3464
rect 4835 -3498 4851 -3464
rect 4899 -3498 4915 -3464
rect 4973 -3498 4989 -3464
rect 5037 -3498 5053 -3464
rect 5111 -3498 5127 -3464
rect 5175 -3498 5191 -3464
rect 5249 -3498 5265 -3464
rect 5313 -3498 5329 -3464
rect 5387 -3498 5403 -3464
rect 5451 -3498 5467 -3464
rect 5525 -3498 5541 -3464
rect 5589 -3498 5605 -3464
rect 5663 -3498 5679 -3464
rect 5727 -3498 5743 -3464
rect 5801 -3498 5817 -3464
rect 5865 -3498 5881 -3464
rect 5939 -3498 5955 -3464
rect 6003 -3498 6019 -3464
rect 6077 -3498 6093 -3464
rect 6141 -3498 6157 -3464
rect 6215 -3498 6231 -3464
rect 6279 -3498 6295 -3464
rect 6353 -3498 6369 -3464
rect 6417 -3498 6433 -3464
rect 6491 -3498 6507 -3464
rect 6555 -3498 6571 -3464
rect 6629 -3498 6645 -3464
rect 6693 -3498 6709 -3464
rect 6767 -3498 6783 -3464
rect 6831 -3498 6847 -3464
rect 6905 -3498 6921 -3464
rect 6969 -3498 6985 -3464
rect 7043 -3498 7059 -3464
rect 7107 -3498 7123 -3464
rect 7181 -3498 7197 -3464
rect 7245 -3498 7261 -3464
rect 7319 -3498 7335 -3464
rect 7383 -3498 7399 -3464
rect 7457 -3498 7473 -3464
rect 7521 -3498 7537 -3464
rect 7595 -3498 7611 -3464
rect 7659 -3498 7675 -3464
rect 7733 -3498 7749 -3464
rect 7797 -3498 7813 -3464
rect 7871 -3498 7887 -3464
rect 7935 -3498 7951 -3464
rect 8009 -3498 8025 -3464
rect 8073 -3498 8089 -3464
rect 8147 -3498 8163 -3464
rect 8211 -3498 8227 -3464
rect 8285 -3498 8301 -3464
rect 8349 -3498 8365 -3464
rect 8423 -3498 8439 -3464
rect 8487 -3498 8503 -3464
rect 8561 -3498 8577 -3464
rect 8625 -3498 8641 -3464
rect 8699 -3498 8715 -3464
rect 8763 -3498 8779 -3464
rect 8837 -3498 8853 -3464
rect 8901 -3498 8917 -3464
rect 8975 -3498 8991 -3464
rect 9039 -3498 9055 -3464
rect 9113 -3498 9129 -3464
rect 9177 -3498 9193 -3464
rect 9251 -3498 9267 -3464
rect 9315 -3498 9331 -3464
rect 9389 -3498 9405 -3464
rect 9453 -3498 9469 -3464
rect 9527 -3498 9543 -3464
rect 9591 -3498 9607 -3464
rect 9665 -3498 9681 -3464
rect 9729 -3498 9745 -3464
rect 9803 -3498 9819 -3464
rect 9867 -3498 9883 -3464
rect 9941 -3498 9957 -3464
rect 10005 -3498 10021 -3464
rect 10079 -3498 10095 -3464
rect 10143 -3498 10159 -3464
rect 10217 -3498 10233 -3464
rect 10281 -3498 10297 -3464
rect 10355 -3498 10371 -3464
rect 10419 -3498 10435 -3464
rect 10493 -3498 10509 -3464
rect 10557 -3498 10573 -3464
rect 10631 -3498 10647 -3464
rect 10695 -3498 10711 -3464
rect 10769 -3498 10785 -3464
rect 10833 -3498 10849 -3464
rect 10907 -3498 10923 -3464
rect 10971 -3498 10987 -3464
rect 11045 -3498 11061 -3464
rect 11109 -3498 11125 -3464
rect 11183 -3498 11199 -3464
rect 11247 -3498 11263 -3464
rect 11321 -3498 11337 -3464
rect 11385 -3498 11401 -3464
rect 11459 -3498 11475 -3464
rect 11523 -3498 11539 -3464
rect 11597 -3498 11613 -3464
rect 11661 -3498 11677 -3464
rect 11735 -3498 11751 -3464
rect 11799 -3498 11815 -3464
rect 11873 -3498 11889 -3464
rect 11937 -3498 11953 -3464
rect 12011 -3498 12027 -3464
rect 12075 -3498 12091 -3464
rect 12149 -3498 12165 -3464
rect 12213 -3498 12229 -3464
rect 12287 -3498 12303 -3464
rect 12351 -3498 12367 -3464
rect 12425 -3498 12441 -3464
rect 12489 -3498 12505 -3464
rect 12563 -3498 12579 -3464
rect 12627 -3498 12643 -3464
rect 12701 -3498 12717 -3464
rect 12765 -3498 12781 -3464
rect 12839 -3498 12855 -3464
rect 12903 -3498 12919 -3464
rect 12977 -3498 12993 -3464
rect 13041 -3498 13057 -3464
rect 13115 -3498 13131 -3464
rect 13179 -3498 13195 -3464
rect 13253 -3498 13269 -3464
rect 13317 -3498 13333 -3464
rect 13391 -3498 13407 -3464
rect 13455 -3498 13471 -3464
rect 13529 -3498 13545 -3464
rect 13593 -3498 13609 -3464
rect 13667 -3498 13683 -3464
rect 13731 -3498 13747 -3464
rect 13805 -3498 13821 -3464
rect 13869 -3498 13885 -3464
rect 14005 -3541 14039 -3479
rect -12 -3575 84 -3541
rect 13943 -3575 14039 -3541
<< viali >>
rect -850 -1551 14344 -970
rect 97 -2519 131 -1743
rect 235 -2519 269 -1743
rect 373 -2519 407 -1743
rect 511 -2519 545 -1743
rect 649 -2519 683 -1743
rect 787 -2519 821 -1743
rect 925 -2519 959 -1743
rect 1063 -2519 1097 -1743
rect 1201 -2519 1235 -1743
rect 1339 -2519 1373 -1743
rect 1477 -2519 1511 -1743
rect 1615 -2519 1649 -1743
rect 1753 -2519 1787 -1743
rect 1891 -2519 1925 -1743
rect 2029 -2519 2063 -1743
rect 2167 -2519 2201 -1743
rect 2305 -2519 2339 -1743
rect 2443 -2519 2477 -1743
rect 2581 -2519 2615 -1743
rect 2719 -2519 2753 -1743
rect 2857 -2519 2891 -1743
rect 2995 -2519 3029 -1743
rect 3133 -2519 3167 -1743
rect 3271 -2519 3305 -1743
rect 3409 -2519 3443 -1743
rect 3547 -2519 3581 -1743
rect 3685 -2519 3719 -1743
rect 3823 -2519 3857 -1743
rect 3961 -2519 3995 -1743
rect 4099 -2519 4133 -1743
rect 4237 -2519 4271 -1743
rect 4375 -2519 4409 -1743
rect 4513 -2519 4547 -1743
rect 4651 -2519 4685 -1743
rect 4789 -2519 4823 -1743
rect 4927 -2519 4961 -1743
rect 5065 -2519 5099 -1743
rect 5203 -2519 5237 -1743
rect 5341 -2519 5375 -1743
rect 5479 -2519 5513 -1743
rect 5617 -2519 5651 -1743
rect 5755 -2519 5789 -1743
rect 5893 -2519 5927 -1743
rect 6031 -2519 6065 -1743
rect 6169 -2519 6203 -1743
rect 6307 -2519 6341 -1743
rect 6445 -2519 6479 -1743
rect 6583 -2519 6617 -1743
rect 6721 -2519 6755 -1743
rect 6859 -2519 6893 -1743
rect 6997 -2519 7031 -1743
rect 7135 -2519 7169 -1743
rect 7273 -2519 7307 -1743
rect 7411 -2519 7445 -1743
rect 7549 -2519 7583 -1743
rect 7687 -2519 7721 -1743
rect 7825 -2519 7859 -1743
rect 7963 -2519 7997 -1743
rect 8101 -2519 8135 -1743
rect 8239 -2519 8273 -1743
rect 8377 -2519 8411 -1743
rect 8515 -2519 8549 -1743
rect 8653 -2519 8687 -1743
rect 8791 -2519 8825 -1743
rect 8929 -2519 8963 -1743
rect 9067 -2519 9101 -1743
rect 9205 -2519 9239 -1743
rect 9343 -2519 9377 -1743
rect 9481 -2519 9515 -1743
rect 9619 -2519 9653 -1743
rect 9757 -2519 9791 -1743
rect 9895 -2519 9929 -1743
rect 10033 -2519 10067 -1743
rect 10171 -2519 10205 -1743
rect 10309 -2519 10343 -1743
rect 10447 -2519 10481 -1743
rect 10585 -2519 10619 -1743
rect 10723 -2519 10757 -1743
rect 10861 -2519 10895 -1743
rect 10999 -2519 11033 -1743
rect 11137 -2519 11171 -1743
rect 11275 -2519 11309 -1743
rect 11413 -2519 11447 -1743
rect 11551 -2519 11585 -1743
rect 11689 -2519 11723 -1743
rect 11827 -2519 11861 -1743
rect 11965 -2519 11999 -1743
rect 12103 -2519 12137 -1743
rect 12241 -2519 12275 -1743
rect 12379 -2519 12413 -1743
rect 12517 -2519 12551 -1743
rect 12655 -2519 12689 -1743
rect 12793 -2519 12827 -1743
rect 12931 -2519 12965 -1743
rect 13069 -2519 13103 -1743
rect 13207 -2519 13241 -1743
rect 13345 -2519 13379 -1743
rect 13483 -2519 13517 -1743
rect 13621 -2519 13655 -1743
rect 13759 -2519 13793 -1743
rect 13897 -2519 13931 -1743
rect 97 -3405 131 -2629
rect 235 -3405 269 -2629
rect 373 -3405 407 -2629
rect 511 -3405 545 -2629
rect 649 -3405 683 -2629
rect 787 -3405 821 -2629
rect 925 -3405 959 -2629
rect 1063 -3405 1097 -2629
rect 1201 -3405 1235 -2629
rect 1339 -3405 1373 -2629
rect 1477 -3405 1511 -2629
rect 1615 -3405 1649 -2629
rect 1753 -3405 1787 -2629
rect 1891 -3405 1925 -2629
rect 2029 -3405 2063 -2629
rect 2167 -3405 2201 -2629
rect 2305 -3405 2339 -2629
rect 2443 -3405 2477 -2629
rect 2581 -3405 2615 -2629
rect 2719 -3405 2753 -2629
rect 2857 -3405 2891 -2629
rect 2995 -3405 3029 -2629
rect 3133 -3405 3167 -2629
rect 3271 -3405 3305 -2629
rect 3409 -3405 3443 -2629
rect 3547 -3405 3581 -2629
rect 3685 -3405 3719 -2629
rect 3823 -3405 3857 -2629
rect 3961 -3405 3995 -2629
rect 4099 -3405 4133 -2629
rect 4237 -3405 4271 -2629
rect 4375 -3405 4409 -2629
rect 4513 -3405 4547 -2629
rect 4651 -3405 4685 -2629
rect 4789 -3405 4823 -2629
rect 4927 -3405 4961 -2629
rect 5065 -3405 5099 -2629
rect 5203 -3405 5237 -2629
rect 5341 -3405 5375 -2629
rect 5479 -3405 5513 -2629
rect 5617 -3405 5651 -2629
rect 5755 -3405 5789 -2629
rect 5893 -3405 5927 -2629
rect 6031 -3405 6065 -2629
rect 6169 -3405 6203 -2629
rect 6307 -3405 6341 -2629
rect 6445 -3405 6479 -2629
rect 6583 -3405 6617 -2629
rect 6721 -3405 6755 -2629
rect 6859 -3405 6893 -2629
rect 6997 -3405 7031 -2629
rect 7135 -3405 7169 -2629
rect 7273 -3405 7307 -2629
rect 7411 -3405 7445 -2629
rect 7549 -3405 7583 -2629
rect 7687 -3405 7721 -2629
rect 7825 -3405 7859 -2629
rect 7963 -3405 7997 -2629
rect 8101 -3405 8135 -2629
rect 8239 -3405 8273 -2629
rect 8377 -3405 8411 -2629
rect 8515 -3405 8549 -2629
rect 8653 -3405 8687 -2629
rect 8791 -3405 8825 -2629
rect 8929 -3405 8963 -2629
rect 9067 -3405 9101 -2629
rect 9205 -3405 9239 -2629
rect 9343 -3405 9377 -2629
rect 9481 -3405 9515 -2629
rect 9619 -3405 9653 -2629
rect 9757 -3405 9791 -2629
rect 9895 -3405 9929 -2629
rect 10033 -3405 10067 -2629
rect 10171 -3405 10205 -2629
rect 10309 -3405 10343 -2629
rect 10447 -3405 10481 -2629
rect 10585 -3405 10619 -2629
rect 10723 -3405 10757 -2629
rect 10861 -3405 10895 -2629
rect 10999 -3405 11033 -2629
rect 11137 -3405 11171 -2629
rect 11275 -3405 11309 -2629
rect 11413 -3405 11447 -2629
rect 11551 -3405 11585 -2629
rect 11689 -3405 11723 -2629
rect 11827 -3405 11861 -2629
rect 11965 -3405 11999 -2629
rect 12103 -3405 12137 -2629
rect 12241 -3405 12275 -2629
rect 12379 -3405 12413 -2629
rect 12517 -3405 12551 -2629
rect 12655 -3405 12689 -2629
rect 12793 -3405 12827 -2629
rect 12931 -3405 12965 -2629
rect 13069 -3405 13103 -2629
rect 13207 -3405 13241 -2629
rect 13345 -3405 13379 -2629
rect 13483 -3405 13517 -2629
rect 13621 -3405 13655 -2629
rect 13759 -3405 13793 -2629
rect 13897 -3405 13931 -2629
rect 159 -3498 207 -3464
rect 297 -3498 345 -3464
rect 435 -3498 483 -3464
rect 573 -3498 621 -3464
rect 711 -3498 759 -3464
rect 849 -3498 897 -3464
rect 987 -3498 1035 -3464
rect 1125 -3498 1173 -3464
rect 1263 -3498 1311 -3464
rect 1401 -3498 1449 -3464
rect 1539 -3498 1587 -3464
rect 1677 -3498 1725 -3464
rect 1815 -3498 1863 -3464
rect 1953 -3498 2001 -3464
rect 2091 -3498 2139 -3464
rect 2229 -3498 2277 -3464
rect 2367 -3498 2415 -3464
rect 2505 -3498 2553 -3464
rect 2643 -3498 2691 -3464
rect 2781 -3498 2829 -3464
rect 2919 -3498 2967 -3464
rect 3057 -3498 3105 -3464
rect 3195 -3498 3243 -3464
rect 3333 -3498 3381 -3464
rect 3471 -3498 3519 -3464
rect 3609 -3498 3657 -3464
rect 3747 -3498 3795 -3464
rect 3885 -3498 3933 -3464
rect 4023 -3498 4071 -3464
rect 4161 -3498 4209 -3464
rect 4299 -3498 4347 -3464
rect 4437 -3498 4485 -3464
rect 4575 -3498 4623 -3464
rect 4713 -3498 4761 -3464
rect 4851 -3498 4899 -3464
rect 4989 -3498 5037 -3464
rect 5127 -3498 5175 -3464
rect 5265 -3498 5313 -3464
rect 5403 -3498 5451 -3464
rect 5541 -3498 5589 -3464
rect 5679 -3498 5727 -3464
rect 5817 -3498 5865 -3464
rect 5955 -3498 6003 -3464
rect 6093 -3498 6141 -3464
rect 6231 -3498 6279 -3464
rect 6369 -3498 6417 -3464
rect 6507 -3498 6555 -3464
rect 6645 -3498 6693 -3464
rect 6783 -3498 6831 -3464
rect 6921 -3498 6969 -3464
rect 7059 -3498 7107 -3464
rect 7197 -3498 7245 -3464
rect 7335 -3498 7383 -3464
rect 7473 -3498 7521 -3464
rect 7611 -3498 7659 -3464
rect 7749 -3498 7797 -3464
rect 7887 -3498 7935 -3464
rect 8025 -3498 8073 -3464
rect 8163 -3498 8211 -3464
rect 8301 -3498 8349 -3464
rect 8439 -3498 8487 -3464
rect 8577 -3498 8625 -3464
rect 8715 -3498 8763 -3464
rect 8853 -3498 8901 -3464
rect 8991 -3498 9039 -3464
rect 9129 -3498 9177 -3464
rect 9267 -3498 9315 -3464
rect 9405 -3498 9453 -3464
rect 9543 -3498 9591 -3464
rect 9681 -3498 9729 -3464
rect 9819 -3498 9867 -3464
rect 9957 -3498 10005 -3464
rect 10095 -3498 10143 -3464
rect 10233 -3498 10281 -3464
rect 10371 -3498 10419 -3464
rect 10509 -3498 10557 -3464
rect 10647 -3498 10695 -3464
rect 10785 -3498 10833 -3464
rect 10923 -3498 10971 -3464
rect 11061 -3498 11109 -3464
rect 11199 -3498 11247 -3464
rect 11337 -3498 11385 -3464
rect 11475 -3498 11523 -3464
rect 11613 -3498 11661 -3464
rect 11751 -3498 11799 -3464
rect 11889 -3498 11937 -3464
rect 12027 -3498 12075 -3464
rect 12165 -3498 12213 -3464
rect 12303 -3498 12351 -3464
rect 12441 -3498 12489 -3464
rect 12579 -3498 12627 -3464
rect 12717 -3498 12765 -3464
rect 12855 -3498 12903 -3464
rect 12993 -3498 13041 -3464
rect 13131 -3498 13179 -3464
rect 13269 -3498 13317 -3464
rect 13407 -3498 13455 -3464
rect 13545 -3498 13593 -3464
rect 13683 -3498 13731 -3464
rect 13821 -3498 13869 -3464
<< metal1 >>
rect 4664 5512 9931 5551
rect 4664 4701 6583 5512
rect 8032 4701 9931 5512
rect 4664 4670 9931 4701
rect 4664 2901 5546 4670
rect 9049 2901 9931 4670
rect 1586 2254 12997 2901
rect 1587 1561 1952 2254
rect 3795 1561 4160 2254
rect 6003 1561 6368 2254
rect 8211 1561 8576 2254
rect 10419 1561 10784 2254
rect 12627 1561 12992 2254
rect 297 1375 13731 1561
rect 297 982 483 1375
rect 849 982 1035 1375
rect 1401 982 1587 1375
rect 1953 982 2139 1375
rect 2505 982 2691 1375
rect 3057 982 3243 1375
rect 3609 982 3795 1375
rect 4161 982 4347 1375
rect 4713 982 4899 1375
rect 5265 982 5451 1375
rect 5817 982 6003 1375
rect 6369 982 6555 1375
rect 6921 982 7107 1375
rect 7473 982 7659 1375
rect 8025 982 8211 1375
rect 8577 982 8763 1375
rect 9129 982 9315 1375
rect 9681 982 9867 1375
rect 10233 982 10419 1375
rect 10785 982 10971 1375
rect 11337 982 11523 1375
rect 11889 982 12075 1375
rect 12441 982 12627 1375
rect 12993 982 13179 1375
rect 13545 982 13731 1375
rect 147 936 13881 982
rect 91 -964 137 895
rect 216 107 226 883
rect 278 107 288 883
rect 216 -771 226 5
rect 278 -771 288 5
rect 367 -964 413 895
rect 492 107 502 883
rect 554 107 564 883
rect 492 -771 502 5
rect 554 -771 564 5
rect 643 -964 689 895
rect 768 107 778 883
rect 830 107 840 883
rect 768 -771 778 5
rect 830 -771 840 5
rect 919 -964 965 895
rect 1044 107 1054 883
rect 1106 107 1116 883
rect 1044 -771 1054 5
rect 1106 -771 1116 5
rect 1195 -964 1241 895
rect 1320 107 1330 883
rect 1382 107 1392 883
rect 1320 -771 1330 5
rect 1382 -771 1392 5
rect 1471 -964 1517 895
rect 1596 107 1606 883
rect 1658 107 1668 883
rect 1596 -771 1606 5
rect 1658 -771 1668 5
rect 1747 -964 1793 895
rect 1872 107 1882 883
rect 1934 107 1944 883
rect 1872 -771 1882 5
rect 1934 -771 1944 5
rect 2023 -964 2069 895
rect 2148 107 2158 883
rect 2210 107 2220 883
rect 2148 -771 2158 5
rect 2210 -771 2220 5
rect 2299 -964 2345 895
rect 2424 107 2434 883
rect 2486 107 2496 883
rect 2424 -771 2434 5
rect 2486 -771 2496 5
rect 2575 -964 2621 895
rect 2700 107 2710 883
rect 2762 107 2772 883
rect 2700 -771 2710 5
rect 2762 -771 2772 5
rect 2851 -964 2897 895
rect 2976 107 2986 883
rect 3038 107 3048 883
rect 2976 -771 2986 5
rect 3038 -771 3048 5
rect 3127 -964 3173 895
rect 3252 107 3262 883
rect 3314 107 3324 883
rect 3252 -771 3262 5
rect 3314 -771 3324 5
rect 3403 -964 3449 895
rect 3528 107 3538 883
rect 3590 107 3600 883
rect 3528 -771 3538 5
rect 3590 -771 3600 5
rect 3679 -964 3725 895
rect 3804 107 3814 883
rect 3866 107 3876 883
rect 3804 -771 3814 5
rect 3866 -771 3876 5
rect 3955 -964 4001 895
rect 4080 107 4090 883
rect 4142 107 4152 883
rect 4080 -771 4090 5
rect 4142 -771 4152 5
rect 4231 -964 4277 895
rect 4356 107 4366 883
rect 4418 107 4428 883
rect 4356 -771 4366 5
rect 4418 -771 4428 5
rect 4507 -964 4553 895
rect 4632 107 4642 883
rect 4694 107 4704 883
rect 4632 -771 4642 5
rect 4694 -771 4704 5
rect 4783 -964 4829 895
rect 4908 107 4918 883
rect 4970 107 4980 883
rect 4908 -771 4918 5
rect 4970 -771 4980 5
rect 5059 -964 5105 895
rect 5184 107 5194 883
rect 5246 107 5256 883
rect 5184 -771 5194 5
rect 5246 -771 5256 5
rect 5335 -964 5381 895
rect 5460 107 5470 883
rect 5522 107 5532 883
rect 5460 -771 5470 5
rect 5522 -771 5532 5
rect 5611 -964 5657 895
rect 5736 107 5746 883
rect 5798 107 5808 883
rect 5736 -771 5746 5
rect 5798 -771 5808 5
rect 5887 -964 5933 895
rect 6012 107 6022 883
rect 6074 107 6084 883
rect 6012 -771 6022 5
rect 6074 -771 6084 5
rect 6163 -964 6209 895
rect 6288 107 6298 883
rect 6350 107 6360 883
rect 6288 -771 6298 5
rect 6350 -771 6360 5
rect 6439 -964 6485 895
rect 6564 107 6574 883
rect 6626 107 6636 883
rect 6564 -771 6574 5
rect 6626 -771 6636 5
rect 6715 -964 6761 895
rect 6840 107 6850 883
rect 6902 107 6912 883
rect 6840 -771 6850 5
rect 6902 -771 6912 5
rect 6991 -964 7037 895
rect 7116 107 7126 883
rect 7178 107 7188 883
rect 7116 -771 7126 5
rect 7178 -771 7188 5
rect 7267 -964 7313 895
rect 7392 107 7402 883
rect 7454 107 7464 883
rect 7392 -771 7402 5
rect 7454 -771 7464 5
rect 7543 -964 7589 895
rect 7668 107 7678 883
rect 7730 107 7740 883
rect 7668 -771 7678 5
rect 7730 -771 7740 5
rect 7819 -964 7865 895
rect 7944 107 7954 883
rect 8006 107 8016 883
rect 7944 -771 7954 5
rect 8006 -771 8016 5
rect 8095 -964 8141 895
rect 8220 107 8230 883
rect 8282 107 8292 883
rect 8220 -771 8230 5
rect 8282 -771 8292 5
rect 8371 -964 8417 895
rect 8496 107 8506 883
rect 8558 107 8568 883
rect 8496 -771 8506 5
rect 8558 -771 8568 5
rect 8647 -964 8693 895
rect 8772 107 8782 883
rect 8834 107 8844 883
rect 8772 -771 8782 5
rect 8834 -771 8844 5
rect 8923 -964 8969 895
rect 9048 107 9058 883
rect 9110 107 9120 883
rect 9048 -771 9058 5
rect 9110 -771 9120 5
rect 9199 -964 9245 895
rect 9324 107 9334 883
rect 9386 107 9396 883
rect 9324 -771 9334 5
rect 9386 -771 9396 5
rect 9475 -964 9521 895
rect 9600 107 9610 883
rect 9662 107 9672 883
rect 9600 -771 9610 5
rect 9662 -771 9672 5
rect 9751 -964 9797 895
rect 9876 107 9886 883
rect 9938 107 9948 883
rect 9876 -771 9886 5
rect 9938 -771 9948 5
rect 10027 -964 10073 895
rect 10152 107 10162 883
rect 10214 107 10224 883
rect 10152 -771 10162 5
rect 10214 -771 10224 5
rect 10303 -964 10349 895
rect 10428 107 10438 883
rect 10490 107 10500 883
rect 10428 -771 10438 5
rect 10490 -771 10500 5
rect 10579 -964 10625 895
rect 10704 107 10714 883
rect 10766 107 10776 883
rect 10704 -771 10714 5
rect 10766 -771 10776 5
rect 10855 -964 10901 895
rect 10980 107 10990 883
rect 11042 107 11052 883
rect 10980 -771 10990 5
rect 11042 -771 11052 5
rect 11131 -964 11177 895
rect 11256 107 11266 883
rect 11318 107 11328 883
rect 11256 -771 11266 5
rect 11318 -771 11328 5
rect 11407 -964 11453 895
rect 11532 107 11542 883
rect 11594 107 11604 883
rect 11532 -771 11542 5
rect 11594 -771 11604 5
rect 11683 -964 11729 895
rect 11808 107 11818 883
rect 11870 107 11880 883
rect 11808 -771 11818 5
rect 11870 -771 11880 5
rect 11959 -964 12005 895
rect 12084 107 12094 883
rect 12146 107 12156 883
rect 12084 -771 12094 5
rect 12146 -771 12156 5
rect 12235 -964 12281 895
rect 12360 107 12370 883
rect 12422 107 12432 883
rect 12360 -771 12370 5
rect 12422 -771 12432 5
rect 12511 -964 12557 895
rect 12636 107 12646 883
rect 12698 107 12708 883
rect 12636 -771 12646 5
rect 12698 -771 12708 5
rect 12787 -964 12833 895
rect 12912 107 12922 883
rect 12974 107 12984 883
rect 12912 -771 12922 5
rect 12974 -771 12984 5
rect 13063 -964 13109 895
rect 13188 107 13198 883
rect 13250 107 13260 883
rect 13188 -771 13198 5
rect 13250 -771 13260 5
rect 13339 -964 13385 895
rect 13464 107 13474 883
rect 13526 107 13536 883
rect 13464 -771 13474 5
rect 13526 -771 13536 5
rect 13615 -964 13661 895
rect 13740 107 13750 883
rect 13802 107 13812 883
rect 13740 -771 13750 5
rect 13802 -771 13812 5
rect 13891 -964 13937 895
rect -862 -970 14356 -964
rect -862 -1551 -850 -970
rect 14344 -1551 14356 -970
rect -862 -1557 14356 -1551
rect 91 -1743 137 -1557
rect 91 -2519 97 -1743
rect 131 -2519 137 -1743
rect 229 -1743 275 -1731
rect 229 -1747 235 -1743
rect 269 -1747 275 -1743
rect 367 -1743 413 -1557
rect 91 -2629 137 -2519
rect 216 -2523 226 -1747
rect 278 -2523 288 -1747
rect 367 -2519 373 -1743
rect 407 -2519 413 -1743
rect 505 -1743 551 -1731
rect 505 -1747 511 -1743
rect 545 -1747 551 -1743
rect 643 -1743 689 -1557
rect 229 -2531 275 -2523
rect 229 -2625 275 -2617
rect 91 -3405 97 -2629
rect 131 -3405 137 -2629
rect 216 -3401 226 -2625
rect 278 -3401 288 -2625
rect 367 -2629 413 -2519
rect 492 -2523 502 -1747
rect 554 -2523 564 -1747
rect 643 -2519 649 -1743
rect 683 -2519 689 -1743
rect 781 -1743 827 -1731
rect 781 -1747 787 -1743
rect 821 -1747 827 -1743
rect 919 -1743 965 -1557
rect 505 -2531 551 -2523
rect 505 -2625 551 -2617
rect 91 -3417 137 -3405
rect 229 -3405 235 -3401
rect 269 -3405 275 -3401
rect 229 -3417 275 -3405
rect 367 -3405 373 -2629
rect 407 -3405 413 -2629
rect 492 -3401 502 -2625
rect 554 -3401 564 -2625
rect 643 -2629 689 -2519
rect 768 -2523 778 -1747
rect 830 -2523 840 -1747
rect 919 -2519 925 -1743
rect 959 -2519 965 -1743
rect 1057 -1743 1103 -1731
rect 1057 -1747 1063 -1743
rect 1097 -1747 1103 -1743
rect 1195 -1743 1241 -1557
rect 781 -2531 827 -2523
rect 781 -2625 827 -2617
rect 367 -3417 413 -3405
rect 505 -3405 511 -3401
rect 545 -3405 551 -3401
rect 505 -3417 551 -3405
rect 643 -3405 649 -2629
rect 683 -3405 689 -2629
rect 768 -3401 778 -2625
rect 830 -3401 840 -2625
rect 919 -2629 965 -2519
rect 1044 -2523 1054 -1747
rect 1106 -2523 1116 -1747
rect 1195 -2519 1201 -1743
rect 1235 -2519 1241 -1743
rect 1333 -1743 1379 -1731
rect 1333 -1747 1339 -1743
rect 1373 -1747 1379 -1743
rect 1471 -1743 1517 -1557
rect 1057 -2531 1103 -2523
rect 1057 -2625 1103 -2617
rect 643 -3417 689 -3405
rect 781 -3405 787 -3401
rect 821 -3405 827 -3401
rect 781 -3417 827 -3405
rect 919 -3405 925 -2629
rect 959 -3405 965 -2629
rect 1044 -3401 1054 -2625
rect 1106 -3401 1116 -2625
rect 1195 -2629 1241 -2519
rect 1320 -2523 1330 -1747
rect 1382 -2523 1392 -1747
rect 1471 -2519 1477 -1743
rect 1511 -2519 1517 -1743
rect 1609 -1743 1655 -1731
rect 1609 -1747 1615 -1743
rect 1649 -1747 1655 -1743
rect 1747 -1743 1793 -1557
rect 1333 -2531 1379 -2523
rect 1333 -2625 1379 -2617
rect 919 -3417 965 -3405
rect 1057 -3405 1063 -3401
rect 1097 -3405 1103 -3401
rect 1057 -3417 1103 -3405
rect 1195 -3405 1201 -2629
rect 1235 -3405 1241 -2629
rect 1320 -3401 1330 -2625
rect 1382 -3401 1392 -2625
rect 1471 -2629 1517 -2519
rect 1596 -2523 1606 -1747
rect 1658 -2523 1668 -1747
rect 1747 -2519 1753 -1743
rect 1787 -2519 1793 -1743
rect 1885 -1743 1931 -1731
rect 1885 -1747 1891 -1743
rect 1925 -1747 1931 -1743
rect 2023 -1743 2069 -1557
rect 1609 -2531 1655 -2523
rect 1609 -2625 1655 -2617
rect 1195 -3417 1241 -3405
rect 1333 -3405 1339 -3401
rect 1373 -3405 1379 -3401
rect 1333 -3417 1379 -3405
rect 1471 -3405 1477 -2629
rect 1511 -3405 1517 -2629
rect 1596 -3401 1606 -2625
rect 1658 -3401 1668 -2625
rect 1747 -2629 1793 -2519
rect 1872 -2523 1882 -1747
rect 1934 -2523 1944 -1747
rect 2023 -2519 2029 -1743
rect 2063 -2519 2069 -1743
rect 2161 -1743 2207 -1731
rect 2161 -1747 2167 -1743
rect 2201 -1747 2207 -1743
rect 2299 -1743 2345 -1557
rect 1885 -2531 1931 -2523
rect 1885 -2625 1931 -2617
rect 1471 -3417 1517 -3405
rect 1609 -3405 1615 -3401
rect 1649 -3405 1655 -3401
rect 1609 -3417 1655 -3405
rect 1747 -3405 1753 -2629
rect 1787 -3405 1793 -2629
rect 1872 -3401 1882 -2625
rect 1934 -3401 1944 -2625
rect 2023 -2629 2069 -2519
rect 2148 -2523 2158 -1747
rect 2210 -2523 2220 -1747
rect 2299 -2519 2305 -1743
rect 2339 -2519 2345 -1743
rect 2437 -1743 2483 -1731
rect 2437 -1747 2443 -1743
rect 2477 -1747 2483 -1743
rect 2575 -1743 2621 -1557
rect 2161 -2531 2207 -2523
rect 2161 -2625 2207 -2617
rect 1747 -3417 1793 -3405
rect 1885 -3405 1891 -3401
rect 1925 -3405 1931 -3401
rect 1885 -3417 1931 -3405
rect 2023 -3405 2029 -2629
rect 2063 -3405 2069 -2629
rect 2148 -3401 2158 -2625
rect 2210 -3401 2220 -2625
rect 2299 -2629 2345 -2519
rect 2424 -2523 2434 -1747
rect 2486 -2523 2496 -1747
rect 2575 -2519 2581 -1743
rect 2615 -2519 2621 -1743
rect 2713 -1743 2759 -1731
rect 2713 -1747 2719 -1743
rect 2753 -1747 2759 -1743
rect 2851 -1743 2897 -1557
rect 2437 -2531 2483 -2523
rect 2437 -2625 2483 -2617
rect 2023 -3417 2069 -3405
rect 2161 -3405 2167 -3401
rect 2201 -3405 2207 -3401
rect 2161 -3417 2207 -3405
rect 2299 -3405 2305 -2629
rect 2339 -3405 2345 -2629
rect 2424 -3401 2434 -2625
rect 2486 -3401 2496 -2625
rect 2575 -2629 2621 -2519
rect 2700 -2523 2710 -1747
rect 2762 -2523 2772 -1747
rect 2851 -2519 2857 -1743
rect 2891 -2519 2897 -1743
rect 2989 -1743 3035 -1731
rect 2989 -1747 2995 -1743
rect 3029 -1747 3035 -1743
rect 3127 -1743 3173 -1557
rect 2713 -2531 2759 -2523
rect 2713 -2625 2759 -2617
rect 2299 -3417 2345 -3405
rect 2437 -3405 2443 -3401
rect 2477 -3405 2483 -3401
rect 2437 -3417 2483 -3405
rect 2575 -3405 2581 -2629
rect 2615 -3405 2621 -2629
rect 2700 -3401 2710 -2625
rect 2762 -3401 2772 -2625
rect 2851 -2629 2897 -2519
rect 2976 -2523 2986 -1747
rect 3038 -2523 3048 -1747
rect 3127 -2519 3133 -1743
rect 3167 -2519 3173 -1743
rect 3265 -1743 3311 -1731
rect 3265 -1747 3271 -1743
rect 3305 -1747 3311 -1743
rect 3403 -1743 3449 -1557
rect 2989 -2531 3035 -2523
rect 2989 -2625 3035 -2617
rect 2575 -3417 2621 -3405
rect 2713 -3405 2719 -3401
rect 2753 -3405 2759 -3401
rect 2713 -3417 2759 -3405
rect 2851 -3405 2857 -2629
rect 2891 -3405 2897 -2629
rect 2976 -3401 2986 -2625
rect 3038 -3401 3048 -2625
rect 3127 -2629 3173 -2519
rect 3252 -2523 3262 -1747
rect 3314 -2523 3324 -1747
rect 3403 -2519 3409 -1743
rect 3443 -2519 3449 -1743
rect 3541 -1743 3587 -1731
rect 3541 -1747 3547 -1743
rect 3581 -1747 3587 -1743
rect 3679 -1743 3725 -1557
rect 3265 -2531 3311 -2523
rect 3265 -2625 3311 -2617
rect 2851 -3417 2897 -3405
rect 2989 -3405 2995 -3401
rect 3029 -3405 3035 -3401
rect 2989 -3417 3035 -3405
rect 3127 -3405 3133 -2629
rect 3167 -3405 3173 -2629
rect 3252 -3401 3262 -2625
rect 3314 -3401 3324 -2625
rect 3403 -2629 3449 -2519
rect 3528 -2523 3538 -1747
rect 3590 -2523 3600 -1747
rect 3679 -2519 3685 -1743
rect 3719 -2519 3725 -1743
rect 3817 -1743 3863 -1731
rect 3817 -1747 3823 -1743
rect 3857 -1747 3863 -1743
rect 3955 -1743 4001 -1557
rect 3541 -2531 3587 -2523
rect 3541 -2625 3587 -2617
rect 3127 -3417 3173 -3405
rect 3265 -3405 3271 -3401
rect 3305 -3405 3311 -3401
rect 3265 -3417 3311 -3405
rect 3403 -3405 3409 -2629
rect 3443 -3405 3449 -2629
rect 3528 -3401 3538 -2625
rect 3590 -3401 3600 -2625
rect 3679 -2629 3725 -2519
rect 3804 -2523 3814 -1747
rect 3866 -2523 3876 -1747
rect 3955 -2519 3961 -1743
rect 3995 -2519 4001 -1743
rect 4093 -1743 4139 -1731
rect 4093 -1747 4099 -1743
rect 4133 -1747 4139 -1743
rect 4231 -1743 4277 -1557
rect 3817 -2531 3863 -2523
rect 3817 -2625 3863 -2617
rect 3403 -3417 3449 -3405
rect 3541 -3405 3547 -3401
rect 3581 -3405 3587 -3401
rect 3541 -3417 3587 -3405
rect 3679 -3405 3685 -2629
rect 3719 -3405 3725 -2629
rect 3804 -3401 3814 -2625
rect 3866 -3401 3876 -2625
rect 3955 -2629 4001 -2519
rect 4080 -2523 4090 -1747
rect 4142 -2523 4152 -1747
rect 4231 -2519 4237 -1743
rect 4271 -2519 4277 -1743
rect 4369 -1743 4415 -1731
rect 4369 -1747 4375 -1743
rect 4409 -1747 4415 -1743
rect 4507 -1743 4553 -1557
rect 4093 -2531 4139 -2523
rect 4093 -2625 4139 -2617
rect 3679 -3417 3725 -3405
rect 3817 -3405 3823 -3401
rect 3857 -3405 3863 -3401
rect 3817 -3417 3863 -3405
rect 3955 -3405 3961 -2629
rect 3995 -3405 4001 -2629
rect 4080 -3401 4090 -2625
rect 4142 -3401 4152 -2625
rect 4231 -2629 4277 -2519
rect 4356 -2523 4366 -1747
rect 4418 -2523 4428 -1747
rect 4507 -2519 4513 -1743
rect 4547 -2519 4553 -1743
rect 4645 -1743 4691 -1731
rect 4645 -1747 4651 -1743
rect 4685 -1747 4691 -1743
rect 4783 -1743 4829 -1557
rect 4369 -2531 4415 -2523
rect 4369 -2625 4415 -2617
rect 3955 -3417 4001 -3405
rect 4093 -3405 4099 -3401
rect 4133 -3405 4139 -3401
rect 4093 -3417 4139 -3405
rect 4231 -3405 4237 -2629
rect 4271 -3405 4277 -2629
rect 4356 -3401 4366 -2625
rect 4418 -3401 4428 -2625
rect 4507 -2629 4553 -2519
rect 4632 -2523 4642 -1747
rect 4694 -2523 4704 -1747
rect 4783 -2519 4789 -1743
rect 4823 -2519 4829 -1743
rect 4921 -1743 4967 -1731
rect 4921 -1747 4927 -1743
rect 4961 -1747 4967 -1743
rect 5059 -1743 5105 -1557
rect 4645 -2531 4691 -2523
rect 4645 -2625 4691 -2617
rect 4231 -3417 4277 -3405
rect 4369 -3405 4375 -3401
rect 4409 -3405 4415 -3401
rect 4369 -3417 4415 -3405
rect 4507 -3405 4513 -2629
rect 4547 -3405 4553 -2629
rect 4632 -3401 4642 -2625
rect 4694 -3401 4704 -2625
rect 4783 -2629 4829 -2519
rect 4908 -2523 4918 -1747
rect 4970 -2523 4980 -1747
rect 5059 -2519 5065 -1743
rect 5099 -2519 5105 -1743
rect 5197 -1743 5243 -1731
rect 5197 -1747 5203 -1743
rect 5237 -1747 5243 -1743
rect 5335 -1743 5381 -1557
rect 4921 -2531 4967 -2523
rect 4921 -2625 4967 -2617
rect 4507 -3417 4553 -3405
rect 4645 -3405 4651 -3401
rect 4685 -3405 4691 -3401
rect 4645 -3417 4691 -3405
rect 4783 -3405 4789 -2629
rect 4823 -3405 4829 -2629
rect 4908 -3401 4918 -2625
rect 4970 -3401 4980 -2625
rect 5059 -2629 5105 -2519
rect 5184 -2523 5194 -1747
rect 5246 -2523 5256 -1747
rect 5335 -2519 5341 -1743
rect 5375 -2519 5381 -1743
rect 5473 -1743 5519 -1731
rect 5473 -1747 5479 -1743
rect 5513 -1747 5519 -1743
rect 5611 -1743 5657 -1557
rect 5197 -2531 5243 -2523
rect 5197 -2625 5243 -2617
rect 4783 -3417 4829 -3405
rect 4921 -3405 4927 -3401
rect 4961 -3405 4967 -3401
rect 4921 -3417 4967 -3405
rect 5059 -3405 5065 -2629
rect 5099 -3405 5105 -2629
rect 5184 -3401 5194 -2625
rect 5246 -3401 5256 -2625
rect 5335 -2629 5381 -2519
rect 5460 -2523 5470 -1747
rect 5522 -2523 5532 -1747
rect 5611 -2519 5617 -1743
rect 5651 -2519 5657 -1743
rect 5749 -1743 5795 -1731
rect 5749 -1747 5755 -1743
rect 5789 -1747 5795 -1743
rect 5887 -1743 5933 -1557
rect 5473 -2531 5519 -2523
rect 5473 -2625 5519 -2617
rect 5059 -3417 5105 -3405
rect 5197 -3405 5203 -3401
rect 5237 -3405 5243 -3401
rect 5197 -3417 5243 -3405
rect 5335 -3405 5341 -2629
rect 5375 -3405 5381 -2629
rect 5460 -3401 5470 -2625
rect 5522 -3401 5532 -2625
rect 5611 -2629 5657 -2519
rect 5736 -2523 5746 -1747
rect 5798 -2523 5808 -1747
rect 5887 -2519 5893 -1743
rect 5927 -2519 5933 -1743
rect 6025 -1743 6071 -1731
rect 6025 -1747 6031 -1743
rect 6065 -1747 6071 -1743
rect 6163 -1743 6209 -1557
rect 5749 -2531 5795 -2523
rect 5749 -2625 5795 -2617
rect 5335 -3417 5381 -3405
rect 5473 -3405 5479 -3401
rect 5513 -3405 5519 -3401
rect 5473 -3417 5519 -3405
rect 5611 -3405 5617 -2629
rect 5651 -3405 5657 -2629
rect 5736 -3401 5746 -2625
rect 5798 -3401 5808 -2625
rect 5887 -2629 5933 -2519
rect 6012 -2523 6022 -1747
rect 6074 -2523 6084 -1747
rect 6163 -2519 6169 -1743
rect 6203 -2519 6209 -1743
rect 6301 -1743 6347 -1731
rect 6301 -1747 6307 -1743
rect 6341 -1747 6347 -1743
rect 6439 -1743 6485 -1557
rect 6025 -2531 6071 -2523
rect 6025 -2625 6071 -2617
rect 5611 -3417 5657 -3405
rect 5749 -3405 5755 -3401
rect 5789 -3405 5795 -3401
rect 5749 -3417 5795 -3405
rect 5887 -3405 5893 -2629
rect 5927 -3405 5933 -2629
rect 6012 -3401 6022 -2625
rect 6074 -3401 6084 -2625
rect 6163 -2629 6209 -2519
rect 6288 -2523 6298 -1747
rect 6350 -2523 6360 -1747
rect 6439 -2519 6445 -1743
rect 6479 -2519 6485 -1743
rect 6577 -1743 6623 -1731
rect 6577 -1747 6583 -1743
rect 6617 -1747 6623 -1743
rect 6715 -1743 6761 -1557
rect 6301 -2531 6347 -2523
rect 6301 -2625 6347 -2617
rect 5887 -3417 5933 -3405
rect 6025 -3405 6031 -3401
rect 6065 -3405 6071 -3401
rect 6025 -3417 6071 -3405
rect 6163 -3405 6169 -2629
rect 6203 -3405 6209 -2629
rect 6288 -3401 6298 -2625
rect 6350 -3401 6360 -2625
rect 6439 -2629 6485 -2519
rect 6564 -2523 6574 -1747
rect 6626 -2523 6636 -1747
rect 6715 -2519 6721 -1743
rect 6755 -2519 6761 -1743
rect 6853 -1743 6899 -1731
rect 6853 -1747 6859 -1743
rect 6893 -1747 6899 -1743
rect 6991 -1743 7037 -1557
rect 6577 -2531 6623 -2523
rect 6577 -2625 6623 -2617
rect 6163 -3417 6209 -3405
rect 6301 -3405 6307 -3401
rect 6341 -3405 6347 -3401
rect 6301 -3417 6347 -3405
rect 6439 -3405 6445 -2629
rect 6479 -3405 6485 -2629
rect 6564 -3401 6574 -2625
rect 6626 -3401 6636 -2625
rect 6715 -2629 6761 -2519
rect 6840 -2523 6850 -1747
rect 6902 -2523 6912 -1747
rect 6991 -2519 6997 -1743
rect 7031 -2519 7037 -1743
rect 7129 -1743 7175 -1731
rect 7129 -1747 7135 -1743
rect 7169 -1747 7175 -1743
rect 7267 -1743 7313 -1557
rect 6853 -2531 6899 -2523
rect 6853 -2625 6899 -2617
rect 6439 -3417 6485 -3405
rect 6577 -3405 6583 -3401
rect 6617 -3405 6623 -3401
rect 6577 -3417 6623 -3405
rect 6715 -3405 6721 -2629
rect 6755 -3405 6761 -2629
rect 6840 -3401 6850 -2625
rect 6902 -3401 6912 -2625
rect 6991 -2629 7037 -2519
rect 7116 -2523 7126 -1747
rect 7178 -2523 7188 -1747
rect 7267 -2519 7273 -1743
rect 7307 -2519 7313 -1743
rect 7405 -1743 7451 -1731
rect 7405 -1747 7411 -1743
rect 7445 -1747 7451 -1743
rect 7543 -1743 7589 -1557
rect 7129 -2531 7175 -2523
rect 7129 -2625 7175 -2617
rect 6715 -3417 6761 -3405
rect 6853 -3405 6859 -3401
rect 6893 -3405 6899 -3401
rect 6853 -3417 6899 -3405
rect 6991 -3405 6997 -2629
rect 7031 -3405 7037 -2629
rect 7116 -3401 7126 -2625
rect 7178 -3401 7188 -2625
rect 7267 -2629 7313 -2519
rect 7392 -2523 7402 -1747
rect 7454 -2523 7464 -1747
rect 7543 -2519 7549 -1743
rect 7583 -2519 7589 -1743
rect 7681 -1743 7727 -1731
rect 7681 -1747 7687 -1743
rect 7721 -1747 7727 -1743
rect 7819 -1743 7865 -1557
rect 7405 -2531 7451 -2523
rect 7405 -2625 7451 -2617
rect 6991 -3417 7037 -3405
rect 7129 -3405 7135 -3401
rect 7169 -3405 7175 -3401
rect 7129 -3417 7175 -3405
rect 7267 -3405 7273 -2629
rect 7307 -3405 7313 -2629
rect 7392 -3401 7402 -2625
rect 7454 -3401 7464 -2625
rect 7543 -2629 7589 -2519
rect 7668 -2523 7678 -1747
rect 7730 -2523 7740 -1747
rect 7819 -2519 7825 -1743
rect 7859 -2519 7865 -1743
rect 7957 -1743 8003 -1731
rect 7957 -1747 7963 -1743
rect 7997 -1747 8003 -1743
rect 8095 -1743 8141 -1557
rect 7681 -2531 7727 -2523
rect 7681 -2625 7727 -2617
rect 7267 -3417 7313 -3405
rect 7405 -3405 7411 -3401
rect 7445 -3405 7451 -3401
rect 7405 -3417 7451 -3405
rect 7543 -3405 7549 -2629
rect 7583 -3405 7589 -2629
rect 7668 -3401 7678 -2625
rect 7730 -3401 7740 -2625
rect 7819 -2629 7865 -2519
rect 7944 -2523 7954 -1747
rect 8006 -2523 8016 -1747
rect 8095 -2519 8101 -1743
rect 8135 -2519 8141 -1743
rect 8233 -1743 8279 -1731
rect 8233 -1747 8239 -1743
rect 8273 -1747 8279 -1743
rect 8371 -1743 8417 -1557
rect 7957 -2531 8003 -2523
rect 7957 -2625 8003 -2617
rect 7543 -3417 7589 -3405
rect 7681 -3405 7687 -3401
rect 7721 -3405 7727 -3401
rect 7681 -3417 7727 -3405
rect 7819 -3405 7825 -2629
rect 7859 -3405 7865 -2629
rect 7944 -3401 7954 -2625
rect 8006 -3401 8016 -2625
rect 8095 -2629 8141 -2519
rect 8220 -2523 8230 -1747
rect 8282 -2523 8292 -1747
rect 8371 -2519 8377 -1743
rect 8411 -2519 8417 -1743
rect 8509 -1743 8555 -1731
rect 8509 -1747 8515 -1743
rect 8549 -1747 8555 -1743
rect 8647 -1743 8693 -1557
rect 8233 -2531 8279 -2523
rect 8233 -2625 8279 -2617
rect 7819 -3417 7865 -3405
rect 7957 -3405 7963 -3401
rect 7997 -3405 8003 -3401
rect 7957 -3417 8003 -3405
rect 8095 -3405 8101 -2629
rect 8135 -3405 8141 -2629
rect 8220 -3401 8230 -2625
rect 8282 -3401 8292 -2625
rect 8371 -2629 8417 -2519
rect 8496 -2523 8506 -1747
rect 8558 -2523 8568 -1747
rect 8647 -2519 8653 -1743
rect 8687 -2519 8693 -1743
rect 8785 -1743 8831 -1731
rect 8785 -1747 8791 -1743
rect 8825 -1747 8831 -1743
rect 8923 -1743 8969 -1557
rect 8509 -2531 8555 -2523
rect 8509 -2625 8555 -2617
rect 8095 -3417 8141 -3405
rect 8233 -3405 8239 -3401
rect 8273 -3405 8279 -3401
rect 8233 -3417 8279 -3405
rect 8371 -3405 8377 -2629
rect 8411 -3405 8417 -2629
rect 8496 -3401 8506 -2625
rect 8558 -3401 8568 -2625
rect 8647 -2629 8693 -2519
rect 8772 -2523 8782 -1747
rect 8834 -2523 8844 -1747
rect 8923 -2519 8929 -1743
rect 8963 -2519 8969 -1743
rect 9061 -1743 9107 -1731
rect 9061 -1747 9067 -1743
rect 9101 -1747 9107 -1743
rect 9199 -1743 9245 -1557
rect 8785 -2531 8831 -2523
rect 8785 -2625 8831 -2617
rect 8371 -3417 8417 -3405
rect 8509 -3405 8515 -3401
rect 8549 -3405 8555 -3401
rect 8509 -3417 8555 -3405
rect 8647 -3405 8653 -2629
rect 8687 -3405 8693 -2629
rect 8772 -3401 8782 -2625
rect 8834 -3401 8844 -2625
rect 8923 -2629 8969 -2519
rect 9048 -2523 9058 -1747
rect 9110 -2523 9120 -1747
rect 9199 -2519 9205 -1743
rect 9239 -2519 9245 -1743
rect 9337 -1743 9383 -1731
rect 9337 -1747 9343 -1743
rect 9377 -1747 9383 -1743
rect 9475 -1743 9521 -1557
rect 9061 -2531 9107 -2523
rect 9061 -2625 9107 -2617
rect 8647 -3417 8693 -3405
rect 8785 -3405 8791 -3401
rect 8825 -3405 8831 -3401
rect 8785 -3417 8831 -3405
rect 8923 -3405 8929 -2629
rect 8963 -3405 8969 -2629
rect 9048 -3401 9058 -2625
rect 9110 -3401 9120 -2625
rect 9199 -2629 9245 -2519
rect 9324 -2523 9334 -1747
rect 9386 -2523 9396 -1747
rect 9475 -2519 9481 -1743
rect 9515 -2519 9521 -1743
rect 9613 -1743 9659 -1731
rect 9613 -1747 9619 -1743
rect 9653 -1747 9659 -1743
rect 9751 -1743 9797 -1557
rect 9337 -2531 9383 -2523
rect 9337 -2625 9383 -2617
rect 8923 -3417 8969 -3405
rect 9061 -3405 9067 -3401
rect 9101 -3405 9107 -3401
rect 9061 -3417 9107 -3405
rect 9199 -3405 9205 -2629
rect 9239 -3405 9245 -2629
rect 9324 -3401 9334 -2625
rect 9386 -3401 9396 -2625
rect 9475 -2629 9521 -2519
rect 9600 -2523 9610 -1747
rect 9662 -2523 9672 -1747
rect 9751 -2519 9757 -1743
rect 9791 -2519 9797 -1743
rect 9889 -1743 9935 -1731
rect 9889 -1747 9895 -1743
rect 9929 -1747 9935 -1743
rect 10027 -1743 10073 -1557
rect 9613 -2531 9659 -2523
rect 9613 -2625 9659 -2617
rect 9199 -3417 9245 -3405
rect 9337 -3405 9343 -3401
rect 9377 -3405 9383 -3401
rect 9337 -3417 9383 -3405
rect 9475 -3405 9481 -2629
rect 9515 -3405 9521 -2629
rect 9600 -3401 9610 -2625
rect 9662 -3401 9672 -2625
rect 9751 -2629 9797 -2519
rect 9876 -2523 9886 -1747
rect 9938 -2523 9948 -1747
rect 10027 -2519 10033 -1743
rect 10067 -2519 10073 -1743
rect 10165 -1743 10211 -1731
rect 10165 -1747 10171 -1743
rect 10205 -1747 10211 -1743
rect 10303 -1743 10349 -1557
rect 9889 -2531 9935 -2523
rect 9889 -2625 9935 -2617
rect 9475 -3417 9521 -3405
rect 9613 -3405 9619 -3401
rect 9653 -3405 9659 -3401
rect 9613 -3417 9659 -3405
rect 9751 -3405 9757 -2629
rect 9791 -3405 9797 -2629
rect 9876 -3401 9886 -2625
rect 9938 -3401 9948 -2625
rect 10027 -2629 10073 -2519
rect 10152 -2523 10162 -1747
rect 10214 -2523 10224 -1747
rect 10303 -2519 10309 -1743
rect 10343 -2519 10349 -1743
rect 10441 -1743 10487 -1731
rect 10441 -1747 10447 -1743
rect 10481 -1747 10487 -1743
rect 10579 -1743 10625 -1557
rect 10165 -2531 10211 -2523
rect 10165 -2625 10211 -2617
rect 9751 -3417 9797 -3405
rect 9889 -3405 9895 -3401
rect 9929 -3405 9935 -3401
rect 9889 -3417 9935 -3405
rect 10027 -3405 10033 -2629
rect 10067 -3405 10073 -2629
rect 10152 -3401 10162 -2625
rect 10214 -3401 10224 -2625
rect 10303 -2629 10349 -2519
rect 10428 -2523 10438 -1747
rect 10490 -2523 10500 -1747
rect 10579 -2519 10585 -1743
rect 10619 -2519 10625 -1743
rect 10717 -1743 10763 -1731
rect 10717 -1747 10723 -1743
rect 10757 -1747 10763 -1743
rect 10855 -1743 10901 -1557
rect 10441 -2531 10487 -2523
rect 10441 -2625 10487 -2617
rect 10027 -3417 10073 -3405
rect 10165 -3405 10171 -3401
rect 10205 -3405 10211 -3401
rect 10165 -3417 10211 -3405
rect 10303 -3405 10309 -2629
rect 10343 -3405 10349 -2629
rect 10428 -3401 10438 -2625
rect 10490 -3401 10500 -2625
rect 10579 -2629 10625 -2519
rect 10704 -2523 10714 -1747
rect 10766 -2523 10776 -1747
rect 10855 -2519 10861 -1743
rect 10895 -2519 10901 -1743
rect 10993 -1743 11039 -1731
rect 10993 -1747 10999 -1743
rect 11033 -1747 11039 -1743
rect 11131 -1743 11177 -1557
rect 10717 -2531 10763 -2523
rect 10717 -2625 10763 -2617
rect 10303 -3417 10349 -3405
rect 10441 -3405 10447 -3401
rect 10481 -3405 10487 -3401
rect 10441 -3417 10487 -3405
rect 10579 -3405 10585 -2629
rect 10619 -3405 10625 -2629
rect 10704 -3401 10714 -2625
rect 10766 -3401 10776 -2625
rect 10855 -2629 10901 -2519
rect 10980 -2523 10990 -1747
rect 11042 -2523 11052 -1747
rect 11131 -2519 11137 -1743
rect 11171 -2519 11177 -1743
rect 11269 -1743 11315 -1731
rect 11269 -1747 11275 -1743
rect 11309 -1747 11315 -1743
rect 11407 -1743 11453 -1557
rect 10993 -2531 11039 -2523
rect 10993 -2625 11039 -2617
rect 10579 -3417 10625 -3405
rect 10717 -3405 10723 -3401
rect 10757 -3405 10763 -3401
rect 10717 -3417 10763 -3405
rect 10855 -3405 10861 -2629
rect 10895 -3405 10901 -2629
rect 10980 -3401 10990 -2625
rect 11042 -3401 11052 -2625
rect 11131 -2629 11177 -2519
rect 11256 -2523 11266 -1747
rect 11318 -2523 11328 -1747
rect 11407 -2519 11413 -1743
rect 11447 -2519 11453 -1743
rect 11545 -1743 11591 -1731
rect 11545 -1747 11551 -1743
rect 11585 -1747 11591 -1743
rect 11683 -1743 11729 -1557
rect 11269 -2531 11315 -2523
rect 11269 -2625 11315 -2617
rect 10855 -3417 10901 -3405
rect 10993 -3405 10999 -3401
rect 11033 -3405 11039 -3401
rect 10993 -3417 11039 -3405
rect 11131 -3405 11137 -2629
rect 11171 -3405 11177 -2629
rect 11256 -3401 11266 -2625
rect 11318 -3401 11328 -2625
rect 11407 -2629 11453 -2519
rect 11532 -2523 11542 -1747
rect 11594 -2523 11604 -1747
rect 11683 -2519 11689 -1743
rect 11723 -2519 11729 -1743
rect 11821 -1743 11867 -1731
rect 11821 -1747 11827 -1743
rect 11861 -1747 11867 -1743
rect 11959 -1743 12005 -1557
rect 11545 -2531 11591 -2523
rect 11545 -2625 11591 -2617
rect 11131 -3417 11177 -3405
rect 11269 -3405 11275 -3401
rect 11309 -3405 11315 -3401
rect 11269 -3417 11315 -3405
rect 11407 -3405 11413 -2629
rect 11447 -3405 11453 -2629
rect 11532 -3401 11542 -2625
rect 11594 -3401 11604 -2625
rect 11683 -2629 11729 -2519
rect 11808 -2523 11818 -1747
rect 11870 -2523 11880 -1747
rect 11959 -2519 11965 -1743
rect 11999 -2519 12005 -1743
rect 12097 -1743 12143 -1731
rect 12097 -1747 12103 -1743
rect 12137 -1747 12143 -1743
rect 12235 -1743 12281 -1557
rect 11821 -2531 11867 -2523
rect 11821 -2625 11867 -2617
rect 11407 -3417 11453 -3405
rect 11545 -3405 11551 -3401
rect 11585 -3405 11591 -3401
rect 11545 -3417 11591 -3405
rect 11683 -3405 11689 -2629
rect 11723 -3405 11729 -2629
rect 11808 -3401 11818 -2625
rect 11870 -3401 11880 -2625
rect 11959 -2629 12005 -2519
rect 12084 -2523 12094 -1747
rect 12146 -2523 12156 -1747
rect 12235 -2519 12241 -1743
rect 12275 -2519 12281 -1743
rect 12373 -1743 12419 -1731
rect 12373 -1747 12379 -1743
rect 12413 -1747 12419 -1743
rect 12511 -1743 12557 -1557
rect 12097 -2531 12143 -2523
rect 12097 -2625 12143 -2617
rect 11683 -3417 11729 -3405
rect 11821 -3405 11827 -3401
rect 11861 -3405 11867 -3401
rect 11821 -3417 11867 -3405
rect 11959 -3405 11965 -2629
rect 11999 -3405 12005 -2629
rect 12084 -3401 12094 -2625
rect 12146 -3401 12156 -2625
rect 12235 -2629 12281 -2519
rect 12360 -2523 12370 -1747
rect 12422 -2523 12432 -1747
rect 12511 -2519 12517 -1743
rect 12551 -2519 12557 -1743
rect 12649 -1743 12695 -1731
rect 12649 -1747 12655 -1743
rect 12689 -1747 12695 -1743
rect 12787 -1743 12833 -1557
rect 12373 -2531 12419 -2523
rect 12373 -2625 12419 -2617
rect 11959 -3417 12005 -3405
rect 12097 -3405 12103 -3401
rect 12137 -3405 12143 -3401
rect 12097 -3417 12143 -3405
rect 12235 -3405 12241 -2629
rect 12275 -3405 12281 -2629
rect 12360 -3401 12370 -2625
rect 12422 -3401 12432 -2625
rect 12511 -2629 12557 -2519
rect 12636 -2523 12646 -1747
rect 12698 -2523 12708 -1747
rect 12787 -2519 12793 -1743
rect 12827 -2519 12833 -1743
rect 12925 -1743 12971 -1731
rect 12925 -1747 12931 -1743
rect 12965 -1747 12971 -1743
rect 13063 -1743 13109 -1557
rect 12649 -2531 12695 -2523
rect 12649 -2625 12695 -2617
rect 12235 -3417 12281 -3405
rect 12373 -3405 12379 -3401
rect 12413 -3405 12419 -3401
rect 12373 -3417 12419 -3405
rect 12511 -3405 12517 -2629
rect 12551 -3405 12557 -2629
rect 12636 -3401 12646 -2625
rect 12698 -3401 12708 -2625
rect 12787 -2629 12833 -2519
rect 12912 -2523 12922 -1747
rect 12974 -2523 12984 -1747
rect 13063 -2519 13069 -1743
rect 13103 -2519 13109 -1743
rect 13201 -1743 13247 -1731
rect 13201 -1747 13207 -1743
rect 13241 -1747 13247 -1743
rect 13339 -1743 13385 -1557
rect 12925 -2531 12971 -2523
rect 12925 -2625 12971 -2617
rect 12511 -3417 12557 -3405
rect 12649 -3405 12655 -3401
rect 12689 -3405 12695 -3401
rect 12649 -3417 12695 -3405
rect 12787 -3405 12793 -2629
rect 12827 -3405 12833 -2629
rect 12912 -3401 12922 -2625
rect 12974 -3401 12984 -2625
rect 13063 -2629 13109 -2519
rect 13188 -2523 13198 -1747
rect 13250 -2523 13260 -1747
rect 13339 -2519 13345 -1743
rect 13379 -2519 13385 -1743
rect 13477 -1743 13523 -1731
rect 13477 -1747 13483 -1743
rect 13517 -1747 13523 -1743
rect 13615 -1743 13661 -1557
rect 13201 -2531 13247 -2523
rect 13201 -2625 13247 -2617
rect 12787 -3417 12833 -3405
rect 12925 -3405 12931 -3401
rect 12965 -3405 12971 -3401
rect 12925 -3417 12971 -3405
rect 13063 -3405 13069 -2629
rect 13103 -3405 13109 -2629
rect 13188 -3401 13198 -2625
rect 13250 -3401 13260 -2625
rect 13339 -2629 13385 -2519
rect 13464 -2523 13474 -1747
rect 13526 -2523 13536 -1747
rect 13615 -2519 13621 -1743
rect 13655 -2519 13661 -1743
rect 13753 -1743 13799 -1731
rect 13753 -1747 13759 -1743
rect 13793 -1747 13799 -1743
rect 13891 -1743 13937 -1557
rect 13477 -2531 13523 -2523
rect 13477 -2625 13523 -2617
rect 13063 -3417 13109 -3405
rect 13201 -3405 13207 -3401
rect 13241 -3405 13247 -3401
rect 13201 -3417 13247 -3405
rect 13339 -3405 13345 -2629
rect 13379 -3405 13385 -2629
rect 13464 -3401 13474 -2625
rect 13526 -3401 13536 -2625
rect 13615 -2629 13661 -2519
rect 13740 -2523 13750 -1747
rect 13802 -2523 13812 -1747
rect 13891 -2519 13897 -1743
rect 13931 -2519 13937 -1743
rect 13753 -2531 13799 -2523
rect 13753 -2625 13799 -2617
rect 13339 -3417 13385 -3405
rect 13477 -3405 13483 -3401
rect 13517 -3405 13523 -3401
rect 13477 -3417 13523 -3405
rect 13615 -3405 13621 -2629
rect 13655 -3405 13661 -2629
rect 13740 -3401 13750 -2625
rect 13802 -3401 13812 -2625
rect 13891 -2629 13937 -2519
rect 13615 -3417 13661 -3405
rect 13753 -3405 13759 -3401
rect 13793 -3405 13799 -3401
rect 13753 -3417 13799 -3405
rect 13891 -3405 13897 -2629
rect 13931 -3405 13937 -2629
rect 13891 -3417 13937 -3405
rect 147 -3464 13881 -3454
rect 147 -3498 159 -3464
rect 207 -3498 297 -3464
rect 345 -3498 435 -3464
rect 483 -3498 573 -3464
rect 621 -3498 711 -3464
rect 759 -3498 849 -3464
rect 897 -3498 987 -3464
rect 1035 -3498 1125 -3464
rect 1173 -3498 1263 -3464
rect 1311 -3498 1401 -3464
rect 1449 -3498 1539 -3464
rect 1587 -3498 1677 -3464
rect 1725 -3498 1815 -3464
rect 1863 -3498 1953 -3464
rect 2001 -3498 2091 -3464
rect 2139 -3498 2229 -3464
rect 2277 -3498 2367 -3464
rect 2415 -3498 2505 -3464
rect 2553 -3498 2643 -3464
rect 2691 -3498 2781 -3464
rect 2829 -3498 2919 -3464
rect 2967 -3498 3057 -3464
rect 3105 -3498 3195 -3464
rect 3243 -3498 3333 -3464
rect 3381 -3498 3471 -3464
rect 3519 -3498 3609 -3464
rect 3657 -3498 3747 -3464
rect 3795 -3498 3885 -3464
rect 3933 -3498 4023 -3464
rect 4071 -3498 4161 -3464
rect 4209 -3498 4299 -3464
rect 4347 -3498 4437 -3464
rect 4485 -3498 4575 -3464
rect 4623 -3498 4713 -3464
rect 4761 -3498 4851 -3464
rect 4899 -3498 4989 -3464
rect 5037 -3498 5127 -3464
rect 5175 -3498 5265 -3464
rect 5313 -3498 5403 -3464
rect 5451 -3498 5541 -3464
rect 5589 -3498 5679 -3464
rect 5727 -3498 5817 -3464
rect 5865 -3498 5955 -3464
rect 6003 -3498 6093 -3464
rect 6141 -3498 6231 -3464
rect 6279 -3498 6369 -3464
rect 6417 -3498 6507 -3464
rect 6555 -3498 6645 -3464
rect 6693 -3498 6783 -3464
rect 6831 -3498 6921 -3464
rect 6969 -3498 7059 -3464
rect 7107 -3498 7197 -3464
rect 7245 -3498 7335 -3464
rect 7383 -3498 7473 -3464
rect 7521 -3498 7611 -3464
rect 7659 -3498 7749 -3464
rect 7797 -3498 7887 -3464
rect 7935 -3498 8025 -3464
rect 8073 -3498 8163 -3464
rect 8211 -3498 8301 -3464
rect 8349 -3498 8439 -3464
rect 8487 -3498 8577 -3464
rect 8625 -3498 8715 -3464
rect 8763 -3498 8853 -3464
rect 8901 -3498 8991 -3464
rect 9039 -3498 9129 -3464
rect 9177 -3498 9267 -3464
rect 9315 -3498 9405 -3464
rect 9453 -3498 9543 -3464
rect 9591 -3498 9681 -3464
rect 9729 -3498 9819 -3464
rect 9867 -3498 9957 -3464
rect 10005 -3498 10095 -3464
rect 10143 -3498 10233 -3464
rect 10281 -3498 10371 -3464
rect 10419 -3498 10509 -3464
rect 10557 -3498 10647 -3464
rect 10695 -3498 10785 -3464
rect 10833 -3498 10923 -3464
rect 10971 -3498 11061 -3464
rect 11109 -3498 11199 -3464
rect 11247 -3498 11337 -3464
rect 11385 -3498 11475 -3464
rect 11523 -3498 11613 -3464
rect 11661 -3498 11751 -3464
rect 11799 -3498 11889 -3464
rect 11937 -3498 12027 -3464
rect 12075 -3498 12165 -3464
rect 12213 -3498 12303 -3464
rect 12351 -3498 12441 -3464
rect 12489 -3498 12579 -3464
rect 12627 -3498 12717 -3464
rect 12765 -3498 12855 -3464
rect 12903 -3498 12993 -3464
rect 13041 -3498 13131 -3464
rect 13179 -3498 13269 -3464
rect 13317 -3498 13407 -3464
rect 13455 -3498 13545 -3464
rect 13593 -3498 13683 -3464
rect 13731 -3498 13821 -3464
rect 13869 -3498 13881 -3464
rect 147 -3500 13881 -3498
rect 147 -3504 219 -3500
rect 285 -3504 495 -3500
rect 561 -3504 633 -3500
rect 699 -3504 771 -3500
rect 837 -3504 1047 -3500
rect 1113 -3504 1185 -3500
rect 1251 -3504 1323 -3500
rect 1389 -3504 1599 -3500
rect 1665 -3504 1737 -3500
rect 1803 -3504 1875 -3500
rect 1941 -3504 2151 -3500
rect 2217 -3504 2289 -3500
rect 2355 -3504 2427 -3500
rect 2493 -3504 2703 -3500
rect 2769 -3504 2841 -3500
rect 2907 -3504 2979 -3500
rect 3045 -3504 3255 -3500
rect 3321 -3504 3393 -3500
rect 3459 -3504 3531 -3500
rect 3597 -3504 3807 -3500
rect 3873 -3504 3945 -3500
rect 4011 -3504 4083 -3500
rect 4149 -3504 4359 -3500
rect 4425 -3504 4497 -3500
rect 4563 -3504 4635 -3500
rect 4701 -3504 4911 -3500
rect 4977 -3504 5049 -3500
rect 5115 -3504 5187 -3500
rect 5253 -3504 5463 -3500
rect 5529 -3504 5601 -3500
rect 5667 -3504 5739 -3500
rect 5805 -3504 6015 -3500
rect 6081 -3504 6153 -3500
rect 6219 -3504 6291 -3500
rect 6357 -3504 6567 -3500
rect 6633 -3504 6705 -3500
rect 6771 -3504 6843 -3500
rect 6909 -3504 7119 -3500
rect 7185 -3504 7257 -3500
rect 7323 -3504 7395 -3500
rect 7461 -3504 7671 -3500
rect 7737 -3504 7809 -3500
rect 7875 -3504 7947 -3500
rect 8013 -3504 8223 -3500
rect 8289 -3504 8361 -3500
rect 8427 -3504 8499 -3500
rect 8565 -3504 8775 -3500
rect 8841 -3504 8913 -3500
rect 8979 -3504 9051 -3500
rect 9117 -3504 9327 -3500
rect 9393 -3504 9465 -3500
rect 9531 -3504 9603 -3500
rect 9669 -3504 9879 -3500
rect 9945 -3504 10017 -3500
rect 10083 -3504 10155 -3500
rect 10221 -3504 10431 -3500
rect 10497 -3504 10569 -3500
rect 10635 -3504 10707 -3500
rect 10773 -3504 10983 -3500
rect 11049 -3504 11121 -3500
rect 11187 -3504 11259 -3500
rect 11325 -3504 11535 -3500
rect 11601 -3504 11673 -3500
rect 11739 -3504 11811 -3500
rect 11877 -3504 12087 -3500
rect 12153 -3504 12225 -3500
rect 12291 -3504 12363 -3500
rect 12429 -3504 12639 -3500
rect 12705 -3504 12777 -3500
rect 12843 -3504 12915 -3500
rect 12981 -3504 13191 -3500
rect 13257 -3504 13329 -3500
rect 13395 -3504 13467 -3500
rect 13533 -3504 13743 -3500
rect 13809 -3504 13881 -3500
rect 297 -3893 483 -3504
rect 849 -3893 1035 -3504
rect 1401 -3893 1587 -3504
rect 1953 -3893 2139 -3504
rect 2505 -3893 2691 -3504
rect 3057 -3893 3243 -3504
rect 3609 -3893 3795 -3504
rect 4161 -3893 4347 -3504
rect 4713 -3893 4899 -3504
rect 5265 -3893 5451 -3504
rect 5817 -3893 6003 -3504
rect 6369 -3893 6555 -3504
rect 6921 -3893 7107 -3504
rect 7473 -3893 7659 -3504
rect 8025 -3893 8211 -3504
rect 8577 -3893 8763 -3504
rect 9129 -3893 9315 -3504
rect 9681 -3893 9867 -3504
rect 10233 -3893 10419 -3504
rect 10785 -3893 10971 -3504
rect 11337 -3893 11523 -3504
rect 11889 -3893 12075 -3504
rect 12441 -3893 12627 -3504
rect 12993 -3893 13179 -3504
rect 13545 -3893 13731 -3504
rect 297 -4079 13731 -3893
rect 1587 -4772 1952 -4079
rect 3795 -4772 4160 -4079
rect 6003 -4772 6368 -4079
rect 8211 -4772 8576 -4079
rect 10419 -4772 10784 -4079
rect 12627 -4772 12992 -4079
rect 1586 -5419 12997 -4772
rect 4664 -7188 5546 -5419
rect 9049 -7188 9931 -5419
rect 4664 -7219 9931 -7188
rect 4664 -8030 6583 -7219
rect 8032 -8030 9931 -7219
rect 4664 -8069 9931 -8030
<< via1 >>
rect 6583 4701 8032 5512
rect 226 107 278 883
rect 226 -771 278 5
rect 502 107 554 883
rect 502 -771 554 5
rect 778 107 830 883
rect 778 -771 830 5
rect 1054 107 1106 883
rect 1054 -771 1106 5
rect 1330 107 1382 883
rect 1330 -771 1382 5
rect 1606 107 1658 883
rect 1606 -771 1658 5
rect 1882 107 1934 883
rect 1882 -771 1934 5
rect 2158 107 2210 883
rect 2158 -771 2210 5
rect 2434 107 2486 883
rect 2434 -771 2486 5
rect 2710 107 2762 883
rect 2710 -771 2762 5
rect 2986 107 3038 883
rect 2986 -771 3038 5
rect 3262 107 3314 883
rect 3262 -771 3314 5
rect 3538 107 3590 883
rect 3538 -771 3590 5
rect 3814 107 3866 883
rect 3814 -771 3866 5
rect 4090 107 4142 883
rect 4090 -771 4142 5
rect 4366 107 4418 883
rect 4366 -771 4418 5
rect 4642 107 4694 883
rect 4642 -771 4694 5
rect 4918 107 4970 883
rect 4918 -771 4970 5
rect 5194 107 5246 883
rect 5194 -771 5246 5
rect 5470 107 5522 883
rect 5470 -771 5522 5
rect 5746 107 5798 883
rect 5746 -771 5798 5
rect 6022 107 6074 883
rect 6022 -771 6074 5
rect 6298 107 6350 883
rect 6298 -771 6350 5
rect 6574 107 6626 883
rect 6574 -771 6626 5
rect 6850 107 6902 883
rect 6850 -771 6902 5
rect 7126 107 7178 883
rect 7126 -771 7178 5
rect 7402 107 7454 883
rect 7402 -771 7454 5
rect 7678 107 7730 883
rect 7678 -771 7730 5
rect 7954 107 8006 883
rect 7954 -771 8006 5
rect 8230 107 8282 883
rect 8230 -771 8282 5
rect 8506 107 8558 883
rect 8506 -771 8558 5
rect 8782 107 8834 883
rect 8782 -771 8834 5
rect 9058 107 9110 883
rect 9058 -771 9110 5
rect 9334 107 9386 883
rect 9334 -771 9386 5
rect 9610 107 9662 883
rect 9610 -771 9662 5
rect 9886 107 9938 883
rect 9886 -771 9938 5
rect 10162 107 10214 883
rect 10162 -771 10214 5
rect 10438 107 10490 883
rect 10438 -771 10490 5
rect 10714 107 10766 883
rect 10714 -771 10766 5
rect 10990 107 11042 883
rect 10990 -771 11042 5
rect 11266 107 11318 883
rect 11266 -771 11318 5
rect 11542 107 11594 883
rect 11542 -771 11594 5
rect 11818 107 11870 883
rect 11818 -771 11870 5
rect 12094 107 12146 883
rect 12094 -771 12146 5
rect 12370 107 12422 883
rect 12370 -771 12422 5
rect 12646 107 12698 883
rect 12646 -771 12698 5
rect 12922 107 12974 883
rect 12922 -771 12974 5
rect 13198 107 13250 883
rect 13198 -771 13250 5
rect 13474 107 13526 883
rect 13474 -771 13526 5
rect 13750 107 13802 883
rect 13750 -771 13802 5
rect -840 -1540 -300 -990
rect 226 -2519 235 -1747
rect 235 -2519 269 -1747
rect 269 -2519 278 -1747
rect 226 -2523 278 -2519
rect 226 -2629 278 -2625
rect 226 -3401 235 -2629
rect 235 -3401 269 -2629
rect 269 -3401 278 -2629
rect 502 -2519 511 -1747
rect 511 -2519 545 -1747
rect 545 -2519 554 -1747
rect 502 -2523 554 -2519
rect 502 -2629 554 -2625
rect 502 -3401 511 -2629
rect 511 -3401 545 -2629
rect 545 -3401 554 -2629
rect 778 -2519 787 -1747
rect 787 -2519 821 -1747
rect 821 -2519 830 -1747
rect 778 -2523 830 -2519
rect 778 -2629 830 -2625
rect 778 -3401 787 -2629
rect 787 -3401 821 -2629
rect 821 -3401 830 -2629
rect 1054 -2519 1063 -1747
rect 1063 -2519 1097 -1747
rect 1097 -2519 1106 -1747
rect 1054 -2523 1106 -2519
rect 1054 -2629 1106 -2625
rect 1054 -3401 1063 -2629
rect 1063 -3401 1097 -2629
rect 1097 -3401 1106 -2629
rect 1330 -2519 1339 -1747
rect 1339 -2519 1373 -1747
rect 1373 -2519 1382 -1747
rect 1330 -2523 1382 -2519
rect 1330 -2629 1382 -2625
rect 1330 -3401 1339 -2629
rect 1339 -3401 1373 -2629
rect 1373 -3401 1382 -2629
rect 1606 -2519 1615 -1747
rect 1615 -2519 1649 -1747
rect 1649 -2519 1658 -1747
rect 1606 -2523 1658 -2519
rect 1606 -2629 1658 -2625
rect 1606 -3401 1615 -2629
rect 1615 -3401 1649 -2629
rect 1649 -3401 1658 -2629
rect 1882 -2519 1891 -1747
rect 1891 -2519 1925 -1747
rect 1925 -2519 1934 -1747
rect 1882 -2523 1934 -2519
rect 1882 -2629 1934 -2625
rect 1882 -3401 1891 -2629
rect 1891 -3401 1925 -2629
rect 1925 -3401 1934 -2629
rect 2158 -2519 2167 -1747
rect 2167 -2519 2201 -1747
rect 2201 -2519 2210 -1747
rect 2158 -2523 2210 -2519
rect 2158 -2629 2210 -2625
rect 2158 -3401 2167 -2629
rect 2167 -3401 2201 -2629
rect 2201 -3401 2210 -2629
rect 2434 -2519 2443 -1747
rect 2443 -2519 2477 -1747
rect 2477 -2519 2486 -1747
rect 2434 -2523 2486 -2519
rect 2434 -2629 2486 -2625
rect 2434 -3401 2443 -2629
rect 2443 -3401 2477 -2629
rect 2477 -3401 2486 -2629
rect 2710 -2519 2719 -1747
rect 2719 -2519 2753 -1747
rect 2753 -2519 2762 -1747
rect 2710 -2523 2762 -2519
rect 2710 -2629 2762 -2625
rect 2710 -3401 2719 -2629
rect 2719 -3401 2753 -2629
rect 2753 -3401 2762 -2629
rect 2986 -2519 2995 -1747
rect 2995 -2519 3029 -1747
rect 3029 -2519 3038 -1747
rect 2986 -2523 3038 -2519
rect 2986 -2629 3038 -2625
rect 2986 -3401 2995 -2629
rect 2995 -3401 3029 -2629
rect 3029 -3401 3038 -2629
rect 3262 -2519 3271 -1747
rect 3271 -2519 3305 -1747
rect 3305 -2519 3314 -1747
rect 3262 -2523 3314 -2519
rect 3262 -2629 3314 -2625
rect 3262 -3401 3271 -2629
rect 3271 -3401 3305 -2629
rect 3305 -3401 3314 -2629
rect 3538 -2519 3547 -1747
rect 3547 -2519 3581 -1747
rect 3581 -2519 3590 -1747
rect 3538 -2523 3590 -2519
rect 3538 -2629 3590 -2625
rect 3538 -3401 3547 -2629
rect 3547 -3401 3581 -2629
rect 3581 -3401 3590 -2629
rect 3814 -2519 3823 -1747
rect 3823 -2519 3857 -1747
rect 3857 -2519 3866 -1747
rect 3814 -2523 3866 -2519
rect 3814 -2629 3866 -2625
rect 3814 -3401 3823 -2629
rect 3823 -3401 3857 -2629
rect 3857 -3401 3866 -2629
rect 4090 -2519 4099 -1747
rect 4099 -2519 4133 -1747
rect 4133 -2519 4142 -1747
rect 4090 -2523 4142 -2519
rect 4090 -2629 4142 -2625
rect 4090 -3401 4099 -2629
rect 4099 -3401 4133 -2629
rect 4133 -3401 4142 -2629
rect 4366 -2519 4375 -1747
rect 4375 -2519 4409 -1747
rect 4409 -2519 4418 -1747
rect 4366 -2523 4418 -2519
rect 4366 -2629 4418 -2625
rect 4366 -3401 4375 -2629
rect 4375 -3401 4409 -2629
rect 4409 -3401 4418 -2629
rect 4642 -2519 4651 -1747
rect 4651 -2519 4685 -1747
rect 4685 -2519 4694 -1747
rect 4642 -2523 4694 -2519
rect 4642 -2629 4694 -2625
rect 4642 -3401 4651 -2629
rect 4651 -3401 4685 -2629
rect 4685 -3401 4694 -2629
rect 4918 -2519 4927 -1747
rect 4927 -2519 4961 -1747
rect 4961 -2519 4970 -1747
rect 4918 -2523 4970 -2519
rect 4918 -2629 4970 -2625
rect 4918 -3401 4927 -2629
rect 4927 -3401 4961 -2629
rect 4961 -3401 4970 -2629
rect 5194 -2519 5203 -1747
rect 5203 -2519 5237 -1747
rect 5237 -2519 5246 -1747
rect 5194 -2523 5246 -2519
rect 5194 -2629 5246 -2625
rect 5194 -3401 5203 -2629
rect 5203 -3401 5237 -2629
rect 5237 -3401 5246 -2629
rect 5470 -2519 5479 -1747
rect 5479 -2519 5513 -1747
rect 5513 -2519 5522 -1747
rect 5470 -2523 5522 -2519
rect 5470 -2629 5522 -2625
rect 5470 -3401 5479 -2629
rect 5479 -3401 5513 -2629
rect 5513 -3401 5522 -2629
rect 5746 -2519 5755 -1747
rect 5755 -2519 5789 -1747
rect 5789 -2519 5798 -1747
rect 5746 -2523 5798 -2519
rect 5746 -2629 5798 -2625
rect 5746 -3401 5755 -2629
rect 5755 -3401 5789 -2629
rect 5789 -3401 5798 -2629
rect 6022 -2519 6031 -1747
rect 6031 -2519 6065 -1747
rect 6065 -2519 6074 -1747
rect 6022 -2523 6074 -2519
rect 6022 -2629 6074 -2625
rect 6022 -3401 6031 -2629
rect 6031 -3401 6065 -2629
rect 6065 -3401 6074 -2629
rect 6298 -2519 6307 -1747
rect 6307 -2519 6341 -1747
rect 6341 -2519 6350 -1747
rect 6298 -2523 6350 -2519
rect 6298 -2629 6350 -2625
rect 6298 -3401 6307 -2629
rect 6307 -3401 6341 -2629
rect 6341 -3401 6350 -2629
rect 6574 -2519 6583 -1747
rect 6583 -2519 6617 -1747
rect 6617 -2519 6626 -1747
rect 6574 -2523 6626 -2519
rect 6574 -2629 6626 -2625
rect 6574 -3401 6583 -2629
rect 6583 -3401 6617 -2629
rect 6617 -3401 6626 -2629
rect 6850 -2519 6859 -1747
rect 6859 -2519 6893 -1747
rect 6893 -2519 6902 -1747
rect 6850 -2523 6902 -2519
rect 6850 -2629 6902 -2625
rect 6850 -3401 6859 -2629
rect 6859 -3401 6893 -2629
rect 6893 -3401 6902 -2629
rect 7126 -2519 7135 -1747
rect 7135 -2519 7169 -1747
rect 7169 -2519 7178 -1747
rect 7126 -2523 7178 -2519
rect 7126 -2629 7178 -2625
rect 7126 -3401 7135 -2629
rect 7135 -3401 7169 -2629
rect 7169 -3401 7178 -2629
rect 7402 -2519 7411 -1747
rect 7411 -2519 7445 -1747
rect 7445 -2519 7454 -1747
rect 7402 -2523 7454 -2519
rect 7402 -2629 7454 -2625
rect 7402 -3401 7411 -2629
rect 7411 -3401 7445 -2629
rect 7445 -3401 7454 -2629
rect 7678 -2519 7687 -1747
rect 7687 -2519 7721 -1747
rect 7721 -2519 7730 -1747
rect 7678 -2523 7730 -2519
rect 7678 -2629 7730 -2625
rect 7678 -3401 7687 -2629
rect 7687 -3401 7721 -2629
rect 7721 -3401 7730 -2629
rect 7954 -2519 7963 -1747
rect 7963 -2519 7997 -1747
rect 7997 -2519 8006 -1747
rect 7954 -2523 8006 -2519
rect 7954 -2629 8006 -2625
rect 7954 -3401 7963 -2629
rect 7963 -3401 7997 -2629
rect 7997 -3401 8006 -2629
rect 8230 -2519 8239 -1747
rect 8239 -2519 8273 -1747
rect 8273 -2519 8282 -1747
rect 8230 -2523 8282 -2519
rect 8230 -2629 8282 -2625
rect 8230 -3401 8239 -2629
rect 8239 -3401 8273 -2629
rect 8273 -3401 8282 -2629
rect 8506 -2519 8515 -1747
rect 8515 -2519 8549 -1747
rect 8549 -2519 8558 -1747
rect 8506 -2523 8558 -2519
rect 8506 -2629 8558 -2625
rect 8506 -3401 8515 -2629
rect 8515 -3401 8549 -2629
rect 8549 -3401 8558 -2629
rect 8782 -2519 8791 -1747
rect 8791 -2519 8825 -1747
rect 8825 -2519 8834 -1747
rect 8782 -2523 8834 -2519
rect 8782 -2629 8834 -2625
rect 8782 -3401 8791 -2629
rect 8791 -3401 8825 -2629
rect 8825 -3401 8834 -2629
rect 9058 -2519 9067 -1747
rect 9067 -2519 9101 -1747
rect 9101 -2519 9110 -1747
rect 9058 -2523 9110 -2519
rect 9058 -2629 9110 -2625
rect 9058 -3401 9067 -2629
rect 9067 -3401 9101 -2629
rect 9101 -3401 9110 -2629
rect 9334 -2519 9343 -1747
rect 9343 -2519 9377 -1747
rect 9377 -2519 9386 -1747
rect 9334 -2523 9386 -2519
rect 9334 -2629 9386 -2625
rect 9334 -3401 9343 -2629
rect 9343 -3401 9377 -2629
rect 9377 -3401 9386 -2629
rect 9610 -2519 9619 -1747
rect 9619 -2519 9653 -1747
rect 9653 -2519 9662 -1747
rect 9610 -2523 9662 -2519
rect 9610 -2629 9662 -2625
rect 9610 -3401 9619 -2629
rect 9619 -3401 9653 -2629
rect 9653 -3401 9662 -2629
rect 9886 -2519 9895 -1747
rect 9895 -2519 9929 -1747
rect 9929 -2519 9938 -1747
rect 9886 -2523 9938 -2519
rect 9886 -2629 9938 -2625
rect 9886 -3401 9895 -2629
rect 9895 -3401 9929 -2629
rect 9929 -3401 9938 -2629
rect 10162 -2519 10171 -1747
rect 10171 -2519 10205 -1747
rect 10205 -2519 10214 -1747
rect 10162 -2523 10214 -2519
rect 10162 -2629 10214 -2625
rect 10162 -3401 10171 -2629
rect 10171 -3401 10205 -2629
rect 10205 -3401 10214 -2629
rect 10438 -2519 10447 -1747
rect 10447 -2519 10481 -1747
rect 10481 -2519 10490 -1747
rect 10438 -2523 10490 -2519
rect 10438 -2629 10490 -2625
rect 10438 -3401 10447 -2629
rect 10447 -3401 10481 -2629
rect 10481 -3401 10490 -2629
rect 10714 -2519 10723 -1747
rect 10723 -2519 10757 -1747
rect 10757 -2519 10766 -1747
rect 10714 -2523 10766 -2519
rect 10714 -2629 10766 -2625
rect 10714 -3401 10723 -2629
rect 10723 -3401 10757 -2629
rect 10757 -3401 10766 -2629
rect 10990 -2519 10999 -1747
rect 10999 -2519 11033 -1747
rect 11033 -2519 11042 -1747
rect 10990 -2523 11042 -2519
rect 10990 -2629 11042 -2625
rect 10990 -3401 10999 -2629
rect 10999 -3401 11033 -2629
rect 11033 -3401 11042 -2629
rect 11266 -2519 11275 -1747
rect 11275 -2519 11309 -1747
rect 11309 -2519 11318 -1747
rect 11266 -2523 11318 -2519
rect 11266 -2629 11318 -2625
rect 11266 -3401 11275 -2629
rect 11275 -3401 11309 -2629
rect 11309 -3401 11318 -2629
rect 11542 -2519 11551 -1747
rect 11551 -2519 11585 -1747
rect 11585 -2519 11594 -1747
rect 11542 -2523 11594 -2519
rect 11542 -2629 11594 -2625
rect 11542 -3401 11551 -2629
rect 11551 -3401 11585 -2629
rect 11585 -3401 11594 -2629
rect 11818 -2519 11827 -1747
rect 11827 -2519 11861 -1747
rect 11861 -2519 11870 -1747
rect 11818 -2523 11870 -2519
rect 11818 -2629 11870 -2625
rect 11818 -3401 11827 -2629
rect 11827 -3401 11861 -2629
rect 11861 -3401 11870 -2629
rect 12094 -2519 12103 -1747
rect 12103 -2519 12137 -1747
rect 12137 -2519 12146 -1747
rect 12094 -2523 12146 -2519
rect 12094 -2629 12146 -2625
rect 12094 -3401 12103 -2629
rect 12103 -3401 12137 -2629
rect 12137 -3401 12146 -2629
rect 12370 -2519 12379 -1747
rect 12379 -2519 12413 -1747
rect 12413 -2519 12422 -1747
rect 12370 -2523 12422 -2519
rect 12370 -2629 12422 -2625
rect 12370 -3401 12379 -2629
rect 12379 -3401 12413 -2629
rect 12413 -3401 12422 -2629
rect 12646 -2519 12655 -1747
rect 12655 -2519 12689 -1747
rect 12689 -2519 12698 -1747
rect 12646 -2523 12698 -2519
rect 12646 -2629 12698 -2625
rect 12646 -3401 12655 -2629
rect 12655 -3401 12689 -2629
rect 12689 -3401 12698 -2629
rect 12922 -2519 12931 -1747
rect 12931 -2519 12965 -1747
rect 12965 -2519 12974 -1747
rect 12922 -2523 12974 -2519
rect 12922 -2629 12974 -2625
rect 12922 -3401 12931 -2629
rect 12931 -3401 12965 -2629
rect 12965 -3401 12974 -2629
rect 13198 -2519 13207 -1747
rect 13207 -2519 13241 -1747
rect 13241 -2519 13250 -1747
rect 13198 -2523 13250 -2519
rect 13198 -2629 13250 -2625
rect 13198 -3401 13207 -2629
rect 13207 -3401 13241 -2629
rect 13241 -3401 13250 -2629
rect 13474 -2519 13483 -1747
rect 13483 -2519 13517 -1747
rect 13517 -2519 13526 -1747
rect 13474 -2523 13526 -2519
rect 13474 -2629 13526 -2625
rect 13474 -3401 13483 -2629
rect 13483 -3401 13517 -2629
rect 13517 -3401 13526 -2629
rect 13750 -2519 13759 -1747
rect 13759 -2519 13793 -1747
rect 13793 -2519 13802 -1747
rect 13750 -2523 13802 -2519
rect 13750 -2629 13802 -2625
rect 13750 -3401 13759 -2629
rect 13759 -3401 13793 -2629
rect 13793 -3401 13802 -2629
rect 6583 -8030 8032 -7219
<< metal2 >>
rect 6583 5512 8032 5522
rect 6583 4691 8032 4701
rect 2434 3997 12148 4040
rect 2434 3217 6579 3997
rect 8000 3217 12148 3997
rect 2434 3158 12148 3217
rect 2434 2015 3316 3158
rect 6850 2015 7732 3158
rect 11266 2015 12148 3158
rect 1106 1670 13474 2015
rect 1106 1263 1330 1670
rect 2210 1263 2434 1670
rect 3314 1263 3538 1670
rect 4418 1263 4642 1670
rect 5522 1263 5746 1670
rect 6626 1263 6850 1670
rect 7730 1263 7954 1670
rect 8834 1263 9058 1670
rect 9938 1263 10162 1670
rect 11042 1263 11266 1670
rect 12146 1263 12370 1670
rect 13250 1263 13474 1670
rect 226 1115 13804 1263
rect 226 883 278 1115
rect 226 5 278 107
rect 226 -786 278 -771
rect 502 883 554 1115
rect 502 5 554 107
rect 502 -786 554 -771
rect 778 883 830 1115
rect 778 5 830 107
rect 778 -786 830 -771
rect 1054 883 1106 1115
rect 1054 5 1106 107
rect 1054 -786 1106 -771
rect 1330 883 1382 1115
rect 1330 5 1382 107
rect 1330 -786 1382 -771
rect 1606 883 1658 1115
rect 1606 5 1658 107
rect 1606 -786 1658 -771
rect 1882 883 1934 1115
rect 1882 5 1934 107
rect 1882 -786 1934 -771
rect 2158 883 2210 1115
rect 2158 5 2210 107
rect 2158 -786 2210 -771
rect 2434 883 2486 1115
rect 2434 5 2486 107
rect 2434 -786 2486 -771
rect 2710 883 2762 1115
rect 2710 5 2762 107
rect 2710 -786 2762 -771
rect 2986 883 3038 1115
rect 2986 5 3038 107
rect 2986 -786 3038 -771
rect 3262 883 3314 1115
rect 3262 5 3314 107
rect 3262 -786 3314 -771
rect 3538 883 3590 1115
rect 3538 5 3590 107
rect 3538 -786 3590 -771
rect 3814 883 3866 1115
rect 3814 5 3866 107
rect 3814 -786 3866 -771
rect 4090 883 4142 1115
rect 4090 5 4142 107
rect 4090 -786 4142 -771
rect 4366 883 4418 1115
rect 4366 5 4418 107
rect 4366 -786 4418 -771
rect 4642 883 4694 1115
rect 4642 5 4694 107
rect 4642 -786 4694 -771
rect 4918 883 4970 1115
rect 4918 5 4970 107
rect 4918 -786 4970 -771
rect 5194 883 5246 1115
rect 5194 5 5246 107
rect 5194 -786 5246 -771
rect 5470 883 5522 1115
rect 5470 5 5522 107
rect 5470 -786 5522 -771
rect 5746 883 5798 1115
rect 5746 5 5798 107
rect 5746 -786 5798 -771
rect 6022 883 6074 1115
rect 6022 5 6074 107
rect 6022 -786 6074 -771
rect 6298 883 6350 1115
rect 6298 5 6350 107
rect 6298 -786 6350 -771
rect 6574 883 6626 1115
rect 6574 5 6626 107
rect 6574 -786 6626 -771
rect 6850 883 6902 1115
rect 6850 5 6902 107
rect 6850 -786 6902 -771
rect 7126 883 7178 1115
rect 7126 5 7178 107
rect 7126 -786 7178 -771
rect 7402 883 7454 1115
rect 7402 5 7454 107
rect 7402 -786 7454 -771
rect 7678 883 7730 1115
rect 7678 5 7730 107
rect 7678 -786 7730 -771
rect 7954 883 8006 1115
rect 7954 5 8006 107
rect 7954 -786 8006 -771
rect 8230 883 8282 1115
rect 8230 5 8282 107
rect 8230 -786 8282 -771
rect 8506 883 8558 1115
rect 8506 5 8558 107
rect 8506 -786 8558 -771
rect 8782 883 8834 1115
rect 8782 5 8834 107
rect 8782 -786 8834 -771
rect 9058 883 9110 1115
rect 9058 5 9110 107
rect 9058 -786 9110 -771
rect 9334 883 9386 1115
rect 9334 5 9386 107
rect 9334 -786 9386 -771
rect 9610 883 9662 1115
rect 9610 5 9662 107
rect 9610 -786 9662 -771
rect 9886 883 9938 1115
rect 9886 5 9938 107
rect 9886 -786 9938 -771
rect 10162 883 10214 1115
rect 10162 5 10214 107
rect 10162 -786 10214 -771
rect 10438 883 10490 1115
rect 10438 5 10490 107
rect 10438 -786 10490 -771
rect 10714 883 10766 1115
rect 10714 5 10766 107
rect 10714 -786 10766 -771
rect 10990 883 11042 1115
rect 10990 5 11042 107
rect 10990 -786 11042 -771
rect 11266 883 11318 1115
rect 11266 5 11318 107
rect 11266 -786 11318 -771
rect 11542 883 11594 1115
rect 11542 5 11594 107
rect 11542 -786 11594 -771
rect 11818 883 11870 1115
rect 11818 5 11870 107
rect 11818 -786 11870 -771
rect 12094 883 12146 1115
rect 12094 5 12146 107
rect 12094 -786 12146 -771
rect 12370 883 12422 1115
rect 12370 5 12422 107
rect 12370 -786 12422 -771
rect 12646 883 12698 1115
rect 12646 5 12698 107
rect 12646 -786 12698 -771
rect 12922 883 12974 1115
rect 12922 5 12974 107
rect 12922 -786 12974 -771
rect 13198 883 13250 1115
rect 13198 5 13250 107
rect 13198 -786 13250 -771
rect 13474 883 13526 1115
rect 13474 5 13526 107
rect 13474 -786 13526 -771
rect 13750 883 13802 1115
rect 13750 5 13802 107
rect 13750 -786 13802 -771
rect -840 -990 -300 -980
rect -840 -1550 -300 -1540
rect 226 -1747 278 -1732
rect 226 -2625 278 -2523
rect 226 -3633 278 -3401
rect 502 -1747 554 -1732
rect 502 -2625 554 -2523
rect 502 -3633 554 -3401
rect 778 -1747 830 -1732
rect 778 -2625 830 -2523
rect 778 -3633 830 -3401
rect 1054 -1747 1106 -1732
rect 1054 -2625 1106 -2523
rect 1054 -3633 1106 -3401
rect 1330 -1747 1382 -1732
rect 1330 -2625 1382 -2523
rect 1330 -3633 1382 -3401
rect 1606 -1747 1658 -1732
rect 1606 -2625 1658 -2523
rect 1606 -3633 1658 -3401
rect 1882 -1747 1934 -1732
rect 1882 -2625 1934 -2523
rect 1882 -3633 1934 -3401
rect 2158 -1747 2210 -1732
rect 2158 -2625 2210 -2523
rect 2158 -3633 2210 -3401
rect 2434 -1747 2486 -1732
rect 2434 -2625 2486 -2523
rect 2434 -3633 2486 -3401
rect 2710 -1747 2762 -1732
rect 2710 -2625 2762 -2523
rect 2710 -3633 2762 -3401
rect 2986 -1747 3038 -1732
rect 2986 -2625 3038 -2523
rect 2986 -3633 3038 -3401
rect 3262 -1747 3314 -1732
rect 3262 -2625 3314 -2523
rect 3262 -3633 3314 -3401
rect 3538 -1747 3590 -1732
rect 3538 -2625 3590 -2523
rect 3538 -3633 3590 -3401
rect 3814 -1747 3866 -1732
rect 3814 -2625 3866 -2523
rect 3814 -3633 3866 -3401
rect 4090 -1747 4142 -1732
rect 4090 -2625 4142 -2523
rect 4090 -3633 4142 -3401
rect 4366 -1747 4418 -1732
rect 4366 -2625 4418 -2523
rect 4366 -3633 4418 -3401
rect 4642 -1747 4694 -1732
rect 4642 -2625 4694 -2523
rect 4642 -3633 4694 -3401
rect 4918 -1747 4970 -1732
rect 4918 -2625 4970 -2523
rect 4918 -3633 4970 -3401
rect 5194 -1747 5246 -1732
rect 5194 -2625 5246 -2523
rect 5194 -3633 5246 -3401
rect 5470 -1747 5522 -1732
rect 5470 -2625 5522 -2523
rect 5470 -3633 5522 -3401
rect 5746 -1747 5798 -1732
rect 5746 -2625 5798 -2523
rect 5746 -3633 5798 -3401
rect 6022 -1747 6074 -1732
rect 6022 -2625 6074 -2523
rect 6022 -3633 6074 -3401
rect 6298 -1747 6350 -1732
rect 6298 -2625 6350 -2523
rect 6298 -3633 6350 -3401
rect 6574 -1747 6626 -1732
rect 6574 -2625 6626 -2523
rect 6574 -3633 6626 -3401
rect 6850 -1747 6902 -1732
rect 6850 -2625 6902 -2523
rect 6850 -3633 6902 -3401
rect 7126 -1747 7178 -1732
rect 7126 -2625 7178 -2523
rect 7126 -3633 7178 -3401
rect 7402 -1747 7454 -1732
rect 7402 -2625 7454 -2523
rect 7402 -3633 7454 -3401
rect 7678 -1747 7730 -1732
rect 7678 -2625 7730 -2523
rect 7678 -3633 7730 -3401
rect 7954 -1747 8006 -1732
rect 7954 -2625 8006 -2523
rect 7954 -3633 8006 -3401
rect 8230 -1747 8282 -1732
rect 8230 -2625 8282 -2523
rect 8230 -3633 8282 -3401
rect 8506 -1747 8558 -1732
rect 8506 -2625 8558 -2523
rect 8506 -3633 8558 -3401
rect 8782 -1747 8834 -1732
rect 8782 -2625 8834 -2523
rect 8782 -3633 8834 -3401
rect 9058 -1747 9110 -1732
rect 9058 -2625 9110 -2523
rect 9058 -3633 9110 -3401
rect 9334 -1747 9386 -1732
rect 9334 -2625 9386 -2523
rect 9334 -3633 9386 -3401
rect 9610 -1747 9662 -1732
rect 9610 -2625 9662 -2523
rect 9610 -3633 9662 -3401
rect 9886 -1747 9938 -1732
rect 9886 -2625 9938 -2523
rect 9886 -3633 9938 -3401
rect 10162 -1747 10214 -1732
rect 10162 -2625 10214 -2523
rect 10162 -3633 10214 -3401
rect 10438 -1747 10490 -1732
rect 10438 -2625 10490 -2523
rect 10438 -3633 10490 -3401
rect 10714 -1747 10766 -1732
rect 10714 -2625 10766 -2523
rect 10714 -3633 10766 -3401
rect 10990 -1747 11042 -1732
rect 10990 -2625 11042 -2523
rect 10990 -3633 11042 -3401
rect 11266 -1747 11318 -1732
rect 11266 -2625 11318 -2523
rect 11266 -3633 11318 -3401
rect 11542 -1747 11594 -1732
rect 11542 -2625 11594 -2523
rect 11542 -3633 11594 -3401
rect 11818 -1747 11870 -1732
rect 11818 -2625 11870 -2523
rect 11818 -3633 11870 -3401
rect 12094 -1747 12146 -1732
rect 12094 -2625 12146 -2523
rect 12094 -3633 12146 -3401
rect 12370 -1747 12422 -1732
rect 12370 -2625 12422 -2523
rect 12370 -3633 12422 -3401
rect 12646 -1747 12698 -1732
rect 12646 -2625 12698 -2523
rect 12646 -3633 12698 -3401
rect 12922 -1747 12974 -1732
rect 12922 -2625 12974 -2523
rect 12922 -3633 12974 -3401
rect 13198 -1747 13250 -1732
rect 13198 -2625 13250 -2523
rect 13198 -3633 13250 -3401
rect 13474 -1747 13526 -1732
rect 13474 -2625 13526 -2523
rect 13474 -3633 13526 -3401
rect 13750 -1747 13802 -1732
rect 13750 -2625 13802 -2523
rect 13750 -3633 13802 -3401
rect 226 -3781 13804 -3633
rect 1106 -4188 1330 -3781
rect 2210 -4188 2434 -3781
rect 3314 -4188 3538 -3781
rect 4418 -4188 4642 -3781
rect 5522 -4188 5746 -3781
rect 6626 -4188 6850 -3781
rect 7730 -4188 7954 -3781
rect 8834 -4188 9058 -3781
rect 9938 -4188 10162 -3781
rect 11042 -4188 11266 -3781
rect 12146 -4188 12370 -3781
rect 13250 -4188 13474 -3781
rect 1106 -4533 13474 -4188
rect 2434 -5676 3316 -4533
rect 6850 -5676 7732 -4533
rect 11266 -5676 12148 -4533
rect 2434 -5735 12148 -5676
rect 2434 -6515 6579 -5735
rect 8000 -6515 12148 -5735
rect 2434 -6558 12148 -6515
rect 6583 -7219 8032 -7209
rect 6583 -8040 8032 -8030
<< via2 >>
rect 6583 4701 8032 5512
rect 6579 3217 8000 3997
rect 6579 -6515 8000 -5735
rect 6583 -8030 8032 -7219
<< metal3 >>
rect -1795 5512 8054 5551
rect -1795 4701 6583 5512
rect 8032 4701 8054 5512
rect -1795 4673 8054 4701
rect 6566 4672 8052 4673
rect 6566 4670 8032 4672
rect 6524 3997 8067 4045
rect 6524 3217 6579 3997
rect 8000 3217 8067 3997
rect 6524 3157 8067 3217
rect 6524 -5735 8067 -5675
rect 6524 -6515 6579 -5735
rect 8000 -6515 8067 -5735
rect 6524 -6563 8067 -6515
rect 6566 -7190 8032 -7188
rect 6566 -7191 8052 -7190
rect -1795 -7219 8054 -7191
rect -1795 -8030 6583 -7219
rect 8032 -8030 8054 -7219
rect -1795 -8069 8054 -8030
use sky130_fd_pr__pfet_01v8_lvt_SNVJWU  sky130_fd_pr__pfet_01v8_lvt_SNVJWU_0
timestamp 1616092564
transform 1 0 7014 0 -1 535
box -6965 -464 6965 498
use sky130_fd_pr__pfet_01v8_lvt_UNVJW6  sky130_fd_pr__pfet_01v8_lvt_UNVJW6_0
timestamp 1616092564
transform 1 0 7014 0 1 -387
box -6965 -462 6965 462
<< end >>
