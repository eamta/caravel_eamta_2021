magic
tech sky130A
magscale 1 2
timestamp 1615911822
<< nwell >>
rect -6302 -3003 6302 3003
<< pmos >>
rect -6208 1541 -6068 2941
rect -6010 1541 -5870 2941
rect -5812 1541 -5672 2941
rect -5614 1541 -5474 2941
rect -5416 1541 -5276 2941
rect -5218 1541 -5078 2941
rect -5020 1541 -4880 2941
rect -4822 1541 -4682 2941
rect -4624 1541 -4484 2941
rect -4426 1541 -4286 2941
rect -4228 1541 -4088 2941
rect -4030 1541 -3890 2941
rect -3832 1541 -3692 2941
rect -3634 1541 -3494 2941
rect -3436 1541 -3296 2941
rect -3238 1541 -3098 2941
rect -3040 1541 -2900 2941
rect -2842 1541 -2702 2941
rect -2644 1541 -2504 2941
rect -2446 1541 -2306 2941
rect -2248 1541 -2108 2941
rect -2050 1541 -1910 2941
rect -1852 1541 -1712 2941
rect -1654 1541 -1514 2941
rect -1456 1541 -1316 2941
rect -1258 1541 -1118 2941
rect -1060 1541 -920 2941
rect -862 1541 -722 2941
rect -664 1541 -524 2941
rect -466 1541 -326 2941
rect -268 1541 -128 2941
rect -70 1541 70 2941
rect 128 1541 268 2941
rect 326 1541 466 2941
rect 524 1541 664 2941
rect 722 1541 862 2941
rect 920 1541 1060 2941
rect 1118 1541 1258 2941
rect 1316 1541 1456 2941
rect 1514 1541 1654 2941
rect 1712 1541 1852 2941
rect 1910 1541 2050 2941
rect 2108 1541 2248 2941
rect 2306 1541 2446 2941
rect 2504 1541 2644 2941
rect 2702 1541 2842 2941
rect 2900 1541 3040 2941
rect 3098 1541 3238 2941
rect 3296 1541 3436 2941
rect 3494 1541 3634 2941
rect 3692 1541 3832 2941
rect 3890 1541 4030 2941
rect 4088 1541 4228 2941
rect 4286 1541 4426 2941
rect 4484 1541 4624 2941
rect 4682 1541 4822 2941
rect 4880 1541 5020 2941
rect 5078 1541 5218 2941
rect 5276 1541 5416 2941
rect 5474 1541 5614 2941
rect 5672 1541 5812 2941
rect 5870 1541 6010 2941
rect 6068 1541 6208 2941
rect -6208 47 -6068 1447
rect -6010 47 -5870 1447
rect -5812 47 -5672 1447
rect -5614 47 -5474 1447
rect -5416 47 -5276 1447
rect -5218 47 -5078 1447
rect -5020 47 -4880 1447
rect -4822 47 -4682 1447
rect -4624 47 -4484 1447
rect -4426 47 -4286 1447
rect -4228 47 -4088 1447
rect -4030 47 -3890 1447
rect -3832 47 -3692 1447
rect -3634 47 -3494 1447
rect -3436 47 -3296 1447
rect -3238 47 -3098 1447
rect -3040 47 -2900 1447
rect -2842 47 -2702 1447
rect -2644 47 -2504 1447
rect -2446 47 -2306 1447
rect -2248 47 -2108 1447
rect -2050 47 -1910 1447
rect -1852 47 -1712 1447
rect -1654 47 -1514 1447
rect -1456 47 -1316 1447
rect -1258 47 -1118 1447
rect -1060 47 -920 1447
rect -862 47 -722 1447
rect -664 47 -524 1447
rect -466 47 -326 1447
rect -268 47 -128 1447
rect -70 47 70 1447
rect 128 47 268 1447
rect 326 47 466 1447
rect 524 47 664 1447
rect 722 47 862 1447
rect 920 47 1060 1447
rect 1118 47 1258 1447
rect 1316 47 1456 1447
rect 1514 47 1654 1447
rect 1712 47 1852 1447
rect 1910 47 2050 1447
rect 2108 47 2248 1447
rect 2306 47 2446 1447
rect 2504 47 2644 1447
rect 2702 47 2842 1447
rect 2900 47 3040 1447
rect 3098 47 3238 1447
rect 3296 47 3436 1447
rect 3494 47 3634 1447
rect 3692 47 3832 1447
rect 3890 47 4030 1447
rect 4088 47 4228 1447
rect 4286 47 4426 1447
rect 4484 47 4624 1447
rect 4682 47 4822 1447
rect 4880 47 5020 1447
rect 5078 47 5218 1447
rect 5276 47 5416 1447
rect 5474 47 5614 1447
rect 5672 47 5812 1447
rect 5870 47 6010 1447
rect 6068 47 6208 1447
rect -6208 -1447 -6068 -47
rect -6010 -1447 -5870 -47
rect -5812 -1447 -5672 -47
rect -5614 -1447 -5474 -47
rect -5416 -1447 -5276 -47
rect -5218 -1447 -5078 -47
rect -5020 -1447 -4880 -47
rect -4822 -1447 -4682 -47
rect -4624 -1447 -4484 -47
rect -4426 -1447 -4286 -47
rect -4228 -1447 -4088 -47
rect -4030 -1447 -3890 -47
rect -3832 -1447 -3692 -47
rect -3634 -1447 -3494 -47
rect -3436 -1447 -3296 -47
rect -3238 -1447 -3098 -47
rect -3040 -1447 -2900 -47
rect -2842 -1447 -2702 -47
rect -2644 -1447 -2504 -47
rect -2446 -1447 -2306 -47
rect -2248 -1447 -2108 -47
rect -2050 -1447 -1910 -47
rect -1852 -1447 -1712 -47
rect -1654 -1447 -1514 -47
rect -1456 -1447 -1316 -47
rect -1258 -1447 -1118 -47
rect -1060 -1447 -920 -47
rect -862 -1447 -722 -47
rect -664 -1447 -524 -47
rect -466 -1447 -326 -47
rect -268 -1447 -128 -47
rect -70 -1447 70 -47
rect 128 -1447 268 -47
rect 326 -1447 466 -47
rect 524 -1447 664 -47
rect 722 -1447 862 -47
rect 920 -1447 1060 -47
rect 1118 -1447 1258 -47
rect 1316 -1447 1456 -47
rect 1514 -1447 1654 -47
rect 1712 -1447 1852 -47
rect 1910 -1447 2050 -47
rect 2108 -1447 2248 -47
rect 2306 -1447 2446 -47
rect 2504 -1447 2644 -47
rect 2702 -1447 2842 -47
rect 2900 -1447 3040 -47
rect 3098 -1447 3238 -47
rect 3296 -1447 3436 -47
rect 3494 -1447 3634 -47
rect 3692 -1447 3832 -47
rect 3890 -1447 4030 -47
rect 4088 -1447 4228 -47
rect 4286 -1447 4426 -47
rect 4484 -1447 4624 -47
rect 4682 -1447 4822 -47
rect 4880 -1447 5020 -47
rect 5078 -1447 5218 -47
rect 5276 -1447 5416 -47
rect 5474 -1447 5614 -47
rect 5672 -1447 5812 -47
rect 5870 -1447 6010 -47
rect 6068 -1447 6208 -47
rect -6208 -2941 -6068 -1541
rect -6010 -2941 -5870 -1541
rect -5812 -2941 -5672 -1541
rect -5614 -2941 -5474 -1541
rect -5416 -2941 -5276 -1541
rect -5218 -2941 -5078 -1541
rect -5020 -2941 -4880 -1541
rect -4822 -2941 -4682 -1541
rect -4624 -2941 -4484 -1541
rect -4426 -2941 -4286 -1541
rect -4228 -2941 -4088 -1541
rect -4030 -2941 -3890 -1541
rect -3832 -2941 -3692 -1541
rect -3634 -2941 -3494 -1541
rect -3436 -2941 -3296 -1541
rect -3238 -2941 -3098 -1541
rect -3040 -2941 -2900 -1541
rect -2842 -2941 -2702 -1541
rect -2644 -2941 -2504 -1541
rect -2446 -2941 -2306 -1541
rect -2248 -2941 -2108 -1541
rect -2050 -2941 -1910 -1541
rect -1852 -2941 -1712 -1541
rect -1654 -2941 -1514 -1541
rect -1456 -2941 -1316 -1541
rect -1258 -2941 -1118 -1541
rect -1060 -2941 -920 -1541
rect -862 -2941 -722 -1541
rect -664 -2941 -524 -1541
rect -466 -2941 -326 -1541
rect -268 -2941 -128 -1541
rect -70 -2941 70 -1541
rect 128 -2941 268 -1541
rect 326 -2941 466 -1541
rect 524 -2941 664 -1541
rect 722 -2941 862 -1541
rect 920 -2941 1060 -1541
rect 1118 -2941 1258 -1541
rect 1316 -2941 1456 -1541
rect 1514 -2941 1654 -1541
rect 1712 -2941 1852 -1541
rect 1910 -2941 2050 -1541
rect 2108 -2941 2248 -1541
rect 2306 -2941 2446 -1541
rect 2504 -2941 2644 -1541
rect 2702 -2941 2842 -1541
rect 2900 -2941 3040 -1541
rect 3098 -2941 3238 -1541
rect 3296 -2941 3436 -1541
rect 3494 -2941 3634 -1541
rect 3692 -2941 3832 -1541
rect 3890 -2941 4030 -1541
rect 4088 -2941 4228 -1541
rect 4286 -2941 4426 -1541
rect 4484 -2941 4624 -1541
rect 4682 -2941 4822 -1541
rect 4880 -2941 5020 -1541
rect 5078 -2941 5218 -1541
rect 5276 -2941 5416 -1541
rect 5474 -2941 5614 -1541
rect 5672 -2941 5812 -1541
rect 5870 -2941 6010 -1541
rect 6068 -2941 6208 -1541
<< pdiff >>
rect -6266 2929 -6208 2941
rect -6266 1553 -6254 2929
rect -6220 1553 -6208 2929
rect -6266 1541 -6208 1553
rect -6068 2929 -6010 2941
rect -6068 1553 -6056 2929
rect -6022 1553 -6010 2929
rect -6068 1541 -6010 1553
rect -5870 2929 -5812 2941
rect -5870 1553 -5858 2929
rect -5824 1553 -5812 2929
rect -5870 1541 -5812 1553
rect -5672 2929 -5614 2941
rect -5672 1553 -5660 2929
rect -5626 1553 -5614 2929
rect -5672 1541 -5614 1553
rect -5474 2929 -5416 2941
rect -5474 1553 -5462 2929
rect -5428 1553 -5416 2929
rect -5474 1541 -5416 1553
rect -5276 2929 -5218 2941
rect -5276 1553 -5264 2929
rect -5230 1553 -5218 2929
rect -5276 1541 -5218 1553
rect -5078 2929 -5020 2941
rect -5078 1553 -5066 2929
rect -5032 1553 -5020 2929
rect -5078 1541 -5020 1553
rect -4880 2929 -4822 2941
rect -4880 1553 -4868 2929
rect -4834 1553 -4822 2929
rect -4880 1541 -4822 1553
rect -4682 2929 -4624 2941
rect -4682 1553 -4670 2929
rect -4636 1553 -4624 2929
rect -4682 1541 -4624 1553
rect -4484 2929 -4426 2941
rect -4484 1553 -4472 2929
rect -4438 1553 -4426 2929
rect -4484 1541 -4426 1553
rect -4286 2929 -4228 2941
rect -4286 1553 -4274 2929
rect -4240 1553 -4228 2929
rect -4286 1541 -4228 1553
rect -4088 2929 -4030 2941
rect -4088 1553 -4076 2929
rect -4042 1553 -4030 2929
rect -4088 1541 -4030 1553
rect -3890 2929 -3832 2941
rect -3890 1553 -3878 2929
rect -3844 1553 -3832 2929
rect -3890 1541 -3832 1553
rect -3692 2929 -3634 2941
rect -3692 1553 -3680 2929
rect -3646 1553 -3634 2929
rect -3692 1541 -3634 1553
rect -3494 2929 -3436 2941
rect -3494 1553 -3482 2929
rect -3448 1553 -3436 2929
rect -3494 1541 -3436 1553
rect -3296 2929 -3238 2941
rect -3296 1553 -3284 2929
rect -3250 1553 -3238 2929
rect -3296 1541 -3238 1553
rect -3098 2929 -3040 2941
rect -3098 1553 -3086 2929
rect -3052 1553 -3040 2929
rect -3098 1541 -3040 1553
rect -2900 2929 -2842 2941
rect -2900 1553 -2888 2929
rect -2854 1553 -2842 2929
rect -2900 1541 -2842 1553
rect -2702 2929 -2644 2941
rect -2702 1553 -2690 2929
rect -2656 1553 -2644 2929
rect -2702 1541 -2644 1553
rect -2504 2929 -2446 2941
rect -2504 1553 -2492 2929
rect -2458 1553 -2446 2929
rect -2504 1541 -2446 1553
rect -2306 2929 -2248 2941
rect -2306 1553 -2294 2929
rect -2260 1553 -2248 2929
rect -2306 1541 -2248 1553
rect -2108 2929 -2050 2941
rect -2108 1553 -2096 2929
rect -2062 1553 -2050 2929
rect -2108 1541 -2050 1553
rect -1910 2929 -1852 2941
rect -1910 1553 -1898 2929
rect -1864 1553 -1852 2929
rect -1910 1541 -1852 1553
rect -1712 2929 -1654 2941
rect -1712 1553 -1700 2929
rect -1666 1553 -1654 2929
rect -1712 1541 -1654 1553
rect -1514 2929 -1456 2941
rect -1514 1553 -1502 2929
rect -1468 1553 -1456 2929
rect -1514 1541 -1456 1553
rect -1316 2929 -1258 2941
rect -1316 1553 -1304 2929
rect -1270 1553 -1258 2929
rect -1316 1541 -1258 1553
rect -1118 2929 -1060 2941
rect -1118 1553 -1106 2929
rect -1072 1553 -1060 2929
rect -1118 1541 -1060 1553
rect -920 2929 -862 2941
rect -920 1553 -908 2929
rect -874 1553 -862 2929
rect -920 1541 -862 1553
rect -722 2929 -664 2941
rect -722 1553 -710 2929
rect -676 1553 -664 2929
rect -722 1541 -664 1553
rect -524 2929 -466 2941
rect -524 1553 -512 2929
rect -478 1553 -466 2929
rect -524 1541 -466 1553
rect -326 2929 -268 2941
rect -326 1553 -314 2929
rect -280 1553 -268 2929
rect -326 1541 -268 1553
rect -128 2929 -70 2941
rect -128 1553 -116 2929
rect -82 1553 -70 2929
rect -128 1541 -70 1553
rect 70 2929 128 2941
rect 70 1553 82 2929
rect 116 1553 128 2929
rect 70 1541 128 1553
rect 268 2929 326 2941
rect 268 1553 280 2929
rect 314 1553 326 2929
rect 268 1541 326 1553
rect 466 2929 524 2941
rect 466 1553 478 2929
rect 512 1553 524 2929
rect 466 1541 524 1553
rect 664 2929 722 2941
rect 664 1553 676 2929
rect 710 1553 722 2929
rect 664 1541 722 1553
rect 862 2929 920 2941
rect 862 1553 874 2929
rect 908 1553 920 2929
rect 862 1541 920 1553
rect 1060 2929 1118 2941
rect 1060 1553 1072 2929
rect 1106 1553 1118 2929
rect 1060 1541 1118 1553
rect 1258 2929 1316 2941
rect 1258 1553 1270 2929
rect 1304 1553 1316 2929
rect 1258 1541 1316 1553
rect 1456 2929 1514 2941
rect 1456 1553 1468 2929
rect 1502 1553 1514 2929
rect 1456 1541 1514 1553
rect 1654 2929 1712 2941
rect 1654 1553 1666 2929
rect 1700 1553 1712 2929
rect 1654 1541 1712 1553
rect 1852 2929 1910 2941
rect 1852 1553 1864 2929
rect 1898 1553 1910 2929
rect 1852 1541 1910 1553
rect 2050 2929 2108 2941
rect 2050 1553 2062 2929
rect 2096 1553 2108 2929
rect 2050 1541 2108 1553
rect 2248 2929 2306 2941
rect 2248 1553 2260 2929
rect 2294 1553 2306 2929
rect 2248 1541 2306 1553
rect 2446 2929 2504 2941
rect 2446 1553 2458 2929
rect 2492 1553 2504 2929
rect 2446 1541 2504 1553
rect 2644 2929 2702 2941
rect 2644 1553 2656 2929
rect 2690 1553 2702 2929
rect 2644 1541 2702 1553
rect 2842 2929 2900 2941
rect 2842 1553 2854 2929
rect 2888 1553 2900 2929
rect 2842 1541 2900 1553
rect 3040 2929 3098 2941
rect 3040 1553 3052 2929
rect 3086 1553 3098 2929
rect 3040 1541 3098 1553
rect 3238 2929 3296 2941
rect 3238 1553 3250 2929
rect 3284 1553 3296 2929
rect 3238 1541 3296 1553
rect 3436 2929 3494 2941
rect 3436 1553 3448 2929
rect 3482 1553 3494 2929
rect 3436 1541 3494 1553
rect 3634 2929 3692 2941
rect 3634 1553 3646 2929
rect 3680 1553 3692 2929
rect 3634 1541 3692 1553
rect 3832 2929 3890 2941
rect 3832 1553 3844 2929
rect 3878 1553 3890 2929
rect 3832 1541 3890 1553
rect 4030 2929 4088 2941
rect 4030 1553 4042 2929
rect 4076 1553 4088 2929
rect 4030 1541 4088 1553
rect 4228 2929 4286 2941
rect 4228 1553 4240 2929
rect 4274 1553 4286 2929
rect 4228 1541 4286 1553
rect 4426 2929 4484 2941
rect 4426 1553 4438 2929
rect 4472 1553 4484 2929
rect 4426 1541 4484 1553
rect 4624 2929 4682 2941
rect 4624 1553 4636 2929
rect 4670 1553 4682 2929
rect 4624 1541 4682 1553
rect 4822 2929 4880 2941
rect 4822 1553 4834 2929
rect 4868 1553 4880 2929
rect 4822 1541 4880 1553
rect 5020 2929 5078 2941
rect 5020 1553 5032 2929
rect 5066 1553 5078 2929
rect 5020 1541 5078 1553
rect 5218 2929 5276 2941
rect 5218 1553 5230 2929
rect 5264 1553 5276 2929
rect 5218 1541 5276 1553
rect 5416 2929 5474 2941
rect 5416 1553 5428 2929
rect 5462 1553 5474 2929
rect 5416 1541 5474 1553
rect 5614 2929 5672 2941
rect 5614 1553 5626 2929
rect 5660 1553 5672 2929
rect 5614 1541 5672 1553
rect 5812 2929 5870 2941
rect 5812 1553 5824 2929
rect 5858 1553 5870 2929
rect 5812 1541 5870 1553
rect 6010 2929 6068 2941
rect 6010 1553 6022 2929
rect 6056 1553 6068 2929
rect 6010 1541 6068 1553
rect 6208 2929 6266 2941
rect 6208 1553 6220 2929
rect 6254 1553 6266 2929
rect 6208 1541 6266 1553
rect -6266 1435 -6208 1447
rect -6266 59 -6254 1435
rect -6220 59 -6208 1435
rect -6266 47 -6208 59
rect -6068 1435 -6010 1447
rect -6068 59 -6056 1435
rect -6022 59 -6010 1435
rect -6068 47 -6010 59
rect -5870 1435 -5812 1447
rect -5870 59 -5858 1435
rect -5824 59 -5812 1435
rect -5870 47 -5812 59
rect -5672 1435 -5614 1447
rect -5672 59 -5660 1435
rect -5626 59 -5614 1435
rect -5672 47 -5614 59
rect -5474 1435 -5416 1447
rect -5474 59 -5462 1435
rect -5428 59 -5416 1435
rect -5474 47 -5416 59
rect -5276 1435 -5218 1447
rect -5276 59 -5264 1435
rect -5230 59 -5218 1435
rect -5276 47 -5218 59
rect -5078 1435 -5020 1447
rect -5078 59 -5066 1435
rect -5032 59 -5020 1435
rect -5078 47 -5020 59
rect -4880 1435 -4822 1447
rect -4880 59 -4868 1435
rect -4834 59 -4822 1435
rect -4880 47 -4822 59
rect -4682 1435 -4624 1447
rect -4682 59 -4670 1435
rect -4636 59 -4624 1435
rect -4682 47 -4624 59
rect -4484 1435 -4426 1447
rect -4484 59 -4472 1435
rect -4438 59 -4426 1435
rect -4484 47 -4426 59
rect -4286 1435 -4228 1447
rect -4286 59 -4274 1435
rect -4240 59 -4228 1435
rect -4286 47 -4228 59
rect -4088 1435 -4030 1447
rect -4088 59 -4076 1435
rect -4042 59 -4030 1435
rect -4088 47 -4030 59
rect -3890 1435 -3832 1447
rect -3890 59 -3878 1435
rect -3844 59 -3832 1435
rect -3890 47 -3832 59
rect -3692 1435 -3634 1447
rect -3692 59 -3680 1435
rect -3646 59 -3634 1435
rect -3692 47 -3634 59
rect -3494 1435 -3436 1447
rect -3494 59 -3482 1435
rect -3448 59 -3436 1435
rect -3494 47 -3436 59
rect -3296 1435 -3238 1447
rect -3296 59 -3284 1435
rect -3250 59 -3238 1435
rect -3296 47 -3238 59
rect -3098 1435 -3040 1447
rect -3098 59 -3086 1435
rect -3052 59 -3040 1435
rect -3098 47 -3040 59
rect -2900 1435 -2842 1447
rect -2900 59 -2888 1435
rect -2854 59 -2842 1435
rect -2900 47 -2842 59
rect -2702 1435 -2644 1447
rect -2702 59 -2690 1435
rect -2656 59 -2644 1435
rect -2702 47 -2644 59
rect -2504 1435 -2446 1447
rect -2504 59 -2492 1435
rect -2458 59 -2446 1435
rect -2504 47 -2446 59
rect -2306 1435 -2248 1447
rect -2306 59 -2294 1435
rect -2260 59 -2248 1435
rect -2306 47 -2248 59
rect -2108 1435 -2050 1447
rect -2108 59 -2096 1435
rect -2062 59 -2050 1435
rect -2108 47 -2050 59
rect -1910 1435 -1852 1447
rect -1910 59 -1898 1435
rect -1864 59 -1852 1435
rect -1910 47 -1852 59
rect -1712 1435 -1654 1447
rect -1712 59 -1700 1435
rect -1666 59 -1654 1435
rect -1712 47 -1654 59
rect -1514 1435 -1456 1447
rect -1514 59 -1502 1435
rect -1468 59 -1456 1435
rect -1514 47 -1456 59
rect -1316 1435 -1258 1447
rect -1316 59 -1304 1435
rect -1270 59 -1258 1435
rect -1316 47 -1258 59
rect -1118 1435 -1060 1447
rect -1118 59 -1106 1435
rect -1072 59 -1060 1435
rect -1118 47 -1060 59
rect -920 1435 -862 1447
rect -920 59 -908 1435
rect -874 59 -862 1435
rect -920 47 -862 59
rect -722 1435 -664 1447
rect -722 59 -710 1435
rect -676 59 -664 1435
rect -722 47 -664 59
rect -524 1435 -466 1447
rect -524 59 -512 1435
rect -478 59 -466 1435
rect -524 47 -466 59
rect -326 1435 -268 1447
rect -326 59 -314 1435
rect -280 59 -268 1435
rect -326 47 -268 59
rect -128 1435 -70 1447
rect -128 59 -116 1435
rect -82 59 -70 1435
rect -128 47 -70 59
rect 70 1435 128 1447
rect 70 59 82 1435
rect 116 59 128 1435
rect 70 47 128 59
rect 268 1435 326 1447
rect 268 59 280 1435
rect 314 59 326 1435
rect 268 47 326 59
rect 466 1435 524 1447
rect 466 59 478 1435
rect 512 59 524 1435
rect 466 47 524 59
rect 664 1435 722 1447
rect 664 59 676 1435
rect 710 59 722 1435
rect 664 47 722 59
rect 862 1435 920 1447
rect 862 59 874 1435
rect 908 59 920 1435
rect 862 47 920 59
rect 1060 1435 1118 1447
rect 1060 59 1072 1435
rect 1106 59 1118 1435
rect 1060 47 1118 59
rect 1258 1435 1316 1447
rect 1258 59 1270 1435
rect 1304 59 1316 1435
rect 1258 47 1316 59
rect 1456 1435 1514 1447
rect 1456 59 1468 1435
rect 1502 59 1514 1435
rect 1456 47 1514 59
rect 1654 1435 1712 1447
rect 1654 59 1666 1435
rect 1700 59 1712 1435
rect 1654 47 1712 59
rect 1852 1435 1910 1447
rect 1852 59 1864 1435
rect 1898 59 1910 1435
rect 1852 47 1910 59
rect 2050 1435 2108 1447
rect 2050 59 2062 1435
rect 2096 59 2108 1435
rect 2050 47 2108 59
rect 2248 1435 2306 1447
rect 2248 59 2260 1435
rect 2294 59 2306 1435
rect 2248 47 2306 59
rect 2446 1435 2504 1447
rect 2446 59 2458 1435
rect 2492 59 2504 1435
rect 2446 47 2504 59
rect 2644 1435 2702 1447
rect 2644 59 2656 1435
rect 2690 59 2702 1435
rect 2644 47 2702 59
rect 2842 1435 2900 1447
rect 2842 59 2854 1435
rect 2888 59 2900 1435
rect 2842 47 2900 59
rect 3040 1435 3098 1447
rect 3040 59 3052 1435
rect 3086 59 3098 1435
rect 3040 47 3098 59
rect 3238 1435 3296 1447
rect 3238 59 3250 1435
rect 3284 59 3296 1435
rect 3238 47 3296 59
rect 3436 1435 3494 1447
rect 3436 59 3448 1435
rect 3482 59 3494 1435
rect 3436 47 3494 59
rect 3634 1435 3692 1447
rect 3634 59 3646 1435
rect 3680 59 3692 1435
rect 3634 47 3692 59
rect 3832 1435 3890 1447
rect 3832 59 3844 1435
rect 3878 59 3890 1435
rect 3832 47 3890 59
rect 4030 1435 4088 1447
rect 4030 59 4042 1435
rect 4076 59 4088 1435
rect 4030 47 4088 59
rect 4228 1435 4286 1447
rect 4228 59 4240 1435
rect 4274 59 4286 1435
rect 4228 47 4286 59
rect 4426 1435 4484 1447
rect 4426 59 4438 1435
rect 4472 59 4484 1435
rect 4426 47 4484 59
rect 4624 1435 4682 1447
rect 4624 59 4636 1435
rect 4670 59 4682 1435
rect 4624 47 4682 59
rect 4822 1435 4880 1447
rect 4822 59 4834 1435
rect 4868 59 4880 1435
rect 4822 47 4880 59
rect 5020 1435 5078 1447
rect 5020 59 5032 1435
rect 5066 59 5078 1435
rect 5020 47 5078 59
rect 5218 1435 5276 1447
rect 5218 59 5230 1435
rect 5264 59 5276 1435
rect 5218 47 5276 59
rect 5416 1435 5474 1447
rect 5416 59 5428 1435
rect 5462 59 5474 1435
rect 5416 47 5474 59
rect 5614 1435 5672 1447
rect 5614 59 5626 1435
rect 5660 59 5672 1435
rect 5614 47 5672 59
rect 5812 1435 5870 1447
rect 5812 59 5824 1435
rect 5858 59 5870 1435
rect 5812 47 5870 59
rect 6010 1435 6068 1447
rect 6010 59 6022 1435
rect 6056 59 6068 1435
rect 6010 47 6068 59
rect 6208 1435 6266 1447
rect 6208 59 6220 1435
rect 6254 59 6266 1435
rect 6208 47 6266 59
rect -6266 -59 -6208 -47
rect -6266 -1435 -6254 -59
rect -6220 -1435 -6208 -59
rect -6266 -1447 -6208 -1435
rect -6068 -59 -6010 -47
rect -6068 -1435 -6056 -59
rect -6022 -1435 -6010 -59
rect -6068 -1447 -6010 -1435
rect -5870 -59 -5812 -47
rect -5870 -1435 -5858 -59
rect -5824 -1435 -5812 -59
rect -5870 -1447 -5812 -1435
rect -5672 -59 -5614 -47
rect -5672 -1435 -5660 -59
rect -5626 -1435 -5614 -59
rect -5672 -1447 -5614 -1435
rect -5474 -59 -5416 -47
rect -5474 -1435 -5462 -59
rect -5428 -1435 -5416 -59
rect -5474 -1447 -5416 -1435
rect -5276 -59 -5218 -47
rect -5276 -1435 -5264 -59
rect -5230 -1435 -5218 -59
rect -5276 -1447 -5218 -1435
rect -5078 -59 -5020 -47
rect -5078 -1435 -5066 -59
rect -5032 -1435 -5020 -59
rect -5078 -1447 -5020 -1435
rect -4880 -59 -4822 -47
rect -4880 -1435 -4868 -59
rect -4834 -1435 -4822 -59
rect -4880 -1447 -4822 -1435
rect -4682 -59 -4624 -47
rect -4682 -1435 -4670 -59
rect -4636 -1435 -4624 -59
rect -4682 -1447 -4624 -1435
rect -4484 -59 -4426 -47
rect -4484 -1435 -4472 -59
rect -4438 -1435 -4426 -59
rect -4484 -1447 -4426 -1435
rect -4286 -59 -4228 -47
rect -4286 -1435 -4274 -59
rect -4240 -1435 -4228 -59
rect -4286 -1447 -4228 -1435
rect -4088 -59 -4030 -47
rect -4088 -1435 -4076 -59
rect -4042 -1435 -4030 -59
rect -4088 -1447 -4030 -1435
rect -3890 -59 -3832 -47
rect -3890 -1435 -3878 -59
rect -3844 -1435 -3832 -59
rect -3890 -1447 -3832 -1435
rect -3692 -59 -3634 -47
rect -3692 -1435 -3680 -59
rect -3646 -1435 -3634 -59
rect -3692 -1447 -3634 -1435
rect -3494 -59 -3436 -47
rect -3494 -1435 -3482 -59
rect -3448 -1435 -3436 -59
rect -3494 -1447 -3436 -1435
rect -3296 -59 -3238 -47
rect -3296 -1435 -3284 -59
rect -3250 -1435 -3238 -59
rect -3296 -1447 -3238 -1435
rect -3098 -59 -3040 -47
rect -3098 -1435 -3086 -59
rect -3052 -1435 -3040 -59
rect -3098 -1447 -3040 -1435
rect -2900 -59 -2842 -47
rect -2900 -1435 -2888 -59
rect -2854 -1435 -2842 -59
rect -2900 -1447 -2842 -1435
rect -2702 -59 -2644 -47
rect -2702 -1435 -2690 -59
rect -2656 -1435 -2644 -59
rect -2702 -1447 -2644 -1435
rect -2504 -59 -2446 -47
rect -2504 -1435 -2492 -59
rect -2458 -1435 -2446 -59
rect -2504 -1447 -2446 -1435
rect -2306 -59 -2248 -47
rect -2306 -1435 -2294 -59
rect -2260 -1435 -2248 -59
rect -2306 -1447 -2248 -1435
rect -2108 -59 -2050 -47
rect -2108 -1435 -2096 -59
rect -2062 -1435 -2050 -59
rect -2108 -1447 -2050 -1435
rect -1910 -59 -1852 -47
rect -1910 -1435 -1898 -59
rect -1864 -1435 -1852 -59
rect -1910 -1447 -1852 -1435
rect -1712 -59 -1654 -47
rect -1712 -1435 -1700 -59
rect -1666 -1435 -1654 -59
rect -1712 -1447 -1654 -1435
rect -1514 -59 -1456 -47
rect -1514 -1435 -1502 -59
rect -1468 -1435 -1456 -59
rect -1514 -1447 -1456 -1435
rect -1316 -59 -1258 -47
rect -1316 -1435 -1304 -59
rect -1270 -1435 -1258 -59
rect -1316 -1447 -1258 -1435
rect -1118 -59 -1060 -47
rect -1118 -1435 -1106 -59
rect -1072 -1435 -1060 -59
rect -1118 -1447 -1060 -1435
rect -920 -59 -862 -47
rect -920 -1435 -908 -59
rect -874 -1435 -862 -59
rect -920 -1447 -862 -1435
rect -722 -59 -664 -47
rect -722 -1435 -710 -59
rect -676 -1435 -664 -59
rect -722 -1447 -664 -1435
rect -524 -59 -466 -47
rect -524 -1435 -512 -59
rect -478 -1435 -466 -59
rect -524 -1447 -466 -1435
rect -326 -59 -268 -47
rect -326 -1435 -314 -59
rect -280 -1435 -268 -59
rect -326 -1447 -268 -1435
rect -128 -59 -70 -47
rect -128 -1435 -116 -59
rect -82 -1435 -70 -59
rect -128 -1447 -70 -1435
rect 70 -59 128 -47
rect 70 -1435 82 -59
rect 116 -1435 128 -59
rect 70 -1447 128 -1435
rect 268 -59 326 -47
rect 268 -1435 280 -59
rect 314 -1435 326 -59
rect 268 -1447 326 -1435
rect 466 -59 524 -47
rect 466 -1435 478 -59
rect 512 -1435 524 -59
rect 466 -1447 524 -1435
rect 664 -59 722 -47
rect 664 -1435 676 -59
rect 710 -1435 722 -59
rect 664 -1447 722 -1435
rect 862 -59 920 -47
rect 862 -1435 874 -59
rect 908 -1435 920 -59
rect 862 -1447 920 -1435
rect 1060 -59 1118 -47
rect 1060 -1435 1072 -59
rect 1106 -1435 1118 -59
rect 1060 -1447 1118 -1435
rect 1258 -59 1316 -47
rect 1258 -1435 1270 -59
rect 1304 -1435 1316 -59
rect 1258 -1447 1316 -1435
rect 1456 -59 1514 -47
rect 1456 -1435 1468 -59
rect 1502 -1435 1514 -59
rect 1456 -1447 1514 -1435
rect 1654 -59 1712 -47
rect 1654 -1435 1666 -59
rect 1700 -1435 1712 -59
rect 1654 -1447 1712 -1435
rect 1852 -59 1910 -47
rect 1852 -1435 1864 -59
rect 1898 -1435 1910 -59
rect 1852 -1447 1910 -1435
rect 2050 -59 2108 -47
rect 2050 -1435 2062 -59
rect 2096 -1435 2108 -59
rect 2050 -1447 2108 -1435
rect 2248 -59 2306 -47
rect 2248 -1435 2260 -59
rect 2294 -1435 2306 -59
rect 2248 -1447 2306 -1435
rect 2446 -59 2504 -47
rect 2446 -1435 2458 -59
rect 2492 -1435 2504 -59
rect 2446 -1447 2504 -1435
rect 2644 -59 2702 -47
rect 2644 -1435 2656 -59
rect 2690 -1435 2702 -59
rect 2644 -1447 2702 -1435
rect 2842 -59 2900 -47
rect 2842 -1435 2854 -59
rect 2888 -1435 2900 -59
rect 2842 -1447 2900 -1435
rect 3040 -59 3098 -47
rect 3040 -1435 3052 -59
rect 3086 -1435 3098 -59
rect 3040 -1447 3098 -1435
rect 3238 -59 3296 -47
rect 3238 -1435 3250 -59
rect 3284 -1435 3296 -59
rect 3238 -1447 3296 -1435
rect 3436 -59 3494 -47
rect 3436 -1435 3448 -59
rect 3482 -1435 3494 -59
rect 3436 -1447 3494 -1435
rect 3634 -59 3692 -47
rect 3634 -1435 3646 -59
rect 3680 -1435 3692 -59
rect 3634 -1447 3692 -1435
rect 3832 -59 3890 -47
rect 3832 -1435 3844 -59
rect 3878 -1435 3890 -59
rect 3832 -1447 3890 -1435
rect 4030 -59 4088 -47
rect 4030 -1435 4042 -59
rect 4076 -1435 4088 -59
rect 4030 -1447 4088 -1435
rect 4228 -59 4286 -47
rect 4228 -1435 4240 -59
rect 4274 -1435 4286 -59
rect 4228 -1447 4286 -1435
rect 4426 -59 4484 -47
rect 4426 -1435 4438 -59
rect 4472 -1435 4484 -59
rect 4426 -1447 4484 -1435
rect 4624 -59 4682 -47
rect 4624 -1435 4636 -59
rect 4670 -1435 4682 -59
rect 4624 -1447 4682 -1435
rect 4822 -59 4880 -47
rect 4822 -1435 4834 -59
rect 4868 -1435 4880 -59
rect 4822 -1447 4880 -1435
rect 5020 -59 5078 -47
rect 5020 -1435 5032 -59
rect 5066 -1435 5078 -59
rect 5020 -1447 5078 -1435
rect 5218 -59 5276 -47
rect 5218 -1435 5230 -59
rect 5264 -1435 5276 -59
rect 5218 -1447 5276 -1435
rect 5416 -59 5474 -47
rect 5416 -1435 5428 -59
rect 5462 -1435 5474 -59
rect 5416 -1447 5474 -1435
rect 5614 -59 5672 -47
rect 5614 -1435 5626 -59
rect 5660 -1435 5672 -59
rect 5614 -1447 5672 -1435
rect 5812 -59 5870 -47
rect 5812 -1435 5824 -59
rect 5858 -1435 5870 -59
rect 5812 -1447 5870 -1435
rect 6010 -59 6068 -47
rect 6010 -1435 6022 -59
rect 6056 -1435 6068 -59
rect 6010 -1447 6068 -1435
rect 6208 -59 6266 -47
rect 6208 -1435 6220 -59
rect 6254 -1435 6266 -59
rect 6208 -1447 6266 -1435
rect -6266 -1553 -6208 -1541
rect -6266 -2929 -6254 -1553
rect -6220 -2929 -6208 -1553
rect -6266 -2941 -6208 -2929
rect -6068 -1553 -6010 -1541
rect -6068 -2929 -6056 -1553
rect -6022 -2929 -6010 -1553
rect -6068 -2941 -6010 -2929
rect -5870 -1553 -5812 -1541
rect -5870 -2929 -5858 -1553
rect -5824 -2929 -5812 -1553
rect -5870 -2941 -5812 -2929
rect -5672 -1553 -5614 -1541
rect -5672 -2929 -5660 -1553
rect -5626 -2929 -5614 -1553
rect -5672 -2941 -5614 -2929
rect -5474 -1553 -5416 -1541
rect -5474 -2929 -5462 -1553
rect -5428 -2929 -5416 -1553
rect -5474 -2941 -5416 -2929
rect -5276 -1553 -5218 -1541
rect -5276 -2929 -5264 -1553
rect -5230 -2929 -5218 -1553
rect -5276 -2941 -5218 -2929
rect -5078 -1553 -5020 -1541
rect -5078 -2929 -5066 -1553
rect -5032 -2929 -5020 -1553
rect -5078 -2941 -5020 -2929
rect -4880 -1553 -4822 -1541
rect -4880 -2929 -4868 -1553
rect -4834 -2929 -4822 -1553
rect -4880 -2941 -4822 -2929
rect -4682 -1553 -4624 -1541
rect -4682 -2929 -4670 -1553
rect -4636 -2929 -4624 -1553
rect -4682 -2941 -4624 -2929
rect -4484 -1553 -4426 -1541
rect -4484 -2929 -4472 -1553
rect -4438 -2929 -4426 -1553
rect -4484 -2941 -4426 -2929
rect -4286 -1553 -4228 -1541
rect -4286 -2929 -4274 -1553
rect -4240 -2929 -4228 -1553
rect -4286 -2941 -4228 -2929
rect -4088 -1553 -4030 -1541
rect -4088 -2929 -4076 -1553
rect -4042 -2929 -4030 -1553
rect -4088 -2941 -4030 -2929
rect -3890 -1553 -3832 -1541
rect -3890 -2929 -3878 -1553
rect -3844 -2929 -3832 -1553
rect -3890 -2941 -3832 -2929
rect -3692 -1553 -3634 -1541
rect -3692 -2929 -3680 -1553
rect -3646 -2929 -3634 -1553
rect -3692 -2941 -3634 -2929
rect -3494 -1553 -3436 -1541
rect -3494 -2929 -3482 -1553
rect -3448 -2929 -3436 -1553
rect -3494 -2941 -3436 -2929
rect -3296 -1553 -3238 -1541
rect -3296 -2929 -3284 -1553
rect -3250 -2929 -3238 -1553
rect -3296 -2941 -3238 -2929
rect -3098 -1553 -3040 -1541
rect -3098 -2929 -3086 -1553
rect -3052 -2929 -3040 -1553
rect -3098 -2941 -3040 -2929
rect -2900 -1553 -2842 -1541
rect -2900 -2929 -2888 -1553
rect -2854 -2929 -2842 -1553
rect -2900 -2941 -2842 -2929
rect -2702 -1553 -2644 -1541
rect -2702 -2929 -2690 -1553
rect -2656 -2929 -2644 -1553
rect -2702 -2941 -2644 -2929
rect -2504 -1553 -2446 -1541
rect -2504 -2929 -2492 -1553
rect -2458 -2929 -2446 -1553
rect -2504 -2941 -2446 -2929
rect -2306 -1553 -2248 -1541
rect -2306 -2929 -2294 -1553
rect -2260 -2929 -2248 -1553
rect -2306 -2941 -2248 -2929
rect -2108 -1553 -2050 -1541
rect -2108 -2929 -2096 -1553
rect -2062 -2929 -2050 -1553
rect -2108 -2941 -2050 -2929
rect -1910 -1553 -1852 -1541
rect -1910 -2929 -1898 -1553
rect -1864 -2929 -1852 -1553
rect -1910 -2941 -1852 -2929
rect -1712 -1553 -1654 -1541
rect -1712 -2929 -1700 -1553
rect -1666 -2929 -1654 -1553
rect -1712 -2941 -1654 -2929
rect -1514 -1553 -1456 -1541
rect -1514 -2929 -1502 -1553
rect -1468 -2929 -1456 -1553
rect -1514 -2941 -1456 -2929
rect -1316 -1553 -1258 -1541
rect -1316 -2929 -1304 -1553
rect -1270 -2929 -1258 -1553
rect -1316 -2941 -1258 -2929
rect -1118 -1553 -1060 -1541
rect -1118 -2929 -1106 -1553
rect -1072 -2929 -1060 -1553
rect -1118 -2941 -1060 -2929
rect -920 -1553 -862 -1541
rect -920 -2929 -908 -1553
rect -874 -2929 -862 -1553
rect -920 -2941 -862 -2929
rect -722 -1553 -664 -1541
rect -722 -2929 -710 -1553
rect -676 -2929 -664 -1553
rect -722 -2941 -664 -2929
rect -524 -1553 -466 -1541
rect -524 -2929 -512 -1553
rect -478 -2929 -466 -1553
rect -524 -2941 -466 -2929
rect -326 -1553 -268 -1541
rect -326 -2929 -314 -1553
rect -280 -2929 -268 -1553
rect -326 -2941 -268 -2929
rect -128 -1553 -70 -1541
rect -128 -2929 -116 -1553
rect -82 -2929 -70 -1553
rect -128 -2941 -70 -2929
rect 70 -1553 128 -1541
rect 70 -2929 82 -1553
rect 116 -2929 128 -1553
rect 70 -2941 128 -2929
rect 268 -1553 326 -1541
rect 268 -2929 280 -1553
rect 314 -2929 326 -1553
rect 268 -2941 326 -2929
rect 466 -1553 524 -1541
rect 466 -2929 478 -1553
rect 512 -2929 524 -1553
rect 466 -2941 524 -2929
rect 664 -1553 722 -1541
rect 664 -2929 676 -1553
rect 710 -2929 722 -1553
rect 664 -2941 722 -2929
rect 862 -1553 920 -1541
rect 862 -2929 874 -1553
rect 908 -2929 920 -1553
rect 862 -2941 920 -2929
rect 1060 -1553 1118 -1541
rect 1060 -2929 1072 -1553
rect 1106 -2929 1118 -1553
rect 1060 -2941 1118 -2929
rect 1258 -1553 1316 -1541
rect 1258 -2929 1270 -1553
rect 1304 -2929 1316 -1553
rect 1258 -2941 1316 -2929
rect 1456 -1553 1514 -1541
rect 1456 -2929 1468 -1553
rect 1502 -2929 1514 -1553
rect 1456 -2941 1514 -2929
rect 1654 -1553 1712 -1541
rect 1654 -2929 1666 -1553
rect 1700 -2929 1712 -1553
rect 1654 -2941 1712 -2929
rect 1852 -1553 1910 -1541
rect 1852 -2929 1864 -1553
rect 1898 -2929 1910 -1553
rect 1852 -2941 1910 -2929
rect 2050 -1553 2108 -1541
rect 2050 -2929 2062 -1553
rect 2096 -2929 2108 -1553
rect 2050 -2941 2108 -2929
rect 2248 -1553 2306 -1541
rect 2248 -2929 2260 -1553
rect 2294 -2929 2306 -1553
rect 2248 -2941 2306 -2929
rect 2446 -1553 2504 -1541
rect 2446 -2929 2458 -1553
rect 2492 -2929 2504 -1553
rect 2446 -2941 2504 -2929
rect 2644 -1553 2702 -1541
rect 2644 -2929 2656 -1553
rect 2690 -2929 2702 -1553
rect 2644 -2941 2702 -2929
rect 2842 -1553 2900 -1541
rect 2842 -2929 2854 -1553
rect 2888 -2929 2900 -1553
rect 2842 -2941 2900 -2929
rect 3040 -1553 3098 -1541
rect 3040 -2929 3052 -1553
rect 3086 -2929 3098 -1553
rect 3040 -2941 3098 -2929
rect 3238 -1553 3296 -1541
rect 3238 -2929 3250 -1553
rect 3284 -2929 3296 -1553
rect 3238 -2941 3296 -2929
rect 3436 -1553 3494 -1541
rect 3436 -2929 3448 -1553
rect 3482 -2929 3494 -1553
rect 3436 -2941 3494 -2929
rect 3634 -1553 3692 -1541
rect 3634 -2929 3646 -1553
rect 3680 -2929 3692 -1553
rect 3634 -2941 3692 -2929
rect 3832 -1553 3890 -1541
rect 3832 -2929 3844 -1553
rect 3878 -2929 3890 -1553
rect 3832 -2941 3890 -2929
rect 4030 -1553 4088 -1541
rect 4030 -2929 4042 -1553
rect 4076 -2929 4088 -1553
rect 4030 -2941 4088 -2929
rect 4228 -1553 4286 -1541
rect 4228 -2929 4240 -1553
rect 4274 -2929 4286 -1553
rect 4228 -2941 4286 -2929
rect 4426 -1553 4484 -1541
rect 4426 -2929 4438 -1553
rect 4472 -2929 4484 -1553
rect 4426 -2941 4484 -2929
rect 4624 -1553 4682 -1541
rect 4624 -2929 4636 -1553
rect 4670 -2929 4682 -1553
rect 4624 -2941 4682 -2929
rect 4822 -1553 4880 -1541
rect 4822 -2929 4834 -1553
rect 4868 -2929 4880 -1553
rect 4822 -2941 4880 -2929
rect 5020 -1553 5078 -1541
rect 5020 -2929 5032 -1553
rect 5066 -2929 5078 -1553
rect 5020 -2941 5078 -2929
rect 5218 -1553 5276 -1541
rect 5218 -2929 5230 -1553
rect 5264 -2929 5276 -1553
rect 5218 -2941 5276 -2929
rect 5416 -1553 5474 -1541
rect 5416 -2929 5428 -1553
rect 5462 -2929 5474 -1553
rect 5416 -2941 5474 -2929
rect 5614 -1553 5672 -1541
rect 5614 -2929 5626 -1553
rect 5660 -2929 5672 -1553
rect 5614 -2941 5672 -2929
rect 5812 -1553 5870 -1541
rect 5812 -2929 5824 -1553
rect 5858 -2929 5870 -1553
rect 5812 -2941 5870 -2929
rect 6010 -1553 6068 -1541
rect 6010 -2929 6022 -1553
rect 6056 -2929 6068 -1553
rect 6010 -2941 6068 -2929
rect 6208 -1553 6266 -1541
rect 6208 -2929 6220 -1553
rect 6254 -2929 6266 -1553
rect 6208 -2941 6266 -2929
<< pdiffc >>
rect -6254 1553 -6220 2929
rect -6056 1553 -6022 2929
rect -5858 1553 -5824 2929
rect -5660 1553 -5626 2929
rect -5462 1553 -5428 2929
rect -5264 1553 -5230 2929
rect -5066 1553 -5032 2929
rect -4868 1553 -4834 2929
rect -4670 1553 -4636 2929
rect -4472 1553 -4438 2929
rect -4274 1553 -4240 2929
rect -4076 1553 -4042 2929
rect -3878 1553 -3844 2929
rect -3680 1553 -3646 2929
rect -3482 1553 -3448 2929
rect -3284 1553 -3250 2929
rect -3086 1553 -3052 2929
rect -2888 1553 -2854 2929
rect -2690 1553 -2656 2929
rect -2492 1553 -2458 2929
rect -2294 1553 -2260 2929
rect -2096 1553 -2062 2929
rect -1898 1553 -1864 2929
rect -1700 1553 -1666 2929
rect -1502 1553 -1468 2929
rect -1304 1553 -1270 2929
rect -1106 1553 -1072 2929
rect -908 1553 -874 2929
rect -710 1553 -676 2929
rect -512 1553 -478 2929
rect -314 1553 -280 2929
rect -116 1553 -82 2929
rect 82 1553 116 2929
rect 280 1553 314 2929
rect 478 1553 512 2929
rect 676 1553 710 2929
rect 874 1553 908 2929
rect 1072 1553 1106 2929
rect 1270 1553 1304 2929
rect 1468 1553 1502 2929
rect 1666 1553 1700 2929
rect 1864 1553 1898 2929
rect 2062 1553 2096 2929
rect 2260 1553 2294 2929
rect 2458 1553 2492 2929
rect 2656 1553 2690 2929
rect 2854 1553 2888 2929
rect 3052 1553 3086 2929
rect 3250 1553 3284 2929
rect 3448 1553 3482 2929
rect 3646 1553 3680 2929
rect 3844 1553 3878 2929
rect 4042 1553 4076 2929
rect 4240 1553 4274 2929
rect 4438 1553 4472 2929
rect 4636 1553 4670 2929
rect 4834 1553 4868 2929
rect 5032 1553 5066 2929
rect 5230 1553 5264 2929
rect 5428 1553 5462 2929
rect 5626 1553 5660 2929
rect 5824 1553 5858 2929
rect 6022 1553 6056 2929
rect 6220 1553 6254 2929
rect -6254 59 -6220 1435
rect -6056 59 -6022 1435
rect -5858 59 -5824 1435
rect -5660 59 -5626 1435
rect -5462 59 -5428 1435
rect -5264 59 -5230 1435
rect -5066 59 -5032 1435
rect -4868 59 -4834 1435
rect -4670 59 -4636 1435
rect -4472 59 -4438 1435
rect -4274 59 -4240 1435
rect -4076 59 -4042 1435
rect -3878 59 -3844 1435
rect -3680 59 -3646 1435
rect -3482 59 -3448 1435
rect -3284 59 -3250 1435
rect -3086 59 -3052 1435
rect -2888 59 -2854 1435
rect -2690 59 -2656 1435
rect -2492 59 -2458 1435
rect -2294 59 -2260 1435
rect -2096 59 -2062 1435
rect -1898 59 -1864 1435
rect -1700 59 -1666 1435
rect -1502 59 -1468 1435
rect -1304 59 -1270 1435
rect -1106 59 -1072 1435
rect -908 59 -874 1435
rect -710 59 -676 1435
rect -512 59 -478 1435
rect -314 59 -280 1435
rect -116 59 -82 1435
rect 82 59 116 1435
rect 280 59 314 1435
rect 478 59 512 1435
rect 676 59 710 1435
rect 874 59 908 1435
rect 1072 59 1106 1435
rect 1270 59 1304 1435
rect 1468 59 1502 1435
rect 1666 59 1700 1435
rect 1864 59 1898 1435
rect 2062 59 2096 1435
rect 2260 59 2294 1435
rect 2458 59 2492 1435
rect 2656 59 2690 1435
rect 2854 59 2888 1435
rect 3052 59 3086 1435
rect 3250 59 3284 1435
rect 3448 59 3482 1435
rect 3646 59 3680 1435
rect 3844 59 3878 1435
rect 4042 59 4076 1435
rect 4240 59 4274 1435
rect 4438 59 4472 1435
rect 4636 59 4670 1435
rect 4834 59 4868 1435
rect 5032 59 5066 1435
rect 5230 59 5264 1435
rect 5428 59 5462 1435
rect 5626 59 5660 1435
rect 5824 59 5858 1435
rect 6022 59 6056 1435
rect 6220 59 6254 1435
rect -6254 -1435 -6220 -59
rect -6056 -1435 -6022 -59
rect -5858 -1435 -5824 -59
rect -5660 -1435 -5626 -59
rect -5462 -1435 -5428 -59
rect -5264 -1435 -5230 -59
rect -5066 -1435 -5032 -59
rect -4868 -1435 -4834 -59
rect -4670 -1435 -4636 -59
rect -4472 -1435 -4438 -59
rect -4274 -1435 -4240 -59
rect -4076 -1435 -4042 -59
rect -3878 -1435 -3844 -59
rect -3680 -1435 -3646 -59
rect -3482 -1435 -3448 -59
rect -3284 -1435 -3250 -59
rect -3086 -1435 -3052 -59
rect -2888 -1435 -2854 -59
rect -2690 -1435 -2656 -59
rect -2492 -1435 -2458 -59
rect -2294 -1435 -2260 -59
rect -2096 -1435 -2062 -59
rect -1898 -1435 -1864 -59
rect -1700 -1435 -1666 -59
rect -1502 -1435 -1468 -59
rect -1304 -1435 -1270 -59
rect -1106 -1435 -1072 -59
rect -908 -1435 -874 -59
rect -710 -1435 -676 -59
rect -512 -1435 -478 -59
rect -314 -1435 -280 -59
rect -116 -1435 -82 -59
rect 82 -1435 116 -59
rect 280 -1435 314 -59
rect 478 -1435 512 -59
rect 676 -1435 710 -59
rect 874 -1435 908 -59
rect 1072 -1435 1106 -59
rect 1270 -1435 1304 -59
rect 1468 -1435 1502 -59
rect 1666 -1435 1700 -59
rect 1864 -1435 1898 -59
rect 2062 -1435 2096 -59
rect 2260 -1435 2294 -59
rect 2458 -1435 2492 -59
rect 2656 -1435 2690 -59
rect 2854 -1435 2888 -59
rect 3052 -1435 3086 -59
rect 3250 -1435 3284 -59
rect 3448 -1435 3482 -59
rect 3646 -1435 3680 -59
rect 3844 -1435 3878 -59
rect 4042 -1435 4076 -59
rect 4240 -1435 4274 -59
rect 4438 -1435 4472 -59
rect 4636 -1435 4670 -59
rect 4834 -1435 4868 -59
rect 5032 -1435 5066 -59
rect 5230 -1435 5264 -59
rect 5428 -1435 5462 -59
rect 5626 -1435 5660 -59
rect 5824 -1435 5858 -59
rect 6022 -1435 6056 -59
rect 6220 -1435 6254 -59
rect -6254 -2929 -6220 -1553
rect -6056 -2929 -6022 -1553
rect -5858 -2929 -5824 -1553
rect -5660 -2929 -5626 -1553
rect -5462 -2929 -5428 -1553
rect -5264 -2929 -5230 -1553
rect -5066 -2929 -5032 -1553
rect -4868 -2929 -4834 -1553
rect -4670 -2929 -4636 -1553
rect -4472 -2929 -4438 -1553
rect -4274 -2929 -4240 -1553
rect -4076 -2929 -4042 -1553
rect -3878 -2929 -3844 -1553
rect -3680 -2929 -3646 -1553
rect -3482 -2929 -3448 -1553
rect -3284 -2929 -3250 -1553
rect -3086 -2929 -3052 -1553
rect -2888 -2929 -2854 -1553
rect -2690 -2929 -2656 -1553
rect -2492 -2929 -2458 -1553
rect -2294 -2929 -2260 -1553
rect -2096 -2929 -2062 -1553
rect -1898 -2929 -1864 -1553
rect -1700 -2929 -1666 -1553
rect -1502 -2929 -1468 -1553
rect -1304 -2929 -1270 -1553
rect -1106 -2929 -1072 -1553
rect -908 -2929 -874 -1553
rect -710 -2929 -676 -1553
rect -512 -2929 -478 -1553
rect -314 -2929 -280 -1553
rect -116 -2929 -82 -1553
rect 82 -2929 116 -1553
rect 280 -2929 314 -1553
rect 478 -2929 512 -1553
rect 676 -2929 710 -1553
rect 874 -2929 908 -1553
rect 1072 -2929 1106 -1553
rect 1270 -2929 1304 -1553
rect 1468 -2929 1502 -1553
rect 1666 -2929 1700 -1553
rect 1864 -2929 1898 -1553
rect 2062 -2929 2096 -1553
rect 2260 -2929 2294 -1553
rect 2458 -2929 2492 -1553
rect 2656 -2929 2690 -1553
rect 2854 -2929 2888 -1553
rect 3052 -2929 3086 -1553
rect 3250 -2929 3284 -1553
rect 3448 -2929 3482 -1553
rect 3646 -2929 3680 -1553
rect 3844 -2929 3878 -1553
rect 4042 -2929 4076 -1553
rect 4240 -2929 4274 -1553
rect 4438 -2929 4472 -1553
rect 4636 -2929 4670 -1553
rect 4834 -2929 4868 -1553
rect 5032 -2929 5066 -1553
rect 5230 -2929 5264 -1553
rect 5428 -2929 5462 -1553
rect 5626 -2929 5660 -1553
rect 5824 -2929 5858 -1553
rect 6022 -2929 6056 -1553
rect 6220 -2929 6254 -1553
<< poly >>
rect -6208 2941 -6068 2967
rect -6010 2941 -5870 2967
rect -5812 2941 -5672 2967
rect -5614 2941 -5474 2967
rect -5416 2941 -5276 2967
rect -5218 2941 -5078 2967
rect -5020 2941 -4880 2967
rect -4822 2941 -4682 2967
rect -4624 2941 -4484 2967
rect -4426 2941 -4286 2967
rect -4228 2941 -4088 2967
rect -4030 2941 -3890 2967
rect -3832 2941 -3692 2967
rect -3634 2941 -3494 2967
rect -3436 2941 -3296 2967
rect -3238 2941 -3098 2967
rect -3040 2941 -2900 2967
rect -2842 2941 -2702 2967
rect -2644 2941 -2504 2967
rect -2446 2941 -2306 2967
rect -2248 2941 -2108 2967
rect -2050 2941 -1910 2967
rect -1852 2941 -1712 2967
rect -1654 2941 -1514 2967
rect -1456 2941 -1316 2967
rect -1258 2941 -1118 2967
rect -1060 2941 -920 2967
rect -862 2941 -722 2967
rect -664 2941 -524 2967
rect -466 2941 -326 2967
rect -268 2941 -128 2967
rect -70 2941 70 2967
rect 128 2941 268 2967
rect 326 2941 466 2967
rect 524 2941 664 2967
rect 722 2941 862 2967
rect 920 2941 1060 2967
rect 1118 2941 1258 2967
rect 1316 2941 1456 2967
rect 1514 2941 1654 2967
rect 1712 2941 1852 2967
rect 1910 2941 2050 2967
rect 2108 2941 2248 2967
rect 2306 2941 2446 2967
rect 2504 2941 2644 2967
rect 2702 2941 2842 2967
rect 2900 2941 3040 2967
rect 3098 2941 3238 2967
rect 3296 2941 3436 2967
rect 3494 2941 3634 2967
rect 3692 2941 3832 2967
rect 3890 2941 4030 2967
rect 4088 2941 4228 2967
rect 4286 2941 4426 2967
rect 4484 2941 4624 2967
rect 4682 2941 4822 2967
rect 4880 2941 5020 2967
rect 5078 2941 5218 2967
rect 5276 2941 5416 2967
rect 5474 2941 5614 2967
rect 5672 2941 5812 2967
rect 5870 2941 6010 2967
rect 6068 2941 6208 2967
rect -6208 1515 -6068 1541
rect -6010 1515 -5870 1541
rect -5812 1515 -5672 1541
rect -5614 1515 -5474 1541
rect -5416 1515 -5276 1541
rect -5218 1515 -5078 1541
rect -5020 1515 -4880 1541
rect -4822 1515 -4682 1541
rect -4624 1515 -4484 1541
rect -4426 1515 -4286 1541
rect -4228 1515 -4088 1541
rect -4030 1515 -3890 1541
rect -3832 1515 -3692 1541
rect -3634 1515 -3494 1541
rect -3436 1515 -3296 1541
rect -3238 1515 -3098 1541
rect -3040 1515 -2900 1541
rect -2842 1515 -2702 1541
rect -2644 1515 -2504 1541
rect -2446 1515 -2306 1541
rect -2248 1515 -2108 1541
rect -2050 1515 -1910 1541
rect -1852 1515 -1712 1541
rect -1654 1515 -1514 1541
rect -1456 1515 -1316 1541
rect -1258 1515 -1118 1541
rect -1060 1515 -920 1541
rect -862 1515 -722 1541
rect -664 1515 -524 1541
rect -466 1515 -326 1541
rect -268 1515 -128 1541
rect -70 1515 70 1541
rect 128 1515 268 1541
rect 326 1515 466 1541
rect 524 1515 664 1541
rect 722 1515 862 1541
rect 920 1515 1060 1541
rect 1118 1515 1258 1541
rect 1316 1515 1456 1541
rect 1514 1515 1654 1541
rect 1712 1515 1852 1541
rect 1910 1515 2050 1541
rect 2108 1515 2248 1541
rect 2306 1515 2446 1541
rect 2504 1515 2644 1541
rect 2702 1515 2842 1541
rect 2900 1515 3040 1541
rect 3098 1515 3238 1541
rect 3296 1515 3436 1541
rect 3494 1515 3634 1541
rect 3692 1515 3832 1541
rect 3890 1515 4030 1541
rect 4088 1515 4228 1541
rect 4286 1515 4426 1541
rect 4484 1515 4624 1541
rect 4682 1515 4822 1541
rect 4880 1515 5020 1541
rect 5078 1515 5218 1541
rect 5276 1515 5416 1541
rect 5474 1515 5614 1541
rect 5672 1515 5812 1541
rect 5870 1515 6010 1541
rect 6068 1515 6208 1541
rect -6208 1447 -6068 1473
rect -6010 1447 -5870 1473
rect -5812 1447 -5672 1473
rect -5614 1447 -5474 1473
rect -5416 1447 -5276 1473
rect -5218 1447 -5078 1473
rect -5020 1447 -4880 1473
rect -4822 1447 -4682 1473
rect -4624 1447 -4484 1473
rect -4426 1447 -4286 1473
rect -4228 1447 -4088 1473
rect -4030 1447 -3890 1473
rect -3832 1447 -3692 1473
rect -3634 1447 -3494 1473
rect -3436 1447 -3296 1473
rect -3238 1447 -3098 1473
rect -3040 1447 -2900 1473
rect -2842 1447 -2702 1473
rect -2644 1447 -2504 1473
rect -2446 1447 -2306 1473
rect -2248 1447 -2108 1473
rect -2050 1447 -1910 1473
rect -1852 1447 -1712 1473
rect -1654 1447 -1514 1473
rect -1456 1447 -1316 1473
rect -1258 1447 -1118 1473
rect -1060 1447 -920 1473
rect -862 1447 -722 1473
rect -664 1447 -524 1473
rect -466 1447 -326 1473
rect -268 1447 -128 1473
rect -70 1447 70 1473
rect 128 1447 268 1473
rect 326 1447 466 1473
rect 524 1447 664 1473
rect 722 1447 862 1473
rect 920 1447 1060 1473
rect 1118 1447 1258 1473
rect 1316 1447 1456 1473
rect 1514 1447 1654 1473
rect 1712 1447 1852 1473
rect 1910 1447 2050 1473
rect 2108 1447 2248 1473
rect 2306 1447 2446 1473
rect 2504 1447 2644 1473
rect 2702 1447 2842 1473
rect 2900 1447 3040 1473
rect 3098 1447 3238 1473
rect 3296 1447 3436 1473
rect 3494 1447 3634 1473
rect 3692 1447 3832 1473
rect 3890 1447 4030 1473
rect 4088 1447 4228 1473
rect 4286 1447 4426 1473
rect 4484 1447 4624 1473
rect 4682 1447 4822 1473
rect 4880 1447 5020 1473
rect 5078 1447 5218 1473
rect 5276 1447 5416 1473
rect 5474 1447 5614 1473
rect 5672 1447 5812 1473
rect 5870 1447 6010 1473
rect 6068 1447 6208 1473
rect -6208 21 -6068 47
rect -6010 21 -5870 47
rect -5812 21 -5672 47
rect -5614 21 -5474 47
rect -5416 21 -5276 47
rect -5218 21 -5078 47
rect -5020 21 -4880 47
rect -4822 21 -4682 47
rect -4624 21 -4484 47
rect -4426 21 -4286 47
rect -4228 21 -4088 47
rect -4030 21 -3890 47
rect -3832 21 -3692 47
rect -3634 21 -3494 47
rect -3436 21 -3296 47
rect -3238 21 -3098 47
rect -3040 21 -2900 47
rect -2842 21 -2702 47
rect -2644 21 -2504 47
rect -2446 21 -2306 47
rect -2248 21 -2108 47
rect -2050 21 -1910 47
rect -1852 21 -1712 47
rect -1654 21 -1514 47
rect -1456 21 -1316 47
rect -1258 21 -1118 47
rect -1060 21 -920 47
rect -862 21 -722 47
rect -664 21 -524 47
rect -466 21 -326 47
rect -268 21 -128 47
rect -70 21 70 47
rect 128 21 268 47
rect 326 21 466 47
rect 524 21 664 47
rect 722 21 862 47
rect 920 21 1060 47
rect 1118 21 1258 47
rect 1316 21 1456 47
rect 1514 21 1654 47
rect 1712 21 1852 47
rect 1910 21 2050 47
rect 2108 21 2248 47
rect 2306 21 2446 47
rect 2504 21 2644 47
rect 2702 21 2842 47
rect 2900 21 3040 47
rect 3098 21 3238 47
rect 3296 21 3436 47
rect 3494 21 3634 47
rect 3692 21 3832 47
rect 3890 21 4030 47
rect 4088 21 4228 47
rect 4286 21 4426 47
rect 4484 21 4624 47
rect 4682 21 4822 47
rect 4880 21 5020 47
rect 5078 21 5218 47
rect 5276 21 5416 47
rect 5474 21 5614 47
rect 5672 21 5812 47
rect 5870 21 6010 47
rect 6068 21 6208 47
rect -6208 -47 -6068 -21
rect -6010 -47 -5870 -21
rect -5812 -47 -5672 -21
rect -5614 -47 -5474 -21
rect -5416 -47 -5276 -21
rect -5218 -47 -5078 -21
rect -5020 -47 -4880 -21
rect -4822 -47 -4682 -21
rect -4624 -47 -4484 -21
rect -4426 -47 -4286 -21
rect -4228 -47 -4088 -21
rect -4030 -47 -3890 -21
rect -3832 -47 -3692 -21
rect -3634 -47 -3494 -21
rect -3436 -47 -3296 -21
rect -3238 -47 -3098 -21
rect -3040 -47 -2900 -21
rect -2842 -47 -2702 -21
rect -2644 -47 -2504 -21
rect -2446 -47 -2306 -21
rect -2248 -47 -2108 -21
rect -2050 -47 -1910 -21
rect -1852 -47 -1712 -21
rect -1654 -47 -1514 -21
rect -1456 -47 -1316 -21
rect -1258 -47 -1118 -21
rect -1060 -47 -920 -21
rect -862 -47 -722 -21
rect -664 -47 -524 -21
rect -466 -47 -326 -21
rect -268 -47 -128 -21
rect -70 -47 70 -21
rect 128 -47 268 -21
rect 326 -47 466 -21
rect 524 -47 664 -21
rect 722 -47 862 -21
rect 920 -47 1060 -21
rect 1118 -47 1258 -21
rect 1316 -47 1456 -21
rect 1514 -47 1654 -21
rect 1712 -47 1852 -21
rect 1910 -47 2050 -21
rect 2108 -47 2248 -21
rect 2306 -47 2446 -21
rect 2504 -47 2644 -21
rect 2702 -47 2842 -21
rect 2900 -47 3040 -21
rect 3098 -47 3238 -21
rect 3296 -47 3436 -21
rect 3494 -47 3634 -21
rect 3692 -47 3832 -21
rect 3890 -47 4030 -21
rect 4088 -47 4228 -21
rect 4286 -47 4426 -21
rect 4484 -47 4624 -21
rect 4682 -47 4822 -21
rect 4880 -47 5020 -21
rect 5078 -47 5218 -21
rect 5276 -47 5416 -21
rect 5474 -47 5614 -21
rect 5672 -47 5812 -21
rect 5870 -47 6010 -21
rect 6068 -47 6208 -21
rect -6208 -1473 -6068 -1447
rect -6010 -1473 -5870 -1447
rect -5812 -1473 -5672 -1447
rect -5614 -1473 -5474 -1447
rect -5416 -1473 -5276 -1447
rect -5218 -1473 -5078 -1447
rect -5020 -1473 -4880 -1447
rect -4822 -1473 -4682 -1447
rect -4624 -1473 -4484 -1447
rect -4426 -1473 -4286 -1447
rect -4228 -1473 -4088 -1447
rect -4030 -1473 -3890 -1447
rect -3832 -1473 -3692 -1447
rect -3634 -1473 -3494 -1447
rect -3436 -1473 -3296 -1447
rect -3238 -1473 -3098 -1447
rect -3040 -1473 -2900 -1447
rect -2842 -1473 -2702 -1447
rect -2644 -1473 -2504 -1447
rect -2446 -1473 -2306 -1447
rect -2248 -1473 -2108 -1447
rect -2050 -1473 -1910 -1447
rect -1852 -1473 -1712 -1447
rect -1654 -1473 -1514 -1447
rect -1456 -1473 -1316 -1447
rect -1258 -1473 -1118 -1447
rect -1060 -1473 -920 -1447
rect -862 -1473 -722 -1447
rect -664 -1473 -524 -1447
rect -466 -1473 -326 -1447
rect -268 -1473 -128 -1447
rect -70 -1473 70 -1447
rect 128 -1473 268 -1447
rect 326 -1473 466 -1447
rect 524 -1473 664 -1447
rect 722 -1473 862 -1447
rect 920 -1473 1060 -1447
rect 1118 -1473 1258 -1447
rect 1316 -1473 1456 -1447
rect 1514 -1473 1654 -1447
rect 1712 -1473 1852 -1447
rect 1910 -1473 2050 -1447
rect 2108 -1473 2248 -1447
rect 2306 -1473 2446 -1447
rect 2504 -1473 2644 -1447
rect 2702 -1473 2842 -1447
rect 2900 -1473 3040 -1447
rect 3098 -1473 3238 -1447
rect 3296 -1473 3436 -1447
rect 3494 -1473 3634 -1447
rect 3692 -1473 3832 -1447
rect 3890 -1473 4030 -1447
rect 4088 -1473 4228 -1447
rect 4286 -1473 4426 -1447
rect 4484 -1473 4624 -1447
rect 4682 -1473 4822 -1447
rect 4880 -1473 5020 -1447
rect 5078 -1473 5218 -1447
rect 5276 -1473 5416 -1447
rect 5474 -1473 5614 -1447
rect 5672 -1473 5812 -1447
rect 5870 -1473 6010 -1447
rect 6068 -1473 6208 -1447
rect -6208 -1541 -6068 -1515
rect -6010 -1541 -5870 -1515
rect -5812 -1541 -5672 -1515
rect -5614 -1541 -5474 -1515
rect -5416 -1541 -5276 -1515
rect -5218 -1541 -5078 -1515
rect -5020 -1541 -4880 -1515
rect -4822 -1541 -4682 -1515
rect -4624 -1541 -4484 -1515
rect -4426 -1541 -4286 -1515
rect -4228 -1541 -4088 -1515
rect -4030 -1541 -3890 -1515
rect -3832 -1541 -3692 -1515
rect -3634 -1541 -3494 -1515
rect -3436 -1541 -3296 -1515
rect -3238 -1541 -3098 -1515
rect -3040 -1541 -2900 -1515
rect -2842 -1541 -2702 -1515
rect -2644 -1541 -2504 -1515
rect -2446 -1541 -2306 -1515
rect -2248 -1541 -2108 -1515
rect -2050 -1541 -1910 -1515
rect -1852 -1541 -1712 -1515
rect -1654 -1541 -1514 -1515
rect -1456 -1541 -1316 -1515
rect -1258 -1541 -1118 -1515
rect -1060 -1541 -920 -1515
rect -862 -1541 -722 -1515
rect -664 -1541 -524 -1515
rect -466 -1541 -326 -1515
rect -268 -1541 -128 -1515
rect -70 -1541 70 -1515
rect 128 -1541 268 -1515
rect 326 -1541 466 -1515
rect 524 -1541 664 -1515
rect 722 -1541 862 -1515
rect 920 -1541 1060 -1515
rect 1118 -1541 1258 -1515
rect 1316 -1541 1456 -1515
rect 1514 -1541 1654 -1515
rect 1712 -1541 1852 -1515
rect 1910 -1541 2050 -1515
rect 2108 -1541 2248 -1515
rect 2306 -1541 2446 -1515
rect 2504 -1541 2644 -1515
rect 2702 -1541 2842 -1515
rect 2900 -1541 3040 -1515
rect 3098 -1541 3238 -1515
rect 3296 -1541 3436 -1515
rect 3494 -1541 3634 -1515
rect 3692 -1541 3832 -1515
rect 3890 -1541 4030 -1515
rect 4088 -1541 4228 -1515
rect 4286 -1541 4426 -1515
rect 4484 -1541 4624 -1515
rect 4682 -1541 4822 -1515
rect 4880 -1541 5020 -1515
rect 5078 -1541 5218 -1515
rect 5276 -1541 5416 -1515
rect 5474 -1541 5614 -1515
rect 5672 -1541 5812 -1515
rect 5870 -1541 6010 -1515
rect 6068 -1541 6208 -1515
rect -6208 -2967 -6068 -2941
rect -6010 -2967 -5870 -2941
rect -5812 -2967 -5672 -2941
rect -5614 -2967 -5474 -2941
rect -5416 -2967 -5276 -2941
rect -5218 -2967 -5078 -2941
rect -5020 -2967 -4880 -2941
rect -4822 -2967 -4682 -2941
rect -4624 -2967 -4484 -2941
rect -4426 -2967 -4286 -2941
rect -4228 -2967 -4088 -2941
rect -4030 -2967 -3890 -2941
rect -3832 -2967 -3692 -2941
rect -3634 -2967 -3494 -2941
rect -3436 -2967 -3296 -2941
rect -3238 -2967 -3098 -2941
rect -3040 -2967 -2900 -2941
rect -2842 -2967 -2702 -2941
rect -2644 -2967 -2504 -2941
rect -2446 -2967 -2306 -2941
rect -2248 -2967 -2108 -2941
rect -2050 -2967 -1910 -2941
rect -1852 -2967 -1712 -2941
rect -1654 -2967 -1514 -2941
rect -1456 -2967 -1316 -2941
rect -1258 -2967 -1118 -2941
rect -1060 -2967 -920 -2941
rect -862 -2967 -722 -2941
rect -664 -2967 -524 -2941
rect -466 -2967 -326 -2941
rect -268 -2967 -128 -2941
rect -70 -2967 70 -2941
rect 128 -2967 268 -2941
rect 326 -2967 466 -2941
rect 524 -2967 664 -2941
rect 722 -2967 862 -2941
rect 920 -2967 1060 -2941
rect 1118 -2967 1258 -2941
rect 1316 -2967 1456 -2941
rect 1514 -2967 1654 -2941
rect 1712 -2967 1852 -2941
rect 1910 -2967 2050 -2941
rect 2108 -2967 2248 -2941
rect 2306 -2967 2446 -2941
rect 2504 -2967 2644 -2941
rect 2702 -2967 2842 -2941
rect 2900 -2967 3040 -2941
rect 3098 -2967 3238 -2941
rect 3296 -2967 3436 -2941
rect 3494 -2967 3634 -2941
rect 3692 -2967 3832 -2941
rect 3890 -2967 4030 -2941
rect 4088 -2967 4228 -2941
rect 4286 -2967 4426 -2941
rect 4484 -2967 4624 -2941
rect 4682 -2967 4822 -2941
rect 4880 -2967 5020 -2941
rect 5078 -2967 5218 -2941
rect 5276 -2967 5416 -2941
rect 5474 -2967 5614 -2941
rect 5672 -2967 5812 -2941
rect 5870 -2967 6010 -2941
rect 6068 -2967 6208 -2941
<< locali >>
rect -6254 2929 -6220 2945
rect -6254 1537 -6220 1553
rect -6056 2929 -6022 2945
rect -6056 1537 -6022 1553
rect -5858 2929 -5824 2945
rect -5858 1537 -5824 1553
rect -5660 2929 -5626 2945
rect -5660 1537 -5626 1553
rect -5462 2929 -5428 2945
rect -5462 1537 -5428 1553
rect -5264 2929 -5230 2945
rect -5264 1537 -5230 1553
rect -5066 2929 -5032 2945
rect -5066 1537 -5032 1553
rect -4868 2929 -4834 2945
rect -4868 1537 -4834 1553
rect -4670 2929 -4636 2945
rect -4670 1537 -4636 1553
rect -4472 2929 -4438 2945
rect -4472 1537 -4438 1553
rect -4274 2929 -4240 2945
rect -4274 1537 -4240 1553
rect -4076 2929 -4042 2945
rect -4076 1537 -4042 1553
rect -3878 2929 -3844 2945
rect -3878 1537 -3844 1553
rect -3680 2929 -3646 2945
rect -3680 1537 -3646 1553
rect -3482 2929 -3448 2945
rect -3482 1537 -3448 1553
rect -3284 2929 -3250 2945
rect -3284 1537 -3250 1553
rect -3086 2929 -3052 2945
rect -3086 1537 -3052 1553
rect -2888 2929 -2854 2945
rect -2888 1537 -2854 1553
rect -2690 2929 -2656 2945
rect -2690 1537 -2656 1553
rect -2492 2929 -2458 2945
rect -2492 1537 -2458 1553
rect -2294 2929 -2260 2945
rect -2294 1537 -2260 1553
rect -2096 2929 -2062 2945
rect -2096 1537 -2062 1553
rect -1898 2929 -1864 2945
rect -1898 1537 -1864 1553
rect -1700 2929 -1666 2945
rect -1700 1537 -1666 1553
rect -1502 2929 -1468 2945
rect -1502 1537 -1468 1553
rect -1304 2929 -1270 2945
rect -1304 1537 -1270 1553
rect -1106 2929 -1072 2945
rect -1106 1537 -1072 1553
rect -908 2929 -874 2945
rect -908 1537 -874 1553
rect -710 2929 -676 2945
rect -710 1537 -676 1553
rect -512 2929 -478 2945
rect -512 1537 -478 1553
rect -314 2929 -280 2945
rect -314 1537 -280 1553
rect -116 2929 -82 2945
rect -116 1537 -82 1553
rect 82 2929 116 2945
rect 82 1537 116 1553
rect 280 2929 314 2945
rect 280 1537 314 1553
rect 478 2929 512 2945
rect 478 1537 512 1553
rect 676 2929 710 2945
rect 676 1537 710 1553
rect 874 2929 908 2945
rect 874 1537 908 1553
rect 1072 2929 1106 2945
rect 1072 1537 1106 1553
rect 1270 2929 1304 2945
rect 1270 1537 1304 1553
rect 1468 2929 1502 2945
rect 1468 1537 1502 1553
rect 1666 2929 1700 2945
rect 1666 1537 1700 1553
rect 1864 2929 1898 2945
rect 1864 1537 1898 1553
rect 2062 2929 2096 2945
rect 2062 1537 2096 1553
rect 2260 2929 2294 2945
rect 2260 1537 2294 1553
rect 2458 2929 2492 2945
rect 2458 1537 2492 1553
rect 2656 2929 2690 2945
rect 2656 1537 2690 1553
rect 2854 2929 2888 2945
rect 2854 1537 2888 1553
rect 3052 2929 3086 2945
rect 3052 1537 3086 1553
rect 3250 2929 3284 2945
rect 3250 1537 3284 1553
rect 3448 2929 3482 2945
rect 3448 1537 3482 1553
rect 3646 2929 3680 2945
rect 3646 1537 3680 1553
rect 3844 2929 3878 2945
rect 3844 1537 3878 1553
rect 4042 2929 4076 2945
rect 4042 1537 4076 1553
rect 4240 2929 4274 2945
rect 4240 1537 4274 1553
rect 4438 2929 4472 2945
rect 4438 1537 4472 1553
rect 4636 2929 4670 2945
rect 4636 1537 4670 1553
rect 4834 2929 4868 2945
rect 4834 1537 4868 1553
rect 5032 2929 5066 2945
rect 5032 1537 5066 1553
rect 5230 2929 5264 2945
rect 5230 1537 5264 1553
rect 5428 2929 5462 2945
rect 5428 1537 5462 1553
rect 5626 2929 5660 2945
rect 5626 1537 5660 1553
rect 5824 2929 5858 2945
rect 5824 1537 5858 1553
rect 6022 2929 6056 2945
rect 6022 1537 6056 1553
rect 6220 2929 6254 2945
rect 6220 1537 6254 1553
rect -6254 1435 -6220 1451
rect -6254 43 -6220 59
rect -6056 1435 -6022 1451
rect -6056 43 -6022 59
rect -5858 1435 -5824 1451
rect -5858 43 -5824 59
rect -5660 1435 -5626 1451
rect -5660 43 -5626 59
rect -5462 1435 -5428 1451
rect -5462 43 -5428 59
rect -5264 1435 -5230 1451
rect -5264 43 -5230 59
rect -5066 1435 -5032 1451
rect -5066 43 -5032 59
rect -4868 1435 -4834 1451
rect -4868 43 -4834 59
rect -4670 1435 -4636 1451
rect -4670 43 -4636 59
rect -4472 1435 -4438 1451
rect -4472 43 -4438 59
rect -4274 1435 -4240 1451
rect -4274 43 -4240 59
rect -4076 1435 -4042 1451
rect -4076 43 -4042 59
rect -3878 1435 -3844 1451
rect -3878 43 -3844 59
rect -3680 1435 -3646 1451
rect -3680 43 -3646 59
rect -3482 1435 -3448 1451
rect -3482 43 -3448 59
rect -3284 1435 -3250 1451
rect -3284 43 -3250 59
rect -3086 1435 -3052 1451
rect -3086 43 -3052 59
rect -2888 1435 -2854 1451
rect -2888 43 -2854 59
rect -2690 1435 -2656 1451
rect -2690 43 -2656 59
rect -2492 1435 -2458 1451
rect -2492 43 -2458 59
rect -2294 1435 -2260 1451
rect -2294 43 -2260 59
rect -2096 1435 -2062 1451
rect -2096 43 -2062 59
rect -1898 1435 -1864 1451
rect -1898 43 -1864 59
rect -1700 1435 -1666 1451
rect -1700 43 -1666 59
rect -1502 1435 -1468 1451
rect -1502 43 -1468 59
rect -1304 1435 -1270 1451
rect -1304 43 -1270 59
rect -1106 1435 -1072 1451
rect -1106 43 -1072 59
rect -908 1435 -874 1451
rect -908 43 -874 59
rect -710 1435 -676 1451
rect -710 43 -676 59
rect -512 1435 -478 1451
rect -512 43 -478 59
rect -314 1435 -280 1451
rect -314 43 -280 59
rect -116 1435 -82 1451
rect -116 43 -82 59
rect 82 1435 116 1451
rect 82 43 116 59
rect 280 1435 314 1451
rect 280 43 314 59
rect 478 1435 512 1451
rect 478 43 512 59
rect 676 1435 710 1451
rect 676 43 710 59
rect 874 1435 908 1451
rect 874 43 908 59
rect 1072 1435 1106 1451
rect 1072 43 1106 59
rect 1270 1435 1304 1451
rect 1270 43 1304 59
rect 1468 1435 1502 1451
rect 1468 43 1502 59
rect 1666 1435 1700 1451
rect 1666 43 1700 59
rect 1864 1435 1898 1451
rect 1864 43 1898 59
rect 2062 1435 2096 1451
rect 2062 43 2096 59
rect 2260 1435 2294 1451
rect 2260 43 2294 59
rect 2458 1435 2492 1451
rect 2458 43 2492 59
rect 2656 1435 2690 1451
rect 2656 43 2690 59
rect 2854 1435 2888 1451
rect 2854 43 2888 59
rect 3052 1435 3086 1451
rect 3052 43 3086 59
rect 3250 1435 3284 1451
rect 3250 43 3284 59
rect 3448 1435 3482 1451
rect 3448 43 3482 59
rect 3646 1435 3680 1451
rect 3646 43 3680 59
rect 3844 1435 3878 1451
rect 3844 43 3878 59
rect 4042 1435 4076 1451
rect 4042 43 4076 59
rect 4240 1435 4274 1451
rect 4240 43 4274 59
rect 4438 1435 4472 1451
rect 4438 43 4472 59
rect 4636 1435 4670 1451
rect 4636 43 4670 59
rect 4834 1435 4868 1451
rect 4834 43 4868 59
rect 5032 1435 5066 1451
rect 5032 43 5066 59
rect 5230 1435 5264 1451
rect 5230 43 5264 59
rect 5428 1435 5462 1451
rect 5428 43 5462 59
rect 5626 1435 5660 1451
rect 5626 43 5660 59
rect 5824 1435 5858 1451
rect 5824 43 5858 59
rect 6022 1435 6056 1451
rect 6022 43 6056 59
rect 6220 1435 6254 1451
rect 6220 43 6254 59
rect -6254 -59 -6220 -43
rect -6254 -1451 -6220 -1435
rect -6056 -59 -6022 -43
rect -6056 -1451 -6022 -1435
rect -5858 -59 -5824 -43
rect -5858 -1451 -5824 -1435
rect -5660 -59 -5626 -43
rect -5660 -1451 -5626 -1435
rect -5462 -59 -5428 -43
rect -5462 -1451 -5428 -1435
rect -5264 -59 -5230 -43
rect -5264 -1451 -5230 -1435
rect -5066 -59 -5032 -43
rect -5066 -1451 -5032 -1435
rect -4868 -59 -4834 -43
rect -4868 -1451 -4834 -1435
rect -4670 -59 -4636 -43
rect -4670 -1451 -4636 -1435
rect -4472 -59 -4438 -43
rect -4472 -1451 -4438 -1435
rect -4274 -59 -4240 -43
rect -4274 -1451 -4240 -1435
rect -4076 -59 -4042 -43
rect -4076 -1451 -4042 -1435
rect -3878 -59 -3844 -43
rect -3878 -1451 -3844 -1435
rect -3680 -59 -3646 -43
rect -3680 -1451 -3646 -1435
rect -3482 -59 -3448 -43
rect -3482 -1451 -3448 -1435
rect -3284 -59 -3250 -43
rect -3284 -1451 -3250 -1435
rect -3086 -59 -3052 -43
rect -3086 -1451 -3052 -1435
rect -2888 -59 -2854 -43
rect -2888 -1451 -2854 -1435
rect -2690 -59 -2656 -43
rect -2690 -1451 -2656 -1435
rect -2492 -59 -2458 -43
rect -2492 -1451 -2458 -1435
rect -2294 -59 -2260 -43
rect -2294 -1451 -2260 -1435
rect -2096 -59 -2062 -43
rect -2096 -1451 -2062 -1435
rect -1898 -59 -1864 -43
rect -1898 -1451 -1864 -1435
rect -1700 -59 -1666 -43
rect -1700 -1451 -1666 -1435
rect -1502 -59 -1468 -43
rect -1502 -1451 -1468 -1435
rect -1304 -59 -1270 -43
rect -1304 -1451 -1270 -1435
rect -1106 -59 -1072 -43
rect -1106 -1451 -1072 -1435
rect -908 -59 -874 -43
rect -908 -1451 -874 -1435
rect -710 -59 -676 -43
rect -710 -1451 -676 -1435
rect -512 -59 -478 -43
rect -512 -1451 -478 -1435
rect -314 -59 -280 -43
rect -314 -1451 -280 -1435
rect -116 -59 -82 -43
rect -116 -1451 -82 -1435
rect 82 -59 116 -43
rect 82 -1451 116 -1435
rect 280 -59 314 -43
rect 280 -1451 314 -1435
rect 478 -59 512 -43
rect 478 -1451 512 -1435
rect 676 -59 710 -43
rect 676 -1451 710 -1435
rect 874 -59 908 -43
rect 874 -1451 908 -1435
rect 1072 -59 1106 -43
rect 1072 -1451 1106 -1435
rect 1270 -59 1304 -43
rect 1270 -1451 1304 -1435
rect 1468 -59 1502 -43
rect 1468 -1451 1502 -1435
rect 1666 -59 1700 -43
rect 1666 -1451 1700 -1435
rect 1864 -59 1898 -43
rect 1864 -1451 1898 -1435
rect 2062 -59 2096 -43
rect 2062 -1451 2096 -1435
rect 2260 -59 2294 -43
rect 2260 -1451 2294 -1435
rect 2458 -59 2492 -43
rect 2458 -1451 2492 -1435
rect 2656 -59 2690 -43
rect 2656 -1451 2690 -1435
rect 2854 -59 2888 -43
rect 2854 -1451 2888 -1435
rect 3052 -59 3086 -43
rect 3052 -1451 3086 -1435
rect 3250 -59 3284 -43
rect 3250 -1451 3284 -1435
rect 3448 -59 3482 -43
rect 3448 -1451 3482 -1435
rect 3646 -59 3680 -43
rect 3646 -1451 3680 -1435
rect 3844 -59 3878 -43
rect 3844 -1451 3878 -1435
rect 4042 -59 4076 -43
rect 4042 -1451 4076 -1435
rect 4240 -59 4274 -43
rect 4240 -1451 4274 -1435
rect 4438 -59 4472 -43
rect 4438 -1451 4472 -1435
rect 4636 -59 4670 -43
rect 4636 -1451 4670 -1435
rect 4834 -59 4868 -43
rect 4834 -1451 4868 -1435
rect 5032 -59 5066 -43
rect 5032 -1451 5066 -1435
rect 5230 -59 5264 -43
rect 5230 -1451 5264 -1435
rect 5428 -59 5462 -43
rect 5428 -1451 5462 -1435
rect 5626 -59 5660 -43
rect 5626 -1451 5660 -1435
rect 5824 -59 5858 -43
rect 5824 -1451 5858 -1435
rect 6022 -59 6056 -43
rect 6022 -1451 6056 -1435
rect 6220 -59 6254 -43
rect 6220 -1451 6254 -1435
rect -6254 -1553 -6220 -1537
rect -6254 -2945 -6220 -2929
rect -6056 -1553 -6022 -1537
rect -6056 -2945 -6022 -2929
rect -5858 -1553 -5824 -1537
rect -5858 -2945 -5824 -2929
rect -5660 -1553 -5626 -1537
rect -5660 -2945 -5626 -2929
rect -5462 -1553 -5428 -1537
rect -5462 -2945 -5428 -2929
rect -5264 -1553 -5230 -1537
rect -5264 -2945 -5230 -2929
rect -5066 -1553 -5032 -1537
rect -5066 -2945 -5032 -2929
rect -4868 -1553 -4834 -1537
rect -4868 -2945 -4834 -2929
rect -4670 -1553 -4636 -1537
rect -4670 -2945 -4636 -2929
rect -4472 -1553 -4438 -1537
rect -4472 -2945 -4438 -2929
rect -4274 -1553 -4240 -1537
rect -4274 -2945 -4240 -2929
rect -4076 -1553 -4042 -1537
rect -4076 -2945 -4042 -2929
rect -3878 -1553 -3844 -1537
rect -3878 -2945 -3844 -2929
rect -3680 -1553 -3646 -1537
rect -3680 -2945 -3646 -2929
rect -3482 -1553 -3448 -1537
rect -3482 -2945 -3448 -2929
rect -3284 -1553 -3250 -1537
rect -3284 -2945 -3250 -2929
rect -3086 -1553 -3052 -1537
rect -3086 -2945 -3052 -2929
rect -2888 -1553 -2854 -1537
rect -2888 -2945 -2854 -2929
rect -2690 -1553 -2656 -1537
rect -2690 -2945 -2656 -2929
rect -2492 -1553 -2458 -1537
rect -2492 -2945 -2458 -2929
rect -2294 -1553 -2260 -1537
rect -2294 -2945 -2260 -2929
rect -2096 -1553 -2062 -1537
rect -2096 -2945 -2062 -2929
rect -1898 -1553 -1864 -1537
rect -1898 -2945 -1864 -2929
rect -1700 -1553 -1666 -1537
rect -1700 -2945 -1666 -2929
rect -1502 -1553 -1468 -1537
rect -1502 -2945 -1468 -2929
rect -1304 -1553 -1270 -1537
rect -1304 -2945 -1270 -2929
rect -1106 -1553 -1072 -1537
rect -1106 -2945 -1072 -2929
rect -908 -1553 -874 -1537
rect -908 -2945 -874 -2929
rect -710 -1553 -676 -1537
rect -710 -2945 -676 -2929
rect -512 -1553 -478 -1537
rect -512 -2945 -478 -2929
rect -314 -1553 -280 -1537
rect -314 -2945 -280 -2929
rect -116 -1553 -82 -1537
rect -116 -2945 -82 -2929
rect 82 -1553 116 -1537
rect 82 -2945 116 -2929
rect 280 -1553 314 -1537
rect 280 -2945 314 -2929
rect 478 -1553 512 -1537
rect 478 -2945 512 -2929
rect 676 -1553 710 -1537
rect 676 -2945 710 -2929
rect 874 -1553 908 -1537
rect 874 -2945 908 -2929
rect 1072 -1553 1106 -1537
rect 1072 -2945 1106 -2929
rect 1270 -1553 1304 -1537
rect 1270 -2945 1304 -2929
rect 1468 -1553 1502 -1537
rect 1468 -2945 1502 -2929
rect 1666 -1553 1700 -1537
rect 1666 -2945 1700 -2929
rect 1864 -1553 1898 -1537
rect 1864 -2945 1898 -2929
rect 2062 -1553 2096 -1537
rect 2062 -2945 2096 -2929
rect 2260 -1553 2294 -1537
rect 2260 -2945 2294 -2929
rect 2458 -1553 2492 -1537
rect 2458 -2945 2492 -2929
rect 2656 -1553 2690 -1537
rect 2656 -2945 2690 -2929
rect 2854 -1553 2888 -1537
rect 2854 -2945 2888 -2929
rect 3052 -1553 3086 -1537
rect 3052 -2945 3086 -2929
rect 3250 -1553 3284 -1537
rect 3250 -2945 3284 -2929
rect 3448 -1553 3482 -1537
rect 3448 -2945 3482 -2929
rect 3646 -1553 3680 -1537
rect 3646 -2945 3680 -2929
rect 3844 -1553 3878 -1537
rect 3844 -2945 3878 -2929
rect 4042 -1553 4076 -1537
rect 4042 -2945 4076 -2929
rect 4240 -1553 4274 -1537
rect 4240 -2945 4274 -2929
rect 4438 -1553 4472 -1537
rect 4438 -2945 4472 -2929
rect 4636 -1553 4670 -1537
rect 4636 -2945 4670 -2929
rect 4834 -1553 4868 -1537
rect 4834 -2945 4868 -2929
rect 5032 -1553 5066 -1537
rect 5032 -2945 5066 -2929
rect 5230 -1553 5264 -1537
rect 5230 -2945 5264 -2929
rect 5428 -1553 5462 -1537
rect 5428 -2945 5462 -2929
rect 5626 -1553 5660 -1537
rect 5626 -2945 5660 -2929
rect 5824 -1553 5858 -1537
rect 5824 -2945 5858 -2929
rect 6022 -1553 6056 -1537
rect 6022 -2945 6056 -2929
rect 6220 -1553 6254 -1537
rect 6220 -2945 6254 -2929
<< viali >>
rect -6254 1553 -6220 2929
rect -6056 1553 -6022 2929
rect -5858 1553 -5824 2929
rect -5660 1553 -5626 2929
rect -5462 1553 -5428 2929
rect -5264 1553 -5230 2929
rect -5066 1553 -5032 2929
rect -4868 1553 -4834 2929
rect -4670 1553 -4636 2929
rect -4472 1553 -4438 2929
rect -4274 1553 -4240 2929
rect -4076 1553 -4042 2929
rect -3878 1553 -3844 2929
rect -3680 1553 -3646 2929
rect -3482 1553 -3448 2929
rect -3284 1553 -3250 2929
rect -3086 1553 -3052 2929
rect -2888 1553 -2854 2929
rect -2690 1553 -2656 2929
rect -2492 1553 -2458 2929
rect -2294 1553 -2260 2929
rect -2096 1553 -2062 2929
rect -1898 1553 -1864 2929
rect -1700 1553 -1666 2929
rect -1502 1553 -1468 2929
rect -1304 1553 -1270 2929
rect -1106 1553 -1072 2929
rect -908 1553 -874 2929
rect -710 1553 -676 2929
rect -512 1553 -478 2929
rect -314 1553 -280 2929
rect -116 1553 -82 2929
rect 82 1553 116 2929
rect 280 1553 314 2929
rect 478 1553 512 2929
rect 676 1553 710 2929
rect 874 1553 908 2929
rect 1072 1553 1106 2929
rect 1270 1553 1304 2929
rect 1468 1553 1502 2929
rect 1666 1553 1700 2929
rect 1864 1553 1898 2929
rect 2062 1553 2096 2929
rect 2260 1553 2294 2929
rect 2458 1553 2492 2929
rect 2656 1553 2690 2929
rect 2854 1553 2888 2929
rect 3052 1553 3086 2929
rect 3250 1553 3284 2929
rect 3448 1553 3482 2929
rect 3646 1553 3680 2929
rect 3844 1553 3878 2929
rect 4042 1553 4076 2929
rect 4240 1553 4274 2929
rect 4438 1553 4472 2929
rect 4636 1553 4670 2929
rect 4834 1553 4868 2929
rect 5032 1553 5066 2929
rect 5230 1553 5264 2929
rect 5428 1553 5462 2929
rect 5626 1553 5660 2929
rect 5824 1553 5858 2929
rect 6022 1553 6056 2929
rect 6220 1553 6254 2929
rect -6254 59 -6220 1435
rect -6056 59 -6022 1435
rect -5858 59 -5824 1435
rect -5660 59 -5626 1435
rect -5462 59 -5428 1435
rect -5264 59 -5230 1435
rect -5066 59 -5032 1435
rect -4868 59 -4834 1435
rect -4670 59 -4636 1435
rect -4472 59 -4438 1435
rect -4274 59 -4240 1435
rect -4076 59 -4042 1435
rect -3878 59 -3844 1435
rect -3680 59 -3646 1435
rect -3482 59 -3448 1435
rect -3284 59 -3250 1435
rect -3086 59 -3052 1435
rect -2888 59 -2854 1435
rect -2690 59 -2656 1435
rect -2492 59 -2458 1435
rect -2294 59 -2260 1435
rect -2096 59 -2062 1435
rect -1898 59 -1864 1435
rect -1700 59 -1666 1435
rect -1502 59 -1468 1435
rect -1304 59 -1270 1435
rect -1106 59 -1072 1435
rect -908 59 -874 1435
rect -710 59 -676 1435
rect -512 59 -478 1435
rect -314 59 -280 1435
rect -116 59 -82 1435
rect 82 59 116 1435
rect 280 59 314 1435
rect 478 59 512 1435
rect 676 59 710 1435
rect 874 59 908 1435
rect 1072 59 1106 1435
rect 1270 59 1304 1435
rect 1468 59 1502 1435
rect 1666 59 1700 1435
rect 1864 59 1898 1435
rect 2062 59 2096 1435
rect 2260 59 2294 1435
rect 2458 59 2492 1435
rect 2656 59 2690 1435
rect 2854 59 2888 1435
rect 3052 59 3086 1435
rect 3250 59 3284 1435
rect 3448 59 3482 1435
rect 3646 59 3680 1435
rect 3844 59 3878 1435
rect 4042 59 4076 1435
rect 4240 59 4274 1435
rect 4438 59 4472 1435
rect 4636 59 4670 1435
rect 4834 59 4868 1435
rect 5032 59 5066 1435
rect 5230 59 5264 1435
rect 5428 59 5462 1435
rect 5626 59 5660 1435
rect 5824 59 5858 1435
rect 6022 59 6056 1435
rect 6220 59 6254 1435
rect -6254 -1435 -6220 -59
rect -6056 -1435 -6022 -59
rect -5858 -1435 -5824 -59
rect -5660 -1435 -5626 -59
rect -5462 -1435 -5428 -59
rect -5264 -1435 -5230 -59
rect -5066 -1435 -5032 -59
rect -4868 -1435 -4834 -59
rect -4670 -1435 -4636 -59
rect -4472 -1435 -4438 -59
rect -4274 -1435 -4240 -59
rect -4076 -1435 -4042 -59
rect -3878 -1435 -3844 -59
rect -3680 -1435 -3646 -59
rect -3482 -1435 -3448 -59
rect -3284 -1435 -3250 -59
rect -3086 -1435 -3052 -59
rect -2888 -1435 -2854 -59
rect -2690 -1435 -2656 -59
rect -2492 -1435 -2458 -59
rect -2294 -1435 -2260 -59
rect -2096 -1435 -2062 -59
rect -1898 -1435 -1864 -59
rect -1700 -1435 -1666 -59
rect -1502 -1435 -1468 -59
rect -1304 -1435 -1270 -59
rect -1106 -1435 -1072 -59
rect -908 -1435 -874 -59
rect -710 -1435 -676 -59
rect -512 -1435 -478 -59
rect -314 -1435 -280 -59
rect -116 -1435 -82 -59
rect 82 -1435 116 -59
rect 280 -1435 314 -59
rect 478 -1435 512 -59
rect 676 -1435 710 -59
rect 874 -1435 908 -59
rect 1072 -1435 1106 -59
rect 1270 -1435 1304 -59
rect 1468 -1435 1502 -59
rect 1666 -1435 1700 -59
rect 1864 -1435 1898 -59
rect 2062 -1435 2096 -59
rect 2260 -1435 2294 -59
rect 2458 -1435 2492 -59
rect 2656 -1435 2690 -59
rect 2854 -1435 2888 -59
rect 3052 -1435 3086 -59
rect 3250 -1435 3284 -59
rect 3448 -1435 3482 -59
rect 3646 -1435 3680 -59
rect 3844 -1435 3878 -59
rect 4042 -1435 4076 -59
rect 4240 -1435 4274 -59
rect 4438 -1435 4472 -59
rect 4636 -1435 4670 -59
rect 4834 -1435 4868 -59
rect 5032 -1435 5066 -59
rect 5230 -1435 5264 -59
rect 5428 -1435 5462 -59
rect 5626 -1435 5660 -59
rect 5824 -1435 5858 -59
rect 6022 -1435 6056 -59
rect 6220 -1435 6254 -59
rect -6254 -2929 -6220 -1553
rect -6056 -2929 -6022 -1553
rect -5858 -2929 -5824 -1553
rect -5660 -2929 -5626 -1553
rect -5462 -2929 -5428 -1553
rect -5264 -2929 -5230 -1553
rect -5066 -2929 -5032 -1553
rect -4868 -2929 -4834 -1553
rect -4670 -2929 -4636 -1553
rect -4472 -2929 -4438 -1553
rect -4274 -2929 -4240 -1553
rect -4076 -2929 -4042 -1553
rect -3878 -2929 -3844 -1553
rect -3680 -2929 -3646 -1553
rect -3482 -2929 -3448 -1553
rect -3284 -2929 -3250 -1553
rect -3086 -2929 -3052 -1553
rect -2888 -2929 -2854 -1553
rect -2690 -2929 -2656 -1553
rect -2492 -2929 -2458 -1553
rect -2294 -2929 -2260 -1553
rect -2096 -2929 -2062 -1553
rect -1898 -2929 -1864 -1553
rect -1700 -2929 -1666 -1553
rect -1502 -2929 -1468 -1553
rect -1304 -2929 -1270 -1553
rect -1106 -2929 -1072 -1553
rect -908 -2929 -874 -1553
rect -710 -2929 -676 -1553
rect -512 -2929 -478 -1553
rect -314 -2929 -280 -1553
rect -116 -2929 -82 -1553
rect 82 -2929 116 -1553
rect 280 -2929 314 -1553
rect 478 -2929 512 -1553
rect 676 -2929 710 -1553
rect 874 -2929 908 -1553
rect 1072 -2929 1106 -1553
rect 1270 -2929 1304 -1553
rect 1468 -2929 1502 -1553
rect 1666 -2929 1700 -1553
rect 1864 -2929 1898 -1553
rect 2062 -2929 2096 -1553
rect 2260 -2929 2294 -1553
rect 2458 -2929 2492 -1553
rect 2656 -2929 2690 -1553
rect 2854 -2929 2888 -1553
rect 3052 -2929 3086 -1553
rect 3250 -2929 3284 -1553
rect 3448 -2929 3482 -1553
rect 3646 -2929 3680 -1553
rect 3844 -2929 3878 -1553
rect 4042 -2929 4076 -1553
rect 4240 -2929 4274 -1553
rect 4438 -2929 4472 -1553
rect 4636 -2929 4670 -1553
rect 4834 -2929 4868 -1553
rect 5032 -2929 5066 -1553
rect 5230 -2929 5264 -1553
rect 5428 -2929 5462 -1553
rect 5626 -2929 5660 -1553
rect 5824 -2929 5858 -1553
rect 6022 -2929 6056 -1553
rect 6220 -2929 6254 -1553
<< metal1 >>
rect -6260 2929 -6214 2941
rect -6260 1553 -6254 2929
rect -6220 1553 -6214 2929
rect -6260 1541 -6214 1553
rect -6062 2929 -6016 2941
rect -6062 1553 -6056 2929
rect -6022 1553 -6016 2929
rect -6062 1541 -6016 1553
rect -5864 2929 -5818 2941
rect -5864 1553 -5858 2929
rect -5824 1553 -5818 2929
rect -5864 1541 -5818 1553
rect -5666 2929 -5620 2941
rect -5666 1553 -5660 2929
rect -5626 1553 -5620 2929
rect -5666 1541 -5620 1553
rect -5468 2929 -5422 2941
rect -5468 1553 -5462 2929
rect -5428 1553 -5422 2929
rect -5468 1541 -5422 1553
rect -5270 2929 -5224 2941
rect -5270 1553 -5264 2929
rect -5230 1553 -5224 2929
rect -5270 1541 -5224 1553
rect -5072 2929 -5026 2941
rect -5072 1553 -5066 2929
rect -5032 1553 -5026 2929
rect -5072 1541 -5026 1553
rect -4874 2929 -4828 2941
rect -4874 1553 -4868 2929
rect -4834 1553 -4828 2929
rect -4874 1541 -4828 1553
rect -4676 2929 -4630 2941
rect -4676 1553 -4670 2929
rect -4636 1553 -4630 2929
rect -4676 1541 -4630 1553
rect -4478 2929 -4432 2941
rect -4478 1553 -4472 2929
rect -4438 1553 -4432 2929
rect -4478 1541 -4432 1553
rect -4280 2929 -4234 2941
rect -4280 1553 -4274 2929
rect -4240 1553 -4234 2929
rect -4280 1541 -4234 1553
rect -4082 2929 -4036 2941
rect -4082 1553 -4076 2929
rect -4042 1553 -4036 2929
rect -4082 1541 -4036 1553
rect -3884 2929 -3838 2941
rect -3884 1553 -3878 2929
rect -3844 1553 -3838 2929
rect -3884 1541 -3838 1553
rect -3686 2929 -3640 2941
rect -3686 1553 -3680 2929
rect -3646 1553 -3640 2929
rect -3686 1541 -3640 1553
rect -3488 2929 -3442 2941
rect -3488 1553 -3482 2929
rect -3448 1553 -3442 2929
rect -3488 1541 -3442 1553
rect -3290 2929 -3244 2941
rect -3290 1553 -3284 2929
rect -3250 1553 -3244 2929
rect -3290 1541 -3244 1553
rect -3092 2929 -3046 2941
rect -3092 1553 -3086 2929
rect -3052 1553 -3046 2929
rect -3092 1541 -3046 1553
rect -2894 2929 -2848 2941
rect -2894 1553 -2888 2929
rect -2854 1553 -2848 2929
rect -2894 1541 -2848 1553
rect -2696 2929 -2650 2941
rect -2696 1553 -2690 2929
rect -2656 1553 -2650 2929
rect -2696 1541 -2650 1553
rect -2498 2929 -2452 2941
rect -2498 1553 -2492 2929
rect -2458 1553 -2452 2929
rect -2498 1541 -2452 1553
rect -2300 2929 -2254 2941
rect -2300 1553 -2294 2929
rect -2260 1553 -2254 2929
rect -2300 1541 -2254 1553
rect -2102 2929 -2056 2941
rect -2102 1553 -2096 2929
rect -2062 1553 -2056 2929
rect -2102 1541 -2056 1553
rect -1904 2929 -1858 2941
rect -1904 1553 -1898 2929
rect -1864 1553 -1858 2929
rect -1904 1541 -1858 1553
rect -1706 2929 -1660 2941
rect -1706 1553 -1700 2929
rect -1666 1553 -1660 2929
rect -1706 1541 -1660 1553
rect -1508 2929 -1462 2941
rect -1508 1553 -1502 2929
rect -1468 1553 -1462 2929
rect -1508 1541 -1462 1553
rect -1310 2929 -1264 2941
rect -1310 1553 -1304 2929
rect -1270 1553 -1264 2929
rect -1310 1541 -1264 1553
rect -1112 2929 -1066 2941
rect -1112 1553 -1106 2929
rect -1072 1553 -1066 2929
rect -1112 1541 -1066 1553
rect -914 2929 -868 2941
rect -914 1553 -908 2929
rect -874 1553 -868 2929
rect -914 1541 -868 1553
rect -716 2929 -670 2941
rect -716 1553 -710 2929
rect -676 1553 -670 2929
rect -716 1541 -670 1553
rect -518 2929 -472 2941
rect -518 1553 -512 2929
rect -478 1553 -472 2929
rect -518 1541 -472 1553
rect -320 2929 -274 2941
rect -320 1553 -314 2929
rect -280 1553 -274 2929
rect -320 1541 -274 1553
rect -122 2929 -76 2941
rect -122 1553 -116 2929
rect -82 1553 -76 2929
rect -122 1541 -76 1553
rect 76 2929 122 2941
rect 76 1553 82 2929
rect 116 1553 122 2929
rect 76 1541 122 1553
rect 274 2929 320 2941
rect 274 1553 280 2929
rect 314 1553 320 2929
rect 274 1541 320 1553
rect 472 2929 518 2941
rect 472 1553 478 2929
rect 512 1553 518 2929
rect 472 1541 518 1553
rect 670 2929 716 2941
rect 670 1553 676 2929
rect 710 1553 716 2929
rect 670 1541 716 1553
rect 868 2929 914 2941
rect 868 1553 874 2929
rect 908 1553 914 2929
rect 868 1541 914 1553
rect 1066 2929 1112 2941
rect 1066 1553 1072 2929
rect 1106 1553 1112 2929
rect 1066 1541 1112 1553
rect 1264 2929 1310 2941
rect 1264 1553 1270 2929
rect 1304 1553 1310 2929
rect 1264 1541 1310 1553
rect 1462 2929 1508 2941
rect 1462 1553 1468 2929
rect 1502 1553 1508 2929
rect 1462 1541 1508 1553
rect 1660 2929 1706 2941
rect 1660 1553 1666 2929
rect 1700 1553 1706 2929
rect 1660 1541 1706 1553
rect 1858 2929 1904 2941
rect 1858 1553 1864 2929
rect 1898 1553 1904 2929
rect 1858 1541 1904 1553
rect 2056 2929 2102 2941
rect 2056 1553 2062 2929
rect 2096 1553 2102 2929
rect 2056 1541 2102 1553
rect 2254 2929 2300 2941
rect 2254 1553 2260 2929
rect 2294 1553 2300 2929
rect 2254 1541 2300 1553
rect 2452 2929 2498 2941
rect 2452 1553 2458 2929
rect 2492 1553 2498 2929
rect 2452 1541 2498 1553
rect 2650 2929 2696 2941
rect 2650 1553 2656 2929
rect 2690 1553 2696 2929
rect 2650 1541 2696 1553
rect 2848 2929 2894 2941
rect 2848 1553 2854 2929
rect 2888 1553 2894 2929
rect 2848 1541 2894 1553
rect 3046 2929 3092 2941
rect 3046 1553 3052 2929
rect 3086 1553 3092 2929
rect 3046 1541 3092 1553
rect 3244 2929 3290 2941
rect 3244 1553 3250 2929
rect 3284 1553 3290 2929
rect 3244 1541 3290 1553
rect 3442 2929 3488 2941
rect 3442 1553 3448 2929
rect 3482 1553 3488 2929
rect 3442 1541 3488 1553
rect 3640 2929 3686 2941
rect 3640 1553 3646 2929
rect 3680 1553 3686 2929
rect 3640 1541 3686 1553
rect 3838 2929 3884 2941
rect 3838 1553 3844 2929
rect 3878 1553 3884 2929
rect 3838 1541 3884 1553
rect 4036 2929 4082 2941
rect 4036 1553 4042 2929
rect 4076 1553 4082 2929
rect 4036 1541 4082 1553
rect 4234 2929 4280 2941
rect 4234 1553 4240 2929
rect 4274 1553 4280 2929
rect 4234 1541 4280 1553
rect 4432 2929 4478 2941
rect 4432 1553 4438 2929
rect 4472 1553 4478 2929
rect 4432 1541 4478 1553
rect 4630 2929 4676 2941
rect 4630 1553 4636 2929
rect 4670 1553 4676 2929
rect 4630 1541 4676 1553
rect 4828 2929 4874 2941
rect 4828 1553 4834 2929
rect 4868 1553 4874 2929
rect 4828 1541 4874 1553
rect 5026 2929 5072 2941
rect 5026 1553 5032 2929
rect 5066 1553 5072 2929
rect 5026 1541 5072 1553
rect 5224 2929 5270 2941
rect 5224 1553 5230 2929
rect 5264 1553 5270 2929
rect 5224 1541 5270 1553
rect 5422 2929 5468 2941
rect 5422 1553 5428 2929
rect 5462 1553 5468 2929
rect 5422 1541 5468 1553
rect 5620 2929 5666 2941
rect 5620 1553 5626 2929
rect 5660 1553 5666 2929
rect 5620 1541 5666 1553
rect 5818 2929 5864 2941
rect 5818 1553 5824 2929
rect 5858 1553 5864 2929
rect 5818 1541 5864 1553
rect 6016 2929 6062 2941
rect 6016 1553 6022 2929
rect 6056 1553 6062 2929
rect 6016 1541 6062 1553
rect 6214 2929 6260 2941
rect 6214 1553 6220 2929
rect 6254 1553 6260 2929
rect 6214 1541 6260 1553
rect -6260 1435 -6214 1447
rect -6260 59 -6254 1435
rect -6220 59 -6214 1435
rect -6260 47 -6214 59
rect -6062 1435 -6016 1447
rect -6062 59 -6056 1435
rect -6022 59 -6016 1435
rect -6062 47 -6016 59
rect -5864 1435 -5818 1447
rect -5864 59 -5858 1435
rect -5824 59 -5818 1435
rect -5864 47 -5818 59
rect -5666 1435 -5620 1447
rect -5666 59 -5660 1435
rect -5626 59 -5620 1435
rect -5666 47 -5620 59
rect -5468 1435 -5422 1447
rect -5468 59 -5462 1435
rect -5428 59 -5422 1435
rect -5468 47 -5422 59
rect -5270 1435 -5224 1447
rect -5270 59 -5264 1435
rect -5230 59 -5224 1435
rect -5270 47 -5224 59
rect -5072 1435 -5026 1447
rect -5072 59 -5066 1435
rect -5032 59 -5026 1435
rect -5072 47 -5026 59
rect -4874 1435 -4828 1447
rect -4874 59 -4868 1435
rect -4834 59 -4828 1435
rect -4874 47 -4828 59
rect -4676 1435 -4630 1447
rect -4676 59 -4670 1435
rect -4636 59 -4630 1435
rect -4676 47 -4630 59
rect -4478 1435 -4432 1447
rect -4478 59 -4472 1435
rect -4438 59 -4432 1435
rect -4478 47 -4432 59
rect -4280 1435 -4234 1447
rect -4280 59 -4274 1435
rect -4240 59 -4234 1435
rect -4280 47 -4234 59
rect -4082 1435 -4036 1447
rect -4082 59 -4076 1435
rect -4042 59 -4036 1435
rect -4082 47 -4036 59
rect -3884 1435 -3838 1447
rect -3884 59 -3878 1435
rect -3844 59 -3838 1435
rect -3884 47 -3838 59
rect -3686 1435 -3640 1447
rect -3686 59 -3680 1435
rect -3646 59 -3640 1435
rect -3686 47 -3640 59
rect -3488 1435 -3442 1447
rect -3488 59 -3482 1435
rect -3448 59 -3442 1435
rect -3488 47 -3442 59
rect -3290 1435 -3244 1447
rect -3290 59 -3284 1435
rect -3250 59 -3244 1435
rect -3290 47 -3244 59
rect -3092 1435 -3046 1447
rect -3092 59 -3086 1435
rect -3052 59 -3046 1435
rect -3092 47 -3046 59
rect -2894 1435 -2848 1447
rect -2894 59 -2888 1435
rect -2854 59 -2848 1435
rect -2894 47 -2848 59
rect -2696 1435 -2650 1447
rect -2696 59 -2690 1435
rect -2656 59 -2650 1435
rect -2696 47 -2650 59
rect -2498 1435 -2452 1447
rect -2498 59 -2492 1435
rect -2458 59 -2452 1435
rect -2498 47 -2452 59
rect -2300 1435 -2254 1447
rect -2300 59 -2294 1435
rect -2260 59 -2254 1435
rect -2300 47 -2254 59
rect -2102 1435 -2056 1447
rect -2102 59 -2096 1435
rect -2062 59 -2056 1435
rect -2102 47 -2056 59
rect -1904 1435 -1858 1447
rect -1904 59 -1898 1435
rect -1864 59 -1858 1435
rect -1904 47 -1858 59
rect -1706 1435 -1660 1447
rect -1706 59 -1700 1435
rect -1666 59 -1660 1435
rect -1706 47 -1660 59
rect -1508 1435 -1462 1447
rect -1508 59 -1502 1435
rect -1468 59 -1462 1435
rect -1508 47 -1462 59
rect -1310 1435 -1264 1447
rect -1310 59 -1304 1435
rect -1270 59 -1264 1435
rect -1310 47 -1264 59
rect -1112 1435 -1066 1447
rect -1112 59 -1106 1435
rect -1072 59 -1066 1435
rect -1112 47 -1066 59
rect -914 1435 -868 1447
rect -914 59 -908 1435
rect -874 59 -868 1435
rect -914 47 -868 59
rect -716 1435 -670 1447
rect -716 59 -710 1435
rect -676 59 -670 1435
rect -716 47 -670 59
rect -518 1435 -472 1447
rect -518 59 -512 1435
rect -478 59 -472 1435
rect -518 47 -472 59
rect -320 1435 -274 1447
rect -320 59 -314 1435
rect -280 59 -274 1435
rect -320 47 -274 59
rect -122 1435 -76 1447
rect -122 59 -116 1435
rect -82 59 -76 1435
rect -122 47 -76 59
rect 76 1435 122 1447
rect 76 59 82 1435
rect 116 59 122 1435
rect 76 47 122 59
rect 274 1435 320 1447
rect 274 59 280 1435
rect 314 59 320 1435
rect 274 47 320 59
rect 472 1435 518 1447
rect 472 59 478 1435
rect 512 59 518 1435
rect 472 47 518 59
rect 670 1435 716 1447
rect 670 59 676 1435
rect 710 59 716 1435
rect 670 47 716 59
rect 868 1435 914 1447
rect 868 59 874 1435
rect 908 59 914 1435
rect 868 47 914 59
rect 1066 1435 1112 1447
rect 1066 59 1072 1435
rect 1106 59 1112 1435
rect 1066 47 1112 59
rect 1264 1435 1310 1447
rect 1264 59 1270 1435
rect 1304 59 1310 1435
rect 1264 47 1310 59
rect 1462 1435 1508 1447
rect 1462 59 1468 1435
rect 1502 59 1508 1435
rect 1462 47 1508 59
rect 1660 1435 1706 1447
rect 1660 59 1666 1435
rect 1700 59 1706 1435
rect 1660 47 1706 59
rect 1858 1435 1904 1447
rect 1858 59 1864 1435
rect 1898 59 1904 1435
rect 1858 47 1904 59
rect 2056 1435 2102 1447
rect 2056 59 2062 1435
rect 2096 59 2102 1435
rect 2056 47 2102 59
rect 2254 1435 2300 1447
rect 2254 59 2260 1435
rect 2294 59 2300 1435
rect 2254 47 2300 59
rect 2452 1435 2498 1447
rect 2452 59 2458 1435
rect 2492 59 2498 1435
rect 2452 47 2498 59
rect 2650 1435 2696 1447
rect 2650 59 2656 1435
rect 2690 59 2696 1435
rect 2650 47 2696 59
rect 2848 1435 2894 1447
rect 2848 59 2854 1435
rect 2888 59 2894 1435
rect 2848 47 2894 59
rect 3046 1435 3092 1447
rect 3046 59 3052 1435
rect 3086 59 3092 1435
rect 3046 47 3092 59
rect 3244 1435 3290 1447
rect 3244 59 3250 1435
rect 3284 59 3290 1435
rect 3244 47 3290 59
rect 3442 1435 3488 1447
rect 3442 59 3448 1435
rect 3482 59 3488 1435
rect 3442 47 3488 59
rect 3640 1435 3686 1447
rect 3640 59 3646 1435
rect 3680 59 3686 1435
rect 3640 47 3686 59
rect 3838 1435 3884 1447
rect 3838 59 3844 1435
rect 3878 59 3884 1435
rect 3838 47 3884 59
rect 4036 1435 4082 1447
rect 4036 59 4042 1435
rect 4076 59 4082 1435
rect 4036 47 4082 59
rect 4234 1435 4280 1447
rect 4234 59 4240 1435
rect 4274 59 4280 1435
rect 4234 47 4280 59
rect 4432 1435 4478 1447
rect 4432 59 4438 1435
rect 4472 59 4478 1435
rect 4432 47 4478 59
rect 4630 1435 4676 1447
rect 4630 59 4636 1435
rect 4670 59 4676 1435
rect 4630 47 4676 59
rect 4828 1435 4874 1447
rect 4828 59 4834 1435
rect 4868 59 4874 1435
rect 4828 47 4874 59
rect 5026 1435 5072 1447
rect 5026 59 5032 1435
rect 5066 59 5072 1435
rect 5026 47 5072 59
rect 5224 1435 5270 1447
rect 5224 59 5230 1435
rect 5264 59 5270 1435
rect 5224 47 5270 59
rect 5422 1435 5468 1447
rect 5422 59 5428 1435
rect 5462 59 5468 1435
rect 5422 47 5468 59
rect 5620 1435 5666 1447
rect 5620 59 5626 1435
rect 5660 59 5666 1435
rect 5620 47 5666 59
rect 5818 1435 5864 1447
rect 5818 59 5824 1435
rect 5858 59 5864 1435
rect 5818 47 5864 59
rect 6016 1435 6062 1447
rect 6016 59 6022 1435
rect 6056 59 6062 1435
rect 6016 47 6062 59
rect 6214 1435 6260 1447
rect 6214 59 6220 1435
rect 6254 59 6260 1435
rect 6214 47 6260 59
rect -6260 -59 -6214 -47
rect -6260 -1435 -6254 -59
rect -6220 -1435 -6214 -59
rect -6260 -1447 -6214 -1435
rect -6062 -59 -6016 -47
rect -6062 -1435 -6056 -59
rect -6022 -1435 -6016 -59
rect -6062 -1447 -6016 -1435
rect -5864 -59 -5818 -47
rect -5864 -1435 -5858 -59
rect -5824 -1435 -5818 -59
rect -5864 -1447 -5818 -1435
rect -5666 -59 -5620 -47
rect -5666 -1435 -5660 -59
rect -5626 -1435 -5620 -59
rect -5666 -1447 -5620 -1435
rect -5468 -59 -5422 -47
rect -5468 -1435 -5462 -59
rect -5428 -1435 -5422 -59
rect -5468 -1447 -5422 -1435
rect -5270 -59 -5224 -47
rect -5270 -1435 -5264 -59
rect -5230 -1435 -5224 -59
rect -5270 -1447 -5224 -1435
rect -5072 -59 -5026 -47
rect -5072 -1435 -5066 -59
rect -5032 -1435 -5026 -59
rect -5072 -1447 -5026 -1435
rect -4874 -59 -4828 -47
rect -4874 -1435 -4868 -59
rect -4834 -1435 -4828 -59
rect -4874 -1447 -4828 -1435
rect -4676 -59 -4630 -47
rect -4676 -1435 -4670 -59
rect -4636 -1435 -4630 -59
rect -4676 -1447 -4630 -1435
rect -4478 -59 -4432 -47
rect -4478 -1435 -4472 -59
rect -4438 -1435 -4432 -59
rect -4478 -1447 -4432 -1435
rect -4280 -59 -4234 -47
rect -4280 -1435 -4274 -59
rect -4240 -1435 -4234 -59
rect -4280 -1447 -4234 -1435
rect -4082 -59 -4036 -47
rect -4082 -1435 -4076 -59
rect -4042 -1435 -4036 -59
rect -4082 -1447 -4036 -1435
rect -3884 -59 -3838 -47
rect -3884 -1435 -3878 -59
rect -3844 -1435 -3838 -59
rect -3884 -1447 -3838 -1435
rect -3686 -59 -3640 -47
rect -3686 -1435 -3680 -59
rect -3646 -1435 -3640 -59
rect -3686 -1447 -3640 -1435
rect -3488 -59 -3442 -47
rect -3488 -1435 -3482 -59
rect -3448 -1435 -3442 -59
rect -3488 -1447 -3442 -1435
rect -3290 -59 -3244 -47
rect -3290 -1435 -3284 -59
rect -3250 -1435 -3244 -59
rect -3290 -1447 -3244 -1435
rect -3092 -59 -3046 -47
rect -3092 -1435 -3086 -59
rect -3052 -1435 -3046 -59
rect -3092 -1447 -3046 -1435
rect -2894 -59 -2848 -47
rect -2894 -1435 -2888 -59
rect -2854 -1435 -2848 -59
rect -2894 -1447 -2848 -1435
rect -2696 -59 -2650 -47
rect -2696 -1435 -2690 -59
rect -2656 -1435 -2650 -59
rect -2696 -1447 -2650 -1435
rect -2498 -59 -2452 -47
rect -2498 -1435 -2492 -59
rect -2458 -1435 -2452 -59
rect -2498 -1447 -2452 -1435
rect -2300 -59 -2254 -47
rect -2300 -1435 -2294 -59
rect -2260 -1435 -2254 -59
rect -2300 -1447 -2254 -1435
rect -2102 -59 -2056 -47
rect -2102 -1435 -2096 -59
rect -2062 -1435 -2056 -59
rect -2102 -1447 -2056 -1435
rect -1904 -59 -1858 -47
rect -1904 -1435 -1898 -59
rect -1864 -1435 -1858 -59
rect -1904 -1447 -1858 -1435
rect -1706 -59 -1660 -47
rect -1706 -1435 -1700 -59
rect -1666 -1435 -1660 -59
rect -1706 -1447 -1660 -1435
rect -1508 -59 -1462 -47
rect -1508 -1435 -1502 -59
rect -1468 -1435 -1462 -59
rect -1508 -1447 -1462 -1435
rect -1310 -59 -1264 -47
rect -1310 -1435 -1304 -59
rect -1270 -1435 -1264 -59
rect -1310 -1447 -1264 -1435
rect -1112 -59 -1066 -47
rect -1112 -1435 -1106 -59
rect -1072 -1435 -1066 -59
rect -1112 -1447 -1066 -1435
rect -914 -59 -868 -47
rect -914 -1435 -908 -59
rect -874 -1435 -868 -59
rect -914 -1447 -868 -1435
rect -716 -59 -670 -47
rect -716 -1435 -710 -59
rect -676 -1435 -670 -59
rect -716 -1447 -670 -1435
rect -518 -59 -472 -47
rect -518 -1435 -512 -59
rect -478 -1435 -472 -59
rect -518 -1447 -472 -1435
rect -320 -59 -274 -47
rect -320 -1435 -314 -59
rect -280 -1435 -274 -59
rect -320 -1447 -274 -1435
rect -122 -59 -76 -47
rect -122 -1435 -116 -59
rect -82 -1435 -76 -59
rect -122 -1447 -76 -1435
rect 76 -59 122 -47
rect 76 -1435 82 -59
rect 116 -1435 122 -59
rect 76 -1447 122 -1435
rect 274 -59 320 -47
rect 274 -1435 280 -59
rect 314 -1435 320 -59
rect 274 -1447 320 -1435
rect 472 -59 518 -47
rect 472 -1435 478 -59
rect 512 -1435 518 -59
rect 472 -1447 518 -1435
rect 670 -59 716 -47
rect 670 -1435 676 -59
rect 710 -1435 716 -59
rect 670 -1447 716 -1435
rect 868 -59 914 -47
rect 868 -1435 874 -59
rect 908 -1435 914 -59
rect 868 -1447 914 -1435
rect 1066 -59 1112 -47
rect 1066 -1435 1072 -59
rect 1106 -1435 1112 -59
rect 1066 -1447 1112 -1435
rect 1264 -59 1310 -47
rect 1264 -1435 1270 -59
rect 1304 -1435 1310 -59
rect 1264 -1447 1310 -1435
rect 1462 -59 1508 -47
rect 1462 -1435 1468 -59
rect 1502 -1435 1508 -59
rect 1462 -1447 1508 -1435
rect 1660 -59 1706 -47
rect 1660 -1435 1666 -59
rect 1700 -1435 1706 -59
rect 1660 -1447 1706 -1435
rect 1858 -59 1904 -47
rect 1858 -1435 1864 -59
rect 1898 -1435 1904 -59
rect 1858 -1447 1904 -1435
rect 2056 -59 2102 -47
rect 2056 -1435 2062 -59
rect 2096 -1435 2102 -59
rect 2056 -1447 2102 -1435
rect 2254 -59 2300 -47
rect 2254 -1435 2260 -59
rect 2294 -1435 2300 -59
rect 2254 -1447 2300 -1435
rect 2452 -59 2498 -47
rect 2452 -1435 2458 -59
rect 2492 -1435 2498 -59
rect 2452 -1447 2498 -1435
rect 2650 -59 2696 -47
rect 2650 -1435 2656 -59
rect 2690 -1435 2696 -59
rect 2650 -1447 2696 -1435
rect 2848 -59 2894 -47
rect 2848 -1435 2854 -59
rect 2888 -1435 2894 -59
rect 2848 -1447 2894 -1435
rect 3046 -59 3092 -47
rect 3046 -1435 3052 -59
rect 3086 -1435 3092 -59
rect 3046 -1447 3092 -1435
rect 3244 -59 3290 -47
rect 3244 -1435 3250 -59
rect 3284 -1435 3290 -59
rect 3244 -1447 3290 -1435
rect 3442 -59 3488 -47
rect 3442 -1435 3448 -59
rect 3482 -1435 3488 -59
rect 3442 -1447 3488 -1435
rect 3640 -59 3686 -47
rect 3640 -1435 3646 -59
rect 3680 -1435 3686 -59
rect 3640 -1447 3686 -1435
rect 3838 -59 3884 -47
rect 3838 -1435 3844 -59
rect 3878 -1435 3884 -59
rect 3838 -1447 3884 -1435
rect 4036 -59 4082 -47
rect 4036 -1435 4042 -59
rect 4076 -1435 4082 -59
rect 4036 -1447 4082 -1435
rect 4234 -59 4280 -47
rect 4234 -1435 4240 -59
rect 4274 -1435 4280 -59
rect 4234 -1447 4280 -1435
rect 4432 -59 4478 -47
rect 4432 -1435 4438 -59
rect 4472 -1435 4478 -59
rect 4432 -1447 4478 -1435
rect 4630 -59 4676 -47
rect 4630 -1435 4636 -59
rect 4670 -1435 4676 -59
rect 4630 -1447 4676 -1435
rect 4828 -59 4874 -47
rect 4828 -1435 4834 -59
rect 4868 -1435 4874 -59
rect 4828 -1447 4874 -1435
rect 5026 -59 5072 -47
rect 5026 -1435 5032 -59
rect 5066 -1435 5072 -59
rect 5026 -1447 5072 -1435
rect 5224 -59 5270 -47
rect 5224 -1435 5230 -59
rect 5264 -1435 5270 -59
rect 5224 -1447 5270 -1435
rect 5422 -59 5468 -47
rect 5422 -1435 5428 -59
rect 5462 -1435 5468 -59
rect 5422 -1447 5468 -1435
rect 5620 -59 5666 -47
rect 5620 -1435 5626 -59
rect 5660 -1435 5666 -59
rect 5620 -1447 5666 -1435
rect 5818 -59 5864 -47
rect 5818 -1435 5824 -59
rect 5858 -1435 5864 -59
rect 5818 -1447 5864 -1435
rect 6016 -59 6062 -47
rect 6016 -1435 6022 -59
rect 6056 -1435 6062 -59
rect 6016 -1447 6062 -1435
rect 6214 -59 6260 -47
rect 6214 -1435 6220 -59
rect 6254 -1435 6260 -59
rect 6214 -1447 6260 -1435
rect -6260 -1553 -6214 -1541
rect -6260 -2929 -6254 -1553
rect -6220 -2929 -6214 -1553
rect -6260 -2941 -6214 -2929
rect -6062 -1553 -6016 -1541
rect -6062 -2929 -6056 -1553
rect -6022 -2929 -6016 -1553
rect -6062 -2941 -6016 -2929
rect -5864 -1553 -5818 -1541
rect -5864 -2929 -5858 -1553
rect -5824 -2929 -5818 -1553
rect -5864 -2941 -5818 -2929
rect -5666 -1553 -5620 -1541
rect -5666 -2929 -5660 -1553
rect -5626 -2929 -5620 -1553
rect -5666 -2941 -5620 -2929
rect -5468 -1553 -5422 -1541
rect -5468 -2929 -5462 -1553
rect -5428 -2929 -5422 -1553
rect -5468 -2941 -5422 -2929
rect -5270 -1553 -5224 -1541
rect -5270 -2929 -5264 -1553
rect -5230 -2929 -5224 -1553
rect -5270 -2941 -5224 -2929
rect -5072 -1553 -5026 -1541
rect -5072 -2929 -5066 -1553
rect -5032 -2929 -5026 -1553
rect -5072 -2941 -5026 -2929
rect -4874 -1553 -4828 -1541
rect -4874 -2929 -4868 -1553
rect -4834 -2929 -4828 -1553
rect -4874 -2941 -4828 -2929
rect -4676 -1553 -4630 -1541
rect -4676 -2929 -4670 -1553
rect -4636 -2929 -4630 -1553
rect -4676 -2941 -4630 -2929
rect -4478 -1553 -4432 -1541
rect -4478 -2929 -4472 -1553
rect -4438 -2929 -4432 -1553
rect -4478 -2941 -4432 -2929
rect -4280 -1553 -4234 -1541
rect -4280 -2929 -4274 -1553
rect -4240 -2929 -4234 -1553
rect -4280 -2941 -4234 -2929
rect -4082 -1553 -4036 -1541
rect -4082 -2929 -4076 -1553
rect -4042 -2929 -4036 -1553
rect -4082 -2941 -4036 -2929
rect -3884 -1553 -3838 -1541
rect -3884 -2929 -3878 -1553
rect -3844 -2929 -3838 -1553
rect -3884 -2941 -3838 -2929
rect -3686 -1553 -3640 -1541
rect -3686 -2929 -3680 -1553
rect -3646 -2929 -3640 -1553
rect -3686 -2941 -3640 -2929
rect -3488 -1553 -3442 -1541
rect -3488 -2929 -3482 -1553
rect -3448 -2929 -3442 -1553
rect -3488 -2941 -3442 -2929
rect -3290 -1553 -3244 -1541
rect -3290 -2929 -3284 -1553
rect -3250 -2929 -3244 -1553
rect -3290 -2941 -3244 -2929
rect -3092 -1553 -3046 -1541
rect -3092 -2929 -3086 -1553
rect -3052 -2929 -3046 -1553
rect -3092 -2941 -3046 -2929
rect -2894 -1553 -2848 -1541
rect -2894 -2929 -2888 -1553
rect -2854 -2929 -2848 -1553
rect -2894 -2941 -2848 -2929
rect -2696 -1553 -2650 -1541
rect -2696 -2929 -2690 -1553
rect -2656 -2929 -2650 -1553
rect -2696 -2941 -2650 -2929
rect -2498 -1553 -2452 -1541
rect -2498 -2929 -2492 -1553
rect -2458 -2929 -2452 -1553
rect -2498 -2941 -2452 -2929
rect -2300 -1553 -2254 -1541
rect -2300 -2929 -2294 -1553
rect -2260 -2929 -2254 -1553
rect -2300 -2941 -2254 -2929
rect -2102 -1553 -2056 -1541
rect -2102 -2929 -2096 -1553
rect -2062 -2929 -2056 -1553
rect -2102 -2941 -2056 -2929
rect -1904 -1553 -1858 -1541
rect -1904 -2929 -1898 -1553
rect -1864 -2929 -1858 -1553
rect -1904 -2941 -1858 -2929
rect -1706 -1553 -1660 -1541
rect -1706 -2929 -1700 -1553
rect -1666 -2929 -1660 -1553
rect -1706 -2941 -1660 -2929
rect -1508 -1553 -1462 -1541
rect -1508 -2929 -1502 -1553
rect -1468 -2929 -1462 -1553
rect -1508 -2941 -1462 -2929
rect -1310 -1553 -1264 -1541
rect -1310 -2929 -1304 -1553
rect -1270 -2929 -1264 -1553
rect -1310 -2941 -1264 -2929
rect -1112 -1553 -1066 -1541
rect -1112 -2929 -1106 -1553
rect -1072 -2929 -1066 -1553
rect -1112 -2941 -1066 -2929
rect -914 -1553 -868 -1541
rect -914 -2929 -908 -1553
rect -874 -2929 -868 -1553
rect -914 -2941 -868 -2929
rect -716 -1553 -670 -1541
rect -716 -2929 -710 -1553
rect -676 -2929 -670 -1553
rect -716 -2941 -670 -2929
rect -518 -1553 -472 -1541
rect -518 -2929 -512 -1553
rect -478 -2929 -472 -1553
rect -518 -2941 -472 -2929
rect -320 -1553 -274 -1541
rect -320 -2929 -314 -1553
rect -280 -2929 -274 -1553
rect -320 -2941 -274 -2929
rect -122 -1553 -76 -1541
rect -122 -2929 -116 -1553
rect -82 -2929 -76 -1553
rect -122 -2941 -76 -2929
rect 76 -1553 122 -1541
rect 76 -2929 82 -1553
rect 116 -2929 122 -1553
rect 76 -2941 122 -2929
rect 274 -1553 320 -1541
rect 274 -2929 280 -1553
rect 314 -2929 320 -1553
rect 274 -2941 320 -2929
rect 472 -1553 518 -1541
rect 472 -2929 478 -1553
rect 512 -2929 518 -1553
rect 472 -2941 518 -2929
rect 670 -1553 716 -1541
rect 670 -2929 676 -1553
rect 710 -2929 716 -1553
rect 670 -2941 716 -2929
rect 868 -1553 914 -1541
rect 868 -2929 874 -1553
rect 908 -2929 914 -1553
rect 868 -2941 914 -2929
rect 1066 -1553 1112 -1541
rect 1066 -2929 1072 -1553
rect 1106 -2929 1112 -1553
rect 1066 -2941 1112 -2929
rect 1264 -1553 1310 -1541
rect 1264 -2929 1270 -1553
rect 1304 -2929 1310 -1553
rect 1264 -2941 1310 -2929
rect 1462 -1553 1508 -1541
rect 1462 -2929 1468 -1553
rect 1502 -2929 1508 -1553
rect 1462 -2941 1508 -2929
rect 1660 -1553 1706 -1541
rect 1660 -2929 1666 -1553
rect 1700 -2929 1706 -1553
rect 1660 -2941 1706 -2929
rect 1858 -1553 1904 -1541
rect 1858 -2929 1864 -1553
rect 1898 -2929 1904 -1553
rect 1858 -2941 1904 -2929
rect 2056 -1553 2102 -1541
rect 2056 -2929 2062 -1553
rect 2096 -2929 2102 -1553
rect 2056 -2941 2102 -2929
rect 2254 -1553 2300 -1541
rect 2254 -2929 2260 -1553
rect 2294 -2929 2300 -1553
rect 2254 -2941 2300 -2929
rect 2452 -1553 2498 -1541
rect 2452 -2929 2458 -1553
rect 2492 -2929 2498 -1553
rect 2452 -2941 2498 -2929
rect 2650 -1553 2696 -1541
rect 2650 -2929 2656 -1553
rect 2690 -2929 2696 -1553
rect 2650 -2941 2696 -2929
rect 2848 -1553 2894 -1541
rect 2848 -2929 2854 -1553
rect 2888 -2929 2894 -1553
rect 2848 -2941 2894 -2929
rect 3046 -1553 3092 -1541
rect 3046 -2929 3052 -1553
rect 3086 -2929 3092 -1553
rect 3046 -2941 3092 -2929
rect 3244 -1553 3290 -1541
rect 3244 -2929 3250 -1553
rect 3284 -2929 3290 -1553
rect 3244 -2941 3290 -2929
rect 3442 -1553 3488 -1541
rect 3442 -2929 3448 -1553
rect 3482 -2929 3488 -1553
rect 3442 -2941 3488 -2929
rect 3640 -1553 3686 -1541
rect 3640 -2929 3646 -1553
rect 3680 -2929 3686 -1553
rect 3640 -2941 3686 -2929
rect 3838 -1553 3884 -1541
rect 3838 -2929 3844 -1553
rect 3878 -2929 3884 -1553
rect 3838 -2941 3884 -2929
rect 4036 -1553 4082 -1541
rect 4036 -2929 4042 -1553
rect 4076 -2929 4082 -1553
rect 4036 -2941 4082 -2929
rect 4234 -1553 4280 -1541
rect 4234 -2929 4240 -1553
rect 4274 -2929 4280 -1553
rect 4234 -2941 4280 -2929
rect 4432 -1553 4478 -1541
rect 4432 -2929 4438 -1553
rect 4472 -2929 4478 -1553
rect 4432 -2941 4478 -2929
rect 4630 -1553 4676 -1541
rect 4630 -2929 4636 -1553
rect 4670 -2929 4676 -1553
rect 4630 -2941 4676 -2929
rect 4828 -1553 4874 -1541
rect 4828 -2929 4834 -1553
rect 4868 -2929 4874 -1553
rect 4828 -2941 4874 -2929
rect 5026 -1553 5072 -1541
rect 5026 -2929 5032 -1553
rect 5066 -2929 5072 -1553
rect 5026 -2941 5072 -2929
rect 5224 -1553 5270 -1541
rect 5224 -2929 5230 -1553
rect 5264 -2929 5270 -1553
rect 5224 -2941 5270 -2929
rect 5422 -1553 5468 -1541
rect 5422 -2929 5428 -1553
rect 5462 -2929 5468 -1553
rect 5422 -2941 5468 -2929
rect 5620 -1553 5666 -1541
rect 5620 -2929 5626 -1553
rect 5660 -2929 5666 -1553
rect 5620 -2941 5666 -2929
rect 5818 -1553 5864 -1541
rect 5818 -2929 5824 -1553
rect 5858 -2929 5864 -1553
rect 5818 -2941 5864 -2929
rect 6016 -1553 6062 -1541
rect 6016 -2929 6022 -1553
rect 6056 -2929 6062 -1553
rect 6016 -2941 6062 -2929
rect 6214 -1553 6260 -1541
rect 6214 -2929 6220 -1553
rect 6254 -2929 6260 -1553
rect 6214 -2941 6260 -2929
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 4 nf 63 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
