magic
tech sky130A
magscale 1 2
timestamp 1616092564
<< nwell >>
rect -6965 -462 6965 462
<< pmoslvt >>
rect -6871 -400 -6791 400
rect -6733 -400 -6653 400
rect -6595 -400 -6515 400
rect -6457 -400 -6377 400
rect -6319 -400 -6239 400
rect -6181 -400 -6101 400
rect -6043 -400 -5963 400
rect -5905 -400 -5825 400
rect -5767 -400 -5687 400
rect -5629 -400 -5549 400
rect -5491 -400 -5411 400
rect -5353 -400 -5273 400
rect -5215 -400 -5135 400
rect -5077 -400 -4997 400
rect -4939 -400 -4859 400
rect -4801 -400 -4721 400
rect -4663 -400 -4583 400
rect -4525 -400 -4445 400
rect -4387 -400 -4307 400
rect -4249 -400 -4169 400
rect -4111 -400 -4031 400
rect -3973 -400 -3893 400
rect -3835 -400 -3755 400
rect -3697 -400 -3617 400
rect -3559 -400 -3479 400
rect -3421 -400 -3341 400
rect -3283 -400 -3203 400
rect -3145 -400 -3065 400
rect -3007 -400 -2927 400
rect -2869 -400 -2789 400
rect -2731 -400 -2651 400
rect -2593 -400 -2513 400
rect -2455 -400 -2375 400
rect -2317 -400 -2237 400
rect -2179 -400 -2099 400
rect -2041 -400 -1961 400
rect -1903 -400 -1823 400
rect -1765 -400 -1685 400
rect -1627 -400 -1547 400
rect -1489 -400 -1409 400
rect -1351 -400 -1271 400
rect -1213 -400 -1133 400
rect -1075 -400 -995 400
rect -937 -400 -857 400
rect -799 -400 -719 400
rect -661 -400 -581 400
rect -523 -400 -443 400
rect -385 -400 -305 400
rect -247 -400 -167 400
rect -109 -400 -29 400
rect 29 -400 109 400
rect 167 -400 247 400
rect 305 -400 385 400
rect 443 -400 523 400
rect 581 -400 661 400
rect 719 -400 799 400
rect 857 -400 937 400
rect 995 -400 1075 400
rect 1133 -400 1213 400
rect 1271 -400 1351 400
rect 1409 -400 1489 400
rect 1547 -400 1627 400
rect 1685 -400 1765 400
rect 1823 -400 1903 400
rect 1961 -400 2041 400
rect 2099 -400 2179 400
rect 2237 -400 2317 400
rect 2375 -400 2455 400
rect 2513 -400 2593 400
rect 2651 -400 2731 400
rect 2789 -400 2869 400
rect 2927 -400 3007 400
rect 3065 -400 3145 400
rect 3203 -400 3283 400
rect 3341 -400 3421 400
rect 3479 -400 3559 400
rect 3617 -400 3697 400
rect 3755 -400 3835 400
rect 3893 -400 3973 400
rect 4031 -400 4111 400
rect 4169 -400 4249 400
rect 4307 -400 4387 400
rect 4445 -400 4525 400
rect 4583 -400 4663 400
rect 4721 -400 4801 400
rect 4859 -400 4939 400
rect 4997 -400 5077 400
rect 5135 -400 5215 400
rect 5273 -400 5353 400
rect 5411 -400 5491 400
rect 5549 -400 5629 400
rect 5687 -400 5767 400
rect 5825 -400 5905 400
rect 5963 -400 6043 400
rect 6101 -400 6181 400
rect 6239 -400 6319 400
rect 6377 -400 6457 400
rect 6515 -400 6595 400
rect 6653 -400 6733 400
rect 6791 -400 6871 400
<< pdiff >>
rect -6929 388 -6871 400
rect -6929 -388 -6917 388
rect -6883 -388 -6871 388
rect -6929 -400 -6871 -388
rect -6791 388 -6733 400
rect -6791 -388 -6779 388
rect -6745 -388 -6733 388
rect -6791 -400 -6733 -388
rect -6653 388 -6595 400
rect -6653 -388 -6641 388
rect -6607 -388 -6595 388
rect -6653 -400 -6595 -388
rect -6515 388 -6457 400
rect -6515 -388 -6503 388
rect -6469 -388 -6457 388
rect -6515 -400 -6457 -388
rect -6377 388 -6319 400
rect -6377 -388 -6365 388
rect -6331 -388 -6319 388
rect -6377 -400 -6319 -388
rect -6239 388 -6181 400
rect -6239 -388 -6227 388
rect -6193 -388 -6181 388
rect -6239 -400 -6181 -388
rect -6101 388 -6043 400
rect -6101 -388 -6089 388
rect -6055 -388 -6043 388
rect -6101 -400 -6043 -388
rect -5963 388 -5905 400
rect -5963 -388 -5951 388
rect -5917 -388 -5905 388
rect -5963 -400 -5905 -388
rect -5825 388 -5767 400
rect -5825 -388 -5813 388
rect -5779 -388 -5767 388
rect -5825 -400 -5767 -388
rect -5687 388 -5629 400
rect -5687 -388 -5675 388
rect -5641 -388 -5629 388
rect -5687 -400 -5629 -388
rect -5549 388 -5491 400
rect -5549 -388 -5537 388
rect -5503 -388 -5491 388
rect -5549 -400 -5491 -388
rect -5411 388 -5353 400
rect -5411 -388 -5399 388
rect -5365 -388 -5353 388
rect -5411 -400 -5353 -388
rect -5273 388 -5215 400
rect -5273 -388 -5261 388
rect -5227 -388 -5215 388
rect -5273 -400 -5215 -388
rect -5135 388 -5077 400
rect -5135 -388 -5123 388
rect -5089 -388 -5077 388
rect -5135 -400 -5077 -388
rect -4997 388 -4939 400
rect -4997 -388 -4985 388
rect -4951 -388 -4939 388
rect -4997 -400 -4939 -388
rect -4859 388 -4801 400
rect -4859 -388 -4847 388
rect -4813 -388 -4801 388
rect -4859 -400 -4801 -388
rect -4721 388 -4663 400
rect -4721 -388 -4709 388
rect -4675 -388 -4663 388
rect -4721 -400 -4663 -388
rect -4583 388 -4525 400
rect -4583 -388 -4571 388
rect -4537 -388 -4525 388
rect -4583 -400 -4525 -388
rect -4445 388 -4387 400
rect -4445 -388 -4433 388
rect -4399 -388 -4387 388
rect -4445 -400 -4387 -388
rect -4307 388 -4249 400
rect -4307 -388 -4295 388
rect -4261 -388 -4249 388
rect -4307 -400 -4249 -388
rect -4169 388 -4111 400
rect -4169 -388 -4157 388
rect -4123 -388 -4111 388
rect -4169 -400 -4111 -388
rect -4031 388 -3973 400
rect -4031 -388 -4019 388
rect -3985 -388 -3973 388
rect -4031 -400 -3973 -388
rect -3893 388 -3835 400
rect -3893 -388 -3881 388
rect -3847 -388 -3835 388
rect -3893 -400 -3835 -388
rect -3755 388 -3697 400
rect -3755 -388 -3743 388
rect -3709 -388 -3697 388
rect -3755 -400 -3697 -388
rect -3617 388 -3559 400
rect -3617 -388 -3605 388
rect -3571 -388 -3559 388
rect -3617 -400 -3559 -388
rect -3479 388 -3421 400
rect -3479 -388 -3467 388
rect -3433 -388 -3421 388
rect -3479 -400 -3421 -388
rect -3341 388 -3283 400
rect -3341 -388 -3329 388
rect -3295 -388 -3283 388
rect -3341 -400 -3283 -388
rect -3203 388 -3145 400
rect -3203 -388 -3191 388
rect -3157 -388 -3145 388
rect -3203 -400 -3145 -388
rect -3065 388 -3007 400
rect -3065 -388 -3053 388
rect -3019 -388 -3007 388
rect -3065 -400 -3007 -388
rect -2927 388 -2869 400
rect -2927 -388 -2915 388
rect -2881 -388 -2869 388
rect -2927 -400 -2869 -388
rect -2789 388 -2731 400
rect -2789 -388 -2777 388
rect -2743 -388 -2731 388
rect -2789 -400 -2731 -388
rect -2651 388 -2593 400
rect -2651 -388 -2639 388
rect -2605 -388 -2593 388
rect -2651 -400 -2593 -388
rect -2513 388 -2455 400
rect -2513 -388 -2501 388
rect -2467 -388 -2455 388
rect -2513 -400 -2455 -388
rect -2375 388 -2317 400
rect -2375 -388 -2363 388
rect -2329 -388 -2317 388
rect -2375 -400 -2317 -388
rect -2237 388 -2179 400
rect -2237 -388 -2225 388
rect -2191 -388 -2179 388
rect -2237 -400 -2179 -388
rect -2099 388 -2041 400
rect -2099 -388 -2087 388
rect -2053 -388 -2041 388
rect -2099 -400 -2041 -388
rect -1961 388 -1903 400
rect -1961 -388 -1949 388
rect -1915 -388 -1903 388
rect -1961 -400 -1903 -388
rect -1823 388 -1765 400
rect -1823 -388 -1811 388
rect -1777 -388 -1765 388
rect -1823 -400 -1765 -388
rect -1685 388 -1627 400
rect -1685 -388 -1673 388
rect -1639 -388 -1627 388
rect -1685 -400 -1627 -388
rect -1547 388 -1489 400
rect -1547 -388 -1535 388
rect -1501 -388 -1489 388
rect -1547 -400 -1489 -388
rect -1409 388 -1351 400
rect -1409 -388 -1397 388
rect -1363 -388 -1351 388
rect -1409 -400 -1351 -388
rect -1271 388 -1213 400
rect -1271 -388 -1259 388
rect -1225 -388 -1213 388
rect -1271 -400 -1213 -388
rect -1133 388 -1075 400
rect -1133 -388 -1121 388
rect -1087 -388 -1075 388
rect -1133 -400 -1075 -388
rect -995 388 -937 400
rect -995 -388 -983 388
rect -949 -388 -937 388
rect -995 -400 -937 -388
rect -857 388 -799 400
rect -857 -388 -845 388
rect -811 -388 -799 388
rect -857 -400 -799 -388
rect -719 388 -661 400
rect -719 -388 -707 388
rect -673 -388 -661 388
rect -719 -400 -661 -388
rect -581 388 -523 400
rect -581 -388 -569 388
rect -535 -388 -523 388
rect -581 -400 -523 -388
rect -443 388 -385 400
rect -443 -388 -431 388
rect -397 -388 -385 388
rect -443 -400 -385 -388
rect -305 388 -247 400
rect -305 -388 -293 388
rect -259 -388 -247 388
rect -305 -400 -247 -388
rect -167 388 -109 400
rect -167 -388 -155 388
rect -121 -388 -109 388
rect -167 -400 -109 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 109 388 167 400
rect 109 -388 121 388
rect 155 -388 167 388
rect 109 -400 167 -388
rect 247 388 305 400
rect 247 -388 259 388
rect 293 -388 305 388
rect 247 -400 305 -388
rect 385 388 443 400
rect 385 -388 397 388
rect 431 -388 443 388
rect 385 -400 443 -388
rect 523 388 581 400
rect 523 -388 535 388
rect 569 -388 581 388
rect 523 -400 581 -388
rect 661 388 719 400
rect 661 -388 673 388
rect 707 -388 719 388
rect 661 -400 719 -388
rect 799 388 857 400
rect 799 -388 811 388
rect 845 -388 857 388
rect 799 -400 857 -388
rect 937 388 995 400
rect 937 -388 949 388
rect 983 -388 995 388
rect 937 -400 995 -388
rect 1075 388 1133 400
rect 1075 -388 1087 388
rect 1121 -388 1133 388
rect 1075 -400 1133 -388
rect 1213 388 1271 400
rect 1213 -388 1225 388
rect 1259 -388 1271 388
rect 1213 -400 1271 -388
rect 1351 388 1409 400
rect 1351 -388 1363 388
rect 1397 -388 1409 388
rect 1351 -400 1409 -388
rect 1489 388 1547 400
rect 1489 -388 1501 388
rect 1535 -388 1547 388
rect 1489 -400 1547 -388
rect 1627 388 1685 400
rect 1627 -388 1639 388
rect 1673 -388 1685 388
rect 1627 -400 1685 -388
rect 1765 388 1823 400
rect 1765 -388 1777 388
rect 1811 -388 1823 388
rect 1765 -400 1823 -388
rect 1903 388 1961 400
rect 1903 -388 1915 388
rect 1949 -388 1961 388
rect 1903 -400 1961 -388
rect 2041 388 2099 400
rect 2041 -388 2053 388
rect 2087 -388 2099 388
rect 2041 -400 2099 -388
rect 2179 388 2237 400
rect 2179 -388 2191 388
rect 2225 -388 2237 388
rect 2179 -400 2237 -388
rect 2317 388 2375 400
rect 2317 -388 2329 388
rect 2363 -388 2375 388
rect 2317 -400 2375 -388
rect 2455 388 2513 400
rect 2455 -388 2467 388
rect 2501 -388 2513 388
rect 2455 -400 2513 -388
rect 2593 388 2651 400
rect 2593 -388 2605 388
rect 2639 -388 2651 388
rect 2593 -400 2651 -388
rect 2731 388 2789 400
rect 2731 -388 2743 388
rect 2777 -388 2789 388
rect 2731 -400 2789 -388
rect 2869 388 2927 400
rect 2869 -388 2881 388
rect 2915 -388 2927 388
rect 2869 -400 2927 -388
rect 3007 388 3065 400
rect 3007 -388 3019 388
rect 3053 -388 3065 388
rect 3007 -400 3065 -388
rect 3145 388 3203 400
rect 3145 -388 3157 388
rect 3191 -388 3203 388
rect 3145 -400 3203 -388
rect 3283 388 3341 400
rect 3283 -388 3295 388
rect 3329 -388 3341 388
rect 3283 -400 3341 -388
rect 3421 388 3479 400
rect 3421 -388 3433 388
rect 3467 -388 3479 388
rect 3421 -400 3479 -388
rect 3559 388 3617 400
rect 3559 -388 3571 388
rect 3605 -388 3617 388
rect 3559 -400 3617 -388
rect 3697 388 3755 400
rect 3697 -388 3709 388
rect 3743 -388 3755 388
rect 3697 -400 3755 -388
rect 3835 388 3893 400
rect 3835 -388 3847 388
rect 3881 -388 3893 388
rect 3835 -400 3893 -388
rect 3973 388 4031 400
rect 3973 -388 3985 388
rect 4019 -388 4031 388
rect 3973 -400 4031 -388
rect 4111 388 4169 400
rect 4111 -388 4123 388
rect 4157 -388 4169 388
rect 4111 -400 4169 -388
rect 4249 388 4307 400
rect 4249 -388 4261 388
rect 4295 -388 4307 388
rect 4249 -400 4307 -388
rect 4387 388 4445 400
rect 4387 -388 4399 388
rect 4433 -388 4445 388
rect 4387 -400 4445 -388
rect 4525 388 4583 400
rect 4525 -388 4537 388
rect 4571 -388 4583 388
rect 4525 -400 4583 -388
rect 4663 388 4721 400
rect 4663 -388 4675 388
rect 4709 -388 4721 388
rect 4663 -400 4721 -388
rect 4801 388 4859 400
rect 4801 -388 4813 388
rect 4847 -388 4859 388
rect 4801 -400 4859 -388
rect 4939 388 4997 400
rect 4939 -388 4951 388
rect 4985 -388 4997 388
rect 4939 -400 4997 -388
rect 5077 388 5135 400
rect 5077 -388 5089 388
rect 5123 -388 5135 388
rect 5077 -400 5135 -388
rect 5215 388 5273 400
rect 5215 -388 5227 388
rect 5261 -388 5273 388
rect 5215 -400 5273 -388
rect 5353 388 5411 400
rect 5353 -388 5365 388
rect 5399 -388 5411 388
rect 5353 -400 5411 -388
rect 5491 388 5549 400
rect 5491 -388 5503 388
rect 5537 -388 5549 388
rect 5491 -400 5549 -388
rect 5629 388 5687 400
rect 5629 -388 5641 388
rect 5675 -388 5687 388
rect 5629 -400 5687 -388
rect 5767 388 5825 400
rect 5767 -388 5779 388
rect 5813 -388 5825 388
rect 5767 -400 5825 -388
rect 5905 388 5963 400
rect 5905 -388 5917 388
rect 5951 -388 5963 388
rect 5905 -400 5963 -388
rect 6043 388 6101 400
rect 6043 -388 6055 388
rect 6089 -388 6101 388
rect 6043 -400 6101 -388
rect 6181 388 6239 400
rect 6181 -388 6193 388
rect 6227 -388 6239 388
rect 6181 -400 6239 -388
rect 6319 388 6377 400
rect 6319 -388 6331 388
rect 6365 -388 6377 388
rect 6319 -400 6377 -388
rect 6457 388 6515 400
rect 6457 -388 6469 388
rect 6503 -388 6515 388
rect 6457 -400 6515 -388
rect 6595 388 6653 400
rect 6595 -388 6607 388
rect 6641 -388 6653 388
rect 6595 -400 6653 -388
rect 6733 388 6791 400
rect 6733 -388 6745 388
rect 6779 -388 6791 388
rect 6733 -400 6791 -388
rect 6871 388 6929 400
rect 6871 -388 6883 388
rect 6917 -388 6929 388
rect 6871 -400 6929 -388
<< pdiffc >>
rect -6917 -388 -6883 388
rect -6779 -388 -6745 388
rect -6641 -388 -6607 388
rect -6503 -388 -6469 388
rect -6365 -388 -6331 388
rect -6227 -388 -6193 388
rect -6089 -388 -6055 388
rect -5951 -388 -5917 388
rect -5813 -388 -5779 388
rect -5675 -388 -5641 388
rect -5537 -388 -5503 388
rect -5399 -388 -5365 388
rect -5261 -388 -5227 388
rect -5123 -388 -5089 388
rect -4985 -388 -4951 388
rect -4847 -388 -4813 388
rect -4709 -388 -4675 388
rect -4571 -388 -4537 388
rect -4433 -388 -4399 388
rect -4295 -388 -4261 388
rect -4157 -388 -4123 388
rect -4019 -388 -3985 388
rect -3881 -388 -3847 388
rect -3743 -388 -3709 388
rect -3605 -388 -3571 388
rect -3467 -388 -3433 388
rect -3329 -388 -3295 388
rect -3191 -388 -3157 388
rect -3053 -388 -3019 388
rect -2915 -388 -2881 388
rect -2777 -388 -2743 388
rect -2639 -388 -2605 388
rect -2501 -388 -2467 388
rect -2363 -388 -2329 388
rect -2225 -388 -2191 388
rect -2087 -388 -2053 388
rect -1949 -388 -1915 388
rect -1811 -388 -1777 388
rect -1673 -388 -1639 388
rect -1535 -388 -1501 388
rect -1397 -388 -1363 388
rect -1259 -388 -1225 388
rect -1121 -388 -1087 388
rect -983 -388 -949 388
rect -845 -388 -811 388
rect -707 -388 -673 388
rect -569 -388 -535 388
rect -431 -388 -397 388
rect -293 -388 -259 388
rect -155 -388 -121 388
rect -17 -388 17 388
rect 121 -388 155 388
rect 259 -388 293 388
rect 397 -388 431 388
rect 535 -388 569 388
rect 673 -388 707 388
rect 811 -388 845 388
rect 949 -388 983 388
rect 1087 -388 1121 388
rect 1225 -388 1259 388
rect 1363 -388 1397 388
rect 1501 -388 1535 388
rect 1639 -388 1673 388
rect 1777 -388 1811 388
rect 1915 -388 1949 388
rect 2053 -388 2087 388
rect 2191 -388 2225 388
rect 2329 -388 2363 388
rect 2467 -388 2501 388
rect 2605 -388 2639 388
rect 2743 -388 2777 388
rect 2881 -388 2915 388
rect 3019 -388 3053 388
rect 3157 -388 3191 388
rect 3295 -388 3329 388
rect 3433 -388 3467 388
rect 3571 -388 3605 388
rect 3709 -388 3743 388
rect 3847 -388 3881 388
rect 3985 -388 4019 388
rect 4123 -388 4157 388
rect 4261 -388 4295 388
rect 4399 -388 4433 388
rect 4537 -388 4571 388
rect 4675 -388 4709 388
rect 4813 -388 4847 388
rect 4951 -388 4985 388
rect 5089 -388 5123 388
rect 5227 -388 5261 388
rect 5365 -388 5399 388
rect 5503 -388 5537 388
rect 5641 -388 5675 388
rect 5779 -388 5813 388
rect 5917 -388 5951 388
rect 6055 -388 6089 388
rect 6193 -388 6227 388
rect 6331 -388 6365 388
rect 6469 -388 6503 388
rect 6607 -388 6641 388
rect 6745 -388 6779 388
rect 6883 -388 6917 388
<< poly >>
rect -6871 400 -6791 426
rect -6733 400 -6653 426
rect -6595 400 -6515 426
rect -6457 400 -6377 426
rect -6319 400 -6239 426
rect -6181 400 -6101 426
rect -6043 400 -5963 426
rect -5905 400 -5825 426
rect -5767 400 -5687 426
rect -5629 400 -5549 426
rect -5491 400 -5411 426
rect -5353 400 -5273 426
rect -5215 400 -5135 426
rect -5077 400 -4997 426
rect -4939 400 -4859 426
rect -4801 400 -4721 426
rect -4663 400 -4583 426
rect -4525 400 -4445 426
rect -4387 400 -4307 426
rect -4249 400 -4169 426
rect -4111 400 -4031 426
rect -3973 400 -3893 426
rect -3835 400 -3755 426
rect -3697 400 -3617 426
rect -3559 400 -3479 426
rect -3421 400 -3341 426
rect -3283 400 -3203 426
rect -3145 400 -3065 426
rect -3007 400 -2927 426
rect -2869 400 -2789 426
rect -2731 400 -2651 426
rect -2593 400 -2513 426
rect -2455 400 -2375 426
rect -2317 400 -2237 426
rect -2179 400 -2099 426
rect -2041 400 -1961 426
rect -1903 400 -1823 426
rect -1765 400 -1685 426
rect -1627 400 -1547 426
rect -1489 400 -1409 426
rect -1351 400 -1271 426
rect -1213 400 -1133 426
rect -1075 400 -995 426
rect -937 400 -857 426
rect -799 400 -719 426
rect -661 400 -581 426
rect -523 400 -443 426
rect -385 400 -305 426
rect -247 400 -167 426
rect -109 400 -29 426
rect 29 400 109 426
rect 167 400 247 426
rect 305 400 385 426
rect 443 400 523 426
rect 581 400 661 426
rect 719 400 799 426
rect 857 400 937 426
rect 995 400 1075 426
rect 1133 400 1213 426
rect 1271 400 1351 426
rect 1409 400 1489 426
rect 1547 400 1627 426
rect 1685 400 1765 426
rect 1823 400 1903 426
rect 1961 400 2041 426
rect 2099 400 2179 426
rect 2237 400 2317 426
rect 2375 400 2455 426
rect 2513 400 2593 426
rect 2651 400 2731 426
rect 2789 400 2869 426
rect 2927 400 3007 426
rect 3065 400 3145 426
rect 3203 400 3283 426
rect 3341 400 3421 426
rect 3479 400 3559 426
rect 3617 400 3697 426
rect 3755 400 3835 426
rect 3893 400 3973 426
rect 4031 400 4111 426
rect 4169 400 4249 426
rect 4307 400 4387 426
rect 4445 400 4525 426
rect 4583 400 4663 426
rect 4721 400 4801 426
rect 4859 400 4939 426
rect 4997 400 5077 426
rect 5135 400 5215 426
rect 5273 400 5353 426
rect 5411 400 5491 426
rect 5549 400 5629 426
rect 5687 400 5767 426
rect 5825 400 5905 426
rect 5963 400 6043 426
rect 6101 400 6181 426
rect 6239 400 6319 426
rect 6377 400 6457 426
rect 6515 400 6595 426
rect 6653 400 6733 426
rect 6791 400 6871 426
rect -6871 -426 -6791 -400
rect -6733 -426 -6653 -400
rect -6595 -426 -6515 -400
rect -6457 -426 -6377 -400
rect -6319 -426 -6239 -400
rect -6181 -426 -6101 -400
rect -6043 -426 -5963 -400
rect -5905 -426 -5825 -400
rect -5767 -426 -5687 -400
rect -5629 -426 -5549 -400
rect -5491 -426 -5411 -400
rect -5353 -426 -5273 -400
rect -5215 -426 -5135 -400
rect -5077 -426 -4997 -400
rect -4939 -426 -4859 -400
rect -4801 -426 -4721 -400
rect -4663 -426 -4583 -400
rect -4525 -426 -4445 -400
rect -4387 -426 -4307 -400
rect -4249 -426 -4169 -400
rect -4111 -426 -4031 -400
rect -3973 -426 -3893 -400
rect -3835 -426 -3755 -400
rect -3697 -426 -3617 -400
rect -3559 -426 -3479 -400
rect -3421 -426 -3341 -400
rect -3283 -426 -3203 -400
rect -3145 -426 -3065 -400
rect -3007 -426 -2927 -400
rect -2869 -426 -2789 -400
rect -2731 -426 -2651 -400
rect -2593 -426 -2513 -400
rect -2455 -426 -2375 -400
rect -2317 -426 -2237 -400
rect -2179 -426 -2099 -400
rect -2041 -426 -1961 -400
rect -1903 -426 -1823 -400
rect -1765 -426 -1685 -400
rect -1627 -426 -1547 -400
rect -1489 -426 -1409 -400
rect -1351 -426 -1271 -400
rect -1213 -426 -1133 -400
rect -1075 -426 -995 -400
rect -937 -426 -857 -400
rect -799 -426 -719 -400
rect -661 -426 -581 -400
rect -523 -426 -443 -400
rect -385 -426 -305 -400
rect -247 -426 -167 -400
rect -109 -426 -29 -400
rect 29 -426 109 -400
rect 167 -426 247 -400
rect 305 -426 385 -400
rect 443 -426 523 -400
rect 581 -426 661 -400
rect 719 -426 799 -400
rect 857 -426 937 -400
rect 995 -426 1075 -400
rect 1133 -426 1213 -400
rect 1271 -426 1351 -400
rect 1409 -426 1489 -400
rect 1547 -426 1627 -400
rect 1685 -426 1765 -400
rect 1823 -426 1903 -400
rect 1961 -426 2041 -400
rect 2099 -426 2179 -400
rect 2237 -426 2317 -400
rect 2375 -426 2455 -400
rect 2513 -426 2593 -400
rect 2651 -426 2731 -400
rect 2789 -426 2869 -400
rect 2927 -426 3007 -400
rect 3065 -426 3145 -400
rect 3203 -426 3283 -400
rect 3341 -426 3421 -400
rect 3479 -426 3559 -400
rect 3617 -426 3697 -400
rect 3755 -426 3835 -400
rect 3893 -426 3973 -400
rect 4031 -426 4111 -400
rect 4169 -426 4249 -400
rect 4307 -426 4387 -400
rect 4445 -426 4525 -400
rect 4583 -426 4663 -400
rect 4721 -426 4801 -400
rect 4859 -426 4939 -400
rect 4997 -426 5077 -400
rect 5135 -426 5215 -400
rect 5273 -426 5353 -400
rect 5411 -426 5491 -400
rect 5549 -426 5629 -400
rect 5687 -426 5767 -400
rect 5825 -426 5905 -400
rect 5963 -426 6043 -400
rect 6101 -426 6181 -400
rect 6239 -426 6319 -400
rect 6377 -426 6457 -400
rect 6515 -426 6595 -400
rect 6653 -426 6733 -400
rect 6791 -426 6871 -400
<< locali >>
rect -6917 388 -6883 404
rect -6917 -404 -6883 -388
rect -6779 388 -6745 404
rect -6779 -404 -6745 -388
rect -6641 388 -6607 404
rect -6641 -404 -6607 -388
rect -6503 388 -6469 404
rect -6503 -404 -6469 -388
rect -6365 388 -6331 404
rect -6365 -404 -6331 -388
rect -6227 388 -6193 404
rect -6227 -404 -6193 -388
rect -6089 388 -6055 404
rect -6089 -404 -6055 -388
rect -5951 388 -5917 404
rect -5951 -404 -5917 -388
rect -5813 388 -5779 404
rect -5813 -404 -5779 -388
rect -5675 388 -5641 404
rect -5675 -404 -5641 -388
rect -5537 388 -5503 404
rect -5537 -404 -5503 -388
rect -5399 388 -5365 404
rect -5399 -404 -5365 -388
rect -5261 388 -5227 404
rect -5261 -404 -5227 -388
rect -5123 388 -5089 404
rect -5123 -404 -5089 -388
rect -4985 388 -4951 404
rect -4985 -404 -4951 -388
rect -4847 388 -4813 404
rect -4847 -404 -4813 -388
rect -4709 388 -4675 404
rect -4709 -404 -4675 -388
rect -4571 388 -4537 404
rect -4571 -404 -4537 -388
rect -4433 388 -4399 404
rect -4433 -404 -4399 -388
rect -4295 388 -4261 404
rect -4295 -404 -4261 -388
rect -4157 388 -4123 404
rect -4157 -404 -4123 -388
rect -4019 388 -3985 404
rect -4019 -404 -3985 -388
rect -3881 388 -3847 404
rect -3881 -404 -3847 -388
rect -3743 388 -3709 404
rect -3743 -404 -3709 -388
rect -3605 388 -3571 404
rect -3605 -404 -3571 -388
rect -3467 388 -3433 404
rect -3467 -404 -3433 -388
rect -3329 388 -3295 404
rect -3329 -404 -3295 -388
rect -3191 388 -3157 404
rect -3191 -404 -3157 -388
rect -3053 388 -3019 404
rect -3053 -404 -3019 -388
rect -2915 388 -2881 404
rect -2915 -404 -2881 -388
rect -2777 388 -2743 404
rect -2777 -404 -2743 -388
rect -2639 388 -2605 404
rect -2639 -404 -2605 -388
rect -2501 388 -2467 404
rect -2501 -404 -2467 -388
rect -2363 388 -2329 404
rect -2363 -404 -2329 -388
rect -2225 388 -2191 404
rect -2225 -404 -2191 -388
rect -2087 388 -2053 404
rect -2087 -404 -2053 -388
rect -1949 388 -1915 404
rect -1949 -404 -1915 -388
rect -1811 388 -1777 404
rect -1811 -404 -1777 -388
rect -1673 388 -1639 404
rect -1673 -404 -1639 -388
rect -1535 388 -1501 404
rect -1535 -404 -1501 -388
rect -1397 388 -1363 404
rect -1397 -404 -1363 -388
rect -1259 388 -1225 404
rect -1259 -404 -1225 -388
rect -1121 388 -1087 404
rect -1121 -404 -1087 -388
rect -983 388 -949 404
rect -983 -404 -949 -388
rect -845 388 -811 404
rect -845 -404 -811 -388
rect -707 388 -673 404
rect -707 -404 -673 -388
rect -569 388 -535 404
rect -569 -404 -535 -388
rect -431 388 -397 404
rect -431 -404 -397 -388
rect -293 388 -259 404
rect -293 -404 -259 -388
rect -155 388 -121 404
rect -155 -404 -121 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 121 388 155 404
rect 121 -404 155 -388
rect 259 388 293 404
rect 259 -404 293 -388
rect 397 388 431 404
rect 397 -404 431 -388
rect 535 388 569 404
rect 535 -404 569 -388
rect 673 388 707 404
rect 673 -404 707 -388
rect 811 388 845 404
rect 811 -404 845 -388
rect 949 388 983 404
rect 949 -404 983 -388
rect 1087 388 1121 404
rect 1087 -404 1121 -388
rect 1225 388 1259 404
rect 1225 -404 1259 -388
rect 1363 388 1397 404
rect 1363 -404 1397 -388
rect 1501 388 1535 404
rect 1501 -404 1535 -388
rect 1639 388 1673 404
rect 1639 -404 1673 -388
rect 1777 388 1811 404
rect 1777 -404 1811 -388
rect 1915 388 1949 404
rect 1915 -404 1949 -388
rect 2053 388 2087 404
rect 2053 -404 2087 -388
rect 2191 388 2225 404
rect 2191 -404 2225 -388
rect 2329 388 2363 404
rect 2329 -404 2363 -388
rect 2467 388 2501 404
rect 2467 -404 2501 -388
rect 2605 388 2639 404
rect 2605 -404 2639 -388
rect 2743 388 2777 404
rect 2743 -404 2777 -388
rect 2881 388 2915 404
rect 2881 -404 2915 -388
rect 3019 388 3053 404
rect 3019 -404 3053 -388
rect 3157 388 3191 404
rect 3157 -404 3191 -388
rect 3295 388 3329 404
rect 3295 -404 3329 -388
rect 3433 388 3467 404
rect 3433 -404 3467 -388
rect 3571 388 3605 404
rect 3571 -404 3605 -388
rect 3709 388 3743 404
rect 3709 -404 3743 -388
rect 3847 388 3881 404
rect 3847 -404 3881 -388
rect 3985 388 4019 404
rect 3985 -404 4019 -388
rect 4123 388 4157 404
rect 4123 -404 4157 -388
rect 4261 388 4295 404
rect 4261 -404 4295 -388
rect 4399 388 4433 404
rect 4399 -404 4433 -388
rect 4537 388 4571 404
rect 4537 -404 4571 -388
rect 4675 388 4709 404
rect 4675 -404 4709 -388
rect 4813 388 4847 404
rect 4813 -404 4847 -388
rect 4951 388 4985 404
rect 4951 -404 4985 -388
rect 5089 388 5123 404
rect 5089 -404 5123 -388
rect 5227 388 5261 404
rect 5227 -404 5261 -388
rect 5365 388 5399 404
rect 5365 -404 5399 -388
rect 5503 388 5537 404
rect 5503 -404 5537 -388
rect 5641 388 5675 404
rect 5641 -404 5675 -388
rect 5779 388 5813 404
rect 5779 -404 5813 -388
rect 5917 388 5951 404
rect 5917 -404 5951 -388
rect 6055 388 6089 404
rect 6055 -404 6089 -388
rect 6193 388 6227 404
rect 6193 -404 6227 -388
rect 6331 388 6365 404
rect 6331 -404 6365 -388
rect 6469 388 6503 404
rect 6469 -404 6503 -388
rect 6607 388 6641 404
rect 6607 -404 6641 -388
rect 6745 388 6779 404
rect 6745 -404 6779 -388
rect 6883 388 6917 404
rect 6883 -404 6917 -388
<< viali >>
rect -6917 -388 -6883 388
rect -6779 -388 -6745 388
rect -6641 -388 -6607 388
rect -6503 -388 -6469 388
rect -6365 -388 -6331 388
rect -6227 -388 -6193 388
rect -6089 -388 -6055 388
rect -5951 -388 -5917 388
rect -5813 -388 -5779 388
rect -5675 -388 -5641 388
rect -5537 -388 -5503 388
rect -5399 -388 -5365 388
rect -5261 -388 -5227 388
rect -5123 -388 -5089 388
rect -4985 -388 -4951 388
rect -4847 -388 -4813 388
rect -4709 -388 -4675 388
rect -4571 -388 -4537 388
rect -4433 -388 -4399 388
rect -4295 -388 -4261 388
rect -4157 -388 -4123 388
rect -4019 -388 -3985 388
rect -3881 -388 -3847 388
rect -3743 -388 -3709 388
rect -3605 -388 -3571 388
rect -3467 -388 -3433 388
rect -3329 -388 -3295 388
rect -3191 -388 -3157 388
rect -3053 -388 -3019 388
rect -2915 -388 -2881 388
rect -2777 -388 -2743 388
rect -2639 -388 -2605 388
rect -2501 -388 -2467 388
rect -2363 -388 -2329 388
rect -2225 -388 -2191 388
rect -2087 -388 -2053 388
rect -1949 -388 -1915 388
rect -1811 -388 -1777 388
rect -1673 -388 -1639 388
rect -1535 -388 -1501 388
rect -1397 -388 -1363 388
rect -1259 -388 -1225 388
rect -1121 -388 -1087 388
rect -983 -388 -949 388
rect -845 -388 -811 388
rect -707 -388 -673 388
rect -569 -388 -535 388
rect -431 -388 -397 388
rect -293 -388 -259 388
rect -155 -388 -121 388
rect -17 -388 17 388
rect 121 -388 155 388
rect 259 -388 293 388
rect 397 -388 431 388
rect 535 -388 569 388
rect 673 -388 707 388
rect 811 -388 845 388
rect 949 -388 983 388
rect 1087 -388 1121 388
rect 1225 -388 1259 388
rect 1363 -388 1397 388
rect 1501 -388 1535 388
rect 1639 -388 1673 388
rect 1777 -388 1811 388
rect 1915 -388 1949 388
rect 2053 -388 2087 388
rect 2191 -388 2225 388
rect 2329 -388 2363 388
rect 2467 -388 2501 388
rect 2605 -388 2639 388
rect 2743 -388 2777 388
rect 2881 -388 2915 388
rect 3019 -388 3053 388
rect 3157 -388 3191 388
rect 3295 -388 3329 388
rect 3433 -388 3467 388
rect 3571 -388 3605 388
rect 3709 -388 3743 388
rect 3847 -388 3881 388
rect 3985 -388 4019 388
rect 4123 -388 4157 388
rect 4261 -388 4295 388
rect 4399 -388 4433 388
rect 4537 -388 4571 388
rect 4675 -388 4709 388
rect 4813 -388 4847 388
rect 4951 -388 4985 388
rect 5089 -388 5123 388
rect 5227 -388 5261 388
rect 5365 -388 5399 388
rect 5503 -388 5537 388
rect 5641 -388 5675 388
rect 5779 -388 5813 388
rect 5917 -388 5951 388
rect 6055 -388 6089 388
rect 6193 -388 6227 388
rect 6331 -388 6365 388
rect 6469 -388 6503 388
rect 6607 -388 6641 388
rect 6745 -388 6779 388
rect 6883 -388 6917 388
<< metal1 >>
rect -6923 388 -6877 400
rect -6923 -388 -6917 388
rect -6883 -388 -6877 388
rect -6923 -400 -6877 -388
rect -6785 388 -6739 400
rect -6785 -388 -6779 388
rect -6745 -388 -6739 388
rect -6785 -400 -6739 -388
rect -6647 388 -6601 400
rect -6647 -388 -6641 388
rect -6607 -388 -6601 388
rect -6647 -400 -6601 -388
rect -6509 388 -6463 400
rect -6509 -388 -6503 388
rect -6469 -388 -6463 388
rect -6509 -400 -6463 -388
rect -6371 388 -6325 400
rect -6371 -388 -6365 388
rect -6331 -388 -6325 388
rect -6371 -400 -6325 -388
rect -6233 388 -6187 400
rect -6233 -388 -6227 388
rect -6193 -388 -6187 388
rect -6233 -400 -6187 -388
rect -6095 388 -6049 400
rect -6095 -388 -6089 388
rect -6055 -388 -6049 388
rect -6095 -400 -6049 -388
rect -5957 388 -5911 400
rect -5957 -388 -5951 388
rect -5917 -388 -5911 388
rect -5957 -400 -5911 -388
rect -5819 388 -5773 400
rect -5819 -388 -5813 388
rect -5779 -388 -5773 388
rect -5819 -400 -5773 -388
rect -5681 388 -5635 400
rect -5681 -388 -5675 388
rect -5641 -388 -5635 388
rect -5681 -400 -5635 -388
rect -5543 388 -5497 400
rect -5543 -388 -5537 388
rect -5503 -388 -5497 388
rect -5543 -400 -5497 -388
rect -5405 388 -5359 400
rect -5405 -388 -5399 388
rect -5365 -388 -5359 388
rect -5405 -400 -5359 -388
rect -5267 388 -5221 400
rect -5267 -388 -5261 388
rect -5227 -388 -5221 388
rect -5267 -400 -5221 -388
rect -5129 388 -5083 400
rect -5129 -388 -5123 388
rect -5089 -388 -5083 388
rect -5129 -400 -5083 -388
rect -4991 388 -4945 400
rect -4991 -388 -4985 388
rect -4951 -388 -4945 388
rect -4991 -400 -4945 -388
rect -4853 388 -4807 400
rect -4853 -388 -4847 388
rect -4813 -388 -4807 388
rect -4853 -400 -4807 -388
rect -4715 388 -4669 400
rect -4715 -388 -4709 388
rect -4675 -388 -4669 388
rect -4715 -400 -4669 -388
rect -4577 388 -4531 400
rect -4577 -388 -4571 388
rect -4537 -388 -4531 388
rect -4577 -400 -4531 -388
rect -4439 388 -4393 400
rect -4439 -388 -4433 388
rect -4399 -388 -4393 388
rect -4439 -400 -4393 -388
rect -4301 388 -4255 400
rect -4301 -388 -4295 388
rect -4261 -388 -4255 388
rect -4301 -400 -4255 -388
rect -4163 388 -4117 400
rect -4163 -388 -4157 388
rect -4123 -388 -4117 388
rect -4163 -400 -4117 -388
rect -4025 388 -3979 400
rect -4025 -388 -4019 388
rect -3985 -388 -3979 388
rect -4025 -400 -3979 -388
rect -3887 388 -3841 400
rect -3887 -388 -3881 388
rect -3847 -388 -3841 388
rect -3887 -400 -3841 -388
rect -3749 388 -3703 400
rect -3749 -388 -3743 388
rect -3709 -388 -3703 388
rect -3749 -400 -3703 -388
rect -3611 388 -3565 400
rect -3611 -388 -3605 388
rect -3571 -388 -3565 388
rect -3611 -400 -3565 -388
rect -3473 388 -3427 400
rect -3473 -388 -3467 388
rect -3433 -388 -3427 388
rect -3473 -400 -3427 -388
rect -3335 388 -3289 400
rect -3335 -388 -3329 388
rect -3295 -388 -3289 388
rect -3335 -400 -3289 -388
rect -3197 388 -3151 400
rect -3197 -388 -3191 388
rect -3157 -388 -3151 388
rect -3197 -400 -3151 -388
rect -3059 388 -3013 400
rect -3059 -388 -3053 388
rect -3019 -388 -3013 388
rect -3059 -400 -3013 -388
rect -2921 388 -2875 400
rect -2921 -388 -2915 388
rect -2881 -388 -2875 388
rect -2921 -400 -2875 -388
rect -2783 388 -2737 400
rect -2783 -388 -2777 388
rect -2743 -388 -2737 388
rect -2783 -400 -2737 -388
rect -2645 388 -2599 400
rect -2645 -388 -2639 388
rect -2605 -388 -2599 388
rect -2645 -400 -2599 -388
rect -2507 388 -2461 400
rect -2507 -388 -2501 388
rect -2467 -388 -2461 388
rect -2507 -400 -2461 -388
rect -2369 388 -2323 400
rect -2369 -388 -2363 388
rect -2329 -388 -2323 388
rect -2369 -400 -2323 -388
rect -2231 388 -2185 400
rect -2231 -388 -2225 388
rect -2191 -388 -2185 388
rect -2231 -400 -2185 -388
rect -2093 388 -2047 400
rect -2093 -388 -2087 388
rect -2053 -388 -2047 388
rect -2093 -400 -2047 -388
rect -1955 388 -1909 400
rect -1955 -388 -1949 388
rect -1915 -388 -1909 388
rect -1955 -400 -1909 -388
rect -1817 388 -1771 400
rect -1817 -388 -1811 388
rect -1777 -388 -1771 388
rect -1817 -400 -1771 -388
rect -1679 388 -1633 400
rect -1679 -388 -1673 388
rect -1639 -388 -1633 388
rect -1679 -400 -1633 -388
rect -1541 388 -1495 400
rect -1541 -388 -1535 388
rect -1501 -388 -1495 388
rect -1541 -400 -1495 -388
rect -1403 388 -1357 400
rect -1403 -388 -1397 388
rect -1363 -388 -1357 388
rect -1403 -400 -1357 -388
rect -1265 388 -1219 400
rect -1265 -388 -1259 388
rect -1225 -388 -1219 388
rect -1265 -400 -1219 -388
rect -1127 388 -1081 400
rect -1127 -388 -1121 388
rect -1087 -388 -1081 388
rect -1127 -400 -1081 -388
rect -989 388 -943 400
rect -989 -388 -983 388
rect -949 -388 -943 388
rect -989 -400 -943 -388
rect -851 388 -805 400
rect -851 -388 -845 388
rect -811 -388 -805 388
rect -851 -400 -805 -388
rect -713 388 -667 400
rect -713 -388 -707 388
rect -673 -388 -667 388
rect -713 -400 -667 -388
rect -575 388 -529 400
rect -575 -388 -569 388
rect -535 -388 -529 388
rect -575 -400 -529 -388
rect -437 388 -391 400
rect -437 -388 -431 388
rect -397 -388 -391 388
rect -437 -400 -391 -388
rect -299 388 -253 400
rect -299 -388 -293 388
rect -259 -388 -253 388
rect -299 -400 -253 -388
rect -161 388 -115 400
rect -161 -388 -155 388
rect -121 -388 -115 388
rect -161 -400 -115 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 115 388 161 400
rect 115 -388 121 388
rect 155 -388 161 388
rect 115 -400 161 -388
rect 253 388 299 400
rect 253 -388 259 388
rect 293 -388 299 388
rect 253 -400 299 -388
rect 391 388 437 400
rect 391 -388 397 388
rect 431 -388 437 388
rect 391 -400 437 -388
rect 529 388 575 400
rect 529 -388 535 388
rect 569 -388 575 388
rect 529 -400 575 -388
rect 667 388 713 400
rect 667 -388 673 388
rect 707 -388 713 388
rect 667 -400 713 -388
rect 805 388 851 400
rect 805 -388 811 388
rect 845 -388 851 388
rect 805 -400 851 -388
rect 943 388 989 400
rect 943 -388 949 388
rect 983 -388 989 388
rect 943 -400 989 -388
rect 1081 388 1127 400
rect 1081 -388 1087 388
rect 1121 -388 1127 388
rect 1081 -400 1127 -388
rect 1219 388 1265 400
rect 1219 -388 1225 388
rect 1259 -388 1265 388
rect 1219 -400 1265 -388
rect 1357 388 1403 400
rect 1357 -388 1363 388
rect 1397 -388 1403 388
rect 1357 -400 1403 -388
rect 1495 388 1541 400
rect 1495 -388 1501 388
rect 1535 -388 1541 388
rect 1495 -400 1541 -388
rect 1633 388 1679 400
rect 1633 -388 1639 388
rect 1673 -388 1679 388
rect 1633 -400 1679 -388
rect 1771 388 1817 400
rect 1771 -388 1777 388
rect 1811 -388 1817 388
rect 1771 -400 1817 -388
rect 1909 388 1955 400
rect 1909 -388 1915 388
rect 1949 -388 1955 388
rect 1909 -400 1955 -388
rect 2047 388 2093 400
rect 2047 -388 2053 388
rect 2087 -388 2093 388
rect 2047 -400 2093 -388
rect 2185 388 2231 400
rect 2185 -388 2191 388
rect 2225 -388 2231 388
rect 2185 -400 2231 -388
rect 2323 388 2369 400
rect 2323 -388 2329 388
rect 2363 -388 2369 388
rect 2323 -400 2369 -388
rect 2461 388 2507 400
rect 2461 -388 2467 388
rect 2501 -388 2507 388
rect 2461 -400 2507 -388
rect 2599 388 2645 400
rect 2599 -388 2605 388
rect 2639 -388 2645 388
rect 2599 -400 2645 -388
rect 2737 388 2783 400
rect 2737 -388 2743 388
rect 2777 -388 2783 388
rect 2737 -400 2783 -388
rect 2875 388 2921 400
rect 2875 -388 2881 388
rect 2915 -388 2921 388
rect 2875 -400 2921 -388
rect 3013 388 3059 400
rect 3013 -388 3019 388
rect 3053 -388 3059 388
rect 3013 -400 3059 -388
rect 3151 388 3197 400
rect 3151 -388 3157 388
rect 3191 -388 3197 388
rect 3151 -400 3197 -388
rect 3289 388 3335 400
rect 3289 -388 3295 388
rect 3329 -388 3335 388
rect 3289 -400 3335 -388
rect 3427 388 3473 400
rect 3427 -388 3433 388
rect 3467 -388 3473 388
rect 3427 -400 3473 -388
rect 3565 388 3611 400
rect 3565 -388 3571 388
rect 3605 -388 3611 388
rect 3565 -400 3611 -388
rect 3703 388 3749 400
rect 3703 -388 3709 388
rect 3743 -388 3749 388
rect 3703 -400 3749 -388
rect 3841 388 3887 400
rect 3841 -388 3847 388
rect 3881 -388 3887 388
rect 3841 -400 3887 -388
rect 3979 388 4025 400
rect 3979 -388 3985 388
rect 4019 -388 4025 388
rect 3979 -400 4025 -388
rect 4117 388 4163 400
rect 4117 -388 4123 388
rect 4157 -388 4163 388
rect 4117 -400 4163 -388
rect 4255 388 4301 400
rect 4255 -388 4261 388
rect 4295 -388 4301 388
rect 4255 -400 4301 -388
rect 4393 388 4439 400
rect 4393 -388 4399 388
rect 4433 -388 4439 388
rect 4393 -400 4439 -388
rect 4531 388 4577 400
rect 4531 -388 4537 388
rect 4571 -388 4577 388
rect 4531 -400 4577 -388
rect 4669 388 4715 400
rect 4669 -388 4675 388
rect 4709 -388 4715 388
rect 4669 -400 4715 -388
rect 4807 388 4853 400
rect 4807 -388 4813 388
rect 4847 -388 4853 388
rect 4807 -400 4853 -388
rect 4945 388 4991 400
rect 4945 -388 4951 388
rect 4985 -388 4991 388
rect 4945 -400 4991 -388
rect 5083 388 5129 400
rect 5083 -388 5089 388
rect 5123 -388 5129 388
rect 5083 -400 5129 -388
rect 5221 388 5267 400
rect 5221 -388 5227 388
rect 5261 -388 5267 388
rect 5221 -400 5267 -388
rect 5359 388 5405 400
rect 5359 -388 5365 388
rect 5399 -388 5405 388
rect 5359 -400 5405 -388
rect 5497 388 5543 400
rect 5497 -388 5503 388
rect 5537 -388 5543 388
rect 5497 -400 5543 -388
rect 5635 388 5681 400
rect 5635 -388 5641 388
rect 5675 -388 5681 388
rect 5635 -400 5681 -388
rect 5773 388 5819 400
rect 5773 -388 5779 388
rect 5813 -388 5819 388
rect 5773 -400 5819 -388
rect 5911 388 5957 400
rect 5911 -388 5917 388
rect 5951 -388 5957 388
rect 5911 -400 5957 -388
rect 6049 388 6095 400
rect 6049 -388 6055 388
rect 6089 -388 6095 388
rect 6049 -400 6095 -388
rect 6187 388 6233 400
rect 6187 -388 6193 388
rect 6227 -388 6233 388
rect 6187 -400 6233 -388
rect 6325 388 6371 400
rect 6325 -388 6331 388
rect 6365 -388 6371 388
rect 6325 -400 6371 -388
rect 6463 388 6509 400
rect 6463 -388 6469 388
rect 6503 -388 6509 388
rect 6463 -400 6509 -388
rect 6601 388 6647 400
rect 6601 -388 6607 388
rect 6641 -388 6647 388
rect 6601 -400 6647 -388
rect 6739 388 6785 400
rect 6739 -388 6745 388
rect 6779 -388 6785 388
rect 6739 -400 6785 -388
rect 6877 388 6923 400
rect 6877 -388 6883 388
rect 6917 -388 6923 388
rect 6877 -400 6923 -388
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 4 l 0.4 m 1 nf 100 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
