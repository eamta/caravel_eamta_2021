magic
tech sky130A
magscale 1 2
timestamp 1623074401
<< pwell >>
rect -1127 -1110 1127 1110
<< nmos >>
rect -927 -900 -897 900
rect -831 -900 -801 900
rect -735 -900 -705 900
rect -639 -900 -609 900
rect -543 -900 -513 900
rect -447 -900 -417 900
rect -351 -900 -321 900
rect -255 -900 -225 900
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
rect 225 -900 255 900
rect 321 -900 351 900
rect 417 -900 447 900
rect 513 -900 543 900
rect 609 -900 639 900
rect 705 -900 735 900
rect 801 -900 831 900
rect 897 -900 927 900
<< ndiff >>
rect -989 888 -927 900
rect -989 -888 -977 888
rect -943 -888 -927 888
rect -989 -900 -927 -888
rect -897 888 -831 900
rect -897 -888 -881 888
rect -847 -888 -831 888
rect -897 -900 -831 -888
rect -801 888 -735 900
rect -801 -888 -785 888
rect -751 -888 -735 888
rect -801 -900 -735 -888
rect -705 888 -639 900
rect -705 -888 -689 888
rect -655 -888 -639 888
rect -705 -900 -639 -888
rect -609 888 -543 900
rect -609 -888 -593 888
rect -559 -888 -543 888
rect -609 -900 -543 -888
rect -513 888 -447 900
rect -513 -888 -497 888
rect -463 -888 -447 888
rect -513 -900 -447 -888
rect -417 888 -351 900
rect -417 -888 -401 888
rect -367 -888 -351 888
rect -417 -900 -351 -888
rect -321 888 -255 900
rect -321 -888 -305 888
rect -271 -888 -255 888
rect -321 -900 -255 -888
rect -225 888 -159 900
rect -225 -888 -209 888
rect -175 -888 -159 888
rect -225 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 225 900
rect 159 -888 175 888
rect 209 -888 225 888
rect 159 -900 225 -888
rect 255 888 321 900
rect 255 -888 271 888
rect 305 -888 321 888
rect 255 -900 321 -888
rect 351 888 417 900
rect 351 -888 367 888
rect 401 -888 417 888
rect 351 -900 417 -888
rect 447 888 513 900
rect 447 -888 463 888
rect 497 -888 513 888
rect 447 -900 513 -888
rect 543 888 609 900
rect 543 -888 559 888
rect 593 -888 609 888
rect 543 -900 609 -888
rect 639 888 705 900
rect 639 -888 655 888
rect 689 -888 705 888
rect 639 -900 705 -888
rect 735 888 801 900
rect 735 -888 751 888
rect 785 -888 801 888
rect 735 -900 801 -888
rect 831 888 897 900
rect 831 -888 847 888
rect 881 -888 897 888
rect 831 -900 897 -888
rect 927 888 989 900
rect 927 -888 943 888
rect 977 -888 989 888
rect 927 -900 989 -888
<< ndiffc >>
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
<< psubdiff >>
rect -1091 1040 -995 1074
rect 995 1040 1091 1074
rect -1091 978 -1057 1040
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1040
rect -1091 -1074 1091 -1040
<< psubdiffcont >>
rect -995 1040 995 1074
rect -1091 -978 -1057 978
<< poly >>
rect -927 985 940 1002
rect -927 949 -910 985
rect 924 949 940 985
rect -927 922 940 949
rect -927 900 -897 922
rect -831 900 -801 922
rect -735 900 -705 922
rect -639 900 -609 922
rect -543 900 -513 922
rect -447 900 -417 922
rect -351 900 -321 922
rect -255 900 -225 922
rect -159 900 -129 922
rect -63 900 -33 922
rect 33 900 63 922
rect 129 900 159 922
rect 225 900 255 922
rect 321 900 351 922
rect 417 900 447 922
rect 513 900 543 922
rect 609 900 639 922
rect 705 900 735 922
rect 801 900 831 922
rect 897 900 927 922
rect -927 -926 -897 -900
rect -831 -926 -801 -900
rect -735 -926 -705 -900
rect -639 -926 -609 -900
rect -543 -926 -513 -900
rect -447 -926 -417 -900
rect -351 -926 -321 -900
rect -255 -926 -225 -900
rect -159 -926 -129 -900
rect -63 -926 -33 -900
rect 33 -926 63 -900
rect 129 -926 159 -900
rect 225 -926 255 -900
rect 321 -926 351 -900
rect 417 -926 447 -900
rect 513 -926 543 -900
rect 609 -926 639 -900
rect 705 -926 735 -900
rect 801 -926 831 -900
rect 897 -926 927 -900
<< polycont >>
rect -910 949 924 985
<< locali >>
rect -1091 1040 -995 1074
rect 995 1040 1091 1074
rect -1091 978 -1057 1040
rect -926 985 940 996
rect -926 949 -910 985
rect 924 949 940 985
rect -926 939 940 949
rect -977 888 -943 904
rect -977 -904 -943 -888
rect -881 888 -847 904
rect -881 -904 -847 -888
rect -785 888 -751 904
rect -785 -904 -751 -888
rect -689 888 -655 904
rect -689 -904 -655 -888
rect -593 888 -559 904
rect -593 -904 -559 -888
rect -497 888 -463 904
rect -497 -904 -463 -888
rect -401 888 -367 904
rect -401 -904 -367 -888
rect -305 888 -271 904
rect -305 -904 -271 -888
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect 271 888 305 904
rect 271 -904 305 -888
rect 367 888 401 904
rect 367 -904 401 -888
rect 463 888 497 904
rect 463 -904 497 -888
rect 559 888 593 904
rect 559 -904 593 -888
rect 655 888 689 904
rect 655 -904 689 -888
rect 751 888 785 904
rect 751 -904 785 -888
rect 847 888 881 904
rect 847 -904 881 -888
rect 943 888 977 904
rect 943 -904 977 -888
rect -1091 -1040 -1057 -978
rect 1057 -1040 1091 1040
rect -1091 -1074 1091 -1040
<< viali >>
rect -910 949 924 985
rect -977 -888 -943 888
rect -881 -888 -847 888
rect -785 -888 -751 888
rect -689 -888 -655 888
rect -593 -888 -559 888
rect -497 -888 -463 888
rect -401 -888 -367 888
rect -305 -888 -271 888
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect 271 -888 305 888
rect 367 -888 401 888
rect 463 -888 497 888
rect 559 -888 593 888
rect 655 -888 689 888
rect 751 -888 785 888
rect 847 -888 881 888
rect 943 -888 977 888
<< metal1 >>
rect -928 1001 940 1004
rect -928 949 -910 1001
rect 924 949 940 1001
rect -928 939 940 949
rect -1002 -904 -992 904
rect -928 -904 -918 904
rect -887 888 -841 900
rect -887 -888 -881 888
rect -847 -888 -841 888
rect -887 -900 -841 -888
rect -810 -904 -800 904
rect -736 -904 -726 904
rect -695 888 -649 900
rect -695 -888 -689 888
rect -655 -888 -649 888
rect -695 -900 -649 -888
rect -618 -904 -608 904
rect -544 -904 -534 904
rect -503 888 -457 900
rect -503 -888 -497 888
rect -463 -888 -457 888
rect -503 -900 -457 -888
rect -426 -904 -416 904
rect -352 -904 -342 904
rect -311 888 -265 900
rect -311 -888 -305 888
rect -271 -888 -265 888
rect -311 -900 -265 -888
rect -234 -904 -224 904
rect -160 -904 -150 904
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -42 -904 -32 904
rect 32 -904 42 904
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 150 -904 160 904
rect 224 -904 234 904
rect 265 888 311 900
rect 265 -888 271 888
rect 305 -888 311 888
rect 265 -900 311 -888
rect 342 -904 352 904
rect 416 -904 426 904
rect 457 888 503 900
rect 457 -888 463 888
rect 497 -888 503 888
rect 457 -900 503 -888
rect 534 -904 544 904
rect 608 -904 618 904
rect 649 888 695 900
rect 649 -888 655 888
rect 689 -888 695 888
rect 649 -900 695 -888
rect 726 -904 736 904
rect 800 -904 810 904
rect 841 888 887 900
rect 841 -888 847 888
rect 881 -888 887 888
rect 841 -900 887 -888
rect 918 -904 928 904
rect 988 -904 998 904
<< via1 >>
rect -910 985 924 1001
rect -910 949 924 985
rect -992 888 -928 904
rect -992 -888 -977 888
rect -977 -888 -943 888
rect -943 -888 -928 888
rect -992 -904 -928 -888
rect -800 888 -736 904
rect -800 -888 -785 888
rect -785 -888 -751 888
rect -751 -888 -736 888
rect -800 -904 -736 -888
rect -608 888 -544 904
rect -608 -888 -593 888
rect -593 -888 -559 888
rect -559 -888 -544 888
rect -608 -904 -544 -888
rect -416 888 -352 904
rect -416 -888 -401 888
rect -401 -888 -367 888
rect -367 -888 -352 888
rect -416 -904 -352 -888
rect -224 888 -160 904
rect -224 -888 -209 888
rect -209 -888 -175 888
rect -175 -888 -160 888
rect -224 -904 -160 -888
rect -32 888 32 904
rect -32 -888 -17 888
rect -17 -888 17 888
rect 17 -888 32 888
rect -32 -904 32 -888
rect 160 888 224 904
rect 160 -888 175 888
rect 175 -888 209 888
rect 209 -888 224 888
rect 160 -904 224 -888
rect 352 888 416 904
rect 352 -888 367 888
rect 367 -888 401 888
rect 401 -888 416 888
rect 352 -904 416 -888
rect 544 888 608 904
rect 544 -888 559 888
rect 559 -888 593 888
rect 593 -888 608 888
rect 544 -904 608 -888
rect 736 888 800 904
rect 736 -888 751 888
rect 751 -888 785 888
rect 785 -888 800 888
rect 736 -904 800 -888
rect 928 888 988 904
rect 928 -888 943 888
rect 943 -888 977 888
rect 977 -888 988 888
rect 928 -904 988 -888
<< metal2 >>
rect -910 1001 924 1011
rect -992 949 -910 1000
rect 924 949 988 1000
rect -992 928 988 949
rect -992 904 -928 928
rect -992 -914 -928 -904
rect -800 904 -736 928
rect -800 -914 -736 -904
rect -608 904 -544 928
rect -608 -914 -544 -904
rect -416 904 -352 928
rect -416 -914 -352 -904
rect -224 904 -160 928
rect -224 -914 -160 -904
rect -32 904 32 928
rect -32 -914 32 -904
rect 160 904 224 928
rect 160 -914 224 -904
rect 352 904 416 928
rect 352 -914 416 -904
rect 544 904 608 928
rect 544 -914 608 -904
rect 736 904 800 928
rect 736 -914 800 -904
rect 928 904 988 928
rect 928 -914 988 -904
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -1057 1074 1057
string parameters w 9 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
