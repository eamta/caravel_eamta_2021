magic
tech sky130A
magscale 1 2
timestamp 1624338677
<< pwell >>
rect -211 -290 211 290
<< nmos >>
rect -15 -142 15 80
<< ndiff >>
rect -73 68 -15 80
rect -73 -130 -61 68
rect -27 -130 -15 68
rect -73 -142 -15 -130
rect 15 68 73 80
rect 15 -130 27 68
rect 61 -130 73 68
rect 15 -142 73 -130
<< ndiffc >>
rect -61 -130 -27 68
rect 27 -130 61 68
<< psubdiff >>
rect -175 220 175 254
rect -175 158 -141 220
rect 141 158 175 220
rect -175 -220 -141 -158
rect 141 -220 175 -158
rect -175 -254 -79 -220
rect 79 -254 175 -220
<< psubdiffcont >>
rect -175 -158 -141 158
rect 141 -158 175 158
rect -79 -254 79 -220
<< poly >>
rect -33 152 33 168
rect -33 118 -17 152
rect 17 118 33 152
rect -33 102 33 118
rect -15 80 15 102
rect -15 -168 15 -142
<< polycont >>
rect -17 118 17 152
<< locali >>
rect -175 220 175 254
rect -175 158 -141 220
rect 141 158 175 220
rect -33 118 -17 152
rect 17 118 33 152
rect -61 68 -27 84
rect -61 -146 -27 -130
rect 27 68 61 84
rect 27 -146 61 -130
rect -175 -220 -141 -158
rect 141 -220 175 -158
rect -175 -254 -79 -220
rect 79 -254 175 -220
<< viali >>
rect -17 118 17 152
rect -61 -130 -27 68
rect 27 -130 61 68
<< metal1 >>
rect -33 152 33 162
rect -33 118 -17 152
rect 17 118 33 152
rect -33 108 33 118
rect -67 68 -21 80
rect -67 -130 -61 68
rect -27 -130 -21 68
rect -67 -142 -21 -130
rect 21 68 67 80
rect 21 -130 27 68
rect 61 -130 67 68
rect 21 -142 67 -130
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -237 158 237
string parameters w 1.11 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
