magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect 667 1042 702 1076
rect 129 919 187 925
rect 129 885 141 919
rect 129 879 187 885
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1042
rect 668 1023 702 1042
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 687 530 702 1023
rect 721 989 756 1023
rect 721 530 755 989
rect 867 921 925 927
rect 867 887 879 921
rect 1037 898 1071 916
rect 867 881 925 887
rect 1037 862 1107 898
rect 1054 828 1125 862
rect 1405 828 1440 862
rect 1828 845 1863 863
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 721 496 736 530
rect 1054 477 1124 828
rect 1406 809 1440 828
rect 1792 830 1863 845
rect 2143 830 2178 864
rect 1236 760 1294 766
rect 1236 726 1248 760
rect 1236 720 1294 726
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1425 424 1440 809
rect 1459 775 1494 809
rect 1459 424 1493 775
rect 1605 707 1663 713
rect 1605 673 1617 707
rect 1605 667 1663 673
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 830
rect 2144 811 2178 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2163 318 2178 811
rect 2197 777 2232 811
rect 2197 318 2231 777
rect 3988 745 4023 779
rect 3989 726 4023 745
rect 2343 709 2401 715
rect 2343 675 2355 709
rect 2513 686 2547 704
rect 2935 686 2970 704
rect 2343 669 2401 675
rect 2513 650 2583 686
rect 2899 671 2970 686
rect 3819 677 3877 683
rect 2530 616 2601 650
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2530 265 2600 616
rect 2712 548 2770 554
rect 2712 514 2724 548
rect 2712 508 2770 514
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
rect 2899 212 2969 671
rect 3819 643 3831 677
rect 3819 637 3877 643
rect 3081 603 3139 609
rect 3081 569 3093 603
rect 3251 580 3285 598
rect 3673 580 3707 598
rect 3081 563 3139 569
rect 3251 544 3321 580
rect 3268 510 3339 544
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2899 176 2952 212
rect 3268 159 3338 510
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3268 123 3321 159
rect 3637 106 3707 580
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3637 70 3690 106
rect 4008 53 4023 726
rect 4042 692 4077 726
rect 4042 53 4076 692
rect 4188 624 4246 630
rect 4188 590 4200 624
rect 4188 584 4246 590
rect 5095 586 5130 620
rect 5096 567 5130 586
rect 4926 518 4984 524
rect 4926 484 4938 518
rect 4926 478 4984 484
rect 4358 421 4392 439
rect 4780 421 4814 439
rect 4358 385 4428 421
rect 4375 351 4446 385
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
rect 4375 0 4445 351
rect 4557 283 4615 289
rect 4557 249 4569 283
rect 4557 243 4615 249
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4375 -36 4428 0
rect 4744 -53 4814 421
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4744 -89 4797 -53
rect 5115 -106 5130 567
rect 5149 533 5184 567
rect 5149 -106 5183 533
rect 5295 465 5353 471
rect 5295 431 5307 465
rect 5295 425 5353 431
rect 5465 262 5499 280
rect 5465 226 5535 262
rect 5482 192 5553 226
rect 5833 192 5868 226
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5149 -140 5164 -106
rect 5482 -159 5552 192
rect 5834 173 5868 192
rect 5664 124 5722 130
rect 5664 90 5676 124
rect 5664 84 5722 90
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5482 -195 5535 -159
rect 5853 -212 5868 173
rect 5887 139 5922 173
rect 6202 139 6237 173
rect 6625 156 6660 174
rect 5887 -212 5921 139
rect 6203 120 6237 139
rect 6589 141 6660 156
rect 6033 71 6091 77
rect 6033 37 6045 71
rect 6033 31 6091 37
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5887 -246 5902 -212
rect 6222 -265 6237 120
rect 6256 86 6291 120
rect 6256 -265 6290 86
rect 6402 18 6460 24
rect 6402 -16 6414 18
rect 6402 -22 6460 -16
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6256 -299 6271 -265
rect 6589 -318 6659 141
rect 6771 73 6829 79
rect 6771 39 6783 73
rect 6941 50 6975 68
rect 6771 33 6829 39
rect 6941 14 7011 50
rect 6958 -20 7029 14
rect 7309 -20 7344 14
rect 7732 -3 7767 15
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6589 -354 6642 -318
rect 6958 -371 7028 -20
rect 7310 -39 7344 -20
rect 7696 -18 7767 -3
rect 7140 -88 7198 -82
rect 7140 -122 7152 -88
rect 7140 -128 7198 -122
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6958 -407 7011 -371
rect 7329 -424 7344 -39
rect 7363 -73 7398 -39
rect 7363 -424 7397 -73
rect 7509 -141 7567 -135
rect 7509 -175 7521 -141
rect 7509 -181 7567 -175
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7363 -458 7378 -424
rect 7696 -477 7766 -18
rect 7878 -86 7936 -80
rect 7878 -120 7890 -86
rect 7878 -126 7936 -120
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7696 -513 7749 -477
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use sky130_fd_pr__pfet_01v8_XSLFBL  XM11
timestamp 1624053917
transform 1 0 2372 0 1 538
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM10
timestamp 1624053917
transform 1 0 2741 0 1 431
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 3110 0 1 432
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM13
timestamp 1624053917
transform 1 0 3848 0 1 416
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM6
timestamp 1624053917
transform 1 0 5324 0 1 204
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM7
timestamp 1624053917
transform 1 0 4955 0 1 257
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM8
timestamp 1624053917
transform 1 0 4586 0 1 166
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM12
timestamp 1624053917
transform 1 0 4217 0 1 363
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XSLFBL  XM19
timestamp 1624053917
transform 1 0 6800 0 1 -98
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM15
timestamp 1624053917
transform 1 0 6431 0 1 -99
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM14
timestamp 1624053917
transform 1 0 6062 0 1 -46
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 5693 0 1 7
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM16
timestamp 1624053917
transform 1 0 7907 0 1 -257
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM17
timestamp 1624053917
transform 1 0 7538 0 1 -258
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM18
timestamp 1624053917
transform 1 0 7169 0 1 -205
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM21
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM20
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM0
timestamp 1624053917
transform 1 0 1265 0 1 643
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM3
timestamp 1624053917
transform 1 0 1634 0 1 590
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Q
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 D
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 CLR
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 CLK
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Qb
port 7 nsew
<< end >>
