magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 1608 1456 1766 1515
rect 1546 1455 1828 1456
rect 1546 1421 1828 1422
rect 1670 1353 1704 1387
rect 129 1291 187 1297
rect 129 1257 141 1291
rect 129 1251 187 1257
rect 867 1185 925 1191
rect 299 1136 333 1154
rect 721 1136 755 1154
rect 867 1151 879 1185
rect 867 1145 925 1151
rect 299 1100 369 1136
rect 316 1066 387 1100
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 625 386 1066
rect 498 998 556 1004
rect 498 964 510 998
rect 498 958 556 964
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect -17 617 17 625
rect 299 617 386 625
rect -17 607 386 617
rect 685 607 755 1136
rect 1037 1030 1071 1048
rect 1037 994 1107 1030
rect 1054 960 1125 994
rect 1512 989 1546 999
rect 1828 989 1862 999
rect 1512 981 1862 989
rect -17 583 755 607
rect 867 613 925 619
rect 867 605 879 613
rect 316 571 755 583
rect 863 579 929 605
rect 867 573 925 579
rect -17 549 738 571
rect 829 565 963 571
rect -343 484 -185 543
rect 316 537 738 549
rect 755 545 963 565
rect 755 537 929 545
rect 316 530 755 537
rect 316 507 738 530
rect 755 509 929 511
rect 755 507 975 509
rect 316 503 975 507
rect 316 494 857 503
rect -405 483 -123 484
rect 721 477 857 494
rect 895 477 975 503
rect 1054 477 1124 960
rect 1476 919 1898 981
rect 1236 892 1294 898
rect 1236 858 1248 892
rect 1236 852 1294 858
rect 1638 629 1658 637
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect -405 449 -123 450
rect 687 443 715 469
rect 757 443 823 469
rect 1054 441 1107 477
rect -281 381 -247 415
rect -439 17 -405 27
rect -123 17 -89 27
rect -439 9 -89 17
rect -475 -53 -53 9
rect 193 -305 200 -200
rect 221 -277 228 -213
rect -313 -343 -293 -335
<< nwell >>
rect -475 579 -53 607
<< pwell >>
rect -53 -584 -1 -53
rect -475 -633 -1 -584
rect 421 -633 525 -53
rect 947 -633 999 -53
<< poly >>
rect 123 419 297 485
rect 649 423 823 489
<< metal1 >>
rect 138 425 148 477
rect 268 425 278 477
rect 388 441 823 493
rect 171 200 181 242
rect 0 178 181 200
rect 239 178 249 242
rect 0 129 200 178
rect 283 129 329 166
rect 0 86 329 129
rect 0 0 200 86
rect 143 -200 189 0
rect 0 -400 200 -200
rect 221 -277 231 -213
rect 289 -277 299 -213
rect 388 -453 440 441
rect 649 423 823 441
rect 697 178 707 242
rect 765 178 775 242
rect 620 170 663 178
rect 617 129 663 170
rect 809 129 855 166
rect 617 86 855 129
rect 669 -204 715 86
rect 747 -277 757 -213
rect 815 -277 825 -213
rect 167 -505 177 -453
rect 236 -505 440 -453
rect 693 -504 703 -452
rect 762 -504 772 -452
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
<< via1 >>
rect 148 425 268 477
rect 181 178 239 242
rect 231 -277 289 -213
rect 707 178 765 242
rect 757 -277 815 -213
rect 177 -505 236 -453
rect 703 -504 762 -452
<< metal2 >>
rect 148 477 268 487
rect -76 425 148 477
rect 268 425 522 477
rect -76 116 -24 425
rect 148 415 268 425
rect 181 242 239 252
rect 181 168 239 178
rect -294 64 -24 116
rect 187 129 233 168
rect 187 83 288 129
rect -294 -27 -242 64
rect -345 -79 -242 -27
rect -105 -79 7 -27
rect -45 -453 7 -79
rect 242 -73 288 83
rect 242 -83 303 -73
rect 242 -165 303 -155
rect 242 -203 288 -165
rect 231 -213 289 -203
rect 231 -287 289 -277
rect 177 -453 236 -443
rect -45 -505 177 -453
rect 470 -450 522 425
rect 707 242 765 252
rect 707 168 765 178
rect 713 129 759 168
rect 713 83 814 129
rect 768 -73 814 83
rect 768 -83 829 -73
rect 768 -165 829 -155
rect 768 -203 814 -165
rect 757 -213 815 -203
rect 757 -287 815 -277
rect 703 -450 762 -442
rect 470 -452 762 -450
rect 470 -502 703 -452
rect 177 -515 236 -505
rect 703 -514 762 -504
<< via2 >>
rect 242 -155 303 -83
rect 768 -155 829 -83
<< metal3 >>
rect 232 -83 313 -78
rect 758 -83 839 -78
rect 232 -155 242 -83
rect 303 -155 768 -83
rect 829 -155 839 -83
rect 232 -160 313 -155
rect 758 -160 839 -155
use sky130_fd_pr__nfet_01v8_HAN8QX  sky130_fd_pr__nfet_01v8_HAN8QX_0
timestamp 1623900471
transform 1 0 210 0 -1 -343
box -211 -290 211 290
use sky130_fd_pr__pfet_01v8_XA7ZMQ  sky130_fd_pr__pfet_01v8_XA7ZMQ_0
timestamp 1623900471
transform 1 0 210 0 1 277
box -263 -330 263 330
use sky130_fd_pr__pfet_01v8_M4ZJ2X  XM5
timestamp 1624053917
transform 1 0 158 0 1 988
box -211 -441 211 441
use sky130_fd_pr__pfet_01v8_XA7ZMQ  sky130_fd_pr__pfet_01v8_XA7ZMQ_1
timestamp 1623900471
transform 1 0 736 0 1 277
box -263 -330 263 330
use sky130_fd_pr__nfet_01v8_HAN8QX  sky130_fd_pr__nfet_01v8_HAN8QX_1
timestamp 1623900471
transform 1 0 736 0 -1 -343
box -211 -290 211 290
use sky130_fd_pr__nfet_01v8_HZDS64  XM6
timestamp 1624053917
transform 1 0 527 0 1 815
box -211 -321 211 321
use sky130_fd_pr__pfet_01v8_M4ZJ2X  XM2
timestamp 1624053917
transform 1 0 896 0 1 882
box -211 -441 211 441
use sky130_fd_pr__nfet_01v8_HZDS64  XM7
timestamp 1624053917
transform 1 0 1265 0 1 709
box -211 -321 211 321
use inverter_min  inverter_min_0
timestamp 1624053917
transform 1 0 -422 0 1 -600
box -53 -1600 369 1179
use inverter_min  x1
timestamp 1624053917
transform 1 0 1529 0 1 372
box -53 -1600 369 1179
<< labels >>
rlabel metal2 -332 -64 -311 -46 1 sel
rlabel metal2 -94 -63 -73 -45 1 sel_b
rlabel metal1 152 -61 173 -43 1 DinA
rlabel metal1 681 -62 702 -44 1 DinB
rlabel via2 786 -132 807 -114 1 out
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd1p8
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 sel
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 avss1p8
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 DinB
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 out
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 DinA
port 6 nsew
<< end >>
