magic
tech sky130A
magscale 1 2
timestamp 1624338677
<< metal1 >>
rect -54 2372 10324 2463
rect -54 2280 -44 2372
rect 28 2326 10324 2372
rect 28 2280 38 2326
rect 9123 2320 10324 2326
rect -54 2186 4 2280
rect 547 1684 557 1756
rect 618 1684 628 1756
rect 1073 1684 1083 1756
rect 1144 1684 1154 1756
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 3495 1684 3505 1756
rect 3566 1684 3576 1756
rect 4021 1684 4031 1756
rect 4092 1684 4102 1756
rect 4969 1684 4979 1756
rect 5040 1684 5050 1756
rect 5495 1684 5505 1756
rect 5566 1684 5576 1756
rect 6443 1684 6453 1756
rect 6514 1684 6524 1756
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 7917 1684 7927 1756
rect 7988 1684 7998 1756
rect 8443 1684 8453 1756
rect 8514 1684 8524 1756
rect 9391 1684 9401 1756
rect 9462 1684 9472 1756
rect 9917 1684 9927 1756
rect 9988 1684 9998 1756
rect 328 1218 9266 1224
rect 0 1136 9266 1218
rect 328 1130 9266 1136
<< via1 >>
rect -44 2280 28 2372
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
<< metal2 >>
rect 62 2537 1547 2538
rect 62 2486 5975 2537
rect -44 2372 28 2382
rect -44 2270 28 2280
rect 15 1812 23 1838
rect 62 1826 114 2486
rect 1495 2485 5975 2486
rect 62 1812 79 1826
rect 1495 1811 1547 2485
rect 2972 2330 3043 2340
rect 2972 2246 3043 2256
rect 2981 1839 3033 2246
rect 2973 1813 3033 1839
rect 4451 1837 4503 2485
rect 2981 1812 3033 1813
rect 4436 1814 4503 1837
rect 5923 1817 5975 2485
rect 7396 2514 7467 2524
rect 7396 2420 7467 2430
rect 7404 1836 7456 2420
rect 4436 1811 4461 1814
rect 5923 1811 5948 1817
rect 7388 1813 7456 1836
rect 7388 1810 7413 1813
rect 8879 1810 8931 2443
rect 557 1756 618 1766
rect 557 1674 618 1684
rect 1083 1756 1144 1766
rect 1083 1674 1144 1684
rect 2031 1756 2092 1766
rect 2031 1674 2092 1684
rect 2557 1756 2618 1766
rect 2557 1674 2618 1684
rect 3505 1756 3566 1766
rect 3505 1674 3566 1684
rect 4031 1756 4092 1766
rect 4031 1674 4092 1684
rect 4979 1756 5040 1766
rect 4979 1674 5040 1684
rect 5505 1756 5566 1766
rect 5505 1674 5566 1684
rect 6453 1756 6514 1766
rect 6453 1674 6514 1684
rect 6979 1756 7040 1766
rect 6979 1674 7040 1684
rect 7927 1756 7988 1766
rect 7927 1674 7988 1684
rect 8453 1756 8514 1766
rect 8453 1674 8514 1684
rect 9401 1756 9462 1766
rect 9401 1674 9462 1684
rect 9927 1756 9988 1766
rect 9927 1674 9988 1684
<< via2 >>
rect 2972 2256 3043 2330
rect 7396 2430 7467 2514
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
<< metal3 >>
rect 2981 2514 7477 2553
rect 2981 2493 7396 2514
rect 2981 2335 3041 2493
rect 7386 2430 7396 2493
rect 7467 2430 7477 2514
rect 7386 2425 7477 2430
rect 2962 2330 3053 2335
rect 2962 2256 2972 2330
rect 3043 2256 3053 2330
rect 2962 2251 3053 2256
rect 4497 2265 7957 2337
rect 1632 2014 3218 2086
rect 1632 1925 1704 2014
rect 1171 1853 1704 1925
rect 2753 1859 2903 1919
rect 2782 1848 2903 1859
rect 525 1756 628 1761
rect 525 1684 557 1756
rect 618 1684 628 1756
rect 525 1679 628 1684
rect 1054 1756 1154 1761
rect 1054 1684 1083 1756
rect 1144 1684 1154 1756
rect 1054 1679 1154 1684
rect 2021 1756 2102 1761
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2021 1679 2102 1684
rect 2547 1756 2628 1761
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 2547 1679 2628 1684
rect 525 1183 585 1679
rect 1054 1173 1114 1679
rect 2031 1072 2091 1679
rect 2564 1072 2624 1679
rect 2843 1536 2903 1848
rect 3146 1769 3218 2014
rect 4497 1925 4569 2265
rect 6173 2039 7718 2111
rect 6173 1925 6245 2039
rect 4119 1853 4569 1925
rect 5593 1853 6245 1925
rect 7067 1853 7366 1925
rect 3146 1761 3560 1769
rect 3146 1756 3576 1761
rect 3146 1697 3505 1756
rect 3495 1684 3505 1697
rect 3566 1684 3576 1756
rect 4021 1756 4102 1761
rect 4021 1734 4031 1756
rect 3495 1679 3576 1684
rect 4020 1684 4031 1734
rect 4092 1684 4102 1756
rect 4020 1679 4102 1684
rect 4969 1756 5050 1761
rect 4969 1684 4979 1756
rect 5040 1748 5050 1756
rect 5495 1756 5576 1761
rect 5040 1684 5060 1748
rect 4969 1679 5060 1684
rect 5495 1684 5505 1756
rect 5566 1743 5576 1756
rect 6443 1756 6524 1761
rect 5566 1684 5585 1743
rect 5495 1679 5585 1684
rect 6443 1684 6453 1756
rect 6514 1734 6524 1756
rect 6969 1756 7050 1761
rect 6514 1684 6525 1734
rect 6443 1679 6525 1684
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 6969 1679 7050 1684
rect 4020 1536 4080 1679
rect 2843 1476 4080 1536
rect 5000 1072 5060 1679
rect 5525 1072 5585 1679
rect 6465 1150 6525 1679
rect 6980 1335 7040 1679
rect 7294 1574 7366 1853
rect 7646 1774 7718 2039
rect 7885 2090 7957 2265
rect 7885 2018 9156 2090
rect 8541 1853 8845 1925
rect 7646 1761 7996 1774
rect 7646 1756 7998 1761
rect 7646 1702 7927 1756
rect 7917 1684 7927 1702
rect 7988 1684 7998 1756
rect 8443 1756 8524 1761
rect 8443 1742 8453 1756
rect 7917 1679 7998 1684
rect 8438 1684 8453 1742
rect 8514 1684 8524 1756
rect 8438 1679 8524 1684
rect 8438 1574 8510 1679
rect 7294 1502 8510 1574
rect 8773 1554 8845 1853
rect 9084 1769 9156 2018
rect 10087 1853 10148 1925
rect 9084 1761 9446 1769
rect 9084 1756 9472 1761
rect 9084 1697 9401 1756
rect 9391 1684 9401 1697
rect 9462 1684 9472 1756
rect 9917 1756 9998 1761
rect 9917 1748 9927 1756
rect 9391 1679 9472 1684
rect 9902 1684 9927 1748
rect 9988 1684 9998 1756
rect 9902 1679 9998 1684
rect 9902 1554 9974 1679
rect 8773 1482 9974 1554
use mux_2to1_logic  mux_2to1_logic_1
timestamp 1624338677
transform 1 0 1949 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_0
timestamp 1624338677
transform 1 0 475 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_2
timestamp 1624338677
transform 1 0 3423 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_3
timestamp 1624338677
transform 1 0 4897 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_4
timestamp 1624338677
transform 1 0 6371 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_5
timestamp 1624338677
transform 1 0 7845 0 -1 1770
box -475 -633 999 607
use mux_2to1_logic  mux_2to1_logic_6
timestamp 1624338677
transform 1 0 9319 0 -1 1770
box -475 -633 999 607
<< labels >>
rlabel metal2 8893 2121 8918 2147 1 reg0
rlabel metal3 6059 2508 6084 2534 1 reg1
rlabel metal2 80 2501 105 2527 1 reg2
rlabel metal3 10087 1853 10148 1925 1 out_mux
rlabel metal3 6980 1335 7040 1684 1 mux_i7
rlabel metal3 6465 1150 6525 1684 1 mux_i6
rlabel metal3 5525 1072 5585 1684 1 mux_i5
rlabel metal3 5000 1072 5060 1684 1 mux_i4
rlabel metal3 1054 1173 1114 1684 1 mux_i1
rlabel metal3 2564 1072 2624 1684 1 mux_i3
rlabel metal3 2031 1072 2091 1684 1 mux_i2
rlabel metal1 28 2326 10324 2463 1 avss1p8
rlabel metal1 0 1136 9266 1218 1 avdd1p8
rlabel metal3 525 1183 585 1684 1 mux_i0
<< end >>
