magic
tech sky130A
magscale 1 2
timestamp 1615997521
<< nwell >>
rect -3517 -884 3517 884
<< pmoslvt >>
rect -3321 -736 -3111 664
rect -3053 -736 -2843 664
rect -2785 -736 -2575 664
rect -2517 -736 -2307 664
rect -2249 -736 -2039 664
rect -1981 -736 -1771 664
rect -1713 -736 -1503 664
rect -1445 -736 -1235 664
rect -1177 -736 -967 664
rect -909 -736 -699 664
rect -641 -736 -431 664
rect -373 -736 -163 664
rect -105 -736 105 664
rect 163 -736 373 664
rect 431 -736 641 664
rect 699 -736 909 664
rect 967 -736 1177 664
rect 1235 -736 1445 664
rect 1503 -736 1713 664
rect 1771 -736 1981 664
rect 2039 -736 2249 664
rect 2307 -736 2517 664
rect 2575 -736 2785 664
rect 2843 -736 3053 664
rect 3111 -736 3321 664
<< pdiff >>
rect -3379 652 -3321 664
rect -3379 -724 -3367 652
rect -3333 -724 -3321 652
rect -3379 -736 -3321 -724
rect -3111 652 -3053 664
rect -3111 -724 -3099 652
rect -3065 -724 -3053 652
rect -3111 -736 -3053 -724
rect -2843 652 -2785 664
rect -2843 -724 -2831 652
rect -2797 -724 -2785 652
rect -2843 -736 -2785 -724
rect -2575 652 -2517 664
rect -2575 -724 -2563 652
rect -2529 -724 -2517 652
rect -2575 -736 -2517 -724
rect -2307 652 -2249 664
rect -2307 -724 -2295 652
rect -2261 -724 -2249 652
rect -2307 -736 -2249 -724
rect -2039 652 -1981 664
rect -2039 -724 -2027 652
rect -1993 -724 -1981 652
rect -2039 -736 -1981 -724
rect -1771 652 -1713 664
rect -1771 -724 -1759 652
rect -1725 -724 -1713 652
rect -1771 -736 -1713 -724
rect -1503 652 -1445 664
rect -1503 -724 -1491 652
rect -1457 -724 -1445 652
rect -1503 -736 -1445 -724
rect -1235 652 -1177 664
rect -1235 -724 -1223 652
rect -1189 -724 -1177 652
rect -1235 -736 -1177 -724
rect -967 652 -909 664
rect -967 -724 -955 652
rect -921 -724 -909 652
rect -967 -736 -909 -724
rect -699 652 -641 664
rect -699 -724 -687 652
rect -653 -724 -641 652
rect -699 -736 -641 -724
rect -431 652 -373 664
rect -431 -724 -419 652
rect -385 -724 -373 652
rect -431 -736 -373 -724
rect -163 652 -105 664
rect -163 -724 -151 652
rect -117 -724 -105 652
rect -163 -736 -105 -724
rect 105 652 163 664
rect 105 -724 117 652
rect 151 -724 163 652
rect 105 -736 163 -724
rect 373 652 431 664
rect 373 -724 385 652
rect 419 -724 431 652
rect 373 -736 431 -724
rect 641 652 699 664
rect 641 -724 653 652
rect 687 -724 699 652
rect 641 -736 699 -724
rect 909 652 967 664
rect 909 -724 921 652
rect 955 -724 967 652
rect 909 -736 967 -724
rect 1177 652 1235 664
rect 1177 -724 1189 652
rect 1223 -724 1235 652
rect 1177 -736 1235 -724
rect 1445 652 1503 664
rect 1445 -724 1457 652
rect 1491 -724 1503 652
rect 1445 -736 1503 -724
rect 1713 652 1771 664
rect 1713 -724 1725 652
rect 1759 -724 1771 652
rect 1713 -736 1771 -724
rect 1981 652 2039 664
rect 1981 -724 1993 652
rect 2027 -724 2039 652
rect 1981 -736 2039 -724
rect 2249 652 2307 664
rect 2249 -724 2261 652
rect 2295 -724 2307 652
rect 2249 -736 2307 -724
rect 2517 652 2575 664
rect 2517 -724 2529 652
rect 2563 -724 2575 652
rect 2517 -736 2575 -724
rect 2785 652 2843 664
rect 2785 -724 2797 652
rect 2831 -724 2843 652
rect 2785 -736 2843 -724
rect 3053 652 3111 664
rect 3053 -724 3065 652
rect 3099 -724 3111 652
rect 3053 -736 3111 -724
rect 3321 652 3379 664
rect 3321 -724 3333 652
rect 3367 -724 3379 652
rect 3321 -736 3379 -724
<< pdiffc >>
rect -3367 -724 -3333 652
rect -3099 -724 -3065 652
rect -2831 -724 -2797 652
rect -2563 -724 -2529 652
rect -2295 -724 -2261 652
rect -2027 -724 -1993 652
rect -1759 -724 -1725 652
rect -1491 -724 -1457 652
rect -1223 -724 -1189 652
rect -955 -724 -921 652
rect -687 -724 -653 652
rect -419 -724 -385 652
rect -151 -724 -117 652
rect 117 -724 151 652
rect 385 -724 419 652
rect 653 -724 687 652
rect 921 -724 955 652
rect 1189 -724 1223 652
rect 1457 -724 1491 652
rect 1725 -724 1759 652
rect 1993 -724 2027 652
rect 2261 -724 2295 652
rect 2529 -724 2563 652
rect 2797 -724 2831 652
rect 3065 -724 3099 652
rect 3333 -724 3367 652
<< nsubdiff >>
rect -3481 814 -3385 848
rect 3385 814 3481 848
rect -3481 751 -3447 814
rect 3447 751 3481 814
rect -3481 -814 -3447 -751
rect 3447 -814 3481 -751
rect -3481 -848 -3385 -814
rect 3385 -848 3481 -814
<< nsubdiffcont >>
rect -3385 814 3385 848
rect -3481 -751 -3447 751
rect 3447 -751 3481 751
rect -3385 -848 3385 -814
<< poly >>
rect -3321 745 -3111 761
rect -3321 711 -3305 745
rect -3127 711 -3111 745
rect -3321 664 -3111 711
rect -3053 745 -2843 761
rect -3053 711 -3037 745
rect -2859 711 -2843 745
rect -3053 664 -2843 711
rect -2785 745 -2575 761
rect -2785 711 -2769 745
rect -2591 711 -2575 745
rect -2785 664 -2575 711
rect -2517 745 -2307 761
rect -2517 711 -2501 745
rect -2323 711 -2307 745
rect -2517 664 -2307 711
rect -2249 745 -2039 761
rect -2249 711 -2233 745
rect -2055 711 -2039 745
rect -2249 664 -2039 711
rect -1981 745 -1771 761
rect -1981 711 -1965 745
rect -1787 711 -1771 745
rect -1981 664 -1771 711
rect -1713 745 -1503 761
rect -1713 711 -1697 745
rect -1519 711 -1503 745
rect -1713 664 -1503 711
rect -1445 745 -1235 761
rect -1445 711 -1429 745
rect -1251 711 -1235 745
rect -1445 664 -1235 711
rect -1177 745 -967 761
rect -1177 711 -1161 745
rect -983 711 -967 745
rect -1177 664 -967 711
rect -909 745 -699 761
rect -909 711 -893 745
rect -715 711 -699 745
rect -909 664 -699 711
rect -641 745 -431 761
rect -641 711 -625 745
rect -447 711 -431 745
rect -641 664 -431 711
rect -373 745 -163 761
rect -373 711 -357 745
rect -179 711 -163 745
rect -373 664 -163 711
rect -105 745 105 761
rect -105 711 -89 745
rect 89 711 105 745
rect -105 664 105 711
rect 163 745 373 761
rect 163 711 179 745
rect 357 711 373 745
rect 163 664 373 711
rect 431 745 641 761
rect 431 711 447 745
rect 625 711 641 745
rect 431 664 641 711
rect 699 745 909 761
rect 699 711 715 745
rect 893 711 909 745
rect 699 664 909 711
rect 967 745 1177 761
rect 967 711 983 745
rect 1161 711 1177 745
rect 967 664 1177 711
rect 1235 745 1445 761
rect 1235 711 1251 745
rect 1429 711 1445 745
rect 1235 664 1445 711
rect 1503 745 1713 761
rect 1503 711 1519 745
rect 1697 711 1713 745
rect 1503 664 1713 711
rect 1771 745 1981 761
rect 1771 711 1787 745
rect 1965 711 1981 745
rect 1771 664 1981 711
rect 2039 745 2249 761
rect 2039 711 2055 745
rect 2233 711 2249 745
rect 2039 664 2249 711
rect 2307 745 2517 761
rect 2307 711 2323 745
rect 2501 711 2517 745
rect 2307 664 2517 711
rect 2575 745 2785 761
rect 2575 711 2591 745
rect 2769 711 2785 745
rect 2575 664 2785 711
rect 2843 745 3053 761
rect 2843 711 2859 745
rect 3037 711 3053 745
rect 2843 664 3053 711
rect 3111 745 3321 761
rect 3111 711 3127 745
rect 3305 711 3321 745
rect 3111 664 3321 711
rect -3321 -762 -3111 -736
rect -3053 -762 -2843 -736
rect -2785 -762 -2575 -736
rect -2517 -762 -2307 -736
rect -2249 -762 -2039 -736
rect -1981 -762 -1771 -736
rect -1713 -762 -1503 -736
rect -1445 -762 -1235 -736
rect -1177 -762 -967 -736
rect -909 -762 -699 -736
rect -641 -762 -431 -736
rect -373 -762 -163 -736
rect -105 -762 105 -736
rect 163 -762 373 -736
rect 431 -762 641 -736
rect 699 -762 909 -736
rect 967 -762 1177 -736
rect 1235 -762 1445 -736
rect 1503 -762 1713 -736
rect 1771 -762 1981 -736
rect 2039 -762 2249 -736
rect 2307 -762 2517 -736
rect 2575 -762 2785 -736
rect 2843 -762 3053 -736
rect 3111 -762 3321 -736
<< polycont >>
rect -3305 711 -3127 745
rect -3037 711 -2859 745
rect -2769 711 -2591 745
rect -2501 711 -2323 745
rect -2233 711 -2055 745
rect -1965 711 -1787 745
rect -1697 711 -1519 745
rect -1429 711 -1251 745
rect -1161 711 -983 745
rect -893 711 -715 745
rect -625 711 -447 745
rect -357 711 -179 745
rect -89 711 89 745
rect 179 711 357 745
rect 447 711 625 745
rect 715 711 893 745
rect 983 711 1161 745
rect 1251 711 1429 745
rect 1519 711 1697 745
rect 1787 711 1965 745
rect 2055 711 2233 745
rect 2323 711 2501 745
rect 2591 711 2769 745
rect 2859 711 3037 745
rect 3127 711 3305 745
<< locali >>
rect -3481 814 -3385 848
rect 3385 814 3481 848
rect -3481 751 -3447 814
rect 3447 751 3481 814
rect -3321 711 -3305 745
rect -3127 711 -3111 745
rect -3053 711 -3037 745
rect -2859 711 -2843 745
rect -2785 711 -2769 745
rect -2591 711 -2575 745
rect -2517 711 -2501 745
rect -2323 711 -2307 745
rect -2249 711 -2233 745
rect -2055 711 -2039 745
rect -1981 711 -1965 745
rect -1787 711 -1771 745
rect -1713 711 -1697 745
rect -1519 711 -1503 745
rect -1445 711 -1429 745
rect -1251 711 -1235 745
rect -1177 711 -1161 745
rect -983 711 -967 745
rect -909 711 -893 745
rect -715 711 -699 745
rect -641 711 -625 745
rect -447 711 -431 745
rect -373 711 -357 745
rect -179 711 -163 745
rect -105 711 -89 745
rect 89 711 105 745
rect 163 711 179 745
rect 357 711 373 745
rect 431 711 447 745
rect 625 711 641 745
rect 699 711 715 745
rect 893 711 909 745
rect 967 711 983 745
rect 1161 711 1177 745
rect 1235 711 1251 745
rect 1429 711 1445 745
rect 1503 711 1519 745
rect 1697 711 1713 745
rect 1771 711 1787 745
rect 1965 711 1981 745
rect 2039 711 2055 745
rect 2233 711 2249 745
rect 2307 711 2323 745
rect 2501 711 2517 745
rect 2575 711 2591 745
rect 2769 711 2785 745
rect 2843 711 2859 745
rect 3037 711 3053 745
rect 3111 711 3127 745
rect 3305 711 3321 745
rect -3367 652 -3333 668
rect -3367 -740 -3333 -724
rect -3099 652 -3065 668
rect -3099 -740 -3065 -724
rect -2831 652 -2797 668
rect -2831 -740 -2797 -724
rect -2563 652 -2529 668
rect -2563 -740 -2529 -724
rect -2295 652 -2261 668
rect -2295 -740 -2261 -724
rect -2027 652 -1993 668
rect -2027 -740 -1993 -724
rect -1759 652 -1725 668
rect -1759 -740 -1725 -724
rect -1491 652 -1457 668
rect -1491 -740 -1457 -724
rect -1223 652 -1189 668
rect -1223 -740 -1189 -724
rect -955 652 -921 668
rect -955 -740 -921 -724
rect -687 652 -653 668
rect -687 -740 -653 -724
rect -419 652 -385 668
rect -419 -740 -385 -724
rect -151 652 -117 668
rect -151 -740 -117 -724
rect 117 652 151 668
rect 117 -740 151 -724
rect 385 652 419 668
rect 385 -740 419 -724
rect 653 652 687 668
rect 653 -740 687 -724
rect 921 652 955 668
rect 921 -740 955 -724
rect 1189 652 1223 668
rect 1189 -740 1223 -724
rect 1457 652 1491 668
rect 1457 -740 1491 -724
rect 1725 652 1759 668
rect 1725 -740 1759 -724
rect 1993 652 2027 668
rect 1993 -740 2027 -724
rect 2261 652 2295 668
rect 2261 -740 2295 -724
rect 2529 652 2563 668
rect 2529 -740 2563 -724
rect 2797 652 2831 668
rect 2797 -740 2831 -724
rect 3065 652 3099 668
rect 3065 -740 3099 -724
rect 3333 652 3367 668
rect 3333 -740 3367 -724
rect -3481 -814 -3447 -751
rect 3447 -814 3481 -751
rect -3481 -848 -3385 -814
rect 3385 -848 3481 -814
<< viali >>
rect -3305 711 -3127 745
rect -3037 711 -2859 745
rect -2769 711 -2591 745
rect -2501 711 -2323 745
rect -2233 711 -2055 745
rect -1965 711 -1787 745
rect -1697 711 -1519 745
rect -1429 711 -1251 745
rect -1161 711 -983 745
rect -893 711 -715 745
rect -625 711 -447 745
rect -357 711 -179 745
rect -89 711 89 745
rect 179 711 357 745
rect 447 711 625 745
rect 715 711 893 745
rect 983 711 1161 745
rect 1251 711 1429 745
rect 1519 711 1697 745
rect 1787 711 1965 745
rect 2055 711 2233 745
rect 2323 711 2501 745
rect 2591 711 2769 745
rect 2859 711 3037 745
rect 3127 711 3305 745
rect -3367 -724 -3333 652
rect -3099 -724 -3065 652
rect -2831 -724 -2797 652
rect -2563 -724 -2529 652
rect -2295 -724 -2261 652
rect -2027 -724 -1993 652
rect -1759 -724 -1725 652
rect -1491 -724 -1457 652
rect -1223 -724 -1189 652
rect -955 -724 -921 652
rect -687 -724 -653 652
rect -419 -724 -385 652
rect -151 -724 -117 652
rect 117 -724 151 652
rect 385 -724 419 652
rect 653 -724 687 652
rect 921 -724 955 652
rect 1189 -724 1223 652
rect 1457 -724 1491 652
rect 1725 -724 1759 652
rect 1993 -724 2027 652
rect 2261 -724 2295 652
rect 2529 -724 2563 652
rect 2797 -724 2831 652
rect 3065 -724 3099 652
rect 3333 -724 3367 652
<< metal1 >>
rect -3317 745 -3115 751
rect -3317 711 -3305 745
rect -3127 711 -3115 745
rect -3317 705 -3115 711
rect -3049 745 -2847 751
rect -3049 711 -3037 745
rect -2859 711 -2847 745
rect -3049 705 -2847 711
rect -2781 745 -2579 751
rect -2781 711 -2769 745
rect -2591 711 -2579 745
rect -2781 705 -2579 711
rect -2513 745 -2311 751
rect -2513 711 -2501 745
rect -2323 711 -2311 745
rect -2513 705 -2311 711
rect -2245 745 -2043 751
rect -2245 711 -2233 745
rect -2055 711 -2043 745
rect -2245 705 -2043 711
rect -1977 745 -1775 751
rect -1977 711 -1965 745
rect -1787 711 -1775 745
rect -1977 705 -1775 711
rect -1709 745 -1507 751
rect -1709 711 -1697 745
rect -1519 711 -1507 745
rect -1709 705 -1507 711
rect -1441 745 -1239 751
rect -1441 711 -1429 745
rect -1251 711 -1239 745
rect -1441 705 -1239 711
rect -1173 745 -971 751
rect -1173 711 -1161 745
rect -983 711 -971 745
rect -1173 705 -971 711
rect -905 745 -703 751
rect -905 711 -893 745
rect -715 711 -703 745
rect -905 705 -703 711
rect -637 745 -435 751
rect -637 711 -625 745
rect -447 711 -435 745
rect -637 705 -435 711
rect -369 745 -167 751
rect -369 711 -357 745
rect -179 711 -167 745
rect -369 705 -167 711
rect -101 745 101 751
rect -101 711 -89 745
rect 89 711 101 745
rect -101 705 101 711
rect 167 745 369 751
rect 167 711 179 745
rect 357 711 369 745
rect 167 705 369 711
rect 435 745 637 751
rect 435 711 447 745
rect 625 711 637 745
rect 435 705 637 711
rect 703 745 905 751
rect 703 711 715 745
rect 893 711 905 745
rect 703 705 905 711
rect 971 745 1173 751
rect 971 711 983 745
rect 1161 711 1173 745
rect 971 705 1173 711
rect 1239 745 1441 751
rect 1239 711 1251 745
rect 1429 711 1441 745
rect 1239 705 1441 711
rect 1507 745 1709 751
rect 1507 711 1519 745
rect 1697 711 1709 745
rect 1507 705 1709 711
rect 1775 745 1977 751
rect 1775 711 1787 745
rect 1965 711 1977 745
rect 1775 705 1977 711
rect 2043 745 2245 751
rect 2043 711 2055 745
rect 2233 711 2245 745
rect 2043 705 2245 711
rect 2311 745 2513 751
rect 2311 711 2323 745
rect 2501 711 2513 745
rect 2311 705 2513 711
rect 2579 745 2781 751
rect 2579 711 2591 745
rect 2769 711 2781 745
rect 2579 705 2781 711
rect 2847 745 3049 751
rect 2847 711 2859 745
rect 3037 711 3049 745
rect 2847 705 3049 711
rect 3115 745 3317 751
rect 3115 711 3127 745
rect 3305 711 3317 745
rect 3115 705 3317 711
rect -3373 652 -3327 664
rect -3373 -724 -3367 652
rect -3333 -724 -3327 652
rect -3373 -736 -3327 -724
rect -3105 652 -3059 664
rect -3105 -724 -3099 652
rect -3065 -724 -3059 652
rect -3105 -736 -3059 -724
rect -2837 652 -2791 664
rect -2837 -724 -2831 652
rect -2797 -724 -2791 652
rect -2837 -736 -2791 -724
rect -2569 652 -2523 664
rect -2569 -724 -2563 652
rect -2529 -724 -2523 652
rect -2569 -736 -2523 -724
rect -2301 652 -2255 664
rect -2301 -724 -2295 652
rect -2261 -724 -2255 652
rect -2301 -736 -2255 -724
rect -2033 652 -1987 664
rect -2033 -724 -2027 652
rect -1993 -724 -1987 652
rect -2033 -736 -1987 -724
rect -1765 652 -1719 664
rect -1765 -724 -1759 652
rect -1725 -724 -1719 652
rect -1765 -736 -1719 -724
rect -1497 652 -1451 664
rect -1497 -724 -1491 652
rect -1457 -724 -1451 652
rect -1497 -736 -1451 -724
rect -1229 652 -1183 664
rect -1229 -724 -1223 652
rect -1189 -724 -1183 652
rect -1229 -736 -1183 -724
rect -961 652 -915 664
rect -961 -724 -955 652
rect -921 -724 -915 652
rect -961 -736 -915 -724
rect -693 652 -647 664
rect -693 -724 -687 652
rect -653 -724 -647 652
rect -693 -736 -647 -724
rect -425 652 -379 664
rect -425 -724 -419 652
rect -385 -724 -379 652
rect -425 -736 -379 -724
rect -157 652 -111 664
rect -157 -724 -151 652
rect -117 -724 -111 652
rect -157 -736 -111 -724
rect 111 652 157 664
rect 111 -724 117 652
rect 151 -724 157 652
rect 111 -736 157 -724
rect 379 652 425 664
rect 379 -724 385 652
rect 419 -724 425 652
rect 379 -736 425 -724
rect 647 652 693 664
rect 647 -724 653 652
rect 687 -724 693 652
rect 647 -736 693 -724
rect 915 652 961 664
rect 915 -724 921 652
rect 955 -724 961 652
rect 915 -736 961 -724
rect 1183 652 1229 664
rect 1183 -724 1189 652
rect 1223 -724 1229 652
rect 1183 -736 1229 -724
rect 1451 652 1497 664
rect 1451 -724 1457 652
rect 1491 -724 1497 652
rect 1451 -736 1497 -724
rect 1719 652 1765 664
rect 1719 -724 1725 652
rect 1759 -724 1765 652
rect 1719 -736 1765 -724
rect 1987 652 2033 664
rect 1987 -724 1993 652
rect 2027 -724 2033 652
rect 1987 -736 2033 -724
rect 2255 652 2301 664
rect 2255 -724 2261 652
rect 2295 -724 2301 652
rect 2255 -736 2301 -724
rect 2523 652 2569 664
rect 2523 -724 2529 652
rect 2563 -724 2569 652
rect 2523 -736 2569 -724
rect 2791 652 2837 664
rect 2791 -724 2797 652
rect 2831 -724 2837 652
rect 2791 -736 2837 -724
rect 3059 652 3105 664
rect 3059 -724 3065 652
rect 3099 -724 3105 652
rect 3059 -736 3105 -724
rect 3327 652 3373 664
rect 3327 -724 3333 652
rect 3367 -724 3373 652
rect 3327 -736 3373 -724
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -3464 -831 3464 831
string parameters w 7 l 1.05 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
