magic
tech sky130A
timestamp 1615558595
<< error_p >>
rect 7 -58 8 58
<< nwell >>
rect -54 -76 54 76
<< pmos >>
rect -7 -45 7 45
<< pdiff >>
rect -36 39 -7 45
rect -36 -39 -30 39
rect -13 -39 -7 39
rect -36 -45 -7 -39
rect 7 39 36 45
rect 7 -39 13 39
rect 30 -39 36 39
rect 7 -45 36 -39
<< pdiffc >>
rect -30 -39 -13 39
rect 13 -39 30 39
<< poly >>
rect -7 45 7 58
rect -7 -58 7 -45
<< locali >>
rect -30 39 -13 47
rect -30 -47 -13 -39
rect 13 39 30 47
rect 13 -47 30 -39
<< viali >>
rect -30 -39 -13 39
rect 13 -39 30 39
<< metal1 >>
rect -33 39 -10 45
rect -33 -39 -30 39
rect -13 -39 -10 39
rect -33 -45 -10 -39
rect 10 39 33 45
rect 10 -39 13 39
rect 30 -39 33 39
rect 10 -45 33 -39
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.9 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
