magic
tech sky130A
magscale 1 2
timestamp 1619042825
<< error_p >>
rect -855 -161 -797 -155
rect -737 -161 -679 -155
rect -619 -161 -561 -155
rect -501 -161 -443 -155
rect -383 -161 -325 -155
rect -265 -161 -207 -155
rect -147 -161 -89 -155
rect -29 -161 29 -155
rect 89 -161 147 -155
rect 207 -161 265 -155
rect 325 -161 383 -155
rect 443 -161 501 -155
rect 561 -161 619 -155
rect 679 -161 737 -155
rect 797 -161 855 -155
rect -855 -195 -843 -161
rect -737 -195 -725 -161
rect -619 -195 -607 -161
rect -501 -195 -489 -161
rect -383 -195 -371 -161
rect -265 -195 -253 -161
rect -147 -195 -135 -161
rect -29 -195 -17 -161
rect 89 -195 101 -161
rect 207 -195 219 -161
rect 325 -195 337 -161
rect 443 -195 455 -161
rect 561 -195 573 -161
rect 679 -195 691 -161
rect 797 -195 809 -161
rect -855 -201 -797 -195
rect -737 -201 -679 -195
rect -619 -201 -561 -195
rect -501 -201 -443 -195
rect -383 -201 -325 -195
rect -265 -201 -207 -195
rect -147 -201 -89 -195
rect -29 -201 29 -195
rect 89 -201 147 -195
rect 207 -201 265 -195
rect 325 -201 383 -195
rect 443 -201 501 -195
rect 561 -201 619 -195
rect 679 -201 737 -195
rect 797 -201 855 -195
<< nwell >>
rect -1052 -334 1052 334
<< pmos >>
rect -856 -114 -796 186
rect -738 -114 -678 186
rect -620 -114 -560 186
rect -502 -114 -442 186
rect -384 -114 -324 186
rect -266 -114 -206 186
rect -148 -114 -88 186
rect -30 -114 30 186
rect 88 -114 148 186
rect 206 -114 266 186
rect 324 -114 384 186
rect 442 -114 502 186
rect 560 -114 620 186
rect 678 -114 738 186
rect 796 -114 856 186
<< pdiff >>
rect -914 174 -856 186
rect -914 -102 -902 174
rect -868 -102 -856 174
rect -914 -114 -856 -102
rect -796 174 -738 186
rect -796 -102 -784 174
rect -750 -102 -738 174
rect -796 -114 -738 -102
rect -678 174 -620 186
rect -678 -102 -666 174
rect -632 -102 -620 174
rect -678 -114 -620 -102
rect -560 174 -502 186
rect -560 -102 -548 174
rect -514 -102 -502 174
rect -560 -114 -502 -102
rect -442 174 -384 186
rect -442 -102 -430 174
rect -396 -102 -384 174
rect -442 -114 -384 -102
rect -324 174 -266 186
rect -324 -102 -312 174
rect -278 -102 -266 174
rect -324 -114 -266 -102
rect -206 174 -148 186
rect -206 -102 -194 174
rect -160 -102 -148 174
rect -206 -114 -148 -102
rect -88 174 -30 186
rect -88 -102 -76 174
rect -42 -102 -30 174
rect -88 -114 -30 -102
rect 30 174 88 186
rect 30 -102 42 174
rect 76 -102 88 174
rect 30 -114 88 -102
rect 148 174 206 186
rect 148 -102 160 174
rect 194 -102 206 174
rect 148 -114 206 -102
rect 266 174 324 186
rect 266 -102 278 174
rect 312 -102 324 174
rect 266 -114 324 -102
rect 384 174 442 186
rect 384 -102 396 174
rect 430 -102 442 174
rect 384 -114 442 -102
rect 502 174 560 186
rect 502 -102 514 174
rect 548 -102 560 174
rect 502 -114 560 -102
rect 620 174 678 186
rect 620 -102 632 174
rect 666 -102 678 174
rect 620 -114 678 -102
rect 738 174 796 186
rect 738 -102 750 174
rect 784 -102 796 174
rect 738 -114 796 -102
rect 856 174 914 186
rect 856 -102 868 174
rect 902 -102 914 174
rect 856 -114 914 -102
<< pdiffc >>
rect -902 -102 -868 174
rect -784 -102 -750 174
rect -666 -102 -632 174
rect -548 -102 -514 174
rect -430 -102 -396 174
rect -312 -102 -278 174
rect -194 -102 -160 174
rect -76 -102 -42 174
rect 42 -102 76 174
rect 160 -102 194 174
rect 278 -102 312 174
rect 396 -102 430 174
rect 514 -102 548 174
rect 632 -102 666 174
rect 750 -102 784 174
rect 868 -102 902 174
<< nsubdiff >>
rect -1016 264 -920 298
rect 920 264 1016 298
rect -1016 201 -982 264
rect 982 201 1016 264
rect -1016 -264 -982 -201
rect 982 -264 1016 -201
rect -1016 -298 -920 -264
rect 920 -298 1016 -264
<< nsubdiffcont >>
rect -920 264 920 298
rect -1016 -201 -982 201
rect 982 -201 1016 201
rect -920 -298 920 -264
<< poly >>
rect -856 186 -796 212
rect -738 186 -678 212
rect -620 186 -560 212
rect -502 186 -442 212
rect -384 186 -324 212
rect -266 186 -206 212
rect -148 186 -88 212
rect -30 186 30 212
rect 88 186 148 212
rect 206 186 266 212
rect 324 186 384 212
rect 442 186 502 212
rect 560 186 620 212
rect 678 186 738 212
rect 796 186 856 212
rect -856 -145 -796 -114
rect -738 -145 -678 -114
rect -620 -145 -560 -114
rect -502 -145 -442 -114
rect -384 -145 -324 -114
rect -266 -145 -206 -114
rect -148 -145 -88 -114
rect -30 -145 30 -114
rect 88 -145 148 -114
rect 206 -145 266 -114
rect 324 -145 384 -114
rect 442 -145 502 -114
rect 560 -145 620 -114
rect 678 -145 738 -114
rect 796 -145 856 -114
rect -859 -161 -793 -145
rect -859 -195 -843 -161
rect -809 -195 -793 -161
rect -859 -211 -793 -195
rect -741 -161 -675 -145
rect -741 -195 -725 -161
rect -691 -195 -675 -161
rect -741 -211 -675 -195
rect -623 -161 -557 -145
rect -623 -195 -607 -161
rect -573 -195 -557 -161
rect -623 -211 -557 -195
rect -505 -161 -439 -145
rect -505 -195 -489 -161
rect -455 -195 -439 -161
rect -505 -211 -439 -195
rect -387 -161 -321 -145
rect -387 -195 -371 -161
rect -337 -195 -321 -161
rect -387 -211 -321 -195
rect -269 -161 -203 -145
rect -269 -195 -253 -161
rect -219 -195 -203 -161
rect -269 -211 -203 -195
rect -151 -161 -85 -145
rect -151 -195 -135 -161
rect -101 -195 -85 -161
rect -151 -211 -85 -195
rect -33 -161 33 -145
rect -33 -195 -17 -161
rect 17 -195 33 -161
rect -33 -211 33 -195
rect 85 -161 151 -145
rect 85 -195 101 -161
rect 135 -195 151 -161
rect 85 -211 151 -195
rect 203 -161 269 -145
rect 203 -195 219 -161
rect 253 -195 269 -161
rect 203 -211 269 -195
rect 321 -161 387 -145
rect 321 -195 337 -161
rect 371 -195 387 -161
rect 321 -211 387 -195
rect 439 -161 505 -145
rect 439 -195 455 -161
rect 489 -195 505 -161
rect 439 -211 505 -195
rect 557 -161 623 -145
rect 557 -195 573 -161
rect 607 -195 623 -161
rect 557 -211 623 -195
rect 675 -161 741 -145
rect 675 -195 691 -161
rect 725 -195 741 -161
rect 675 -211 741 -195
rect 793 -161 859 -145
rect 793 -195 809 -161
rect 843 -195 859 -161
rect 793 -211 859 -195
<< polycont >>
rect -843 -195 -809 -161
rect -725 -195 -691 -161
rect -607 -195 -573 -161
rect -489 -195 -455 -161
rect -371 -195 -337 -161
rect -253 -195 -219 -161
rect -135 -195 -101 -161
rect -17 -195 17 -161
rect 101 -195 135 -161
rect 219 -195 253 -161
rect 337 -195 371 -161
rect 455 -195 489 -161
rect 573 -195 607 -161
rect 691 -195 725 -161
rect 809 -195 843 -161
<< locali >>
rect -1016 264 -920 298
rect 920 264 1016 298
rect -1016 201 -982 264
rect 982 201 1016 264
rect -902 174 -868 190
rect -902 -118 -868 -102
rect -784 174 -750 190
rect -784 -118 -750 -102
rect -666 174 -632 190
rect -666 -118 -632 -102
rect -548 174 -514 190
rect -548 -118 -514 -102
rect -430 174 -396 190
rect -430 -118 -396 -102
rect -312 174 -278 190
rect -312 -118 -278 -102
rect -194 174 -160 190
rect -194 -118 -160 -102
rect -76 174 -42 190
rect -76 -118 -42 -102
rect 42 174 76 190
rect 42 -118 76 -102
rect 160 174 194 190
rect 160 -118 194 -102
rect 278 174 312 190
rect 278 -118 312 -102
rect 396 174 430 190
rect 396 -118 430 -102
rect 514 174 548 190
rect 514 -118 548 -102
rect 632 174 666 190
rect 632 -118 666 -102
rect 750 174 784 190
rect 750 -118 784 -102
rect 868 174 902 190
rect 868 -118 902 -102
rect -859 -195 -843 -161
rect -809 -195 -793 -161
rect -741 -195 -725 -161
rect -691 -195 -675 -161
rect -623 -195 -607 -161
rect -573 -195 -557 -161
rect -505 -195 -489 -161
rect -455 -195 -439 -161
rect -387 -195 -371 -161
rect -337 -195 -321 -161
rect -269 -195 -253 -161
rect -219 -195 -203 -161
rect -151 -195 -135 -161
rect -101 -195 -85 -161
rect -33 -195 -17 -161
rect 17 -195 33 -161
rect 85 -195 101 -161
rect 135 -195 151 -161
rect 203 -195 219 -161
rect 253 -195 269 -161
rect 321 -195 337 -161
rect 371 -195 387 -161
rect 439 -195 455 -161
rect 489 -195 505 -161
rect 557 -195 573 -161
rect 607 -195 623 -161
rect 675 -195 691 -161
rect 725 -195 741 -161
rect 793 -195 809 -161
rect 843 -195 859 -161
rect -1016 -264 -982 -201
rect 982 -264 1016 -201
rect -1016 -298 -920 -264
rect 920 -298 1016 -264
<< viali >>
rect -902 -102 -868 174
rect -784 -102 -750 174
rect -666 -102 -632 174
rect -548 -102 -514 174
rect -430 -102 -396 174
rect -312 -102 -278 174
rect -194 -102 -160 174
rect -76 -102 -42 174
rect 42 -102 76 174
rect 160 -102 194 174
rect 278 -102 312 174
rect 396 -102 430 174
rect 514 -102 548 174
rect 632 -102 666 174
rect 750 -102 784 174
rect 868 -102 902 174
rect -843 -195 -809 -161
rect -725 -195 -691 -161
rect -607 -195 -573 -161
rect -489 -195 -455 -161
rect -371 -195 -337 -161
rect -253 -195 -219 -161
rect -135 -195 -101 -161
rect -17 -195 17 -161
rect 101 -195 135 -161
rect 219 -195 253 -161
rect 337 -195 371 -161
rect 455 -195 489 -161
rect 573 -195 607 -161
rect 691 -195 725 -161
rect 809 -195 843 -161
<< metal1 >>
rect -908 174 -862 186
rect -908 -102 -902 174
rect -868 -102 -862 174
rect -908 -114 -862 -102
rect -790 174 -744 186
rect -790 -102 -784 174
rect -750 -102 -744 174
rect -790 -114 -744 -102
rect -672 174 -626 186
rect -672 -102 -666 174
rect -632 -102 -626 174
rect -672 -114 -626 -102
rect -554 174 -508 186
rect -554 -102 -548 174
rect -514 -102 -508 174
rect -554 -114 -508 -102
rect -436 174 -390 186
rect -436 -102 -430 174
rect -396 -102 -390 174
rect -436 -114 -390 -102
rect -318 174 -272 186
rect -318 -102 -312 174
rect -278 -102 -272 174
rect -318 -114 -272 -102
rect -200 174 -154 186
rect -200 -102 -194 174
rect -160 -102 -154 174
rect -200 -114 -154 -102
rect -82 174 -36 186
rect -82 -102 -76 174
rect -42 -102 -36 174
rect -82 -114 -36 -102
rect 36 174 82 186
rect 36 -102 42 174
rect 76 -102 82 174
rect 36 -114 82 -102
rect 154 174 200 186
rect 154 -102 160 174
rect 194 -102 200 174
rect 154 -114 200 -102
rect 272 174 318 186
rect 272 -102 278 174
rect 312 -102 318 174
rect 272 -114 318 -102
rect 390 174 436 186
rect 390 -102 396 174
rect 430 -102 436 174
rect 390 -114 436 -102
rect 508 174 554 186
rect 508 -102 514 174
rect 548 -102 554 174
rect 508 -114 554 -102
rect 626 174 672 186
rect 626 -102 632 174
rect 666 -102 672 174
rect 626 -114 672 -102
rect 744 174 790 186
rect 744 -102 750 174
rect 784 -102 790 174
rect 744 -114 790 -102
rect 862 174 908 186
rect 862 -102 868 174
rect 902 -102 908 174
rect 862 -114 908 -102
rect -855 -161 -797 -155
rect -855 -195 -843 -161
rect -809 -195 -797 -161
rect -855 -201 -797 -195
rect -737 -161 -679 -155
rect -737 -195 -725 -161
rect -691 -195 -679 -161
rect -737 -201 -679 -195
rect -619 -161 -561 -155
rect -619 -195 -607 -161
rect -573 -195 -561 -161
rect -619 -201 -561 -195
rect -501 -161 -443 -155
rect -501 -195 -489 -161
rect -455 -195 -443 -161
rect -501 -201 -443 -195
rect -383 -161 -325 -155
rect -383 -195 -371 -161
rect -337 -195 -325 -161
rect -383 -201 -325 -195
rect -265 -161 -207 -155
rect -265 -195 -253 -161
rect -219 -195 -207 -161
rect -265 -201 -207 -195
rect -147 -161 -89 -155
rect -147 -195 -135 -161
rect -101 -195 -89 -161
rect -147 -201 -89 -195
rect -29 -161 29 -155
rect -29 -195 -17 -161
rect 17 -195 29 -161
rect -29 -201 29 -195
rect 89 -161 147 -155
rect 89 -195 101 -161
rect 135 -195 147 -161
rect 89 -201 147 -195
rect 207 -161 265 -155
rect 207 -195 219 -161
rect 253 -195 265 -161
rect 207 -201 265 -195
rect 325 -161 383 -155
rect 325 -195 337 -161
rect 371 -195 383 -161
rect 325 -201 383 -195
rect 443 -161 501 -155
rect 443 -195 455 -161
rect 489 -195 501 -161
rect 443 -201 501 -195
rect 561 -161 619 -155
rect 561 -195 573 -161
rect 607 -195 619 -161
rect 561 -201 619 -195
rect 679 -161 737 -155
rect 679 -195 691 -161
rect 725 -195 737 -161
rect 679 -201 737 -195
rect 797 -161 855 -155
rect 797 -195 809 -161
rect 843 -195 855 -161
rect 797 -201 855 -195
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -999 -281 999 281
string parameters w 1.5 l 0.3 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
