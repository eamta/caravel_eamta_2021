magic
tech sky130A
magscale 1 2
timestamp 1619550847
<< viali >>
rect 0 8960 16400 9020
rect 0 7600 40 8960
rect 3180 7600 3340 8960
rect 6480 7600 6620 8960
rect 9780 7600 9920 8960
rect 13060 7600 13200 8960
rect 16360 7600 16400 8960
rect 0 7460 16400 7600
rect 0 6080 40 7460
rect 3180 6080 3340 7460
rect 6480 6080 6620 7460
rect 9780 6080 9920 7460
rect 13060 6080 13200 7460
rect 16360 6080 16400 7460
rect 0 5940 16400 6080
rect 0 4560 40 5940
rect 3180 4560 3340 5940
rect 6480 4560 6620 5940
rect 9780 4560 9920 5940
rect 13060 4560 13200 5940
rect 16360 4560 16400 5940
rect 0 4420 16400 4560
rect 0 3040 40 4420
rect 3180 3040 3340 4420
rect 6480 3040 6620 4420
rect 9780 3040 9920 4420
rect 13060 3040 13200 4420
rect 16360 3040 16400 4420
rect 0 2900 16400 3040
rect 0 1520 40 2900
rect 3180 1520 3340 2900
rect 6480 1520 6620 2900
rect 9780 1520 9920 2900
rect 13060 1520 13200 2900
rect 16360 1520 16400 2900
rect 0 1380 16400 1520
rect 0 20 40 1380
rect 3180 20 3340 1380
rect 6480 20 6620 1380
rect 9780 20 9920 1380
rect 13060 20 13200 1380
rect 16360 20 16400 1380
rect 0 -40 16400 20
<< metal1 >>
rect -6 9026 46 9032
rect 3174 9026 3346 9032
rect 6474 9026 6626 9032
rect 9774 9026 9926 9032
rect 13054 9026 13206 9032
rect 16354 9026 16406 9032
rect -12 9020 16412 9026
rect -12 8954 0 9020
rect -6 7606 0 8954
rect -12 7454 0 7606
rect 40 8954 3180 8960
rect 40 7606 46 8954
rect 150 8860 160 8920
rect 3060 8860 3070 8920
rect 90 8610 100 8790
rect 160 8610 170 8790
rect 390 8610 400 8790
rect 460 8610 470 8790
rect 680 8610 690 8790
rect 750 8610 760 8790
rect 980 8610 990 8790
rect 1050 8610 1060 8790
rect 1280 8610 1290 8790
rect 1350 8610 1360 8790
rect 1580 8610 1590 8790
rect 1650 8610 1660 8790
rect 1870 8610 1880 8790
rect 1940 8610 1950 8790
rect 2160 8610 2170 8790
rect 2230 8610 2240 8790
rect 2460 8610 2470 8790
rect 2530 8610 2540 8790
rect 2750 8610 2760 8790
rect 2820 8610 2830 8790
rect 3050 8610 3060 8790
rect 3120 8610 3130 8790
rect 240 8350 250 8530
rect 310 8350 320 8530
rect 540 8350 550 8530
rect 610 8350 620 8530
rect 830 8350 840 8530
rect 900 8350 910 8530
rect 1130 8350 1140 8530
rect 1200 8350 1210 8530
rect 1430 8350 1440 8530
rect 1500 8350 1510 8530
rect 1720 8350 1730 8530
rect 1790 8350 1800 8530
rect 2020 8350 2030 8530
rect 2090 8350 2100 8530
rect 2310 8350 2320 8530
rect 2380 8350 2390 8530
rect 2610 8350 2620 8530
rect 2680 8350 2690 8530
rect 2910 8350 2920 8530
rect 2980 8350 2990 8530
rect 90 8090 100 8270
rect 160 8090 170 8270
rect 390 8090 400 8270
rect 460 8090 470 8270
rect 680 8090 690 8270
rect 750 8090 760 8270
rect 980 8090 990 8270
rect 1050 8090 1060 8270
rect 1280 8090 1290 8270
rect 1350 8090 1360 8270
rect 1580 8090 1590 8270
rect 1650 8090 1660 8270
rect 1870 8090 1880 8270
rect 1940 8090 1950 8270
rect 2160 8090 2170 8270
rect 2230 8090 2240 8270
rect 2460 8090 2470 8270
rect 2530 8090 2540 8270
rect 2760 8090 2770 8270
rect 2830 8090 2840 8270
rect 3050 8090 3060 8270
rect 3120 8090 3130 8270
rect 240 7830 250 8010
rect 310 7830 320 8010
rect 530 7830 540 8010
rect 600 7830 610 8010
rect 830 7830 840 8010
rect 900 7830 910 8010
rect 1120 7830 1130 8010
rect 1190 7830 1200 8010
rect 1420 7830 1430 8010
rect 1490 7830 1500 8010
rect 1720 7830 1730 8010
rect 1790 7830 1800 8010
rect 2020 7830 2030 8010
rect 2090 7830 2100 8010
rect 2320 7830 2330 8010
rect 2390 7830 2400 8010
rect 2610 7830 2620 8010
rect 2680 7830 2690 8010
rect 2910 7830 2920 8010
rect 2980 7830 2990 8010
rect 150 7650 160 7710
rect 3060 7650 3070 7710
rect 3174 7606 3180 8954
rect 40 7600 3180 7606
rect 3340 8954 6480 8960
rect 3340 7606 3346 8954
rect 3450 8860 3460 8920
rect 6360 8860 6370 8920
rect 3390 8620 3400 8800
rect 3460 8620 3470 8800
rect 3670 8620 3680 8800
rect 3740 8620 3750 8800
rect 3970 8620 3980 8800
rect 4040 8620 4050 8800
rect 4270 8620 4280 8800
rect 4340 8620 4350 8800
rect 4570 8620 4580 8800
rect 4640 8620 4650 8800
rect 4870 8620 4880 8800
rect 4940 8620 4950 8800
rect 5150 8620 5160 8800
rect 5220 8620 5230 8800
rect 5450 8620 5460 8800
rect 5520 8620 5530 8800
rect 5750 8620 5760 8800
rect 5820 8620 5830 8800
rect 6050 8620 6060 8800
rect 6120 8620 6130 8800
rect 6330 8620 6340 8800
rect 6400 8620 6410 8800
rect 3530 8360 3540 8520
rect 3600 8360 3610 8520
rect 3830 8360 3840 8520
rect 3900 8360 3910 8520
rect 4130 8360 4140 8520
rect 4200 8360 4210 8520
rect 4430 8360 4440 8520
rect 4500 8360 4510 8520
rect 4710 8360 4720 8520
rect 4780 8360 4790 8520
rect 5010 8360 5020 8520
rect 5080 8360 5090 8520
rect 5310 8360 5320 8520
rect 5380 8360 5390 8520
rect 5590 8360 5600 8520
rect 5660 8360 5670 8520
rect 5910 8360 5920 8520
rect 5980 8360 5990 8520
rect 6190 8360 6200 8520
rect 6260 8360 6270 8520
rect 3390 8100 3400 8260
rect 3460 8100 3470 8260
rect 3690 8100 3700 8260
rect 3760 8100 3770 8260
rect 3970 8100 3980 8260
rect 4040 8100 4050 8260
rect 4270 8100 4280 8260
rect 4340 8100 4350 8260
rect 4550 8100 4560 8260
rect 4620 8100 4630 8260
rect 4870 8100 4880 8260
rect 4940 8100 4950 8260
rect 5150 8100 5160 8260
rect 5220 8100 5230 8260
rect 5450 8100 5460 8260
rect 5520 8100 5530 8260
rect 5750 8100 5760 8260
rect 5820 8100 5830 8260
rect 6050 8100 6060 8260
rect 6120 8100 6130 8260
rect 6350 8100 6360 8260
rect 6420 8100 6430 8260
rect 3530 7840 3540 8000
rect 3600 7840 3610 8000
rect 3830 7840 3840 8000
rect 3900 7840 3910 8000
rect 4130 7840 4140 8000
rect 4200 7840 4210 8000
rect 4410 7840 4420 8000
rect 4480 7840 4490 8000
rect 4710 7840 4720 8000
rect 4780 7840 4790 8000
rect 5010 7840 5020 8000
rect 5080 7840 5090 8000
rect 5310 7840 5320 8000
rect 5380 7840 5390 8000
rect 5610 7840 5620 8000
rect 5680 7840 5690 8000
rect 5910 7840 5920 8000
rect 5980 7840 5990 8000
rect 6190 7840 6200 8000
rect 6260 7840 6270 8000
rect 3450 7650 3460 7710
rect 6360 7650 6370 7710
rect 6474 7606 6480 8954
rect 3340 7600 6480 7606
rect 6620 8954 9780 8960
rect 6620 7606 6626 8954
rect 6740 8860 6750 8920
rect 9650 8860 9660 8920
rect 6670 8640 6680 8800
rect 6740 8640 6750 8800
rect 6970 8640 6980 8800
rect 7040 8640 7050 8800
rect 7270 8640 7280 8800
rect 7340 8640 7350 8800
rect 7570 8640 7580 8800
rect 7640 8640 7650 8800
rect 7870 8640 7880 8800
rect 7940 8640 7950 8800
rect 8150 8640 8160 8800
rect 8220 8640 8230 8800
rect 8450 8620 8460 8780
rect 8520 8620 8530 8780
rect 8750 8620 8760 8780
rect 8820 8620 8830 8780
rect 9030 8620 9040 8780
rect 9100 8620 9110 8780
rect 9330 8620 9340 8780
rect 9400 8620 9410 8780
rect 9630 8620 9640 8780
rect 9700 8620 9710 8780
rect 6810 8360 6820 8520
rect 6880 8360 6890 8520
rect 7110 8360 7120 8520
rect 7180 8360 7190 8520
rect 7410 8360 7420 8520
rect 7480 8360 7490 8520
rect 7710 8360 7720 8520
rect 7780 8360 7790 8520
rect 8010 8360 8020 8520
rect 8080 8360 8090 8520
rect 8310 8360 8320 8520
rect 8380 8360 8390 8520
rect 8610 8360 8620 8520
rect 8680 8360 8690 8520
rect 8910 8360 8920 8520
rect 8980 8360 8990 8520
rect 9190 8360 9200 8520
rect 9260 8360 9270 8520
rect 9490 8360 9500 8520
rect 9560 8360 9570 8520
rect 6670 8100 6680 8260
rect 6740 8100 6750 8260
rect 6970 8100 6980 8260
rect 7040 8100 7050 8260
rect 7270 8100 7280 8260
rect 7340 8100 7350 8260
rect 7570 8100 7580 8260
rect 7640 8100 7650 8260
rect 7850 8100 7860 8260
rect 7920 8100 7930 8260
rect 8150 8100 8160 8260
rect 8220 8100 8230 8260
rect 8450 8100 8460 8260
rect 8520 8100 8530 8260
rect 8750 8100 8760 8260
rect 8820 8100 8830 8260
rect 9050 8100 9060 8260
rect 9120 8100 9130 8260
rect 9330 8100 9340 8260
rect 9400 8100 9410 8260
rect 9630 8100 9640 8260
rect 9700 8100 9710 8260
rect 6830 7840 6840 8000
rect 6900 7840 6910 8000
rect 7130 7840 7140 8000
rect 7200 7840 7210 8000
rect 7410 7840 7420 8000
rect 7480 7840 7490 8000
rect 7710 7840 7720 8000
rect 7780 7840 7790 8000
rect 8010 7840 8020 8000
rect 8080 7840 8090 8000
rect 8290 7840 8300 8000
rect 8360 7840 8370 8000
rect 8610 7840 8620 8000
rect 8680 7840 8690 8000
rect 8890 7840 8900 8000
rect 8960 7840 8970 8000
rect 9190 7840 9200 8000
rect 9260 7840 9270 8000
rect 9490 7840 9500 8000
rect 9560 7840 9570 8000
rect 6740 7650 6750 7710
rect 9650 7650 9660 7710
rect 9774 7606 9780 8954
rect 6620 7600 9780 7606
rect 9920 8954 13060 8960
rect 9920 7606 9926 8954
rect 10030 8860 10040 8920
rect 12940 8860 12950 8920
rect 9970 8640 9980 8800
rect 10040 8640 10050 8800
rect 10270 8640 10280 8800
rect 10340 8640 10350 8800
rect 10570 8640 10580 8800
rect 10640 8640 10650 8800
rect 10870 8640 10880 8800
rect 10940 8640 10950 8800
rect 11150 8620 11160 8780
rect 11220 8620 11230 8780
rect 11450 8620 11460 8780
rect 11520 8620 11530 8780
rect 11750 8620 11760 8780
rect 11820 8620 11830 8780
rect 12030 8620 12040 8780
rect 12100 8620 12110 8780
rect 12350 8620 12360 8780
rect 12420 8620 12430 8780
rect 12630 8620 12640 8780
rect 12700 8620 12710 8780
rect 12930 8620 12940 8780
rect 13000 8620 13010 8780
rect 10130 8360 10140 8520
rect 10200 8360 10210 8520
rect 10410 8360 10420 8520
rect 10480 8360 10490 8520
rect 10710 8360 10720 8520
rect 10780 8360 10790 8520
rect 11010 8360 11020 8520
rect 11080 8360 11090 8520
rect 11310 8360 11320 8520
rect 11380 8360 11390 8520
rect 11590 8360 11600 8520
rect 11660 8360 11670 8520
rect 11890 8360 11900 8520
rect 11960 8360 11970 8520
rect 12190 8360 12200 8520
rect 12260 8360 12270 8520
rect 12490 8360 12500 8520
rect 12560 8360 12570 8520
rect 12790 8360 12800 8520
rect 12860 8360 12870 8520
rect 9970 8100 9980 8260
rect 10040 8100 10050 8260
rect 10270 8100 10280 8260
rect 10340 8100 10350 8260
rect 10570 8100 10580 8260
rect 10640 8100 10650 8260
rect 10850 8100 10860 8260
rect 10920 8100 10930 8260
rect 11170 8100 11180 8260
rect 11240 8100 11250 8260
rect 11450 8100 11460 8260
rect 11520 8100 11530 8260
rect 11750 8100 11760 8260
rect 11820 8100 11830 8260
rect 12050 8100 12060 8260
rect 12120 8100 12130 8260
rect 12330 8100 12340 8260
rect 12400 8100 12410 8260
rect 12630 8100 12640 8260
rect 12700 8100 12710 8260
rect 12930 8100 12940 8260
rect 13000 8100 13010 8260
rect 10130 7840 10140 8000
rect 10200 7840 10210 8000
rect 10430 7840 10440 8000
rect 10500 7840 10510 8000
rect 10710 7840 10720 8000
rect 10780 7840 10790 8000
rect 11010 7840 11020 8000
rect 11080 7840 11090 8000
rect 11310 7840 11320 8000
rect 11380 7840 11390 8000
rect 11590 7840 11600 8000
rect 11660 7840 11670 8000
rect 11890 7840 11900 8000
rect 11960 7840 11970 8000
rect 12190 7840 12200 8000
rect 12260 7840 12270 8000
rect 12490 7840 12500 8000
rect 12560 7840 12570 8000
rect 12790 7840 12800 8000
rect 12860 7840 12870 8000
rect 10030 7650 10040 7710
rect 12940 7650 12950 7710
rect 13054 7606 13060 8954
rect 9920 7600 13060 7606
rect 13200 8954 16360 8960
rect 13200 7606 13206 8954
rect 13330 8860 13340 8920
rect 16240 8860 16250 8920
rect 13270 8620 13280 8780
rect 13340 8620 13350 8780
rect 13570 8620 13580 8780
rect 13640 8620 13650 8780
rect 13850 8620 13860 8780
rect 13920 8620 13930 8780
rect 14170 8620 14180 8780
rect 14240 8620 14250 8780
rect 14450 8620 14460 8780
rect 14520 8620 14530 8780
rect 14750 8620 14760 8780
rect 14820 8620 14830 8780
rect 15030 8620 15040 8780
rect 15100 8620 15110 8780
rect 15330 8620 15340 8780
rect 15400 8620 15410 8780
rect 15630 8620 15640 8780
rect 15700 8620 15710 8780
rect 15930 8620 15940 8780
rect 16000 8620 16010 8780
rect 16230 8620 16240 8780
rect 16300 8620 16310 8780
rect 13410 8360 13420 8520
rect 13480 8360 13490 8520
rect 13710 8360 13720 8520
rect 13780 8360 13790 8520
rect 13990 8360 14000 8520
rect 14060 8360 14070 8520
rect 14310 8360 14320 8520
rect 14380 8360 14390 8520
rect 14590 8360 14600 8520
rect 14660 8360 14670 8520
rect 14890 8360 14900 8520
rect 14960 8360 14970 8520
rect 15190 8360 15200 8520
rect 15260 8360 15270 8520
rect 15490 8360 15500 8520
rect 15560 8360 15570 8520
rect 15770 8360 15780 8520
rect 15840 8360 15850 8520
rect 16070 8360 16080 8520
rect 16140 8360 16150 8520
rect 13270 8100 13280 8260
rect 13340 8100 13350 8260
rect 13570 8100 13580 8260
rect 13640 8100 13650 8260
rect 13850 8100 13860 8260
rect 13920 8100 13930 8260
rect 14170 8100 14180 8260
rect 14240 8100 14250 8260
rect 14450 8100 14460 8260
rect 14520 8100 14530 8260
rect 14750 8100 14760 8260
rect 14820 8100 14830 8260
rect 15050 8100 15060 8260
rect 15120 8100 15130 8260
rect 15350 8100 15360 8260
rect 15420 8100 15430 8260
rect 15630 8100 15640 8260
rect 15700 8100 15710 8260
rect 15930 8100 15940 8260
rect 16000 8100 16010 8260
rect 16230 8100 16240 8260
rect 16300 8100 16310 8260
rect 13410 7840 13420 8000
rect 13480 7840 13490 8000
rect 13710 7840 13720 8000
rect 13780 7840 13790 8000
rect 14010 7840 14020 8000
rect 14080 7840 14090 8000
rect 14310 7840 14320 8000
rect 14380 7840 14390 8000
rect 14590 7840 14600 8000
rect 14660 7840 14670 8000
rect 14890 7840 14900 8000
rect 14960 7840 14970 8000
rect 15190 7840 15200 8000
rect 15260 7840 15270 8000
rect 15490 7840 15500 8000
rect 15560 7840 15570 8000
rect 15790 7840 15800 8000
rect 15860 7840 15870 8000
rect 16070 7840 16080 8000
rect 16140 7840 16150 8000
rect 13330 7650 13340 7710
rect 16240 7650 16250 7710
rect 16354 7606 16360 8954
rect 13200 7600 16360 7606
rect 16400 8954 16412 9020
rect 16400 7606 16406 8954
rect 16400 7600 16412 7606
rect 16780 7460 16800 7600
rect -6 6086 0 7454
rect -12 5934 0 6086
rect 40 7454 3180 7460
rect 40 6086 46 7454
rect 150 7340 160 7400
rect 3060 7340 3070 7400
rect 90 7120 100 7280
rect 160 7120 170 7280
rect 390 7120 400 7280
rect 460 7120 470 7280
rect 690 7120 700 7280
rect 760 7120 770 7280
rect 970 7120 980 7280
rect 1040 7120 1050 7280
rect 1270 7120 1280 7280
rect 1340 7120 1350 7280
rect 1570 7120 1580 7280
rect 1640 7120 1650 7280
rect 1870 7120 1880 7280
rect 1940 7120 1950 7280
rect 2170 7120 2180 7280
rect 2240 7120 2250 7280
rect 2450 7120 2460 7280
rect 2520 7120 2530 7280
rect 2770 7120 2780 7280
rect 2840 7120 2850 7280
rect 3050 7120 3060 7280
rect 3120 7120 3130 7280
rect 250 6860 260 7020
rect 320 6860 330 7020
rect 550 6860 560 7020
rect 620 6860 630 7020
rect 830 6860 840 7020
rect 900 6860 910 7020
rect 1130 6860 1140 7020
rect 1200 6860 1210 7020
rect 1410 6860 1420 7020
rect 1480 6860 1490 7020
rect 1710 6860 1720 7020
rect 1780 6860 1790 7020
rect 2030 6860 2040 7020
rect 2100 6860 2110 7020
rect 2310 6860 2320 7020
rect 2380 6860 2390 7020
rect 2610 6860 2620 7020
rect 2680 6860 2690 7020
rect 2890 6860 2900 7020
rect 2960 6860 2970 7020
rect 90 6340 100 6500
rect 160 6340 170 6500
rect 370 6340 380 6500
rect 440 6340 450 6500
rect 690 6340 700 6500
rect 760 6340 770 6500
rect 990 6340 1000 6500
rect 1060 6340 1070 6500
rect 1270 6340 1280 6500
rect 1340 6340 1350 6500
rect 1570 6340 1580 6500
rect 1640 6340 1650 6500
rect 1870 6340 1880 6500
rect 1940 6340 1950 6500
rect 2170 6340 2180 6500
rect 2240 6340 2250 6500
rect 2470 6340 2480 6500
rect 2540 6340 2550 6500
rect 2750 6340 2760 6500
rect 2820 6340 2830 6500
rect 3050 6340 3060 6500
rect 3120 6340 3130 6500
rect 150 6130 160 6190
rect 3060 6130 3070 6190
rect 3174 6086 3180 7454
rect 40 6080 3180 6086
rect 3340 7454 6480 7460
rect 3340 6086 3346 7454
rect 3450 7340 3460 7400
rect 6360 7340 6370 7400
rect 3390 7120 3400 7280
rect 3460 7120 3470 7280
rect 3670 7120 3680 7280
rect 3740 7120 3750 7280
rect 3970 7120 3980 7280
rect 4040 7120 4050 7280
rect 4270 7120 4280 7280
rect 4340 7120 4350 7280
rect 4570 7120 4580 7280
rect 4640 7120 4650 7280
rect 4870 7120 4880 7280
rect 4940 7120 4950 7280
rect 5170 7120 5180 7280
rect 5240 7120 5250 7280
rect 5450 7120 5460 7280
rect 5520 7120 5530 7280
rect 5750 7120 5760 7280
rect 5820 7120 5830 7280
rect 6050 7120 6060 7280
rect 6120 7120 6130 7280
rect 6350 7120 6360 7280
rect 6420 7120 6430 7280
rect 3530 6860 3540 7020
rect 3600 6860 3610 7020
rect 3830 6860 3840 7020
rect 3900 6860 3910 7020
rect 4110 6860 4120 7020
rect 4180 6860 4190 7020
rect 4410 6860 4420 7020
rect 4480 6860 4490 7020
rect 4710 6860 4720 7020
rect 4780 6860 4790 7020
rect 5010 6860 5020 7020
rect 5080 6860 5090 7020
rect 5310 6860 5320 7020
rect 5380 6860 5390 7020
rect 5610 6860 5620 7020
rect 5680 6860 5690 7020
rect 5890 6860 5900 7020
rect 5960 6860 5970 7020
rect 6210 6860 6220 7020
rect 6280 6860 6290 7020
rect 3390 6340 3400 6500
rect 3460 6340 3470 6500
rect 3670 6340 3680 6500
rect 3740 6340 3750 6500
rect 3970 6340 3980 6500
rect 4040 6340 4050 6500
rect 4270 6340 4280 6500
rect 4340 6340 4350 6500
rect 4570 6340 4580 6500
rect 4640 6340 4650 6500
rect 4870 6340 4880 6500
rect 4940 6340 4950 6500
rect 5150 6340 5160 6500
rect 5220 6340 5230 6500
rect 5450 6340 5460 6500
rect 5520 6340 5530 6500
rect 5750 6340 5760 6500
rect 5820 6340 5830 6500
rect 6050 6340 6060 6500
rect 6120 6340 6130 6500
rect 6350 6340 6360 6500
rect 6420 6340 6430 6500
rect 3450 6130 3460 6190
rect 6360 6130 6370 6190
rect 6474 6086 6480 7454
rect 3340 6080 6480 6086
rect 6620 7454 9780 7460
rect 6620 6086 6626 7454
rect 6740 7340 6750 7400
rect 9650 7340 9660 7400
rect 6670 7120 6680 7280
rect 6740 7120 6750 7280
rect 6970 7120 6980 7280
rect 7040 7120 7050 7280
rect 7270 7120 7280 7280
rect 7340 7120 7350 7280
rect 7570 7120 7580 7280
rect 7640 7120 7650 7280
rect 7870 7120 7880 7280
rect 7940 7120 7950 7280
rect 8150 7120 8160 7280
rect 8220 7120 8230 7280
rect 8450 7120 8460 7280
rect 8520 7120 8530 7280
rect 8750 7120 8760 7280
rect 8820 7120 8830 7280
rect 9050 7120 9060 7280
rect 9120 7120 9130 7280
rect 9330 7120 9340 7280
rect 9400 7120 9410 7280
rect 9630 7120 9640 7280
rect 9700 7120 9710 7280
rect 6830 6600 6840 6760
rect 6900 6600 6910 6760
rect 7130 6600 7140 6760
rect 7200 6600 7210 6760
rect 7410 6600 7420 6760
rect 7480 6600 7490 6760
rect 7710 6600 7720 6760
rect 7780 6600 7790 6760
rect 8010 6600 8020 6760
rect 8080 6600 8090 6760
rect 8310 6600 8320 6760
rect 8380 6600 8390 6760
rect 8610 6600 8620 6760
rect 8680 6600 8690 6760
rect 8910 6600 8920 6760
rect 8980 6600 8990 6760
rect 9190 6600 9200 6760
rect 9260 6600 9270 6760
rect 9490 6600 9500 6760
rect 9560 6600 9570 6760
rect 6670 6340 6680 6500
rect 6740 6340 6750 6500
rect 6970 6340 6980 6500
rect 7040 6340 7050 6500
rect 7270 6340 7280 6500
rect 7340 6340 7350 6500
rect 7570 6340 7580 6500
rect 7640 6340 7650 6500
rect 7870 6340 7880 6500
rect 7940 6340 7950 6500
rect 8170 6340 8180 6500
rect 8240 6340 8250 6500
rect 8450 6340 8460 6500
rect 8520 6340 8530 6500
rect 8750 6340 8760 6500
rect 8820 6340 8830 6500
rect 9050 6340 9060 6500
rect 9120 6340 9130 6500
rect 9350 6340 9360 6500
rect 9420 6340 9430 6500
rect 9630 6340 9640 6500
rect 9700 6340 9710 6500
rect 6740 6130 6750 6190
rect 9650 6130 9660 6190
rect 9774 6086 9780 7454
rect 6620 6080 9780 6086
rect 9920 7454 13060 7460
rect 9920 6086 9926 7454
rect 10030 7340 10040 7400
rect 12940 7340 12950 7400
rect 9970 7120 9980 7280
rect 10040 7120 10050 7280
rect 10270 7120 10280 7280
rect 10340 7120 10350 7280
rect 10570 7120 10580 7280
rect 10640 7120 10650 7280
rect 10870 7120 10880 7280
rect 10940 7120 10950 7280
rect 11150 7120 11160 7280
rect 11220 7120 11230 7280
rect 11450 7120 11460 7280
rect 11520 7120 11530 7280
rect 11750 7120 11760 7280
rect 11820 7120 11830 7280
rect 12050 7120 12060 7280
rect 12120 7120 12130 7280
rect 12330 7120 12340 7280
rect 12400 7120 12410 7280
rect 12650 7120 12660 7280
rect 12720 7120 12730 7280
rect 12930 7120 12940 7280
rect 13000 7120 13010 7280
rect 10130 6860 10140 7020
rect 10200 6860 10210 7020
rect 10410 6860 10420 7020
rect 10480 6860 10490 7020
rect 10710 6860 10720 7020
rect 10780 6860 10790 7020
rect 11010 6860 11020 7020
rect 11080 6860 11090 7020
rect 11310 6860 11320 7020
rect 11380 6860 11390 7020
rect 11610 6860 11620 7020
rect 11680 6860 11690 7020
rect 11910 6860 11920 7020
rect 11980 6860 11990 7020
rect 12190 6860 12200 7020
rect 12260 6860 12270 7020
rect 12490 6860 12500 7020
rect 12560 6860 12570 7020
rect 12790 6860 12800 7020
rect 12860 6860 12870 7020
rect 9990 6340 10000 6500
rect 10060 6340 10070 6500
rect 10270 6340 10280 6500
rect 10340 6340 10350 6500
rect 10550 6340 10560 6500
rect 10620 6340 10630 6500
rect 10850 6340 10860 6500
rect 10920 6340 10930 6500
rect 11150 6340 11160 6500
rect 11220 6340 11230 6500
rect 11450 6340 11460 6500
rect 11520 6340 11530 6500
rect 11750 6340 11760 6500
rect 11820 6340 11830 6500
rect 12050 6340 12060 6500
rect 12120 6340 12130 6500
rect 12330 6340 12340 6500
rect 12400 6340 12410 6500
rect 12630 6340 12640 6500
rect 12700 6340 12710 6500
rect 12930 6340 12940 6500
rect 13000 6340 13010 6500
rect 10030 6130 10040 6190
rect 12940 6130 12950 6190
rect 13054 6086 13060 7454
rect 9920 6080 13060 6086
rect 13200 7454 16360 7460
rect 13200 6086 13206 7454
rect 13330 7340 13340 7400
rect 16240 7340 16250 7400
rect 13270 7120 13280 7280
rect 13340 7120 13350 7280
rect 13550 7120 13560 7280
rect 13620 7120 13630 7280
rect 13870 7120 13880 7280
rect 13940 7120 13950 7280
rect 14150 7120 14160 7280
rect 14220 7120 14230 7280
rect 14470 7120 14480 7280
rect 14540 7120 14550 7280
rect 14750 7120 14760 7280
rect 14820 7120 14830 7280
rect 15050 7120 15060 7280
rect 15120 7120 15130 7280
rect 15330 7120 15340 7280
rect 15400 7120 15410 7280
rect 15630 7120 15640 7280
rect 15700 7120 15710 7280
rect 15930 7120 15940 7280
rect 16000 7120 16010 7280
rect 16230 7120 16240 7280
rect 16300 7120 16310 7280
rect 13430 6860 13440 7020
rect 13500 6860 13510 7020
rect 13710 6860 13720 7020
rect 13780 6860 13790 7020
rect 14010 6860 14020 7020
rect 14080 6860 14090 7020
rect 14290 6860 14300 7020
rect 14360 6860 14370 7020
rect 14610 6860 14620 7020
rect 14680 6860 14690 7020
rect 14910 6860 14920 7020
rect 14980 6860 14990 7020
rect 15190 6860 15200 7020
rect 15260 6860 15270 7020
rect 15490 6860 15500 7020
rect 15560 6860 15570 7020
rect 15770 6860 15780 7020
rect 15840 6860 15850 7020
rect 16070 6860 16080 7020
rect 16140 6860 16150 7020
rect 13250 6340 13260 6500
rect 13320 6340 13330 6500
rect 13550 6340 13560 6500
rect 13620 6340 13630 6500
rect 13870 6340 13880 6500
rect 13940 6340 13950 6500
rect 14150 6340 14160 6500
rect 14220 6340 14230 6500
rect 14450 6340 14460 6500
rect 14520 6340 14530 6500
rect 14730 6340 14740 6500
rect 14800 6340 14810 6500
rect 15050 6340 15060 6500
rect 15120 6340 15130 6500
rect 15330 6340 15340 6500
rect 15400 6340 15410 6500
rect 15650 6340 15660 6500
rect 15720 6340 15730 6500
rect 15930 6340 15940 6500
rect 16000 6340 16010 6500
rect 16230 6340 16240 6500
rect 16300 6340 16310 6500
rect 13330 6130 13340 6190
rect 16240 6130 16250 6190
rect 16354 6086 16360 7454
rect 13200 6080 16360 6086
rect 16400 7454 16412 7460
rect 16400 6086 16406 7454
rect 16400 6080 16412 6086
rect 16780 5940 16800 6080
rect -6 4566 0 5934
rect -12 4414 0 4566
rect 40 5934 3180 5940
rect 40 4566 46 5934
rect 150 5820 160 5880
rect 3060 5820 3070 5880
rect 90 5600 100 5760
rect 160 5600 170 5760
rect 390 5600 400 5760
rect 460 5600 470 5760
rect 670 5600 680 5760
rect 740 5600 750 5760
rect 990 5600 1000 5760
rect 1060 5600 1070 5760
rect 1270 5600 1280 5760
rect 1340 5600 1350 5760
rect 1570 5600 1580 5760
rect 1640 5600 1650 5760
rect 1870 5600 1880 5760
rect 1940 5600 1950 5760
rect 2170 5600 2180 5760
rect 2240 5600 2250 5760
rect 2470 5600 2480 5760
rect 2540 5600 2550 5760
rect 2750 5600 2760 5760
rect 2820 5600 2830 5760
rect 3050 5600 3060 5760
rect 3120 5600 3130 5760
rect 250 5340 260 5500
rect 320 5340 330 5500
rect 550 5340 560 5500
rect 620 5340 630 5500
rect 830 5340 840 5500
rect 900 5340 910 5500
rect 1130 5340 1140 5500
rect 1200 5340 1210 5500
rect 1430 5340 1440 5500
rect 1500 5340 1510 5500
rect 1710 5340 1720 5500
rect 1780 5340 1790 5500
rect 2030 5340 2040 5500
rect 2100 5340 2110 5500
rect 2310 5340 2320 5500
rect 2380 5340 2390 5500
rect 2610 5340 2620 5500
rect 2680 5340 2690 5500
rect 2910 5340 2920 5500
rect 2980 5340 2990 5500
rect 150 4610 160 4670
rect 3060 4610 3070 4670
rect 3174 4566 3180 5934
rect 40 4560 3180 4566
rect 3340 5934 6480 5940
rect 3340 4566 3346 5934
rect 3450 5820 3460 5880
rect 6360 5820 6370 5880
rect 3390 5600 3400 5760
rect 3460 5600 3470 5760
rect 3670 5600 3680 5760
rect 3740 5600 3750 5760
rect 3970 5600 3980 5760
rect 4040 5600 4050 5760
rect 4270 5600 4280 5760
rect 4340 5600 4350 5760
rect 4570 5600 4580 5760
rect 4640 5600 4650 5760
rect 4850 5600 4860 5760
rect 4920 5600 4930 5760
rect 5150 5600 5160 5760
rect 5220 5600 5230 5760
rect 5450 5600 5460 5760
rect 5520 5600 5530 5760
rect 5750 5600 5760 5760
rect 5820 5600 5830 5760
rect 6050 5600 6060 5760
rect 6120 5600 6130 5760
rect 6350 5600 6360 5760
rect 6420 5600 6430 5760
rect 3550 5080 3560 5240
rect 3620 5080 3630 5240
rect 3830 5080 3840 5240
rect 3900 5080 3910 5240
rect 4130 5080 4140 5240
rect 4200 5080 4210 5240
rect 4410 5080 4420 5240
rect 4480 5080 4490 5240
rect 4730 5080 4740 5240
rect 4800 5080 4810 5240
rect 5010 5080 5020 5240
rect 5080 5080 5090 5240
rect 5310 5080 5320 5240
rect 5380 5080 5390 5240
rect 5610 5080 5620 5240
rect 5680 5080 5690 5240
rect 5890 5080 5900 5240
rect 5960 5080 5970 5240
rect 6190 5080 6200 5240
rect 6260 5080 6270 5240
rect 3450 4610 3460 4670
rect 6360 4610 6370 4670
rect 6474 4566 6480 5934
rect 3340 4560 6480 4566
rect 6620 5934 9780 5940
rect 6620 4566 6626 5934
rect 6740 5820 6750 5880
rect 9650 5820 9660 5880
rect 6670 5600 6680 5760
rect 6740 5600 6750 5760
rect 6970 5600 6980 5760
rect 7040 5600 7050 5760
rect 7270 5600 7280 5760
rect 7340 5600 7350 5760
rect 7570 5600 7580 5760
rect 7640 5600 7650 5760
rect 7870 5600 7880 5760
rect 7940 5600 7950 5760
rect 8170 5600 8180 5760
rect 8240 5600 8250 5760
rect 8450 5600 8460 5760
rect 8520 5600 8530 5760
rect 8750 5600 8760 5760
rect 8820 5600 8830 5760
rect 9050 5600 9060 5760
rect 9120 5600 9130 5760
rect 9350 5600 9360 5760
rect 9420 5600 9430 5760
rect 9650 5600 9660 5760
rect 9720 5600 9730 5760
rect 6830 4820 6840 4980
rect 6900 4820 6910 4980
rect 7130 4820 7140 4980
rect 7200 4820 7210 4980
rect 7430 4820 7440 4980
rect 7500 4820 7510 4980
rect 7710 4820 7720 4980
rect 7780 4820 7790 4980
rect 8010 4820 8020 4980
rect 8080 4820 8090 4980
rect 8310 4820 8320 4980
rect 8380 4820 8390 4980
rect 8590 4820 8600 4980
rect 8660 4820 8670 4980
rect 8890 4820 8900 4980
rect 8960 4820 8970 4980
rect 9190 4820 9200 4980
rect 9260 4820 9270 4980
rect 9490 4820 9500 4980
rect 9560 4820 9570 4980
rect 6740 4610 6750 4670
rect 9650 4610 9660 4670
rect 9774 4566 9780 5934
rect 6620 4560 9780 4566
rect 9920 5934 13060 5940
rect 9920 4566 9926 5934
rect 10030 5820 10040 5880
rect 12940 5820 12950 5880
rect 9970 5600 9980 5760
rect 10040 5600 10050 5760
rect 10270 5600 10280 5760
rect 10340 5600 10350 5760
rect 10570 5600 10580 5760
rect 10640 5600 10650 5760
rect 10870 5600 10880 5760
rect 10940 5600 10950 5760
rect 11150 5600 11160 5760
rect 11220 5600 11230 5760
rect 11450 5600 11460 5760
rect 11520 5600 11530 5760
rect 11750 5600 11760 5760
rect 11820 5600 11830 5760
rect 12050 5600 12060 5760
rect 12120 5600 12130 5760
rect 12330 5600 12340 5760
rect 12400 5600 12410 5760
rect 12630 5600 12640 5760
rect 12700 5600 12710 5760
rect 12930 5600 12940 5760
rect 13000 5600 13010 5760
rect 10110 5080 10120 5240
rect 10180 5080 10190 5240
rect 10410 5080 10420 5240
rect 10480 5080 10490 5240
rect 10730 5080 10740 5240
rect 10800 5080 10810 5240
rect 11010 5080 11020 5240
rect 11080 5080 11090 5240
rect 11310 5080 11320 5240
rect 11380 5080 11390 5240
rect 11590 5080 11600 5240
rect 11660 5080 11670 5240
rect 11910 5080 11920 5240
rect 11980 5080 11990 5240
rect 12190 5080 12200 5240
rect 12260 5080 12270 5240
rect 12490 5080 12500 5240
rect 12560 5080 12570 5240
rect 12790 5080 12800 5240
rect 12860 5080 12870 5240
rect 10030 4610 10040 4670
rect 12940 4610 12950 4670
rect 13054 4566 13060 5934
rect 9920 4560 13060 4566
rect 13200 5934 16360 5940
rect 13200 4566 13206 5934
rect 13330 5820 13340 5880
rect 16240 5820 16250 5880
rect 13270 5600 13280 5760
rect 13340 5600 13350 5760
rect 13550 5600 13560 5760
rect 13620 5600 13630 5760
rect 13870 5600 13880 5760
rect 13940 5600 13950 5760
rect 14150 5600 14160 5760
rect 14220 5600 14230 5760
rect 14450 5600 14460 5760
rect 14520 5600 14530 5760
rect 14730 5600 14740 5760
rect 14800 5600 14810 5760
rect 15050 5600 15060 5760
rect 15120 5600 15130 5760
rect 15350 5600 15360 5760
rect 15420 5600 15430 5760
rect 15630 5600 15640 5760
rect 15700 5600 15710 5760
rect 15930 5600 15940 5760
rect 16000 5600 16010 5760
rect 16230 5600 16240 5760
rect 16300 5600 16310 5760
rect 13430 5340 13440 5500
rect 13500 5340 13510 5500
rect 13710 5340 13720 5500
rect 13780 5340 13790 5500
rect 14010 5340 14020 5500
rect 14080 5340 14090 5500
rect 14310 5340 14320 5500
rect 14380 5340 14390 5500
rect 14590 5340 14600 5500
rect 14660 5340 14670 5500
rect 14890 5340 14900 5500
rect 14960 5340 14970 5500
rect 15190 5340 15200 5500
rect 15260 5340 15270 5500
rect 15490 5340 15500 5500
rect 15560 5340 15570 5500
rect 15790 5340 15800 5500
rect 15860 5340 15870 5500
rect 16070 5340 16080 5500
rect 16140 5340 16150 5500
rect 13330 4610 13340 4670
rect 16240 4610 16250 4670
rect 16354 4566 16360 5934
rect 13200 4560 16360 4566
rect 16400 5934 16412 5940
rect 16400 4566 16406 5934
rect 16400 4560 16412 4566
rect 16780 4420 16800 4560
rect -6 3046 0 4414
rect -12 2894 0 3046
rect 40 4414 3180 4420
rect 40 3046 46 4414
rect 150 4300 160 4360
rect 3060 4300 3070 4360
rect 90 4080 100 4240
rect 160 4080 170 4240
rect 390 4080 400 4240
rect 460 4080 470 4240
rect 670 4080 680 4240
rect 740 4080 750 4240
rect 970 4080 980 4240
rect 1040 4080 1050 4240
rect 1270 4080 1280 4240
rect 1340 4080 1350 4240
rect 1570 4080 1580 4240
rect 1640 4080 1650 4240
rect 1870 4080 1880 4240
rect 1940 4080 1950 4240
rect 2170 4080 2180 4240
rect 2240 4080 2250 4240
rect 2450 4080 2460 4240
rect 2520 4080 2530 4240
rect 2750 4080 2760 4240
rect 2820 4080 2830 4240
rect 3050 4080 3060 4240
rect 3120 4080 3130 4240
rect 230 3820 240 3980
rect 300 3820 310 3980
rect 530 3820 540 3980
rect 600 3820 610 3980
rect 830 3820 840 3980
rect 900 3820 910 3980
rect 1130 3820 1140 3980
rect 1200 3820 1210 3980
rect 1430 3820 1440 3980
rect 1500 3820 1510 3980
rect 1730 3820 1740 3980
rect 1800 3820 1810 3980
rect 2010 3820 2020 3980
rect 2080 3820 2090 3980
rect 2310 3820 2320 3980
rect 2380 3820 2390 3980
rect 2610 3820 2620 3980
rect 2680 3820 2690 3980
rect 2890 3820 2900 3980
rect 2960 3820 2970 3980
rect 90 3300 100 3460
rect 160 3300 170 3460
rect 390 3300 400 3460
rect 460 3300 470 3460
rect 670 3300 680 3460
rect 740 3300 750 3460
rect 970 3300 980 3460
rect 1040 3300 1050 3460
rect 1270 3300 1280 3460
rect 1340 3300 1350 3460
rect 1570 3300 1580 3460
rect 1640 3300 1650 3460
rect 1850 3300 1860 3460
rect 1920 3300 1930 3460
rect 2150 3300 2160 3460
rect 2220 3300 2230 3460
rect 2470 3300 2480 3460
rect 2540 3300 2550 3460
rect 2750 3300 2760 3460
rect 2820 3300 2830 3460
rect 3050 3300 3060 3460
rect 3120 3300 3130 3460
rect 150 3100 160 3160
rect 3060 3100 3070 3160
rect 3174 3046 3180 4414
rect 40 3040 3180 3046
rect 3340 4414 6480 4420
rect 3340 3046 3346 4414
rect 3450 4300 3460 4360
rect 6360 4300 6370 4360
rect 3390 4080 3400 4240
rect 3460 4080 3470 4240
rect 3670 4080 3680 4240
rect 3740 4080 3750 4240
rect 3970 4080 3980 4240
rect 4040 4080 4050 4240
rect 4270 4080 4280 4240
rect 4340 4080 4350 4240
rect 4550 4080 4560 4240
rect 4620 4080 4630 4240
rect 4850 4080 4860 4240
rect 4920 4080 4930 4240
rect 5150 4080 5160 4240
rect 5220 4080 5230 4240
rect 5450 4080 5460 4240
rect 5520 4080 5530 4240
rect 5770 4080 5780 4240
rect 5840 4080 5850 4240
rect 6050 4080 6060 4240
rect 6120 4080 6130 4240
rect 6350 4080 6360 4240
rect 6420 4080 6430 4240
rect 3530 3560 3540 3720
rect 3600 3560 3610 3720
rect 3830 3560 3840 3720
rect 3900 3560 3910 3720
rect 4130 3560 4140 3720
rect 4200 3560 4210 3720
rect 4410 3560 4420 3720
rect 4480 3560 4490 3720
rect 4710 3560 4720 3720
rect 4780 3560 4790 3720
rect 5010 3560 5020 3720
rect 5080 3560 5090 3720
rect 5310 3560 5320 3720
rect 5380 3560 5390 3720
rect 5610 3560 5620 3720
rect 5680 3560 5690 3720
rect 5910 3560 5920 3720
rect 5980 3560 5990 3720
rect 6190 3560 6200 3720
rect 6260 3560 6270 3720
rect 3390 3300 3400 3460
rect 3460 3300 3470 3460
rect 3670 3300 3680 3460
rect 3740 3300 3750 3460
rect 3990 3300 4000 3460
rect 4060 3300 4070 3460
rect 4270 3300 4280 3460
rect 4340 3300 4350 3460
rect 4570 3300 4580 3460
rect 4640 3300 4650 3460
rect 4850 3300 4860 3460
rect 4920 3300 4930 3460
rect 5150 3300 5160 3460
rect 5220 3300 5230 3460
rect 5450 3300 5460 3460
rect 5520 3300 5530 3460
rect 5750 3300 5760 3460
rect 5820 3300 5830 3460
rect 6050 3300 6060 3460
rect 6120 3300 6130 3460
rect 6350 3300 6360 3460
rect 6420 3300 6430 3460
rect 3450 3100 3460 3160
rect 6360 3100 6370 3160
rect 6474 3046 6480 4414
rect 3340 3040 6480 3046
rect 6620 4414 9780 4420
rect 6620 3046 6626 4414
rect 6740 4300 6750 4360
rect 9650 4300 9660 4360
rect 6690 4080 6700 4240
rect 6760 4080 6770 4240
rect 6970 4080 6980 4240
rect 7040 4080 7050 4240
rect 7270 4080 7280 4240
rect 7340 4080 7350 4240
rect 7570 4080 7580 4240
rect 7640 4080 7650 4240
rect 7870 4080 7880 4240
rect 7940 4080 7950 4240
rect 8150 4080 8160 4240
rect 8220 4080 8230 4240
rect 8450 4080 8460 4240
rect 8520 4080 8530 4240
rect 8750 4080 8760 4240
rect 8820 4080 8830 4240
rect 9050 4080 9060 4240
rect 9120 4080 9130 4240
rect 9330 4080 9340 4240
rect 9400 4080 9410 4240
rect 9630 4080 9640 4240
rect 9700 4080 9710 4240
rect 6830 3560 6840 3720
rect 6900 3560 6910 3720
rect 7130 3560 7140 3720
rect 7200 3560 7210 3720
rect 7430 3560 7440 3720
rect 7500 3560 7510 3720
rect 7710 3560 7720 3720
rect 7780 3560 7790 3720
rect 8010 3560 8020 3720
rect 8080 3560 8090 3720
rect 8310 3560 8320 3720
rect 8380 3560 8390 3720
rect 8610 3560 8620 3720
rect 8680 3560 8690 3720
rect 8890 3560 8900 3720
rect 8960 3560 8970 3720
rect 9190 3560 9200 3720
rect 9260 3560 9270 3720
rect 9490 3560 9500 3720
rect 9560 3560 9570 3720
rect 6670 3300 6680 3460
rect 6740 3300 6750 3460
rect 6970 3300 6980 3460
rect 7040 3300 7050 3460
rect 7270 3300 7280 3460
rect 7340 3300 7350 3460
rect 7570 3300 7580 3460
rect 7640 3300 7650 3460
rect 7870 3300 7880 3460
rect 7940 3300 7950 3460
rect 8150 3300 8160 3460
rect 8220 3300 8230 3460
rect 8450 3300 8460 3460
rect 8520 3300 8530 3460
rect 8770 3300 8780 3460
rect 8840 3300 8850 3460
rect 9050 3300 9060 3460
rect 9120 3300 9130 3460
rect 9350 3300 9360 3460
rect 9420 3300 9430 3460
rect 9650 3300 9660 3460
rect 9720 3300 9730 3460
rect 6740 3100 6750 3160
rect 9650 3100 9660 3160
rect 9774 3046 9780 4414
rect 6620 3040 9780 3046
rect 9920 4414 13060 4420
rect 9920 3046 9926 4414
rect 10030 4300 10040 4360
rect 12940 4300 12950 4360
rect 9970 4080 9980 4240
rect 10040 4080 10050 4240
rect 10270 4080 10280 4240
rect 10340 4080 10350 4240
rect 10550 4080 10560 4240
rect 10620 4080 10630 4240
rect 10850 4080 10860 4240
rect 10920 4080 10930 4240
rect 11150 4080 11160 4240
rect 11220 4080 11230 4240
rect 11450 4080 11460 4240
rect 11520 4080 11530 4240
rect 11750 4080 11760 4240
rect 11820 4080 11830 4240
rect 12050 4080 12060 4240
rect 12120 4080 12130 4240
rect 12330 4080 12340 4240
rect 12400 4080 12410 4240
rect 12630 4080 12640 4240
rect 12700 4080 12710 4240
rect 12930 4080 12940 4240
rect 13000 4080 13010 4240
rect 10130 3560 10140 3720
rect 10200 3560 10210 3720
rect 10410 3560 10420 3720
rect 10480 3560 10490 3720
rect 10710 3560 10720 3720
rect 10780 3560 10790 3720
rect 11010 3560 11020 3720
rect 11080 3560 11090 3720
rect 11310 3560 11320 3720
rect 11380 3560 11390 3720
rect 11590 3560 11600 3720
rect 11660 3560 11670 3720
rect 11890 3560 11900 3720
rect 11960 3560 11970 3720
rect 12190 3560 12200 3720
rect 12260 3560 12270 3720
rect 12490 3560 12500 3720
rect 12560 3560 12570 3720
rect 12790 3560 12800 3720
rect 12860 3560 12870 3720
rect 9990 3300 10000 3460
rect 10060 3300 10070 3460
rect 10270 3300 10280 3460
rect 10340 3300 10350 3460
rect 10570 3300 10580 3460
rect 10640 3300 10650 3460
rect 10850 3300 10860 3460
rect 10920 3300 10930 3460
rect 11170 3300 11180 3460
rect 11240 3300 11250 3460
rect 11450 3300 11460 3460
rect 11520 3300 11530 3460
rect 11750 3300 11760 3460
rect 11820 3300 11830 3460
rect 12050 3300 12060 3460
rect 12120 3300 12130 3460
rect 12350 3300 12360 3460
rect 12420 3300 12430 3460
rect 12630 3300 12640 3460
rect 12700 3300 12710 3460
rect 12930 3300 12940 3460
rect 13000 3300 13010 3460
rect 10030 3100 10040 3160
rect 12940 3100 12950 3160
rect 13054 3046 13060 4414
rect 9920 3040 13060 3046
rect 13200 4414 16360 4420
rect 13200 3046 13206 4414
rect 13330 4300 13340 4360
rect 16240 4300 16250 4360
rect 13270 4080 13280 4240
rect 13340 4080 13350 4240
rect 13550 4080 13560 4240
rect 13620 4080 13630 4240
rect 13850 4080 13860 4240
rect 13920 4080 13930 4240
rect 14150 4080 14160 4240
rect 14220 4080 14230 4240
rect 14450 4080 14460 4240
rect 14520 4080 14530 4240
rect 14750 4080 14760 4240
rect 14820 4080 14830 4240
rect 15050 4080 15060 4240
rect 15120 4080 15130 4240
rect 15350 4080 15360 4240
rect 15420 4080 15430 4240
rect 15630 4080 15640 4240
rect 15700 4080 15710 4240
rect 15930 4080 15940 4240
rect 16000 4080 16010 4240
rect 16210 4080 16220 4240
rect 16280 4080 16290 4240
rect 13430 3820 13440 3980
rect 13500 3820 13510 3980
rect 13710 3820 13720 3980
rect 13780 3820 13790 3980
rect 14010 3820 14020 3980
rect 14080 3820 14090 3980
rect 14310 3820 14320 3980
rect 14380 3820 14390 3980
rect 14590 3820 14600 3980
rect 14660 3820 14670 3980
rect 14890 3820 14900 3980
rect 14960 3820 14970 3980
rect 15190 3820 15200 3980
rect 15260 3820 15270 3980
rect 15490 3820 15500 3980
rect 15560 3820 15570 3980
rect 15770 3820 15780 3980
rect 15840 3820 15850 3980
rect 16070 3820 16080 3980
rect 16140 3820 16150 3980
rect 13270 3300 13280 3460
rect 13340 3300 13350 3460
rect 13550 3300 13560 3460
rect 13620 3300 13630 3460
rect 13870 3300 13880 3460
rect 13940 3300 13950 3460
rect 14170 3300 14180 3460
rect 14240 3300 14250 3460
rect 14450 3300 14460 3460
rect 14520 3300 14530 3460
rect 14730 3300 14740 3460
rect 14800 3300 14810 3460
rect 15030 3300 15040 3460
rect 15100 3300 15110 3460
rect 15350 3300 15360 3460
rect 15420 3300 15430 3460
rect 15630 3300 15640 3460
rect 15700 3300 15710 3460
rect 15930 3300 15940 3460
rect 16000 3300 16010 3460
rect 16230 3300 16240 3460
rect 16300 3300 16310 3460
rect 13330 3100 13340 3160
rect 16240 3100 16250 3160
rect 16354 3046 16360 4414
rect 13200 3040 16360 3046
rect 16400 4414 16412 4420
rect 16400 3046 16406 4414
rect 16400 3040 16412 3046
rect 16780 2900 16800 3040
rect -6 1526 0 2894
rect -12 1374 0 1526
rect 40 2894 3180 2900
rect 40 1526 46 2894
rect 140 2780 150 2840
rect 3050 2834 3060 2840
rect 3050 2800 3066 2834
rect 3050 2780 3060 2800
rect 90 2560 100 2720
rect 160 2560 170 2720
rect 390 2560 400 2720
rect 460 2560 470 2720
rect 670 2560 680 2720
rect 740 2560 750 2720
rect 970 2560 980 2720
rect 1040 2560 1050 2720
rect 1290 2560 1300 2720
rect 1360 2560 1370 2720
rect 1590 2560 1600 2720
rect 1660 2560 1670 2720
rect 1870 2560 1880 2720
rect 1940 2560 1950 2720
rect 2170 2560 2180 2720
rect 2240 2560 2250 2720
rect 2450 2560 2460 2720
rect 2520 2560 2530 2720
rect 2750 2560 2760 2720
rect 2820 2560 2830 2720
rect 3050 2560 3060 2720
rect 3120 2560 3130 2720
rect 250 2300 260 2460
rect 320 2300 330 2460
rect 530 2300 540 2460
rect 600 2300 610 2460
rect 830 2300 840 2460
rect 900 2300 910 2460
rect 1130 2300 1140 2460
rect 1200 2300 1210 2460
rect 1430 2300 1440 2460
rect 1500 2300 1510 2460
rect 1730 2300 1740 2460
rect 1800 2300 1810 2460
rect 2010 2300 2020 2460
rect 2080 2300 2090 2460
rect 2310 2300 2320 2460
rect 2380 2300 2390 2460
rect 2610 2300 2620 2460
rect 2680 2300 2690 2460
rect 2890 2300 2900 2460
rect 2960 2300 2970 2460
rect 90 1780 100 1940
rect 160 1780 170 1940
rect 390 1780 400 1940
rect 460 1780 470 1940
rect 670 1780 680 1940
rect 740 1780 750 1940
rect 990 1780 1000 1940
rect 1060 1780 1070 1940
rect 1290 1780 1300 1940
rect 1360 1780 1370 1940
rect 1590 1780 1600 1940
rect 1660 1780 1670 1940
rect 1870 1780 1880 1940
rect 1940 1780 1950 1940
rect 2170 1780 2180 1940
rect 2240 1780 2250 1940
rect 2450 1780 2460 1940
rect 2520 1780 2530 1940
rect 2750 1780 2760 1940
rect 2820 1780 2830 1940
rect 3050 1780 3060 1940
rect 3120 1780 3130 1940
rect 140 1570 150 1630
rect 3050 1624 3060 1630
rect 3050 1590 3063 1624
rect 3050 1570 3060 1590
rect 3174 1526 3180 2894
rect 40 1520 3180 1526
rect 3340 2894 6480 2900
rect 3340 1526 3346 2894
rect 3440 2780 3450 2840
rect 6350 2780 6360 2840
rect 3390 2560 3400 2720
rect 3460 2560 3470 2720
rect 3670 2560 3680 2720
rect 3740 2560 3750 2720
rect 3970 2560 3980 2720
rect 4040 2560 4050 2720
rect 4270 2560 4280 2720
rect 4340 2560 4350 2720
rect 4570 2560 4580 2720
rect 4640 2560 4650 2720
rect 4870 2560 4880 2720
rect 4940 2560 4950 2720
rect 5150 2560 5160 2720
rect 5220 2560 5230 2720
rect 5450 2560 5460 2720
rect 5520 2560 5530 2720
rect 5750 2560 5760 2720
rect 5820 2560 5830 2720
rect 6050 2560 6060 2720
rect 6120 2560 6130 2720
rect 6350 2560 6360 2720
rect 6420 2560 6430 2720
rect 3530 2000 3540 2460
rect 3620 2000 3630 2460
rect 3810 2000 3820 2460
rect 3900 2000 3910 2460
rect 4110 2000 4120 2460
rect 4200 2000 4210 2460
rect 4410 2000 4420 2460
rect 4500 2000 4510 2460
rect 4710 2000 4720 2460
rect 4800 2000 4810 2460
rect 5010 2000 5020 2460
rect 5100 2000 5110 2460
rect 5310 2000 5320 2460
rect 5400 2000 5410 2460
rect 5590 2000 5600 2460
rect 5680 2000 5690 2460
rect 5890 2000 5900 2460
rect 5980 2000 5990 2460
rect 6190 2000 6200 2460
rect 6280 2000 6290 2460
rect 3390 1780 3400 1940
rect 3460 1780 3470 1940
rect 3670 1780 3680 1940
rect 3740 1780 3750 1940
rect 3970 1780 3980 1940
rect 4040 1780 4050 1940
rect 4270 1780 4280 1940
rect 4340 1780 4350 1940
rect 4570 1780 4580 1940
rect 4640 1780 4650 1940
rect 4870 1780 4880 1940
rect 4940 1780 4950 1940
rect 5150 1780 5160 1940
rect 5220 1780 5230 1940
rect 5450 1780 5460 1940
rect 5520 1780 5530 1940
rect 5770 1780 5780 1940
rect 5840 1780 5850 1940
rect 6050 1780 6060 1940
rect 6120 1780 6130 1940
rect 6330 1780 6340 1940
rect 6400 1780 6410 1940
rect 3440 1570 3450 1630
rect 6350 1570 6360 1630
rect 6474 1526 6480 2894
rect 3340 1520 6480 1526
rect 6620 2894 9780 2900
rect 6620 1526 6626 2894
rect 6730 2780 6740 2840
rect 9640 2835 9650 2840
rect 9640 2801 9655 2835
rect 9640 2780 9650 2801
rect 6670 2560 6680 2720
rect 6740 2560 6750 2720
rect 6970 2560 6980 2720
rect 7040 2560 7050 2720
rect 7270 2560 7280 2720
rect 7340 2560 7350 2720
rect 7570 2560 7580 2720
rect 7640 2560 7650 2720
rect 7870 2560 7880 2720
rect 7940 2560 7950 2720
rect 8150 2560 8160 2720
rect 8220 2560 8230 2720
rect 8450 2560 8460 2720
rect 8520 2560 8530 2720
rect 8750 2560 8760 2720
rect 8820 2560 8830 2720
rect 9030 2560 9040 2720
rect 9100 2560 9110 2720
rect 9330 2560 9340 2720
rect 9400 2560 9410 2720
rect 9630 2560 9640 2720
rect 9700 2560 9710 2720
rect 6830 2040 6840 2200
rect 6900 2040 6910 2200
rect 7130 2040 7140 2200
rect 7200 2040 7210 2200
rect 7430 2040 7440 2200
rect 7500 2040 7510 2200
rect 7710 2040 7720 2200
rect 7780 2040 7790 2200
rect 8010 2040 8020 2200
rect 8080 2040 8090 2200
rect 8310 2040 8320 2200
rect 8380 2040 8390 2200
rect 8590 2040 8600 2200
rect 8660 2040 8670 2200
rect 8890 2040 8900 2200
rect 8960 2040 8970 2200
rect 9190 2040 9200 2200
rect 9260 2040 9270 2200
rect 9490 2040 9500 2200
rect 9560 2040 9570 2200
rect 6670 1780 6680 1940
rect 6740 1780 6750 1940
rect 6990 1780 7000 1940
rect 7060 1780 7070 1940
rect 7270 1780 7280 1940
rect 7340 1780 7350 1940
rect 7570 1780 7580 1940
rect 7640 1780 7650 1940
rect 7850 1780 7860 1940
rect 7920 1780 7930 1940
rect 8170 1780 8180 1940
rect 8240 1780 8250 1940
rect 8450 1780 8460 1940
rect 8520 1780 8530 1940
rect 8750 1780 8760 1940
rect 8820 1780 8830 1940
rect 9050 1780 9060 1940
rect 9120 1780 9130 1940
rect 9330 1780 9340 1940
rect 9400 1780 9410 1940
rect 9630 1780 9640 1940
rect 9700 1780 9710 1940
rect 6730 1570 6740 1630
rect 9640 1624 9650 1630
rect 9640 1590 9652 1624
rect 9640 1570 9650 1590
rect 9774 1526 9780 2894
rect 6620 1520 9780 1526
rect 9920 2894 13060 2900
rect 9920 1526 9926 2894
rect 10020 2780 10030 2840
rect 12930 2833 12940 2840
rect 12930 2799 12946 2833
rect 12930 2780 12940 2799
rect 9970 2560 9980 2720
rect 10040 2560 10050 2720
rect 10270 2560 10280 2720
rect 10340 2560 10350 2720
rect 10550 2560 10560 2720
rect 10620 2560 10630 2720
rect 10850 2560 10860 2720
rect 10920 2560 10930 2720
rect 11150 2560 11160 2720
rect 11220 2560 11230 2720
rect 11450 2560 11460 2720
rect 11520 2560 11530 2720
rect 11750 2560 11760 2720
rect 11820 2560 11830 2720
rect 12030 2560 12040 2720
rect 12100 2560 12110 2720
rect 12330 2560 12340 2720
rect 12400 2560 12410 2720
rect 12630 2560 12640 2720
rect 12700 2560 12710 2720
rect 12930 2560 12940 2720
rect 13000 2560 13010 2720
rect 10130 2300 10140 2460
rect 10200 2300 10210 2460
rect 10410 2300 10420 2460
rect 10480 2300 10490 2460
rect 10710 2300 10720 2460
rect 10780 2300 10790 2460
rect 11010 2300 11020 2460
rect 11080 2300 11090 2460
rect 11310 2300 11320 2460
rect 11380 2300 11390 2460
rect 11590 2300 11600 2460
rect 11660 2300 11670 2460
rect 11910 2300 11920 2460
rect 11980 2300 11990 2460
rect 12190 2300 12200 2460
rect 12260 2300 12270 2460
rect 12490 2300 12500 2460
rect 12560 2300 12570 2460
rect 12790 2300 12800 2460
rect 12860 2300 12870 2460
rect 9990 1780 10000 1940
rect 10060 1780 10070 1940
rect 10270 1780 10280 1940
rect 10340 1780 10350 1940
rect 10570 1780 10580 1940
rect 10640 1780 10650 1940
rect 10870 1780 10880 1940
rect 10940 1780 10950 1940
rect 11150 1780 11160 1940
rect 11220 1780 11230 1940
rect 11450 1780 11460 1940
rect 11520 1780 11530 1940
rect 11750 1780 11760 1940
rect 11820 1780 11830 1940
rect 12050 1780 12060 1940
rect 12120 1780 12130 1940
rect 12350 1780 12360 1940
rect 12420 1780 12430 1940
rect 12630 1780 12640 1940
rect 12700 1780 12710 1940
rect 12930 1780 12940 1940
rect 13000 1780 13010 1940
rect 10020 1570 10030 1630
rect 12930 1626 12940 1630
rect 12930 1592 12947 1626
rect 12930 1570 12940 1592
rect 13054 1526 13060 2894
rect 9920 1520 13060 1526
rect 13200 2894 16360 2900
rect 13200 1526 13206 2894
rect 13320 2780 13330 2840
rect 16230 2780 16240 2840
rect 13270 2560 13280 2720
rect 13340 2560 13350 2720
rect 13570 2560 13580 2720
rect 13640 2560 13650 2720
rect 13850 2560 13860 2720
rect 13920 2560 13930 2720
rect 14150 2560 14160 2720
rect 14220 2560 14230 2720
rect 14450 2560 14460 2720
rect 14520 2560 14530 2720
rect 14750 2560 14760 2720
rect 14820 2560 14830 2720
rect 15050 2560 15060 2720
rect 15120 2560 15130 2720
rect 15330 2560 15340 2720
rect 15400 2560 15410 2720
rect 15630 2560 15640 2720
rect 15700 2560 15710 2720
rect 15930 2560 15940 2720
rect 16000 2560 16010 2720
rect 16230 2560 16240 2720
rect 16300 2560 16310 2720
rect 13430 2300 13440 2460
rect 13500 2300 13510 2460
rect 13710 2300 13720 2460
rect 13780 2300 13790 2460
rect 14010 2300 14020 2460
rect 14080 2300 14090 2460
rect 14310 2300 14320 2460
rect 14380 2300 14390 2460
rect 14610 2300 14620 2460
rect 14680 2300 14690 2460
rect 14890 2300 14900 2460
rect 14960 2300 14970 2460
rect 15190 2300 15200 2460
rect 15260 2300 15270 2460
rect 15490 2300 15500 2460
rect 15560 2300 15570 2460
rect 15790 2300 15800 2460
rect 15860 2300 15870 2460
rect 16090 2300 16100 2460
rect 16160 2300 16170 2460
rect 13270 1780 13280 1940
rect 13340 1780 13350 1940
rect 13550 1780 13560 1940
rect 13620 1780 13630 1940
rect 13870 1780 13880 1940
rect 13940 1780 13950 1940
rect 14150 1780 14160 1940
rect 14220 1780 14230 1940
rect 14450 1780 14460 1940
rect 14520 1780 14530 1940
rect 14750 1780 14760 1940
rect 14820 1780 14830 1940
rect 15050 1780 15060 1940
rect 15120 1780 15130 1940
rect 15330 1780 15340 1940
rect 15400 1780 15410 1940
rect 15630 1780 15640 1940
rect 15700 1780 15710 1940
rect 15930 1780 15940 1940
rect 16000 1780 16010 1940
rect 16230 1780 16240 1940
rect 16300 1780 16310 1940
rect 13320 1570 13330 1630
rect 16230 1624 16240 1630
rect 16230 1590 16241 1624
rect 16230 1570 16240 1590
rect 16354 1526 16360 2894
rect 13200 1520 16360 1526
rect 16400 2894 16412 2900
rect 16400 1526 16406 2894
rect 16400 1520 16412 1526
rect 16780 1380 16800 1520
rect -6 26 0 1374
rect -12 -40 0 26
rect 40 1374 3180 1380
rect 40 26 46 1374
rect 140 1270 150 1330
rect 3050 1316 3060 1330
rect 3050 1282 3066 1316
rect 3050 1270 3060 1282
rect 90 1030 100 1210
rect 160 1030 170 1210
rect 390 1030 400 1210
rect 460 1030 470 1210
rect 690 1030 700 1210
rect 760 1030 770 1210
rect 990 1030 1000 1210
rect 1060 1030 1070 1210
rect 1270 1030 1280 1210
rect 1340 1030 1350 1210
rect 1570 1030 1580 1210
rect 1640 1030 1650 1210
rect 1870 1030 1880 1210
rect 1940 1030 1950 1210
rect 2170 1030 2180 1210
rect 2240 1030 2250 1210
rect 2470 1030 2480 1210
rect 2540 1030 2550 1210
rect 2750 1030 2760 1210
rect 2820 1030 2830 1210
rect 3050 1030 3060 1210
rect 3120 1030 3130 1210
rect 230 770 240 950
rect 300 770 310 950
rect 530 770 540 950
rect 600 770 610 950
rect 830 770 840 950
rect 900 770 910 950
rect 1130 770 1140 950
rect 1200 770 1210 950
rect 1430 770 1440 950
rect 1500 770 1510 950
rect 1730 770 1740 950
rect 1800 770 1810 950
rect 2010 770 2020 950
rect 2080 770 2090 950
rect 2310 770 2320 950
rect 2380 770 2390 950
rect 2610 770 2620 950
rect 2680 770 2690 950
rect 2910 770 2920 950
rect 2980 770 2990 950
rect 110 510 120 690
rect 180 510 190 690
rect 390 510 400 690
rect 460 510 470 690
rect 670 510 680 690
rect 740 510 750 690
rect 970 510 980 690
rect 1040 510 1050 690
rect 1290 510 1300 690
rect 1360 510 1370 690
rect 1590 510 1600 690
rect 1660 510 1670 690
rect 1870 510 1880 690
rect 1940 510 1950 690
rect 2150 510 2160 690
rect 2220 510 2230 690
rect 2470 510 2480 690
rect 2540 510 2550 690
rect 2750 510 2760 690
rect 2820 510 2830 690
rect 3050 510 3060 690
rect 3120 510 3130 690
rect 230 250 240 430
rect 300 250 310 430
rect 530 250 540 430
rect 600 250 610 430
rect 830 250 840 430
rect 900 250 910 430
rect 1130 250 1140 430
rect 1200 250 1210 430
rect 1430 250 1440 430
rect 1500 250 1510 430
rect 1730 250 1740 430
rect 1800 250 1810 430
rect 2010 250 2020 430
rect 2080 250 2090 430
rect 2330 250 2340 430
rect 2400 250 2410 430
rect 2610 250 2620 430
rect 2680 250 2690 430
rect 2910 250 2920 430
rect 2980 250 2990 430
rect 140 60 150 120
rect 3050 107 3060 120
rect 3050 73 3066 107
rect 3050 60 3060 73
rect 3174 26 3180 1374
rect 40 20 3180 26
rect 3340 1374 6480 1380
rect 3340 26 3346 1374
rect 3440 1270 3450 1330
rect 6350 1316 6360 1330
rect 6350 1282 6361 1316
rect 6350 1270 6360 1282
rect 3390 1030 3400 1210
rect 3460 1030 3470 1210
rect 3670 1030 3680 1210
rect 3740 1030 3750 1210
rect 3990 1030 4000 1210
rect 4060 1030 4070 1210
rect 4270 1030 4280 1210
rect 4340 1030 4350 1210
rect 4570 1030 4580 1210
rect 4640 1030 4650 1210
rect 4870 1030 4880 1210
rect 4940 1030 4950 1210
rect 5150 1030 5160 1210
rect 5220 1030 5230 1210
rect 5450 1030 5460 1210
rect 5520 1030 5530 1210
rect 5750 1030 5760 1210
rect 5820 1030 5830 1210
rect 6050 1030 6060 1210
rect 6120 1030 6130 1210
rect 6350 1030 6360 1210
rect 6420 1030 6430 1210
rect 3530 770 3540 950
rect 3600 770 3610 950
rect 3830 770 3840 950
rect 3900 770 3910 950
rect 4130 770 4140 950
rect 4200 770 4210 950
rect 4430 770 4440 950
rect 4500 770 4510 950
rect 4710 770 4720 950
rect 4780 770 4790 950
rect 5010 770 5020 950
rect 5080 770 5090 950
rect 5310 770 5320 950
rect 5380 770 5390 950
rect 5610 770 5620 950
rect 5680 770 5690 950
rect 5890 770 5900 950
rect 5960 770 5970 950
rect 6210 770 6220 950
rect 6280 770 6290 950
rect 3390 510 3400 690
rect 3460 510 3470 690
rect 3690 510 3700 690
rect 3760 510 3770 690
rect 3990 510 4000 690
rect 4060 510 4070 690
rect 4270 510 4280 690
rect 4340 510 4350 690
rect 4570 510 4580 690
rect 4640 510 4650 690
rect 4870 510 4880 690
rect 4940 510 4950 690
rect 5170 510 5180 690
rect 5240 510 5250 690
rect 5450 510 5460 690
rect 5520 510 5530 690
rect 5750 510 5760 690
rect 5820 510 5830 690
rect 6050 510 6060 690
rect 6120 510 6130 690
rect 6350 510 6360 690
rect 6420 510 6430 690
rect 3530 250 3540 430
rect 3600 250 3610 430
rect 3830 250 3840 430
rect 3900 250 3910 430
rect 4130 250 4140 430
rect 4200 250 4210 430
rect 4430 250 4440 430
rect 4500 250 4510 430
rect 4710 250 4720 430
rect 4780 250 4790 430
rect 5010 250 5020 430
rect 5080 250 5090 430
rect 5310 250 5320 430
rect 5380 250 5390 430
rect 5610 250 5620 430
rect 5680 250 5690 430
rect 5890 250 5900 430
rect 5960 250 5970 430
rect 6210 250 6220 430
rect 6280 250 6290 430
rect 3440 60 3450 120
rect 6350 60 6360 120
rect 6474 26 6480 1374
rect 3340 20 6480 26
rect 6620 1374 9780 1380
rect 6620 26 6626 1374
rect 6730 1270 6740 1330
rect 9640 1314 9650 1330
rect 9640 1280 9655 1314
rect 9640 1270 9650 1280
rect 6690 1030 6700 1210
rect 6760 1030 6770 1210
rect 6970 1030 6980 1210
rect 7040 1030 7050 1210
rect 7270 1030 7280 1210
rect 7340 1030 7350 1210
rect 7570 1030 7580 1210
rect 7640 1030 7650 1210
rect 7870 1030 7880 1210
rect 7940 1030 7950 1210
rect 8170 1030 8180 1210
rect 8240 1030 8250 1210
rect 8450 1030 8460 1210
rect 8520 1030 8530 1210
rect 8750 1030 8760 1210
rect 8820 1030 8830 1210
rect 9050 1030 9060 1210
rect 9120 1030 9130 1210
rect 9350 1030 9360 1210
rect 9420 1030 9430 1210
rect 9630 1030 9640 1210
rect 9700 1030 9710 1210
rect 6830 770 6840 950
rect 6900 770 6910 950
rect 7130 770 7140 950
rect 7200 770 7210 950
rect 7410 770 7420 950
rect 7480 770 7490 950
rect 7710 770 7720 950
rect 7780 770 7790 950
rect 8010 770 8020 950
rect 8080 770 8090 950
rect 8290 770 8300 950
rect 8360 770 8370 950
rect 8610 770 8620 950
rect 8680 770 8690 950
rect 8910 770 8920 950
rect 8980 770 8990 950
rect 9210 770 9220 950
rect 9280 770 9290 950
rect 9510 770 9520 950
rect 9580 770 9590 950
rect 6690 510 6700 690
rect 6760 510 6770 690
rect 6990 510 7000 690
rect 7060 510 7070 690
rect 7270 510 7280 690
rect 7340 510 7350 690
rect 7570 510 7580 690
rect 7640 510 7650 690
rect 7850 510 7860 690
rect 7920 510 7930 690
rect 8170 510 8180 690
rect 8240 510 8250 690
rect 8470 510 8480 690
rect 8540 510 8550 690
rect 8750 510 8760 690
rect 8820 510 8830 690
rect 9050 510 9060 690
rect 9120 510 9130 690
rect 9350 510 9360 690
rect 9420 510 9430 690
rect 9650 510 9660 690
rect 9720 510 9730 690
rect 6830 250 6840 430
rect 6900 250 6910 430
rect 7130 250 7140 430
rect 7200 250 7210 430
rect 7430 250 7440 430
rect 7500 250 7510 430
rect 7710 250 7720 430
rect 7780 250 7790 430
rect 8010 250 8020 430
rect 8080 250 8090 430
rect 8310 250 8320 430
rect 8380 250 8390 430
rect 8610 250 8620 430
rect 8680 250 8690 430
rect 8910 250 8920 430
rect 8980 250 8990 430
rect 9190 250 9200 430
rect 9260 250 9270 430
rect 9510 250 9520 430
rect 9580 250 9590 430
rect 6730 60 6740 120
rect 9640 107 9650 120
rect 9640 73 9652 107
rect 9640 60 9650 73
rect 9774 26 9780 1374
rect 6620 20 9780 26
rect 9920 1374 13060 1380
rect 9920 26 9926 1374
rect 10020 1270 10030 1330
rect 12930 1315 12940 1330
rect 12930 1281 12945 1315
rect 12930 1270 12940 1281
rect 9970 1030 9980 1210
rect 10040 1030 10050 1210
rect 10270 1030 10280 1210
rect 10340 1030 10350 1210
rect 10550 1030 10560 1210
rect 10620 1030 10630 1210
rect 10850 1030 10860 1210
rect 10920 1030 10930 1210
rect 11150 1030 11160 1210
rect 11220 1030 11230 1210
rect 11450 1030 11460 1210
rect 11520 1030 11530 1210
rect 11750 1030 11760 1210
rect 11820 1030 11830 1210
rect 12050 1030 12060 1210
rect 12120 1030 12130 1210
rect 12350 1030 12360 1210
rect 12420 1030 12430 1210
rect 12650 1030 12660 1210
rect 12720 1030 12730 1210
rect 12930 1030 12940 1210
rect 13000 1030 13010 1210
rect 10130 770 10140 950
rect 10200 770 10210 950
rect 10410 770 10420 950
rect 10480 770 10490 950
rect 10730 770 10740 950
rect 10800 770 10810 950
rect 11010 770 11020 950
rect 11080 770 11090 950
rect 11310 770 11320 950
rect 11380 770 11390 950
rect 11610 770 11620 950
rect 11680 770 11690 950
rect 11910 770 11920 950
rect 11980 770 11990 950
rect 12210 770 12220 950
rect 12280 770 12290 950
rect 12490 770 12500 950
rect 12560 770 12570 950
rect 12790 770 12800 950
rect 12860 770 12870 950
rect 9990 510 10000 690
rect 10060 510 10070 690
rect 10270 510 10280 690
rect 10340 510 10350 690
rect 10570 510 10580 690
rect 10640 510 10650 690
rect 10850 510 10860 690
rect 10920 510 10930 690
rect 11150 510 11160 690
rect 11220 510 11230 690
rect 11470 510 11480 690
rect 11540 510 11550 690
rect 11750 510 11760 690
rect 11820 510 11830 690
rect 12050 510 12060 690
rect 12120 510 12130 690
rect 12350 510 12360 690
rect 12420 510 12430 690
rect 12650 510 12660 690
rect 12720 510 12730 690
rect 12930 510 12940 690
rect 13000 510 13010 690
rect 10130 250 10140 430
rect 10200 250 10210 430
rect 10430 250 10440 430
rect 10500 250 10510 430
rect 10730 250 10740 430
rect 10800 250 10810 430
rect 11010 250 11020 430
rect 11080 250 11090 430
rect 11290 250 11300 430
rect 11360 250 11370 430
rect 11590 250 11600 430
rect 11660 250 11670 430
rect 11890 250 11900 430
rect 11960 250 11970 430
rect 12210 250 12220 430
rect 12280 250 12290 430
rect 12490 250 12500 430
rect 12560 250 12570 430
rect 12790 250 12800 430
rect 12860 250 12870 430
rect 10020 60 10030 120
rect 12930 106 12940 120
rect 12930 72 12948 106
rect 12930 60 12940 72
rect 13054 26 13060 1374
rect 9920 20 13060 26
rect 13200 1374 16360 1380
rect 13200 26 13206 1374
rect 13320 1270 13330 1330
rect 16230 1316 16240 1330
rect 16230 1282 16242 1316
rect 16230 1270 16240 1282
rect 13270 1030 13280 1210
rect 13340 1030 13350 1210
rect 13570 1030 13580 1210
rect 13640 1030 13650 1210
rect 13870 1030 13880 1210
rect 13940 1030 13950 1210
rect 14170 1030 14180 1210
rect 14240 1030 14250 1210
rect 14450 1030 14460 1210
rect 14520 1030 14530 1210
rect 14750 1030 14760 1210
rect 14820 1030 14830 1210
rect 15050 1030 15060 1210
rect 15120 1030 15130 1210
rect 15350 1030 15360 1210
rect 15420 1030 15430 1210
rect 15630 1030 15640 1210
rect 15700 1030 15710 1210
rect 15950 1030 15960 1210
rect 16020 1030 16030 1210
rect 16230 1030 16240 1210
rect 16300 1030 16310 1210
rect 13410 770 13420 950
rect 13480 770 13490 950
rect 13730 770 13740 950
rect 13800 770 13810 950
rect 14010 770 14020 950
rect 14080 770 14090 950
rect 14290 770 14300 950
rect 14360 770 14370 950
rect 14610 770 14620 950
rect 14680 770 14690 950
rect 14910 770 14920 950
rect 14980 770 14990 950
rect 15190 770 15200 950
rect 15260 770 15270 950
rect 15490 770 15500 950
rect 15560 770 15570 950
rect 15770 770 15780 950
rect 15840 770 15850 950
rect 16090 770 16100 950
rect 16160 770 16170 950
rect 13270 510 13280 690
rect 13340 510 13350 690
rect 13570 510 13580 690
rect 13640 510 13650 690
rect 13870 510 13880 690
rect 13940 510 13950 690
rect 14150 510 14160 690
rect 14220 510 14230 690
rect 14450 510 14460 690
rect 14520 510 14530 690
rect 14750 510 14760 690
rect 14820 510 14830 690
rect 15050 510 15060 690
rect 15120 510 15130 690
rect 15350 510 15360 690
rect 15420 510 15430 690
rect 15630 510 15640 690
rect 15700 510 15710 690
rect 15930 510 15940 690
rect 16000 510 16010 690
rect 16230 510 16240 690
rect 16300 510 16310 690
rect 13430 250 13440 430
rect 13500 250 13510 430
rect 13730 250 13740 430
rect 13800 250 13810 430
rect 14010 250 14020 430
rect 14080 250 14090 430
rect 14310 250 14320 430
rect 14380 250 14390 430
rect 14590 250 14600 430
rect 14660 250 14670 430
rect 14890 250 14900 430
rect 14960 250 14970 430
rect 15190 250 15200 430
rect 15260 250 15270 430
rect 15490 250 15500 430
rect 15560 250 15570 430
rect 15770 250 15780 430
rect 15840 250 15850 430
rect 16090 250 16100 430
rect 16160 250 16170 430
rect 13320 60 13330 120
rect 16230 60 16240 120
rect 16354 26 16360 1374
rect 13200 20 16360 26
rect 16400 1374 16412 1380
rect 16400 26 16406 1374
rect 16400 -40 16412 26
rect -12 -46 16412 -40
rect -6 -52 46 -46
rect 3174 -52 3346 -46
rect 6474 -52 6626 -46
rect 9774 -52 9926 -46
rect 13054 -52 13206 -46
rect 16354 -52 16406 -46
<< via1 >>
rect 160 8860 3060 8920
rect 100 8610 160 8790
rect 400 8610 460 8790
rect 690 8610 750 8790
rect 990 8610 1050 8790
rect 1290 8610 1350 8790
rect 1590 8610 1650 8790
rect 1880 8610 1940 8790
rect 2170 8610 2230 8790
rect 2470 8610 2530 8790
rect 2760 8610 2820 8790
rect 3060 8610 3120 8790
rect 250 8350 310 8530
rect 550 8350 610 8530
rect 840 8350 900 8530
rect 1140 8350 1200 8530
rect 1440 8350 1500 8530
rect 1730 8350 1790 8530
rect 2030 8350 2090 8530
rect 2320 8350 2380 8530
rect 2620 8350 2680 8530
rect 2920 8350 2980 8530
rect 100 8090 160 8270
rect 400 8090 460 8270
rect 690 8090 750 8270
rect 990 8090 1050 8270
rect 1290 8090 1350 8270
rect 1590 8090 1650 8270
rect 1880 8090 1940 8270
rect 2170 8090 2230 8270
rect 2470 8090 2530 8270
rect 2770 8090 2830 8270
rect 3060 8090 3120 8270
rect 250 7830 310 8010
rect 540 7830 600 8010
rect 840 7830 900 8010
rect 1130 7830 1190 8010
rect 1430 7830 1490 8010
rect 1730 7830 1790 8010
rect 2030 7830 2090 8010
rect 2330 7830 2390 8010
rect 2620 7830 2680 8010
rect 2920 7830 2980 8010
rect 160 7650 3060 7710
rect 3460 8860 6360 8920
rect 3400 8620 3460 8800
rect 3680 8620 3740 8800
rect 3980 8620 4040 8800
rect 4280 8620 4340 8800
rect 4580 8620 4640 8800
rect 4880 8620 4940 8800
rect 5160 8620 5220 8800
rect 5460 8620 5520 8800
rect 5760 8620 5820 8800
rect 6060 8620 6120 8800
rect 6340 8620 6400 8800
rect 3540 8360 3600 8520
rect 3840 8360 3900 8520
rect 4140 8360 4200 8520
rect 4440 8360 4500 8520
rect 4720 8360 4780 8520
rect 5020 8360 5080 8520
rect 5320 8360 5380 8520
rect 5600 8360 5660 8520
rect 5920 8360 5980 8520
rect 6200 8360 6260 8520
rect 3400 8100 3460 8260
rect 3700 8100 3760 8260
rect 3980 8100 4040 8260
rect 4280 8100 4340 8260
rect 4560 8100 4620 8260
rect 4880 8100 4940 8260
rect 5160 8100 5220 8260
rect 5460 8100 5520 8260
rect 5760 8100 5820 8260
rect 6060 8100 6120 8260
rect 6360 8100 6420 8260
rect 3540 7840 3600 8000
rect 3840 7840 3900 8000
rect 4140 7840 4200 8000
rect 4420 7840 4480 8000
rect 4720 7840 4780 8000
rect 5020 7840 5080 8000
rect 5320 7840 5380 8000
rect 5620 7840 5680 8000
rect 5920 7840 5980 8000
rect 6200 7840 6260 8000
rect 3460 7650 6360 7710
rect 6750 8860 9650 8920
rect 6680 8640 6740 8800
rect 6980 8640 7040 8800
rect 7280 8640 7340 8800
rect 7580 8640 7640 8800
rect 7880 8640 7940 8800
rect 8160 8640 8220 8800
rect 8460 8620 8520 8780
rect 8760 8620 8820 8780
rect 9040 8620 9100 8780
rect 9340 8620 9400 8780
rect 9640 8620 9700 8780
rect 6820 8360 6880 8520
rect 7120 8360 7180 8520
rect 7420 8360 7480 8520
rect 7720 8360 7780 8520
rect 8020 8360 8080 8520
rect 8320 8360 8380 8520
rect 8620 8360 8680 8520
rect 8920 8360 8980 8520
rect 9200 8360 9260 8520
rect 9500 8360 9560 8520
rect 6680 8100 6740 8260
rect 6980 8100 7040 8260
rect 7280 8100 7340 8260
rect 7580 8100 7640 8260
rect 7860 8100 7920 8260
rect 8160 8100 8220 8260
rect 8460 8100 8520 8260
rect 8760 8100 8820 8260
rect 9060 8100 9120 8260
rect 9340 8100 9400 8260
rect 9640 8100 9700 8260
rect 6840 7840 6900 8000
rect 7140 7840 7200 8000
rect 7420 7840 7480 8000
rect 7720 7840 7780 8000
rect 8020 7840 8080 8000
rect 8300 7840 8360 8000
rect 8620 7840 8680 8000
rect 8900 7840 8960 8000
rect 9200 7840 9260 8000
rect 9500 7840 9560 8000
rect 6750 7650 9650 7710
rect 10040 8860 12940 8920
rect 9980 8640 10040 8800
rect 10280 8640 10340 8800
rect 10580 8640 10640 8800
rect 10880 8640 10940 8800
rect 11160 8620 11220 8780
rect 11460 8620 11520 8780
rect 11760 8620 11820 8780
rect 12040 8620 12100 8780
rect 12360 8620 12420 8780
rect 12640 8620 12700 8780
rect 12940 8620 13000 8780
rect 10140 8360 10200 8520
rect 10420 8360 10480 8520
rect 10720 8360 10780 8520
rect 11020 8360 11080 8520
rect 11320 8360 11380 8520
rect 11600 8360 11660 8520
rect 11900 8360 11960 8520
rect 12200 8360 12260 8520
rect 12500 8360 12560 8520
rect 12800 8360 12860 8520
rect 9980 8100 10040 8260
rect 10280 8100 10340 8260
rect 10580 8100 10640 8260
rect 10860 8100 10920 8260
rect 11180 8100 11240 8260
rect 11460 8100 11520 8260
rect 11760 8100 11820 8260
rect 12060 8100 12120 8260
rect 12340 8100 12400 8260
rect 12640 8100 12700 8260
rect 12940 8100 13000 8260
rect 10140 7840 10200 8000
rect 10440 7840 10500 8000
rect 10720 7840 10780 8000
rect 11020 7840 11080 8000
rect 11320 7840 11380 8000
rect 11600 7840 11660 8000
rect 11900 7840 11960 8000
rect 12200 7840 12260 8000
rect 12500 7840 12560 8000
rect 12800 7840 12860 8000
rect 10040 7650 12940 7710
rect 13340 8860 16240 8920
rect 13280 8620 13340 8780
rect 13580 8620 13640 8780
rect 13860 8620 13920 8780
rect 14180 8620 14240 8780
rect 14460 8620 14520 8780
rect 14760 8620 14820 8780
rect 15040 8620 15100 8780
rect 15340 8620 15400 8780
rect 15640 8620 15700 8780
rect 15940 8620 16000 8780
rect 16240 8620 16300 8780
rect 13420 8360 13480 8520
rect 13720 8360 13780 8520
rect 14000 8360 14060 8520
rect 14320 8360 14380 8520
rect 14600 8360 14660 8520
rect 14900 8360 14960 8520
rect 15200 8360 15260 8520
rect 15500 8360 15560 8520
rect 15780 8360 15840 8520
rect 16080 8360 16140 8520
rect 13280 8100 13340 8260
rect 13580 8100 13640 8260
rect 13860 8100 13920 8260
rect 14180 8100 14240 8260
rect 14460 8100 14520 8260
rect 14760 8100 14820 8260
rect 15060 8100 15120 8260
rect 15360 8100 15420 8260
rect 15640 8100 15700 8260
rect 15940 8100 16000 8260
rect 16240 8100 16300 8260
rect 13420 7840 13480 8000
rect 13720 7840 13780 8000
rect 14020 7840 14080 8000
rect 14320 7840 14380 8000
rect 14600 7840 14660 8000
rect 14900 7840 14960 8000
rect 15200 7840 15260 8000
rect 15500 7840 15560 8000
rect 15800 7840 15860 8000
rect 16080 7840 16140 8000
rect 13340 7650 16240 7710
rect 16400 7460 16780 7600
rect 160 7340 3060 7400
rect 100 7120 160 7280
rect 400 7120 460 7280
rect 700 7120 760 7280
rect 980 7120 1040 7280
rect 1280 7120 1340 7280
rect 1580 7120 1640 7280
rect 1880 7120 1940 7280
rect 2180 7120 2240 7280
rect 2460 7120 2520 7280
rect 2780 7120 2840 7280
rect 3060 7120 3120 7280
rect 260 6860 320 7020
rect 560 6860 620 7020
rect 840 6860 900 7020
rect 1140 6860 1200 7020
rect 1420 6860 1480 7020
rect 1720 6860 1780 7020
rect 2040 6860 2100 7020
rect 2320 6860 2380 7020
rect 2620 6860 2680 7020
rect 2900 6860 2960 7020
rect 100 6340 160 6500
rect 380 6340 440 6500
rect 700 6340 760 6500
rect 1000 6340 1060 6500
rect 1280 6340 1340 6500
rect 1580 6340 1640 6500
rect 1880 6340 1940 6500
rect 2180 6340 2240 6500
rect 2480 6340 2540 6500
rect 2760 6340 2820 6500
rect 3060 6340 3120 6500
rect 160 6130 3060 6190
rect 3460 7340 6360 7400
rect 3400 7120 3460 7280
rect 3680 7120 3740 7280
rect 3980 7120 4040 7280
rect 4280 7120 4340 7280
rect 4580 7120 4640 7280
rect 4880 7120 4940 7280
rect 5180 7120 5240 7280
rect 5460 7120 5520 7280
rect 5760 7120 5820 7280
rect 6060 7120 6120 7280
rect 6360 7120 6420 7280
rect 3540 6860 3600 7020
rect 3840 6860 3900 7020
rect 4120 6860 4180 7020
rect 4420 6860 4480 7020
rect 4720 6860 4780 7020
rect 5020 6860 5080 7020
rect 5320 6860 5380 7020
rect 5620 6860 5680 7020
rect 5900 6860 5960 7020
rect 6220 6860 6280 7020
rect 3400 6340 3460 6500
rect 3680 6340 3740 6500
rect 3980 6340 4040 6500
rect 4280 6340 4340 6500
rect 4580 6340 4640 6500
rect 4880 6340 4940 6500
rect 5160 6340 5220 6500
rect 5460 6340 5520 6500
rect 5760 6340 5820 6500
rect 6060 6340 6120 6500
rect 6360 6340 6420 6500
rect 3460 6130 6360 6190
rect 6750 7340 9650 7400
rect 6680 7120 6740 7280
rect 6980 7120 7040 7280
rect 7280 7120 7340 7280
rect 7580 7120 7640 7280
rect 7880 7120 7940 7280
rect 8160 7120 8220 7280
rect 8460 7120 8520 7280
rect 8760 7120 8820 7280
rect 9060 7120 9120 7280
rect 9340 7120 9400 7280
rect 9640 7120 9700 7280
rect 6840 6600 6900 6760
rect 7140 6600 7200 6760
rect 7420 6600 7480 6760
rect 7720 6600 7780 6760
rect 8020 6600 8080 6760
rect 8320 6600 8380 6760
rect 8620 6600 8680 6760
rect 8920 6600 8980 6760
rect 9200 6600 9260 6760
rect 9500 6600 9560 6760
rect 6680 6340 6740 6500
rect 6980 6340 7040 6500
rect 7280 6340 7340 6500
rect 7580 6340 7640 6500
rect 7880 6340 7940 6500
rect 8180 6340 8240 6500
rect 8460 6340 8520 6500
rect 8760 6340 8820 6500
rect 9060 6340 9120 6500
rect 9360 6340 9420 6500
rect 9640 6340 9700 6500
rect 6750 6130 9650 6190
rect 10040 7340 12940 7400
rect 9980 7120 10040 7280
rect 10280 7120 10340 7280
rect 10580 7120 10640 7280
rect 10880 7120 10940 7280
rect 11160 7120 11220 7280
rect 11460 7120 11520 7280
rect 11760 7120 11820 7280
rect 12060 7120 12120 7280
rect 12340 7120 12400 7280
rect 12660 7120 12720 7280
rect 12940 7120 13000 7280
rect 10140 6860 10200 7020
rect 10420 6860 10480 7020
rect 10720 6860 10780 7020
rect 11020 6860 11080 7020
rect 11320 6860 11380 7020
rect 11620 6860 11680 7020
rect 11920 6860 11980 7020
rect 12200 6860 12260 7020
rect 12500 6860 12560 7020
rect 12800 6860 12860 7020
rect 10000 6340 10060 6500
rect 10280 6340 10340 6500
rect 10560 6340 10620 6500
rect 10860 6340 10920 6500
rect 11160 6340 11220 6500
rect 11460 6340 11520 6500
rect 11760 6340 11820 6500
rect 12060 6340 12120 6500
rect 12340 6340 12400 6500
rect 12640 6340 12700 6500
rect 12940 6340 13000 6500
rect 10040 6130 12940 6190
rect 13340 7340 16240 7400
rect 13280 7120 13340 7280
rect 13560 7120 13620 7280
rect 13880 7120 13940 7280
rect 14160 7120 14220 7280
rect 14480 7120 14540 7280
rect 14760 7120 14820 7280
rect 15060 7120 15120 7280
rect 15340 7120 15400 7280
rect 15640 7120 15700 7280
rect 15940 7120 16000 7280
rect 16240 7120 16300 7280
rect 13440 6860 13500 7020
rect 13720 6860 13780 7020
rect 14020 6860 14080 7020
rect 14300 6860 14360 7020
rect 14620 6860 14680 7020
rect 14920 6860 14980 7020
rect 15200 6860 15260 7020
rect 15500 6860 15560 7020
rect 15780 6860 15840 7020
rect 16080 6860 16140 7020
rect 13260 6340 13320 6500
rect 13560 6340 13620 6500
rect 13880 6340 13940 6500
rect 14160 6340 14220 6500
rect 14460 6340 14520 6500
rect 14740 6340 14800 6500
rect 15060 6340 15120 6500
rect 15340 6340 15400 6500
rect 15660 6340 15720 6500
rect 15940 6340 16000 6500
rect 16240 6340 16300 6500
rect 13340 6130 16240 6190
rect 16400 5940 16780 6080
rect 160 5820 3060 5880
rect 100 5600 160 5760
rect 400 5600 460 5760
rect 680 5600 740 5760
rect 1000 5600 1060 5760
rect 1280 5600 1340 5760
rect 1580 5600 1640 5760
rect 1880 5600 1940 5760
rect 2180 5600 2240 5760
rect 2480 5600 2540 5760
rect 2760 5600 2820 5760
rect 3060 5600 3120 5760
rect 260 5340 320 5500
rect 560 5340 620 5500
rect 840 5340 900 5500
rect 1140 5340 1200 5500
rect 1440 5340 1500 5500
rect 1720 5340 1780 5500
rect 2040 5340 2100 5500
rect 2320 5340 2380 5500
rect 2620 5340 2680 5500
rect 2920 5340 2980 5500
rect 160 4610 3060 4670
rect 3460 5820 6360 5880
rect 3400 5600 3460 5760
rect 3680 5600 3740 5760
rect 3980 5600 4040 5760
rect 4280 5600 4340 5760
rect 4580 5600 4640 5760
rect 4860 5600 4920 5760
rect 5160 5600 5220 5760
rect 5460 5600 5520 5760
rect 5760 5600 5820 5760
rect 6060 5600 6120 5760
rect 6360 5600 6420 5760
rect 3560 5080 3620 5240
rect 3840 5080 3900 5240
rect 4140 5080 4200 5240
rect 4420 5080 4480 5240
rect 4740 5080 4800 5240
rect 5020 5080 5080 5240
rect 5320 5080 5380 5240
rect 5620 5080 5680 5240
rect 5900 5080 5960 5240
rect 6200 5080 6260 5240
rect 3460 4610 6360 4670
rect 6750 5820 9650 5880
rect 6680 5600 6740 5760
rect 6980 5600 7040 5760
rect 7280 5600 7340 5760
rect 7580 5600 7640 5760
rect 7880 5600 7940 5760
rect 8180 5600 8240 5760
rect 8460 5600 8520 5760
rect 8760 5600 8820 5760
rect 9060 5600 9120 5760
rect 9360 5600 9420 5760
rect 9660 5600 9720 5760
rect 6840 4820 6900 4980
rect 7140 4820 7200 4980
rect 7440 4820 7500 4980
rect 7720 4820 7780 4980
rect 8020 4820 8080 4980
rect 8320 4820 8380 4980
rect 8600 4820 8660 4980
rect 8900 4820 8960 4980
rect 9200 4820 9260 4980
rect 9500 4820 9560 4980
rect 6750 4610 9650 4670
rect 10040 5820 12940 5880
rect 9980 5600 10040 5760
rect 10280 5600 10340 5760
rect 10580 5600 10640 5760
rect 10880 5600 10940 5760
rect 11160 5600 11220 5760
rect 11460 5600 11520 5760
rect 11760 5600 11820 5760
rect 12060 5600 12120 5760
rect 12340 5600 12400 5760
rect 12640 5600 12700 5760
rect 12940 5600 13000 5760
rect 10120 5080 10180 5240
rect 10420 5080 10480 5240
rect 10740 5080 10800 5240
rect 11020 5080 11080 5240
rect 11320 5080 11380 5240
rect 11600 5080 11660 5240
rect 11920 5080 11980 5240
rect 12200 5080 12260 5240
rect 12500 5080 12560 5240
rect 12800 5080 12860 5240
rect 10040 4610 12940 4670
rect 13340 5820 16240 5880
rect 13280 5600 13340 5760
rect 13560 5600 13620 5760
rect 13880 5600 13940 5760
rect 14160 5600 14220 5760
rect 14460 5600 14520 5760
rect 14740 5600 14800 5760
rect 15060 5600 15120 5760
rect 15360 5600 15420 5760
rect 15640 5600 15700 5760
rect 15940 5600 16000 5760
rect 16240 5600 16300 5760
rect 13440 5340 13500 5500
rect 13720 5340 13780 5500
rect 14020 5340 14080 5500
rect 14320 5340 14380 5500
rect 14600 5340 14660 5500
rect 14900 5340 14960 5500
rect 15200 5340 15260 5500
rect 15500 5340 15560 5500
rect 15800 5340 15860 5500
rect 16080 5340 16140 5500
rect 13340 4610 16240 4670
rect 16400 4420 16780 4560
rect 160 4300 3060 4360
rect 100 4080 160 4240
rect 400 4080 460 4240
rect 680 4080 740 4240
rect 980 4080 1040 4240
rect 1280 4080 1340 4240
rect 1580 4080 1640 4240
rect 1880 4080 1940 4240
rect 2180 4080 2240 4240
rect 2460 4080 2520 4240
rect 2760 4080 2820 4240
rect 3060 4080 3120 4240
rect 240 3820 300 3980
rect 540 3820 600 3980
rect 840 3820 900 3980
rect 1140 3820 1200 3980
rect 1440 3820 1500 3980
rect 1740 3820 1800 3980
rect 2020 3820 2080 3980
rect 2320 3820 2380 3980
rect 2620 3820 2680 3980
rect 2900 3820 2960 3980
rect 100 3300 160 3460
rect 400 3300 460 3460
rect 680 3300 740 3460
rect 980 3300 1040 3460
rect 1280 3300 1340 3460
rect 1580 3300 1640 3460
rect 1860 3300 1920 3460
rect 2160 3300 2220 3460
rect 2480 3300 2540 3460
rect 2760 3300 2820 3460
rect 3060 3300 3120 3460
rect 160 3100 3060 3160
rect 3460 4300 6360 4360
rect 3400 4080 3460 4240
rect 3680 4080 3740 4240
rect 3980 4080 4040 4240
rect 4280 4080 4340 4240
rect 4560 4080 4620 4240
rect 4860 4080 4920 4240
rect 5160 4080 5220 4240
rect 5460 4080 5520 4240
rect 5780 4080 5840 4240
rect 6060 4080 6120 4240
rect 6360 4080 6420 4240
rect 3540 3560 3600 3720
rect 3840 3560 3900 3720
rect 4140 3560 4200 3720
rect 4420 3560 4480 3720
rect 4720 3560 4780 3720
rect 5020 3560 5080 3720
rect 5320 3560 5380 3720
rect 5620 3560 5680 3720
rect 5920 3560 5980 3720
rect 6200 3560 6260 3720
rect 3400 3300 3460 3460
rect 3680 3300 3740 3460
rect 4000 3300 4060 3460
rect 4280 3300 4340 3460
rect 4580 3300 4640 3460
rect 4860 3300 4920 3460
rect 5160 3300 5220 3460
rect 5460 3300 5520 3460
rect 5760 3300 5820 3460
rect 6060 3300 6120 3460
rect 6360 3300 6420 3460
rect 3460 3100 6360 3160
rect 6750 4300 9650 4360
rect 6700 4080 6760 4240
rect 6980 4080 7040 4240
rect 7280 4080 7340 4240
rect 7580 4080 7640 4240
rect 7880 4080 7940 4240
rect 8160 4080 8220 4240
rect 8460 4080 8520 4240
rect 8760 4080 8820 4240
rect 9060 4080 9120 4240
rect 9340 4080 9400 4240
rect 9640 4080 9700 4240
rect 6840 3560 6900 3720
rect 7140 3560 7200 3720
rect 7440 3560 7500 3720
rect 7720 3560 7780 3720
rect 8020 3560 8080 3720
rect 8320 3560 8380 3720
rect 8620 3560 8680 3720
rect 8900 3560 8960 3720
rect 9200 3560 9260 3720
rect 9500 3560 9560 3720
rect 6680 3300 6740 3460
rect 6980 3300 7040 3460
rect 7280 3300 7340 3460
rect 7580 3300 7640 3460
rect 7880 3300 7940 3460
rect 8160 3300 8220 3460
rect 8460 3300 8520 3460
rect 8780 3300 8840 3460
rect 9060 3300 9120 3460
rect 9360 3300 9420 3460
rect 9660 3300 9720 3460
rect 6750 3100 9650 3160
rect 10040 4300 12940 4360
rect 9980 4080 10040 4240
rect 10280 4080 10340 4240
rect 10560 4080 10620 4240
rect 10860 4080 10920 4240
rect 11160 4080 11220 4240
rect 11460 4080 11520 4240
rect 11760 4080 11820 4240
rect 12060 4080 12120 4240
rect 12340 4080 12400 4240
rect 12640 4080 12700 4240
rect 12940 4080 13000 4240
rect 10140 3560 10200 3720
rect 10420 3560 10480 3720
rect 10720 3560 10780 3720
rect 11020 3560 11080 3720
rect 11320 3560 11380 3720
rect 11600 3560 11660 3720
rect 11900 3560 11960 3720
rect 12200 3560 12260 3720
rect 12500 3560 12560 3720
rect 12800 3560 12860 3720
rect 10000 3300 10060 3460
rect 10280 3300 10340 3460
rect 10580 3300 10640 3460
rect 10860 3300 10920 3460
rect 11180 3300 11240 3460
rect 11460 3300 11520 3460
rect 11760 3300 11820 3460
rect 12060 3300 12120 3460
rect 12360 3300 12420 3460
rect 12640 3300 12700 3460
rect 12940 3300 13000 3460
rect 10040 3100 12940 3160
rect 13340 4300 16240 4360
rect 13280 4080 13340 4240
rect 13560 4080 13620 4240
rect 13860 4080 13920 4240
rect 14160 4080 14220 4240
rect 14460 4080 14520 4240
rect 14760 4080 14820 4240
rect 15060 4080 15120 4240
rect 15360 4080 15420 4240
rect 15640 4080 15700 4240
rect 15940 4080 16000 4240
rect 16220 4080 16280 4240
rect 13440 3820 13500 3980
rect 13720 3820 13780 3980
rect 14020 3820 14080 3980
rect 14320 3820 14380 3980
rect 14600 3820 14660 3980
rect 14900 3820 14960 3980
rect 15200 3820 15260 3980
rect 15500 3820 15560 3980
rect 15780 3820 15840 3980
rect 16080 3820 16140 3980
rect 13280 3300 13340 3460
rect 13560 3300 13620 3460
rect 13880 3300 13940 3460
rect 14180 3300 14240 3460
rect 14460 3300 14520 3460
rect 14740 3300 14800 3460
rect 15040 3300 15100 3460
rect 15360 3300 15420 3460
rect 15640 3300 15700 3460
rect 15940 3300 16000 3460
rect 16240 3300 16300 3460
rect 13340 3100 16240 3160
rect 16400 2900 16780 3040
rect 150 2780 3050 2840
rect 100 2560 160 2720
rect 400 2560 460 2720
rect 680 2560 740 2720
rect 980 2560 1040 2720
rect 1300 2560 1360 2720
rect 1600 2560 1660 2720
rect 1880 2560 1940 2720
rect 2180 2560 2240 2720
rect 2460 2560 2520 2720
rect 2760 2560 2820 2720
rect 3060 2560 3120 2720
rect 260 2300 320 2460
rect 540 2300 600 2460
rect 840 2300 900 2460
rect 1140 2300 1200 2460
rect 1440 2300 1500 2460
rect 1740 2300 1800 2460
rect 2020 2300 2080 2460
rect 2320 2300 2380 2460
rect 2620 2300 2680 2460
rect 2900 2300 2960 2460
rect 100 1780 160 1940
rect 400 1780 460 1940
rect 680 1780 740 1940
rect 1000 1780 1060 1940
rect 1300 1780 1360 1940
rect 1600 1780 1660 1940
rect 1880 1780 1940 1940
rect 2180 1780 2240 1940
rect 2460 1780 2520 1940
rect 2760 1780 2820 1940
rect 3060 1780 3120 1940
rect 150 1570 3050 1630
rect 3450 2780 6350 2840
rect 3400 2560 3460 2720
rect 3680 2560 3740 2720
rect 3980 2560 4040 2720
rect 4280 2560 4340 2720
rect 4580 2560 4640 2720
rect 4880 2560 4940 2720
rect 5160 2560 5220 2720
rect 5460 2560 5520 2720
rect 5760 2560 5820 2720
rect 6060 2560 6120 2720
rect 6360 2560 6420 2720
rect 3540 2000 3620 2460
rect 3820 2000 3900 2460
rect 4120 2000 4200 2460
rect 4420 2000 4500 2460
rect 4720 2000 4800 2460
rect 5020 2000 5100 2460
rect 5320 2000 5400 2460
rect 5600 2000 5680 2460
rect 5900 2000 5980 2460
rect 6200 2000 6280 2460
rect 3400 1780 3460 1940
rect 3680 1780 3740 1940
rect 3980 1780 4040 1940
rect 4280 1780 4340 1940
rect 4580 1780 4640 1940
rect 4880 1780 4940 1940
rect 5160 1780 5220 1940
rect 5460 1780 5520 1940
rect 5780 1780 5840 1940
rect 6060 1780 6120 1940
rect 6340 1780 6400 1940
rect 3450 1570 6350 1630
rect 6740 2780 9640 2840
rect 6680 2560 6740 2720
rect 6980 2560 7040 2720
rect 7280 2560 7340 2720
rect 7580 2560 7640 2720
rect 7880 2560 7940 2720
rect 8160 2560 8220 2720
rect 8460 2560 8520 2720
rect 8760 2560 8820 2720
rect 9040 2560 9100 2720
rect 9340 2560 9400 2720
rect 9640 2560 9700 2720
rect 6840 2040 6900 2200
rect 7140 2040 7200 2200
rect 7440 2040 7500 2200
rect 7720 2040 7780 2200
rect 8020 2040 8080 2200
rect 8320 2040 8380 2200
rect 8600 2040 8660 2200
rect 8900 2040 8960 2200
rect 9200 2040 9260 2200
rect 9500 2040 9560 2200
rect 6680 1780 6740 1940
rect 7000 1780 7060 1940
rect 7280 1780 7340 1940
rect 7580 1780 7640 1940
rect 7860 1780 7920 1940
rect 8180 1780 8240 1940
rect 8460 1780 8520 1940
rect 8760 1780 8820 1940
rect 9060 1780 9120 1940
rect 9340 1780 9400 1940
rect 9640 1780 9700 1940
rect 6740 1570 9640 1630
rect 10030 2780 12930 2840
rect 9980 2560 10040 2720
rect 10280 2560 10340 2720
rect 10560 2560 10620 2720
rect 10860 2560 10920 2720
rect 11160 2560 11220 2720
rect 11460 2560 11520 2720
rect 11760 2560 11820 2720
rect 12040 2560 12100 2720
rect 12340 2560 12400 2720
rect 12640 2560 12700 2720
rect 12940 2560 13000 2720
rect 10140 2300 10200 2460
rect 10420 2300 10480 2460
rect 10720 2300 10780 2460
rect 11020 2300 11080 2460
rect 11320 2300 11380 2460
rect 11600 2300 11660 2460
rect 11920 2300 11980 2460
rect 12200 2300 12260 2460
rect 12500 2300 12560 2460
rect 12800 2300 12860 2460
rect 10000 1780 10060 1940
rect 10280 1780 10340 1940
rect 10580 1780 10640 1940
rect 10880 1780 10940 1940
rect 11160 1780 11220 1940
rect 11460 1780 11520 1940
rect 11760 1780 11820 1940
rect 12060 1780 12120 1940
rect 12360 1780 12420 1940
rect 12640 1780 12700 1940
rect 12940 1780 13000 1940
rect 10030 1570 12930 1630
rect 13330 2780 16230 2840
rect 13280 2560 13340 2720
rect 13580 2560 13640 2720
rect 13860 2560 13920 2720
rect 14160 2560 14220 2720
rect 14460 2560 14520 2720
rect 14760 2560 14820 2720
rect 15060 2560 15120 2720
rect 15340 2560 15400 2720
rect 15640 2560 15700 2720
rect 15940 2560 16000 2720
rect 16240 2560 16300 2720
rect 13440 2300 13500 2460
rect 13720 2300 13780 2460
rect 14020 2300 14080 2460
rect 14320 2300 14380 2460
rect 14620 2300 14680 2460
rect 14900 2300 14960 2460
rect 15200 2300 15260 2460
rect 15500 2300 15560 2460
rect 15800 2300 15860 2460
rect 16100 2300 16160 2460
rect 13280 1780 13340 1940
rect 13560 1780 13620 1940
rect 13880 1780 13940 1940
rect 14160 1780 14220 1940
rect 14460 1780 14520 1940
rect 14760 1780 14820 1940
rect 15060 1780 15120 1940
rect 15340 1780 15400 1940
rect 15640 1780 15700 1940
rect 15940 1780 16000 1940
rect 16240 1780 16300 1940
rect 13330 1570 16230 1630
rect 16400 1380 16780 1520
rect 150 1270 3050 1330
rect 100 1030 160 1210
rect 400 1030 460 1210
rect 700 1030 760 1210
rect 1000 1030 1060 1210
rect 1280 1030 1340 1210
rect 1580 1030 1640 1210
rect 1880 1030 1940 1210
rect 2180 1030 2240 1210
rect 2480 1030 2540 1210
rect 2760 1030 2820 1210
rect 3060 1030 3120 1210
rect 240 770 300 950
rect 540 770 600 950
rect 840 770 900 950
rect 1140 770 1200 950
rect 1440 770 1500 950
rect 1740 770 1800 950
rect 2020 770 2080 950
rect 2320 770 2380 950
rect 2620 770 2680 950
rect 2920 770 2980 950
rect 120 510 180 690
rect 400 510 460 690
rect 680 510 740 690
rect 980 510 1040 690
rect 1300 510 1360 690
rect 1600 510 1660 690
rect 1880 510 1940 690
rect 2160 510 2220 690
rect 2480 510 2540 690
rect 2760 510 2820 690
rect 3060 510 3120 690
rect 240 250 300 430
rect 540 250 600 430
rect 840 250 900 430
rect 1140 250 1200 430
rect 1440 250 1500 430
rect 1740 250 1800 430
rect 2020 250 2080 430
rect 2340 250 2400 430
rect 2620 250 2680 430
rect 2920 250 2980 430
rect 150 60 3050 120
rect 3450 1270 6350 1330
rect 3400 1030 3460 1210
rect 3680 1030 3740 1210
rect 4000 1030 4060 1210
rect 4280 1030 4340 1210
rect 4580 1030 4640 1210
rect 4880 1030 4940 1210
rect 5160 1030 5220 1210
rect 5460 1030 5520 1210
rect 5760 1030 5820 1210
rect 6060 1030 6120 1210
rect 6360 1030 6420 1210
rect 3540 770 3600 950
rect 3840 770 3900 950
rect 4140 770 4200 950
rect 4440 770 4500 950
rect 4720 770 4780 950
rect 5020 770 5080 950
rect 5320 770 5380 950
rect 5620 770 5680 950
rect 5900 770 5960 950
rect 6220 770 6280 950
rect 3400 510 3460 690
rect 3700 510 3760 690
rect 4000 510 4060 690
rect 4280 510 4340 690
rect 4580 510 4640 690
rect 4880 510 4940 690
rect 5180 510 5240 690
rect 5460 510 5520 690
rect 5760 510 5820 690
rect 6060 510 6120 690
rect 6360 510 6420 690
rect 3540 250 3600 430
rect 3840 250 3900 430
rect 4140 250 4200 430
rect 4440 250 4500 430
rect 4720 250 4780 430
rect 5020 250 5080 430
rect 5320 250 5380 430
rect 5620 250 5680 430
rect 5900 250 5960 430
rect 6220 250 6280 430
rect 3450 60 6350 120
rect 6740 1270 9640 1330
rect 6700 1030 6760 1210
rect 6980 1030 7040 1210
rect 7280 1030 7340 1210
rect 7580 1030 7640 1210
rect 7880 1030 7940 1210
rect 8180 1030 8240 1210
rect 8460 1030 8520 1210
rect 8760 1030 8820 1210
rect 9060 1030 9120 1210
rect 9360 1030 9420 1210
rect 9640 1030 9700 1210
rect 6840 770 6900 950
rect 7140 770 7200 950
rect 7420 770 7480 950
rect 7720 770 7780 950
rect 8020 770 8080 950
rect 8300 770 8360 950
rect 8620 770 8680 950
rect 8920 770 8980 950
rect 9220 770 9280 950
rect 9520 770 9580 950
rect 6700 510 6760 690
rect 7000 510 7060 690
rect 7280 510 7340 690
rect 7580 510 7640 690
rect 7860 510 7920 690
rect 8180 510 8240 690
rect 8480 510 8540 690
rect 8760 510 8820 690
rect 9060 510 9120 690
rect 9360 510 9420 690
rect 9660 510 9720 690
rect 6840 250 6900 430
rect 7140 250 7200 430
rect 7440 250 7500 430
rect 7720 250 7780 430
rect 8020 250 8080 430
rect 8320 250 8380 430
rect 8620 250 8680 430
rect 8920 250 8980 430
rect 9200 250 9260 430
rect 9520 250 9580 430
rect 6740 60 9640 120
rect 10030 1270 12930 1330
rect 9980 1030 10040 1210
rect 10280 1030 10340 1210
rect 10560 1030 10620 1210
rect 10860 1030 10920 1210
rect 11160 1030 11220 1210
rect 11460 1030 11520 1210
rect 11760 1030 11820 1210
rect 12060 1030 12120 1210
rect 12360 1030 12420 1210
rect 12660 1030 12720 1210
rect 12940 1030 13000 1210
rect 10140 770 10200 950
rect 10420 770 10480 950
rect 10740 770 10800 950
rect 11020 770 11080 950
rect 11320 770 11380 950
rect 11620 770 11680 950
rect 11920 770 11980 950
rect 12220 770 12280 950
rect 12500 770 12560 950
rect 12800 770 12860 950
rect 10000 510 10060 690
rect 10280 510 10340 690
rect 10580 510 10640 690
rect 10860 510 10920 690
rect 11160 510 11220 690
rect 11480 510 11540 690
rect 11760 510 11820 690
rect 12060 510 12120 690
rect 12360 510 12420 690
rect 12660 510 12720 690
rect 12940 510 13000 690
rect 10140 250 10200 430
rect 10440 250 10500 430
rect 10740 250 10800 430
rect 11020 250 11080 430
rect 11300 250 11360 430
rect 11600 250 11660 430
rect 11900 250 11960 430
rect 12220 250 12280 430
rect 12500 250 12560 430
rect 12800 250 12860 430
rect 10030 60 12930 120
rect 13330 1270 16230 1330
rect 13280 1030 13340 1210
rect 13580 1030 13640 1210
rect 13880 1030 13940 1210
rect 14180 1030 14240 1210
rect 14460 1030 14520 1210
rect 14760 1030 14820 1210
rect 15060 1030 15120 1210
rect 15360 1030 15420 1210
rect 15640 1030 15700 1210
rect 15960 1030 16020 1210
rect 16240 1030 16300 1210
rect 13420 770 13480 950
rect 13740 770 13800 950
rect 14020 770 14080 950
rect 14300 770 14360 950
rect 14620 770 14680 950
rect 14920 770 14980 950
rect 15200 770 15260 950
rect 15500 770 15560 950
rect 15780 770 15840 950
rect 16100 770 16160 950
rect 13280 510 13340 690
rect 13580 510 13640 690
rect 13880 510 13940 690
rect 14160 510 14220 690
rect 14460 510 14520 690
rect 14760 510 14820 690
rect 15060 510 15120 690
rect 15360 510 15420 690
rect 15640 510 15700 690
rect 15940 510 16000 690
rect 16240 510 16300 690
rect 13440 250 13500 430
rect 13740 250 13800 430
rect 14020 250 14080 430
rect 14320 250 14380 430
rect 14600 250 14660 430
rect 14900 250 14960 430
rect 15200 250 15260 430
rect 15500 250 15560 430
rect 15780 250 15840 430
rect 16100 250 16160 430
rect 13330 60 16230 120
<< metal2 >>
rect 160 8920 3060 8930
rect 3180 8920 3340 9020
rect 3460 8920 6360 8930
rect 6480 8920 6620 9030
rect 6750 8920 9650 8930
rect 9780 8920 9920 9030
rect 10040 8920 12940 8930
rect 13060 8920 13200 9030
rect 13340 8920 16240 8930
rect 3060 8860 3460 8920
rect 6360 8860 6750 8920
rect 9650 8860 10040 8920
rect 12940 8860 13340 8920
rect 160 8850 3060 8860
rect 100 8790 160 8800
rect 100 8600 160 8610
rect 400 8790 460 8800
rect 400 8600 460 8610
rect 690 8790 750 8800
rect 690 8600 750 8610
rect 990 8790 1050 8800
rect 990 8600 1050 8610
rect 1290 8790 1350 8800
rect 1290 8600 1350 8610
rect 1590 8790 1650 8800
rect 1590 8600 1650 8610
rect 1880 8790 1940 8800
rect 1880 8600 1940 8610
rect 2170 8790 2230 8800
rect 2170 8600 2230 8610
rect 2470 8790 2530 8800
rect 2470 8600 2530 8610
rect 2760 8790 2820 8800
rect 2760 8600 2820 8610
rect 3060 8790 3120 8800
rect 3060 8600 3120 8610
rect 250 8530 310 8540
rect 250 8340 310 8350
rect 550 8530 610 8540
rect 550 8340 610 8350
rect 840 8530 900 8540
rect 840 8340 900 8350
rect 1140 8530 1200 8540
rect 1140 8340 1200 8350
rect 1440 8530 1500 8540
rect 1440 8340 1500 8350
rect 1730 8530 1790 8540
rect 1730 8340 1790 8350
rect 2030 8530 2090 8540
rect 2030 8340 2090 8350
rect 2320 8530 2380 8540
rect 2320 8340 2380 8350
rect 2620 8530 2680 8540
rect 2620 8340 2680 8350
rect 2920 8530 2980 8540
rect 2920 8340 2980 8350
rect 100 8270 160 8280
rect 100 8080 160 8090
rect 400 8270 460 8280
rect 400 8080 460 8090
rect 690 8270 750 8280
rect 690 8080 750 8090
rect 990 8270 1050 8280
rect 990 8080 1050 8090
rect 1290 8270 1350 8280
rect 1290 8080 1350 8090
rect 1590 8270 1650 8280
rect 1590 8080 1650 8090
rect 1880 8270 1940 8280
rect 1880 8080 1940 8090
rect 2170 8270 2230 8280
rect 2170 8080 2230 8090
rect 2470 8270 2530 8280
rect 2470 8080 2530 8090
rect 2770 8270 2830 8280
rect 2770 8080 2830 8090
rect 3060 8270 3120 8280
rect 3060 8080 3120 8090
rect 250 8010 310 8020
rect 250 7820 310 7830
rect 540 8010 600 8020
rect 540 7820 600 7830
rect 840 8010 900 8020
rect 840 7820 900 7830
rect 1130 8010 1190 8020
rect 1130 7820 1190 7830
rect 1430 8010 1490 8020
rect 1430 7820 1490 7830
rect 1730 8010 1790 8020
rect 1730 7820 1790 7830
rect 2030 8010 2090 8020
rect 2030 7820 2090 7830
rect 2330 8010 2390 8020
rect 2330 7820 2390 7830
rect 2620 8010 2680 8020
rect 2620 7820 2680 7830
rect 2920 8010 2980 8020
rect 2920 7820 2980 7830
rect 160 7710 3060 7720
rect 3180 7710 3340 8860
rect 3460 8850 6360 8860
rect 3400 8800 3460 8810
rect 3400 8610 3460 8620
rect 3680 8800 3740 8810
rect 3680 8610 3740 8620
rect 3980 8800 4040 8810
rect 3980 8610 4040 8620
rect 4280 8800 4340 8810
rect 4280 8610 4340 8620
rect 4580 8800 4640 8810
rect 4580 8610 4640 8620
rect 4880 8800 4940 8810
rect 4880 8610 4940 8620
rect 5160 8800 5220 8810
rect 5160 8610 5220 8620
rect 5460 8800 5520 8810
rect 5460 8610 5520 8620
rect 5760 8800 5820 8810
rect 5760 8610 5820 8620
rect 6060 8800 6120 8810
rect 6060 8610 6120 8620
rect 6340 8800 6400 8810
rect 6340 8610 6400 8620
rect 3540 8520 3600 8530
rect 3540 8350 3600 8360
rect 3840 8520 3900 8530
rect 3840 8350 3900 8360
rect 4140 8520 4200 8530
rect 4140 8350 4200 8360
rect 4440 8520 4500 8530
rect 4440 8350 4500 8360
rect 4720 8520 4780 8530
rect 4720 8350 4780 8360
rect 5020 8520 5080 8530
rect 5020 8350 5080 8360
rect 5320 8520 5380 8530
rect 5320 8350 5380 8360
rect 5600 8520 5660 8530
rect 5600 8350 5660 8360
rect 5920 8520 5980 8530
rect 5920 8350 5980 8360
rect 6200 8520 6260 8530
rect 6200 8350 6260 8360
rect 3400 8260 3460 8270
rect 3400 8090 3460 8100
rect 3700 8260 3760 8270
rect 3700 8090 3760 8100
rect 3980 8260 4040 8270
rect 3980 8090 4040 8100
rect 4280 8260 4340 8270
rect 4280 8090 4340 8100
rect 4560 8260 4620 8270
rect 4560 8090 4620 8100
rect 4880 8260 4940 8270
rect 4880 8090 4940 8100
rect 5160 8260 5220 8270
rect 5160 8090 5220 8100
rect 5460 8260 5520 8270
rect 5460 8090 5520 8100
rect 5760 8260 5820 8270
rect 5760 8090 5820 8100
rect 6060 8260 6120 8270
rect 6060 8090 6120 8100
rect 6360 8260 6420 8270
rect 6360 8090 6420 8100
rect 3540 8000 3600 8010
rect 3540 7830 3600 7840
rect 3840 8000 3900 8010
rect 3840 7830 3900 7840
rect 4140 8000 4200 8010
rect 4140 7830 4200 7840
rect 4420 8000 4480 8010
rect 4420 7830 4480 7840
rect 4720 8000 4780 8010
rect 4720 7830 4780 7840
rect 5020 8000 5080 8010
rect 5020 7830 5080 7840
rect 5320 8000 5380 8010
rect 5320 7830 5380 7840
rect 5620 8000 5680 8010
rect 5620 7830 5680 7840
rect 5920 8000 5980 8010
rect 5920 7830 5980 7840
rect 6200 8000 6260 8010
rect 6200 7830 6260 7840
rect 3460 7710 6360 7720
rect 6480 7710 6620 8860
rect 6750 8850 9650 8860
rect 6680 8800 6740 8810
rect 6680 8630 6740 8640
rect 6980 8800 7040 8810
rect 6980 8630 7040 8640
rect 7280 8800 7340 8810
rect 7280 8630 7340 8640
rect 7580 8800 7640 8810
rect 7580 8630 7640 8640
rect 7880 8800 7940 8810
rect 7880 8630 7940 8640
rect 8160 8800 8220 8810
rect 8160 8630 8220 8640
rect 8460 8780 8520 8790
rect 8460 8610 8520 8620
rect 8760 8780 8820 8790
rect 8760 8610 8820 8620
rect 9040 8780 9100 8790
rect 9040 8610 9100 8620
rect 9340 8780 9400 8790
rect 9340 8610 9400 8620
rect 9640 8780 9700 8790
rect 9640 8610 9700 8620
rect 6820 8520 6880 8530
rect 6820 8350 6880 8360
rect 7120 8520 7180 8530
rect 7120 8350 7180 8360
rect 7420 8520 7480 8530
rect 7420 8350 7480 8360
rect 7720 8520 7780 8530
rect 7720 8350 7780 8360
rect 8020 8520 8080 8530
rect 8020 8350 8080 8360
rect 8320 8520 8380 8530
rect 8320 8350 8380 8360
rect 8620 8520 8680 8530
rect 8620 8350 8680 8360
rect 8920 8520 8980 8530
rect 8920 8350 8980 8360
rect 9200 8520 9260 8530
rect 9200 8350 9260 8360
rect 9500 8520 9560 8530
rect 9500 8350 9560 8360
rect 6680 8260 6740 8270
rect 6680 8090 6740 8100
rect 6980 8260 7040 8270
rect 6980 8090 7040 8100
rect 7280 8260 7340 8270
rect 7280 8090 7340 8100
rect 7580 8260 7640 8270
rect 7580 8090 7640 8100
rect 7860 8260 7920 8270
rect 7860 8090 7920 8100
rect 8160 8260 8220 8270
rect 8160 8090 8220 8100
rect 8460 8260 8520 8270
rect 8460 8090 8520 8100
rect 8760 8260 8820 8270
rect 8760 8090 8820 8100
rect 9060 8260 9120 8270
rect 9060 8090 9120 8100
rect 9340 8260 9400 8270
rect 9340 8090 9400 8100
rect 9640 8260 9700 8270
rect 9640 8090 9700 8100
rect 6840 8000 6900 8010
rect 6840 7830 6900 7840
rect 7140 8000 7200 8010
rect 7140 7830 7200 7840
rect 7420 8000 7480 8010
rect 7420 7830 7480 7840
rect 7720 8000 7780 8010
rect 7720 7830 7780 7840
rect 8020 8000 8080 8010
rect 8020 7830 8080 7840
rect 8300 8000 8360 8010
rect 8300 7830 8360 7840
rect 8620 8000 8680 8010
rect 8620 7830 8680 7840
rect 8900 8000 8960 8010
rect 8900 7830 8960 7840
rect 9200 8000 9260 8010
rect 9200 7830 9260 7840
rect 9500 8000 9560 8010
rect 9500 7830 9560 7840
rect 6750 7710 9650 7720
rect 9780 7710 9920 8860
rect 10040 8850 12940 8860
rect 9980 8800 10040 8810
rect 9980 8630 10040 8640
rect 10280 8800 10340 8810
rect 10280 8630 10340 8640
rect 10580 8800 10640 8810
rect 10580 8630 10640 8640
rect 10880 8800 10940 8810
rect 10880 8630 10940 8640
rect 11160 8780 11220 8790
rect 11160 8610 11220 8620
rect 11460 8780 11520 8790
rect 11460 8610 11520 8620
rect 11760 8780 11820 8790
rect 11760 8610 11820 8620
rect 12040 8780 12100 8790
rect 12040 8610 12100 8620
rect 12360 8780 12420 8790
rect 12360 8610 12420 8620
rect 12640 8780 12700 8790
rect 12640 8610 12700 8620
rect 12940 8780 13000 8790
rect 12940 8610 13000 8620
rect 10140 8520 10200 8530
rect 10140 8350 10200 8360
rect 10420 8520 10480 8530
rect 10420 8350 10480 8360
rect 10720 8520 10780 8530
rect 10720 8350 10780 8360
rect 11020 8520 11080 8530
rect 11020 8350 11080 8360
rect 11320 8520 11380 8530
rect 11320 8350 11380 8360
rect 11600 8520 11660 8530
rect 11600 8350 11660 8360
rect 11900 8520 11960 8530
rect 11900 8350 11960 8360
rect 12200 8520 12260 8530
rect 12200 8350 12260 8360
rect 12500 8520 12560 8530
rect 12500 8350 12560 8360
rect 12800 8520 12860 8530
rect 12800 8350 12860 8360
rect 9980 8260 10040 8270
rect 9980 8090 10040 8100
rect 10280 8260 10340 8270
rect 10280 8090 10340 8100
rect 10580 8260 10640 8270
rect 10580 8090 10640 8100
rect 10860 8260 10920 8270
rect 10860 8090 10920 8100
rect 11180 8260 11240 8270
rect 11180 8090 11240 8100
rect 11460 8260 11520 8270
rect 11460 8090 11520 8100
rect 11760 8260 11820 8270
rect 11760 8090 11820 8100
rect 12060 8260 12120 8270
rect 12060 8090 12120 8100
rect 12340 8260 12400 8270
rect 12340 8090 12400 8100
rect 12640 8260 12700 8270
rect 12640 8090 12700 8100
rect 12940 8260 13000 8270
rect 12940 8090 13000 8100
rect 10140 8000 10200 8010
rect 10140 7830 10200 7840
rect 10440 8000 10500 8010
rect 10440 7830 10500 7840
rect 10720 8000 10780 8010
rect 10720 7830 10780 7840
rect 11020 8000 11080 8010
rect 11020 7830 11080 7840
rect 11320 8000 11380 8010
rect 11320 7830 11380 7840
rect 11600 8000 11660 8010
rect 11600 7830 11660 7840
rect 11900 8000 11960 8010
rect 11900 7830 11960 7840
rect 12200 8000 12260 8010
rect 12200 7830 12260 7840
rect 12500 8000 12560 8010
rect 12500 7830 12560 7840
rect 12800 8000 12860 8010
rect 12800 7830 12860 7840
rect 10040 7710 12940 7720
rect 13060 7710 13200 8860
rect 13340 8850 16240 8860
rect 13280 8780 13340 8790
rect 13280 8610 13340 8620
rect 13580 8780 13640 8790
rect 13580 8610 13640 8620
rect 13860 8780 13920 8790
rect 13860 8610 13920 8620
rect 14180 8780 14240 8790
rect 14180 8610 14240 8620
rect 14460 8780 14520 8790
rect 14460 8610 14520 8620
rect 14760 8780 14820 8790
rect 14760 8610 14820 8620
rect 15040 8780 15100 8790
rect 15040 8610 15100 8620
rect 15340 8780 15400 8790
rect 15340 8610 15400 8620
rect 15640 8780 15700 8790
rect 15640 8610 15700 8620
rect 15940 8780 16000 8790
rect 15940 8610 16000 8620
rect 16240 8780 16300 8790
rect 16240 8610 16300 8620
rect 16400 8780 16800 8800
rect 16400 8620 16420 8780
rect 16780 8620 16800 8780
rect 13420 8520 13480 8530
rect 13420 8350 13480 8360
rect 13720 8520 13780 8530
rect 13720 8350 13780 8360
rect 14000 8520 14060 8530
rect 14000 8350 14060 8360
rect 14320 8520 14380 8530
rect 14320 8350 14380 8360
rect 14600 8520 14660 8530
rect 14600 8350 14660 8360
rect 14900 8520 14960 8530
rect 14900 8350 14960 8360
rect 15200 8520 15260 8530
rect 15200 8350 15260 8360
rect 15500 8520 15560 8530
rect 15500 8350 15560 8360
rect 15780 8520 15840 8530
rect 15780 8350 15840 8360
rect 16080 8520 16140 8530
rect 16080 8350 16140 8360
rect 13280 8260 13340 8270
rect 13280 8090 13340 8100
rect 13580 8260 13640 8270
rect 13580 8090 13640 8100
rect 13860 8260 13920 8270
rect 13860 8090 13920 8100
rect 14180 8260 14240 8270
rect 14180 8090 14240 8100
rect 14460 8260 14520 8270
rect 14460 8090 14520 8100
rect 14760 8260 14820 8270
rect 14760 8090 14820 8100
rect 15060 8260 15120 8270
rect 15060 8090 15120 8100
rect 15360 8260 15420 8270
rect 15360 8090 15420 8100
rect 15640 8260 15700 8270
rect 15640 8090 15700 8100
rect 15940 8260 16000 8270
rect 15940 8090 16000 8100
rect 16240 8260 16300 8270
rect 16240 8090 16300 8100
rect 16400 8260 16800 8620
rect 16400 8100 16420 8260
rect 16780 8100 16800 8260
rect 13420 8000 13480 8010
rect 13420 7830 13480 7840
rect 13720 8000 13780 8010
rect 13720 7830 13780 7840
rect 14020 8000 14080 8010
rect 14020 7830 14080 7840
rect 14320 8000 14380 8010
rect 14320 7830 14380 7840
rect 14600 8000 14660 8010
rect 14600 7830 14660 7840
rect 14900 8000 14960 8010
rect 14900 7830 14960 7840
rect 15200 8000 15260 8010
rect 15200 7830 15260 7840
rect 15500 8000 15560 8010
rect 15500 7830 15560 7840
rect 15800 8000 15860 8010
rect 15800 7830 15860 7840
rect 16080 8000 16140 8010
rect 16080 7830 16140 7840
rect 13340 7710 16240 7720
rect 3060 7650 3460 7710
rect 6360 7650 6750 7710
rect 9650 7650 10040 7710
rect 12940 7650 13340 7710
rect 160 7640 3060 7650
rect 160 7400 3060 7410
rect 3180 7400 3340 7650
rect 3460 7640 6360 7650
rect 3460 7400 6360 7410
rect 6480 7400 6620 7650
rect 6750 7640 9650 7650
rect 6750 7400 9650 7410
rect 9780 7400 9920 7650
rect 10040 7640 12940 7650
rect 10040 7400 12940 7410
rect 13060 7400 13200 7650
rect 13340 7640 16240 7650
rect 16400 7600 16800 8100
rect 16780 7460 16800 7600
rect 13340 7400 16240 7410
rect 3060 7340 3460 7400
rect 6360 7340 6750 7400
rect 9650 7340 10040 7400
rect 12940 7340 13340 7400
rect 160 7330 3060 7340
rect 100 7280 160 7290
rect 100 7110 160 7120
rect 400 7280 460 7290
rect 400 7110 460 7120
rect 700 7280 760 7290
rect 700 7110 760 7120
rect 980 7280 1040 7290
rect 980 7110 1040 7120
rect 1280 7280 1340 7290
rect 1280 7110 1340 7120
rect 1580 7280 1640 7290
rect 1580 7110 1640 7120
rect 1880 7280 1940 7290
rect 1880 7110 1940 7120
rect 2180 7280 2240 7290
rect 2180 7110 2240 7120
rect 2460 7280 2520 7290
rect 2460 7110 2520 7120
rect 2780 7280 2840 7290
rect 2780 7110 2840 7120
rect 3060 7280 3120 7290
rect 3060 7110 3120 7120
rect 260 7020 320 7030
rect 260 6850 320 6860
rect 560 7020 620 7030
rect 560 6850 620 6860
rect 840 7020 900 7030
rect 840 6850 900 6860
rect 1140 7020 1200 7030
rect 1140 6850 1200 6860
rect 1420 7020 1480 7030
rect 1420 6850 1480 6860
rect 1720 7020 1780 7030
rect 1720 6850 1780 6860
rect 2040 7020 2100 7030
rect 2040 6850 2100 6860
rect 2320 7020 2380 7030
rect 2320 6850 2380 6860
rect 2620 7020 2680 7030
rect 2620 6850 2680 6860
rect 2900 7020 2960 7030
rect 2900 6850 2960 6860
rect 100 6500 160 6510
rect 100 6330 160 6340
rect 380 6500 440 6510
rect 380 6330 440 6340
rect 700 6500 760 6510
rect 700 6330 760 6340
rect 1000 6500 1060 6510
rect 1000 6330 1060 6340
rect 1280 6500 1340 6510
rect 1280 6330 1340 6340
rect 1580 6500 1640 6510
rect 1580 6330 1640 6340
rect 1880 6500 1940 6510
rect 1880 6330 1940 6340
rect 2180 6500 2240 6510
rect 2180 6330 2240 6340
rect 2480 6500 2540 6510
rect 2480 6330 2540 6340
rect 2760 6500 2820 6510
rect 2760 6330 2820 6340
rect 3060 6500 3120 6510
rect 3060 6330 3120 6340
rect 160 6190 3060 6200
rect 3180 6190 3340 7340
rect 3460 7330 6360 7340
rect 3400 7280 3460 7290
rect 3400 7110 3460 7120
rect 3680 7280 3740 7290
rect 3680 7110 3740 7120
rect 3980 7280 4040 7290
rect 3980 7110 4040 7120
rect 4280 7280 4340 7290
rect 4280 7110 4340 7120
rect 4580 7280 4640 7290
rect 4580 7110 4640 7120
rect 4880 7280 4940 7290
rect 4880 7110 4940 7120
rect 5180 7280 5240 7290
rect 5180 7110 5240 7120
rect 5460 7280 5520 7290
rect 5460 7110 5520 7120
rect 5760 7280 5820 7290
rect 5760 7110 5820 7120
rect 6060 7280 6120 7290
rect 6060 7110 6120 7120
rect 6360 7280 6420 7290
rect 6360 7110 6420 7120
rect 3540 7020 3600 7030
rect 3540 6850 3600 6860
rect 3840 7020 3900 7030
rect 3840 6850 3900 6860
rect 4120 7020 4180 7030
rect 4120 6850 4180 6860
rect 4420 7020 4480 7030
rect 4420 6850 4480 6860
rect 4720 7020 4780 7030
rect 4720 6850 4780 6860
rect 5020 7020 5080 7030
rect 5020 6850 5080 6860
rect 5320 7020 5380 7030
rect 5320 6850 5380 6860
rect 5620 7020 5680 7030
rect 5620 6850 5680 6860
rect 5900 7020 5960 7030
rect 5900 6850 5960 6860
rect 6220 7020 6280 7030
rect 6220 6850 6280 6860
rect 3400 6500 3460 6510
rect 3400 6330 3460 6340
rect 3680 6500 3740 6510
rect 3680 6330 3740 6340
rect 3980 6500 4040 6510
rect 3980 6330 4040 6340
rect 4280 6500 4340 6510
rect 4280 6330 4340 6340
rect 4580 6500 4640 6510
rect 4580 6330 4640 6340
rect 4880 6500 4940 6510
rect 4880 6330 4940 6340
rect 5160 6500 5220 6510
rect 5160 6330 5220 6340
rect 5460 6500 5520 6510
rect 5460 6330 5520 6340
rect 5760 6500 5820 6510
rect 5760 6330 5820 6340
rect 6060 6500 6120 6510
rect 6060 6330 6120 6340
rect 6360 6500 6420 6510
rect 6360 6330 6420 6340
rect 3460 6190 6360 6200
rect 6480 6190 6620 7340
rect 6750 7330 9650 7340
rect 6680 7280 6740 7290
rect 6680 7110 6740 7120
rect 6980 7280 7040 7290
rect 6980 7110 7040 7120
rect 7280 7280 7340 7290
rect 7280 7110 7340 7120
rect 7580 7280 7640 7290
rect 7580 7110 7640 7120
rect 7880 7280 7940 7290
rect 7880 7110 7940 7120
rect 8160 7280 8220 7290
rect 8160 7110 8220 7120
rect 8460 7280 8520 7290
rect 8460 7110 8520 7120
rect 8760 7280 8820 7290
rect 8760 7110 8820 7120
rect 9060 7280 9120 7290
rect 9060 7110 9120 7120
rect 9340 7280 9400 7290
rect 9340 7110 9400 7120
rect 9640 7280 9700 7290
rect 9640 7110 9700 7120
rect 6840 6760 6900 6770
rect 6840 6590 6900 6600
rect 7140 6760 7200 6770
rect 7140 6590 7200 6600
rect 7420 6760 7480 6770
rect 7420 6590 7480 6600
rect 7720 6760 7780 6770
rect 7720 6590 7780 6600
rect 8020 6760 8080 6770
rect 8020 6590 8080 6600
rect 8320 6760 8380 6770
rect 8320 6590 8380 6600
rect 8620 6760 8680 6770
rect 8620 6590 8680 6600
rect 8920 6760 8980 6770
rect 8920 6590 8980 6600
rect 9200 6760 9260 6770
rect 9200 6590 9260 6600
rect 9500 6760 9560 6770
rect 9500 6590 9560 6600
rect 6680 6500 6740 6510
rect 6680 6330 6740 6340
rect 6980 6500 7040 6510
rect 6980 6330 7040 6340
rect 7280 6500 7340 6510
rect 7280 6330 7340 6340
rect 7580 6500 7640 6510
rect 7580 6330 7640 6340
rect 7880 6500 7940 6510
rect 7880 6330 7940 6340
rect 8180 6500 8240 6510
rect 8180 6330 8240 6340
rect 8460 6500 8520 6510
rect 8460 6330 8520 6340
rect 8760 6500 8820 6510
rect 8760 6330 8820 6340
rect 9060 6500 9120 6510
rect 9060 6330 9120 6340
rect 9360 6500 9420 6510
rect 9360 6330 9420 6340
rect 9640 6500 9700 6510
rect 9640 6330 9700 6340
rect 6750 6190 9650 6200
rect 9780 6190 9920 7340
rect 10040 7330 12940 7340
rect 9980 7280 10040 7290
rect 9980 7110 10040 7120
rect 10280 7280 10340 7290
rect 10280 7110 10340 7120
rect 10580 7280 10640 7290
rect 10580 7110 10640 7120
rect 10880 7280 10940 7290
rect 10880 7110 10940 7120
rect 11160 7280 11220 7290
rect 11160 7110 11220 7120
rect 11460 7280 11520 7290
rect 11460 7110 11520 7120
rect 11760 7280 11820 7290
rect 11760 7110 11820 7120
rect 12060 7280 12120 7290
rect 12060 7110 12120 7120
rect 12340 7280 12400 7290
rect 12340 7110 12400 7120
rect 12660 7280 12720 7290
rect 12660 7110 12720 7120
rect 12940 7280 13000 7290
rect 12940 7110 13000 7120
rect 10140 7020 10200 7030
rect 10140 6850 10200 6860
rect 10420 7020 10480 7030
rect 10420 6850 10480 6860
rect 10720 7020 10780 7030
rect 10720 6850 10780 6860
rect 11020 7020 11080 7030
rect 11020 6850 11080 6860
rect 11320 7020 11380 7030
rect 11320 6850 11380 6860
rect 11620 7020 11680 7030
rect 11620 6850 11680 6860
rect 11920 7020 11980 7030
rect 11920 6850 11980 6860
rect 12200 7020 12260 7030
rect 12200 6850 12260 6860
rect 12500 7020 12560 7030
rect 12500 6850 12560 6860
rect 12800 7020 12860 7030
rect 12800 6850 12860 6860
rect 10000 6500 10060 6510
rect 10000 6330 10060 6340
rect 10280 6500 10340 6510
rect 10280 6330 10340 6340
rect 10560 6500 10620 6510
rect 10560 6330 10620 6340
rect 10860 6500 10920 6510
rect 10860 6330 10920 6340
rect 11160 6500 11220 6510
rect 11160 6330 11220 6340
rect 11460 6500 11520 6510
rect 11460 6330 11520 6340
rect 11760 6500 11820 6510
rect 11760 6330 11820 6340
rect 12060 6500 12120 6510
rect 12060 6330 12120 6340
rect 12340 6500 12400 6510
rect 12340 6330 12400 6340
rect 12640 6500 12700 6510
rect 12640 6330 12700 6340
rect 12940 6500 13000 6510
rect 12940 6330 13000 6340
rect 10040 6190 12940 6200
rect 13060 6190 13200 7340
rect 13340 7330 16240 7340
rect 13280 7280 13340 7290
rect 13280 7110 13340 7120
rect 13560 7280 13620 7290
rect 13560 7110 13620 7120
rect 13880 7280 13940 7290
rect 13880 7110 13940 7120
rect 14160 7280 14220 7290
rect 14160 7110 14220 7120
rect 14480 7280 14540 7290
rect 14480 7110 14540 7120
rect 14760 7280 14820 7290
rect 14760 7110 14820 7120
rect 15060 7280 15120 7290
rect 15060 7110 15120 7120
rect 15340 7280 15400 7290
rect 15340 7110 15400 7120
rect 15640 7280 15700 7290
rect 15640 7110 15700 7120
rect 15940 7280 16000 7290
rect 15940 7110 16000 7120
rect 16240 7280 16300 7290
rect 16240 7110 16300 7120
rect 16400 7280 16800 7460
rect 16400 7120 16420 7280
rect 16780 7120 16800 7280
rect 13440 7020 13500 7030
rect 13440 6850 13500 6860
rect 13720 7020 13780 7030
rect 13720 6850 13780 6860
rect 14020 7020 14080 7030
rect 14020 6850 14080 6860
rect 14300 7020 14360 7030
rect 14300 6850 14360 6860
rect 14620 7020 14680 7030
rect 14620 6850 14680 6860
rect 14920 7020 14980 7030
rect 14920 6850 14980 6860
rect 15200 7020 15260 7030
rect 15200 6850 15260 6860
rect 15500 7020 15560 7030
rect 15500 6850 15560 6860
rect 15780 7020 15840 7030
rect 15780 6850 15840 6860
rect 16080 7020 16140 7030
rect 16080 6850 16140 6860
rect 13260 6500 13320 6510
rect 13260 6330 13320 6340
rect 13560 6500 13620 6510
rect 13560 6330 13620 6340
rect 13880 6500 13940 6510
rect 13880 6330 13940 6340
rect 14160 6500 14220 6510
rect 14160 6330 14220 6340
rect 14460 6500 14520 6510
rect 14460 6330 14520 6340
rect 14740 6500 14800 6510
rect 14740 6330 14800 6340
rect 15060 6500 15120 6510
rect 15060 6330 15120 6340
rect 15340 6500 15400 6510
rect 15340 6330 15400 6340
rect 15660 6500 15720 6510
rect 15660 6330 15720 6340
rect 15940 6500 16000 6510
rect 15940 6330 16000 6340
rect 16240 6500 16300 6510
rect 16240 6330 16300 6340
rect 16400 6500 16800 7120
rect 16400 6340 16420 6500
rect 16780 6340 16800 6500
rect 13340 6190 16240 6200
rect 3060 6130 3460 6190
rect 6360 6130 6750 6190
rect 9650 6130 10040 6190
rect 12940 6130 13340 6190
rect 160 6120 3060 6130
rect 160 5880 3060 5890
rect 3180 5880 3340 6130
rect 3460 6120 6360 6130
rect 3460 5880 6360 5890
rect 6480 5880 6620 6130
rect 6750 6120 9650 6130
rect 6750 5880 9650 5890
rect 9780 5880 9920 6130
rect 10040 6120 12940 6130
rect 10040 5880 12940 5890
rect 13060 5880 13200 6130
rect 13340 6120 16240 6130
rect 16400 6080 16800 6340
rect 16780 5940 16800 6080
rect 13340 5880 16240 5890
rect 3060 5820 3460 5880
rect 6360 5820 6750 5880
rect 9650 5820 10040 5880
rect 12940 5820 13340 5880
rect 160 5810 3060 5820
rect 100 5760 160 5770
rect 100 5590 160 5600
rect 400 5760 460 5770
rect 400 5590 460 5600
rect 680 5760 740 5770
rect 680 5590 740 5600
rect 1000 5760 1060 5770
rect 1000 5590 1060 5600
rect 1280 5760 1340 5770
rect 1280 5590 1340 5600
rect 1580 5760 1640 5770
rect 1580 5590 1640 5600
rect 1880 5760 1940 5770
rect 1880 5590 1940 5600
rect 2180 5760 2240 5770
rect 2180 5590 2240 5600
rect 2480 5760 2540 5770
rect 2480 5590 2540 5600
rect 2760 5760 2820 5770
rect 2760 5590 2820 5600
rect 3060 5760 3120 5770
rect 3060 5590 3120 5600
rect 260 5500 320 5510
rect 260 5330 320 5340
rect 560 5500 620 5510
rect 560 5330 620 5340
rect 840 5500 900 5510
rect 840 5330 900 5340
rect 1140 5500 1200 5510
rect 1140 5330 1200 5340
rect 1440 5500 1500 5510
rect 1440 5330 1500 5340
rect 1720 5500 1780 5510
rect 1720 5330 1780 5340
rect 2040 5500 2100 5510
rect 2040 5330 2100 5340
rect 2320 5500 2380 5510
rect 2320 5330 2380 5340
rect 2620 5500 2680 5510
rect 2620 5330 2680 5340
rect 2920 5500 2980 5510
rect 2920 5330 2980 5340
rect 3180 4980 3340 5820
rect 3460 5810 6360 5820
rect 3400 5760 3460 5770
rect 3400 5590 3460 5600
rect 3680 5760 3740 5770
rect 3680 5590 3740 5600
rect 3980 5760 4040 5770
rect 3980 5590 4040 5600
rect 4280 5760 4340 5770
rect 4280 5590 4340 5600
rect 4580 5760 4640 5770
rect 4580 5590 4640 5600
rect 4860 5760 4920 5770
rect 4860 5590 4920 5600
rect 5160 5760 5220 5770
rect 5160 5590 5220 5600
rect 5460 5760 5520 5770
rect 5460 5590 5520 5600
rect 5760 5760 5820 5770
rect 5760 5590 5820 5600
rect 6060 5760 6120 5770
rect 6060 5590 6120 5600
rect 6360 5760 6420 5770
rect 6360 5590 6420 5600
rect 3560 5240 3620 5250
rect 3560 5070 3620 5080
rect 3840 5240 3900 5250
rect 3840 5070 3900 5080
rect 4140 5240 4200 5250
rect 4140 5070 4200 5080
rect 4420 5240 4480 5250
rect 4420 5070 4480 5080
rect 4740 5240 4800 5250
rect 4740 5070 4800 5080
rect 5020 5240 5080 5250
rect 5020 5070 5080 5080
rect 5320 5240 5380 5250
rect 5320 5070 5380 5080
rect 5620 5240 5680 5250
rect 5620 5070 5680 5080
rect 5900 5240 5960 5250
rect 5900 5070 5960 5080
rect 6200 5240 6260 5250
rect 6200 5070 6260 5080
rect 3180 4820 3200 4980
rect 3320 4820 3340 4980
rect 160 4670 3060 4680
rect 3180 4670 3340 4820
rect 6480 4980 6620 5820
rect 6750 5810 9650 5820
rect 6680 5760 6740 5770
rect 6680 5590 6740 5600
rect 6980 5760 7040 5770
rect 6980 5590 7040 5600
rect 7280 5760 7340 5770
rect 7280 5590 7340 5600
rect 7580 5760 7640 5770
rect 7580 5590 7640 5600
rect 7880 5760 7940 5770
rect 7880 5590 7940 5600
rect 8180 5760 8240 5770
rect 8180 5590 8240 5600
rect 8460 5760 8520 5770
rect 8460 5590 8520 5600
rect 8760 5760 8820 5770
rect 8760 5590 8820 5600
rect 9060 5760 9120 5770
rect 9060 5590 9120 5600
rect 9360 5760 9420 5770
rect 9360 5590 9420 5600
rect 9660 5760 9720 5770
rect 9660 5590 9720 5600
rect 6480 4820 6500 4980
rect 6600 4820 6620 4980
rect 3460 4670 6360 4680
rect 6480 4670 6620 4820
rect 6840 4980 6900 4990
rect 6840 4810 6900 4820
rect 7140 4980 7200 4990
rect 7140 4810 7200 4820
rect 7440 4980 7500 4990
rect 7440 4810 7500 4820
rect 7720 4980 7780 4990
rect 7720 4810 7780 4820
rect 8020 4980 8080 4990
rect 8020 4810 8080 4820
rect 8320 4980 8380 4990
rect 8320 4810 8380 4820
rect 8600 4980 8660 4990
rect 8600 4810 8660 4820
rect 8900 4980 8960 4990
rect 8900 4810 8960 4820
rect 9200 4980 9260 4990
rect 9200 4810 9260 4820
rect 9500 4980 9560 4990
rect 9500 4810 9560 4820
rect 9780 4980 9920 5820
rect 10040 5810 12940 5820
rect 9980 5760 10040 5770
rect 9980 5590 10040 5600
rect 10280 5760 10340 5770
rect 10280 5590 10340 5600
rect 10580 5760 10640 5770
rect 10580 5590 10640 5600
rect 10880 5760 10940 5770
rect 10880 5590 10940 5600
rect 11160 5760 11220 5770
rect 11160 5590 11220 5600
rect 11460 5760 11520 5770
rect 11460 5590 11520 5600
rect 11760 5760 11820 5770
rect 11760 5590 11820 5600
rect 12060 5760 12120 5770
rect 12060 5590 12120 5600
rect 12340 5760 12400 5770
rect 12340 5590 12400 5600
rect 12640 5760 12700 5770
rect 12640 5590 12700 5600
rect 12940 5760 13000 5770
rect 12940 5590 13000 5600
rect 10120 5240 10180 5250
rect 10120 5070 10180 5080
rect 10420 5240 10480 5250
rect 10420 5070 10480 5080
rect 10740 5240 10800 5250
rect 10740 5070 10800 5080
rect 11020 5240 11080 5250
rect 11020 5070 11080 5080
rect 11320 5240 11380 5250
rect 11320 5070 11380 5080
rect 11600 5240 11660 5250
rect 11600 5070 11660 5080
rect 11920 5240 11980 5250
rect 11920 5070 11980 5080
rect 12200 5240 12260 5250
rect 12200 5070 12260 5080
rect 12500 5240 12560 5250
rect 12500 5070 12560 5080
rect 12800 5240 12860 5250
rect 12800 5070 12860 5080
rect 9780 4820 9800 4980
rect 9900 4820 9920 4980
rect 6750 4670 9650 4680
rect 9780 4670 9920 4820
rect 13060 4980 13200 5820
rect 13340 5810 16240 5820
rect 13280 5760 13340 5770
rect 13280 5590 13340 5600
rect 13560 5760 13620 5770
rect 13560 5590 13620 5600
rect 13880 5760 13940 5770
rect 13880 5590 13940 5600
rect 14160 5760 14220 5770
rect 14160 5590 14220 5600
rect 14460 5760 14520 5770
rect 14460 5590 14520 5600
rect 14740 5760 14800 5770
rect 14740 5590 14800 5600
rect 15060 5760 15120 5770
rect 15060 5590 15120 5600
rect 15360 5760 15420 5770
rect 15360 5590 15420 5600
rect 15640 5760 15700 5770
rect 15640 5590 15700 5600
rect 15940 5760 16000 5770
rect 15940 5590 16000 5600
rect 16240 5760 16300 5770
rect 16240 5590 16300 5600
rect 16400 5760 16800 5940
rect 16400 5600 16420 5760
rect 16780 5600 16800 5760
rect 13440 5500 13500 5510
rect 13440 5330 13500 5340
rect 13720 5500 13780 5510
rect 13720 5330 13780 5340
rect 14020 5500 14080 5510
rect 14020 5330 14080 5340
rect 14320 5500 14380 5510
rect 14320 5330 14380 5340
rect 14600 5500 14660 5510
rect 14600 5330 14660 5340
rect 14900 5500 14960 5510
rect 14900 5330 14960 5340
rect 15200 5500 15260 5510
rect 15200 5330 15260 5340
rect 15500 5500 15560 5510
rect 15500 5330 15560 5340
rect 15800 5500 15860 5510
rect 15800 5330 15860 5340
rect 16080 5500 16140 5510
rect 16080 5330 16140 5340
rect 13060 4820 13080 4980
rect 13180 4820 13200 4980
rect 10040 4670 12940 4680
rect 13060 4670 13200 4820
rect 13340 4670 16240 4680
rect 3060 4610 3460 4670
rect 6360 4610 6750 4670
rect 9650 4610 10040 4670
rect 12940 4610 13340 4670
rect 160 4600 3060 4610
rect 160 4360 3060 4370
rect 3180 4360 3340 4610
rect 3460 4600 6360 4610
rect 3460 4360 6360 4370
rect 6480 4360 6620 4610
rect 6750 4600 9650 4610
rect 6750 4360 9650 4370
rect 9780 4360 9920 4610
rect 10040 4600 12940 4610
rect 10040 4360 12940 4370
rect 13060 4360 13200 4610
rect 13340 4600 16240 4610
rect 16400 4560 16800 5600
rect 16780 4420 16800 4560
rect 13340 4360 16240 4370
rect 3060 4300 3460 4360
rect 6360 4300 6750 4360
rect 9650 4300 10040 4360
rect 12940 4300 13340 4360
rect 160 4290 3060 4300
rect 100 4240 160 4250
rect 100 4070 160 4080
rect 400 4240 460 4250
rect 400 4070 460 4080
rect 680 4240 740 4250
rect 680 4070 740 4080
rect 980 4240 1040 4250
rect 980 4070 1040 4080
rect 1280 4240 1340 4250
rect 1280 4070 1340 4080
rect 1580 4240 1640 4250
rect 1580 4070 1640 4080
rect 1880 4240 1940 4250
rect 1880 4070 1940 4080
rect 2180 4240 2240 4250
rect 2180 4070 2240 4080
rect 2460 4240 2520 4250
rect 2460 4070 2520 4080
rect 2760 4240 2820 4250
rect 2760 4070 2820 4080
rect 3060 4240 3120 4250
rect 3060 4070 3120 4080
rect 240 3980 300 3990
rect 240 3810 300 3820
rect 540 3980 600 3990
rect 540 3810 600 3820
rect 840 3980 900 3990
rect 840 3810 900 3820
rect 1140 3980 1200 3990
rect 1140 3810 1200 3820
rect 1440 3980 1500 3990
rect 1440 3810 1500 3820
rect 1740 3980 1800 3990
rect 1740 3810 1800 3820
rect 2020 3980 2080 3990
rect 2020 3810 2080 3820
rect 2320 3980 2380 3990
rect 2320 3810 2380 3820
rect 2620 3980 2680 3990
rect 2620 3810 2680 3820
rect 2900 3980 2960 3990
rect 2900 3810 2960 3820
rect 100 3460 160 3470
rect 100 3290 160 3300
rect 400 3460 460 3470
rect 400 3290 460 3300
rect 680 3460 740 3470
rect 680 3290 740 3300
rect 980 3460 1040 3470
rect 980 3290 1040 3300
rect 1280 3460 1340 3470
rect 1280 3290 1340 3300
rect 1580 3460 1640 3470
rect 1580 3290 1640 3300
rect 1860 3460 1920 3470
rect 1860 3290 1920 3300
rect 2160 3460 2220 3470
rect 2160 3290 2220 3300
rect 2480 3460 2540 3470
rect 2480 3290 2540 3300
rect 2760 3460 2820 3470
rect 2760 3290 2820 3300
rect 3060 3460 3120 3470
rect 3060 3290 3120 3300
rect 160 3160 3060 3170
rect 3180 3160 3340 4300
rect 3460 4290 6360 4300
rect 3400 4240 3460 4250
rect 3400 4070 3460 4080
rect 3680 4240 3740 4250
rect 3680 4070 3740 4080
rect 3980 4240 4040 4250
rect 3980 4070 4040 4080
rect 4280 4240 4340 4250
rect 4280 4070 4340 4080
rect 4560 4240 4620 4250
rect 4560 4070 4620 4080
rect 4860 4240 4920 4250
rect 4860 4070 4920 4080
rect 5160 4240 5220 4250
rect 5160 4070 5220 4080
rect 5460 4240 5520 4250
rect 5460 4070 5520 4080
rect 5780 4240 5840 4250
rect 5780 4070 5840 4080
rect 6060 4240 6120 4250
rect 6060 4070 6120 4080
rect 6360 4240 6420 4250
rect 6360 4070 6420 4080
rect 3540 3720 3600 3730
rect 3540 3550 3600 3560
rect 3840 3720 3900 3730
rect 3840 3550 3900 3560
rect 4140 3720 4200 3730
rect 4140 3550 4200 3560
rect 4420 3720 4480 3730
rect 4420 3550 4480 3560
rect 4720 3720 4780 3730
rect 4720 3550 4780 3560
rect 5020 3720 5080 3730
rect 5020 3550 5080 3560
rect 5320 3720 5380 3730
rect 5320 3550 5380 3560
rect 5620 3720 5680 3730
rect 5620 3550 5680 3560
rect 5920 3720 5980 3730
rect 5920 3550 5980 3560
rect 6200 3720 6260 3730
rect 6200 3550 6260 3560
rect 3400 3460 3460 3470
rect 3400 3290 3460 3300
rect 3680 3460 3740 3470
rect 3680 3290 3740 3300
rect 4000 3460 4060 3470
rect 4000 3290 4060 3300
rect 4280 3460 4340 3470
rect 4280 3290 4340 3300
rect 4580 3460 4640 3470
rect 4580 3290 4640 3300
rect 4860 3460 4920 3470
rect 4860 3290 4920 3300
rect 5160 3460 5220 3470
rect 5160 3290 5220 3300
rect 5460 3460 5520 3470
rect 5460 3290 5520 3300
rect 5760 3460 5820 3470
rect 5760 3290 5820 3300
rect 6060 3460 6120 3470
rect 6060 3290 6120 3300
rect 6360 3460 6420 3470
rect 6360 3290 6420 3300
rect 3460 3160 6360 3170
rect 6480 3160 6620 4300
rect 6750 4290 9650 4300
rect 6700 4240 6760 4250
rect 6700 4070 6760 4080
rect 6980 4240 7040 4250
rect 6980 4070 7040 4080
rect 7280 4240 7340 4250
rect 7280 4070 7340 4080
rect 7580 4240 7640 4250
rect 7580 4070 7640 4080
rect 7880 4240 7940 4250
rect 7880 4070 7940 4080
rect 8160 4240 8220 4250
rect 8160 4070 8220 4080
rect 8460 4240 8520 4250
rect 8460 4070 8520 4080
rect 8760 4240 8820 4250
rect 8760 4070 8820 4080
rect 9060 4240 9120 4250
rect 9060 4070 9120 4080
rect 9340 4240 9400 4250
rect 9340 4070 9400 4080
rect 9640 4240 9700 4250
rect 9640 4070 9700 4080
rect 6840 3720 6900 3730
rect 6840 3550 6900 3560
rect 7140 3720 7200 3730
rect 7140 3550 7200 3560
rect 7440 3720 7500 3730
rect 7440 3550 7500 3560
rect 7720 3720 7780 3730
rect 7720 3550 7780 3560
rect 8020 3720 8080 3730
rect 8020 3550 8080 3560
rect 8320 3720 8380 3730
rect 8320 3550 8380 3560
rect 8620 3720 8680 3730
rect 8620 3550 8680 3560
rect 8900 3720 8960 3730
rect 8900 3550 8960 3560
rect 9200 3720 9260 3730
rect 9200 3550 9260 3560
rect 9500 3720 9560 3730
rect 9500 3550 9560 3560
rect 6680 3460 6740 3470
rect 6680 3290 6740 3300
rect 6980 3460 7040 3470
rect 6980 3290 7040 3300
rect 7280 3460 7340 3470
rect 7280 3290 7340 3300
rect 7580 3460 7640 3470
rect 7580 3290 7640 3300
rect 7880 3460 7940 3470
rect 7880 3290 7940 3300
rect 8160 3460 8220 3470
rect 8160 3290 8220 3300
rect 8460 3460 8520 3470
rect 8460 3290 8520 3300
rect 8780 3460 8840 3470
rect 8780 3290 8840 3300
rect 9060 3460 9120 3470
rect 9060 3290 9120 3300
rect 9360 3460 9420 3470
rect 9360 3290 9420 3300
rect 9660 3460 9720 3470
rect 9660 3290 9720 3300
rect 6750 3160 9650 3170
rect 9780 3160 9920 4300
rect 10040 4290 12940 4300
rect 9980 4240 10040 4250
rect 9980 4070 10040 4080
rect 10280 4240 10340 4250
rect 10280 4070 10340 4080
rect 10560 4240 10620 4250
rect 10560 4070 10620 4080
rect 10860 4240 10920 4250
rect 10860 4070 10920 4080
rect 11160 4240 11220 4250
rect 11160 4070 11220 4080
rect 11460 4240 11520 4250
rect 11460 4070 11520 4080
rect 11760 4240 11820 4250
rect 11760 4070 11820 4080
rect 12060 4240 12120 4250
rect 12060 4070 12120 4080
rect 12340 4240 12400 4250
rect 12340 4070 12400 4080
rect 12640 4240 12700 4250
rect 12640 4070 12700 4080
rect 12940 4240 13000 4250
rect 12940 4070 13000 4080
rect 10140 3720 10200 3730
rect 10140 3550 10200 3560
rect 10420 3720 10480 3730
rect 10420 3550 10480 3560
rect 10720 3720 10780 3730
rect 10720 3550 10780 3560
rect 11020 3720 11080 3730
rect 11020 3550 11080 3560
rect 11320 3720 11380 3730
rect 11320 3550 11380 3560
rect 11600 3720 11660 3730
rect 11600 3550 11660 3560
rect 11900 3720 11960 3730
rect 11900 3550 11960 3560
rect 12200 3720 12260 3730
rect 12200 3550 12260 3560
rect 12500 3720 12560 3730
rect 12500 3550 12560 3560
rect 12800 3720 12860 3730
rect 12800 3550 12860 3560
rect 10000 3460 10060 3470
rect 10000 3290 10060 3300
rect 10280 3460 10340 3470
rect 10280 3290 10340 3300
rect 10580 3460 10640 3470
rect 10580 3290 10640 3300
rect 10860 3460 10920 3470
rect 10860 3290 10920 3300
rect 11180 3460 11240 3470
rect 11180 3290 11240 3300
rect 11460 3460 11520 3470
rect 11460 3290 11520 3300
rect 11760 3460 11820 3470
rect 11760 3290 11820 3300
rect 12060 3460 12120 3470
rect 12060 3290 12120 3300
rect 12360 3460 12420 3470
rect 12360 3290 12420 3300
rect 12640 3460 12700 3470
rect 12640 3290 12700 3300
rect 12940 3460 13000 3470
rect 12940 3290 13000 3300
rect 10040 3160 12940 3170
rect 13060 3160 13200 4300
rect 13340 4290 16240 4300
rect 13280 4240 13340 4250
rect 13280 4070 13340 4080
rect 13560 4240 13620 4250
rect 13560 4070 13620 4080
rect 13860 4240 13920 4250
rect 13860 4070 13920 4080
rect 14160 4240 14220 4250
rect 14160 4070 14220 4080
rect 14460 4240 14520 4250
rect 14460 4070 14520 4080
rect 14760 4240 14820 4250
rect 14760 4070 14820 4080
rect 15060 4240 15120 4250
rect 15060 4070 15120 4080
rect 15360 4240 15420 4250
rect 15360 4070 15420 4080
rect 15640 4240 15700 4250
rect 15640 4070 15700 4080
rect 15940 4240 16000 4250
rect 15940 4070 16000 4080
rect 16220 4240 16280 4250
rect 16220 4070 16280 4080
rect 16400 4240 16800 4420
rect 16400 4080 16420 4240
rect 16780 4080 16800 4240
rect 13440 3980 13500 3990
rect 13440 3810 13500 3820
rect 13720 3980 13780 3990
rect 13720 3810 13780 3820
rect 14020 3980 14080 3990
rect 14020 3810 14080 3820
rect 14320 3980 14380 3990
rect 14320 3810 14380 3820
rect 14600 3980 14660 3990
rect 14600 3810 14660 3820
rect 14900 3980 14960 3990
rect 14900 3810 14960 3820
rect 15200 3980 15260 3990
rect 15200 3810 15260 3820
rect 15500 3980 15560 3990
rect 15500 3810 15560 3820
rect 15780 3980 15840 3990
rect 15780 3810 15840 3820
rect 16080 3980 16140 3990
rect 16080 3810 16140 3820
rect 13280 3460 13340 3470
rect 13280 3290 13340 3300
rect 13560 3460 13620 3470
rect 13560 3290 13620 3300
rect 13880 3460 13940 3470
rect 13880 3290 13940 3300
rect 14180 3460 14240 3470
rect 14180 3290 14240 3300
rect 14460 3460 14520 3470
rect 14460 3290 14520 3300
rect 14740 3460 14800 3470
rect 14740 3290 14800 3300
rect 15040 3460 15100 3470
rect 15040 3290 15100 3300
rect 15360 3460 15420 3470
rect 15360 3290 15420 3300
rect 15640 3460 15700 3470
rect 15640 3290 15700 3300
rect 15940 3460 16000 3470
rect 15940 3290 16000 3300
rect 16240 3460 16300 3470
rect 16240 3290 16300 3300
rect 16400 3460 16800 4080
rect 16400 3300 16420 3460
rect 16780 3300 16800 3460
rect 13340 3160 16240 3170
rect 3060 3100 3460 3160
rect 6360 3100 6750 3160
rect 9650 3100 10040 3160
rect 12940 3100 13340 3160
rect 160 3090 3060 3100
rect 150 2840 3050 2850
rect 3180 2840 3340 3100
rect 3460 3090 6360 3100
rect 3450 2840 6350 2850
rect 6480 2840 6620 3100
rect 6750 3090 9650 3100
rect 6740 2840 9640 2850
rect 9780 2840 9920 3100
rect 10040 3090 12940 3100
rect 10030 2840 12930 2850
rect 13060 2840 13200 3100
rect 13340 3090 16240 3100
rect 16400 3040 16800 3300
rect 16780 2900 16800 3040
rect 13330 2840 16230 2850
rect 3050 2780 3450 2840
rect 6350 2780 6740 2840
rect 9640 2780 10030 2840
rect 12930 2780 13330 2840
rect 150 2770 3050 2780
rect 100 2720 160 2730
rect 100 2550 160 2560
rect 400 2720 460 2730
rect 400 2550 460 2560
rect 680 2720 740 2730
rect 680 2550 740 2560
rect 980 2720 1040 2730
rect 980 2550 1040 2560
rect 1300 2720 1360 2730
rect 1300 2550 1360 2560
rect 1600 2720 1660 2730
rect 1600 2550 1660 2560
rect 1880 2720 1940 2730
rect 1880 2550 1940 2560
rect 2180 2720 2240 2730
rect 2180 2550 2240 2560
rect 2460 2720 2520 2730
rect 2460 2550 2520 2560
rect 2760 2720 2820 2730
rect 2760 2550 2820 2560
rect 3060 2720 3120 2730
rect 3060 2550 3120 2560
rect 260 2460 320 2470
rect 260 2290 320 2300
rect 540 2460 600 2470
rect 540 2290 600 2300
rect 840 2460 900 2470
rect 840 2290 900 2300
rect 1140 2460 1200 2470
rect 1140 2290 1200 2300
rect 1440 2460 1500 2470
rect 1440 2290 1500 2300
rect 1740 2460 1800 2470
rect 1740 2290 1800 2300
rect 2020 2460 2080 2470
rect 2020 2290 2080 2300
rect 2320 2460 2380 2470
rect 2320 2290 2380 2300
rect 2620 2460 2680 2470
rect 2620 2290 2680 2300
rect 2900 2460 2960 2470
rect 2900 2290 2960 2300
rect 100 1940 160 1950
rect 100 1770 160 1780
rect 400 1940 460 1950
rect 400 1770 460 1780
rect 680 1940 740 1950
rect 680 1770 740 1780
rect 1000 1940 1060 1950
rect 1000 1770 1060 1780
rect 1300 1940 1360 1950
rect 1300 1770 1360 1780
rect 1600 1940 1660 1950
rect 1600 1770 1660 1780
rect 1880 1940 1940 1950
rect 1880 1770 1940 1780
rect 2180 1940 2240 1950
rect 2180 1770 2240 1780
rect 2460 1940 2520 1950
rect 2460 1770 2520 1780
rect 2760 1940 2820 1950
rect 2760 1770 2820 1780
rect 3060 1940 3120 1950
rect 3060 1770 3120 1780
rect 150 1630 3050 1640
rect 3180 1630 3340 2780
rect 3450 2770 6350 2780
rect 3400 2720 3460 2730
rect 3680 2720 3740 2730
rect 3460 2560 3680 2600
rect 3980 2720 4040 2730
rect 3740 2560 3980 2600
rect 4280 2720 4340 2730
rect 4040 2560 4280 2600
rect 4580 2720 4640 2730
rect 4340 2560 4580 2600
rect 4880 2720 4940 2730
rect 4640 2560 4880 2600
rect 5160 2720 5220 2730
rect 4940 2560 5160 2600
rect 5460 2720 5520 2730
rect 5220 2560 5460 2600
rect 5760 2720 5820 2730
rect 5520 2560 5760 2600
rect 6060 2720 6120 2730
rect 5820 2560 6060 2600
rect 6360 2720 6420 2730
rect 6120 2560 6360 2600
rect 3400 2550 6420 2560
rect 3440 2460 6360 2550
rect 3440 2000 3540 2460
rect 3620 2000 3820 2460
rect 3900 2000 4120 2460
rect 4200 2000 4420 2460
rect 4500 2000 4720 2460
rect 4800 2000 5020 2460
rect 5100 2000 5320 2460
rect 5400 2000 5600 2460
rect 5680 2000 5900 2460
rect 5980 2000 6200 2460
rect 6280 2000 6360 2460
rect 3440 1950 6360 2000
rect 3400 1940 6400 1950
rect 3460 1920 3680 1940
rect 3400 1770 3460 1780
rect 3740 1920 3980 1940
rect 3680 1770 3740 1780
rect 4040 1920 4280 1940
rect 3980 1770 4040 1780
rect 4340 1920 4580 1940
rect 4280 1770 4340 1780
rect 4640 1920 4880 1940
rect 4580 1770 4640 1780
rect 4940 1920 5160 1940
rect 4880 1770 4940 1780
rect 5220 1920 5460 1940
rect 5160 1770 5220 1780
rect 5520 1920 5780 1940
rect 5460 1770 5520 1780
rect 5840 1920 6060 1940
rect 5780 1770 5840 1780
rect 6120 1920 6340 1940
rect 6060 1770 6120 1780
rect 6340 1770 6400 1780
rect 3450 1630 6350 1640
rect 6480 1630 6620 2780
rect 6740 2770 9640 2780
rect 6680 2720 6740 2730
rect 6680 2550 6740 2560
rect 6980 2720 7040 2730
rect 6980 2550 7040 2560
rect 7280 2720 7340 2730
rect 7280 2550 7340 2560
rect 7580 2720 7640 2730
rect 7580 2550 7640 2560
rect 7880 2720 7940 2730
rect 7880 2550 7940 2560
rect 8160 2720 8220 2730
rect 8160 2550 8220 2560
rect 8460 2720 8520 2730
rect 8460 2550 8520 2560
rect 8760 2720 8820 2730
rect 8760 2550 8820 2560
rect 9040 2720 9100 2730
rect 9040 2550 9100 2560
rect 9340 2720 9400 2730
rect 9340 2550 9400 2560
rect 9640 2720 9700 2730
rect 9640 2550 9700 2560
rect 6840 2200 6900 2210
rect 6840 2030 6900 2040
rect 7140 2200 7200 2210
rect 7140 2030 7200 2040
rect 7440 2200 7500 2210
rect 7440 2030 7500 2040
rect 7720 2200 7780 2210
rect 7720 2030 7780 2040
rect 8020 2200 8080 2210
rect 8020 2030 8080 2040
rect 8320 2200 8380 2210
rect 8320 2030 8380 2040
rect 8600 2200 8660 2210
rect 8600 2030 8660 2040
rect 8900 2200 8960 2210
rect 8900 2030 8960 2040
rect 9200 2200 9260 2210
rect 9200 2030 9260 2040
rect 9500 2200 9560 2210
rect 9500 2030 9560 2040
rect 6680 1940 6740 1950
rect 6680 1770 6740 1780
rect 7000 1940 7060 1950
rect 7000 1770 7060 1780
rect 7280 1940 7340 1950
rect 7280 1770 7340 1780
rect 7580 1940 7640 1950
rect 7580 1770 7640 1780
rect 7860 1940 7920 1950
rect 7860 1770 7920 1780
rect 8180 1940 8240 1950
rect 8180 1770 8240 1780
rect 8460 1940 8520 1950
rect 8460 1770 8520 1780
rect 8760 1940 8820 1950
rect 8760 1770 8820 1780
rect 9060 1940 9120 1950
rect 9060 1770 9120 1780
rect 9340 1940 9400 1950
rect 9340 1770 9400 1780
rect 9640 1940 9700 1950
rect 9640 1770 9700 1780
rect 6740 1630 9640 1640
rect 9780 1630 9920 2780
rect 10030 2770 12930 2780
rect 9980 2720 10040 2730
rect 9980 2550 10040 2560
rect 10280 2720 10340 2730
rect 10280 2550 10340 2560
rect 10560 2720 10620 2730
rect 10560 2550 10620 2560
rect 10860 2720 10920 2730
rect 10860 2550 10920 2560
rect 11160 2720 11220 2730
rect 11160 2550 11220 2560
rect 11460 2720 11520 2730
rect 11460 2550 11520 2560
rect 11760 2720 11820 2730
rect 11760 2550 11820 2560
rect 12040 2720 12100 2730
rect 12040 2550 12100 2560
rect 12340 2720 12400 2730
rect 12340 2550 12400 2560
rect 12640 2720 12700 2730
rect 12640 2550 12700 2560
rect 12940 2720 13000 2730
rect 12940 2550 13000 2560
rect 10140 2460 10200 2470
rect 10140 2290 10200 2300
rect 10420 2460 10480 2470
rect 10420 2290 10480 2300
rect 10720 2460 10780 2470
rect 10720 2290 10780 2300
rect 11020 2460 11080 2470
rect 11020 2290 11080 2300
rect 11320 2460 11380 2470
rect 11320 2290 11380 2300
rect 11600 2460 11660 2470
rect 11600 2290 11660 2300
rect 11920 2460 11980 2470
rect 11920 2290 11980 2300
rect 12200 2460 12260 2470
rect 12200 2290 12260 2300
rect 12500 2460 12560 2470
rect 12500 2290 12560 2300
rect 12800 2460 12860 2470
rect 12800 2290 12860 2300
rect 10000 1940 10060 1950
rect 10000 1770 10060 1780
rect 10280 1940 10340 1950
rect 10280 1770 10340 1780
rect 10580 1940 10640 1950
rect 10580 1770 10640 1780
rect 10880 1940 10940 1950
rect 10880 1770 10940 1780
rect 11160 1940 11220 1950
rect 11160 1770 11220 1780
rect 11460 1940 11520 1950
rect 11460 1770 11520 1780
rect 11760 1940 11820 1950
rect 11760 1770 11820 1780
rect 12060 1940 12120 1950
rect 12060 1770 12120 1780
rect 12360 1940 12420 1950
rect 12360 1770 12420 1780
rect 12640 1940 12700 1950
rect 12640 1770 12700 1780
rect 12940 1940 13000 1950
rect 12940 1770 13000 1780
rect 10030 1630 12930 1640
rect 13060 1630 13200 2780
rect 13330 2770 16230 2780
rect 13280 2720 13340 2730
rect 13280 2550 13340 2560
rect 13580 2720 13640 2730
rect 13580 2550 13640 2560
rect 13860 2720 13920 2730
rect 13860 2550 13920 2560
rect 14160 2720 14220 2730
rect 14160 2550 14220 2560
rect 14460 2720 14520 2730
rect 14460 2550 14520 2560
rect 14760 2720 14820 2730
rect 14760 2550 14820 2560
rect 15060 2720 15120 2730
rect 15060 2550 15120 2560
rect 15340 2720 15400 2730
rect 15340 2550 15400 2560
rect 15640 2720 15700 2730
rect 15640 2550 15700 2560
rect 15940 2720 16000 2730
rect 15940 2550 16000 2560
rect 16240 2720 16300 2730
rect 16240 2550 16300 2560
rect 16400 2720 16800 2900
rect 16400 2560 16420 2720
rect 16780 2560 16800 2720
rect 13440 2460 13500 2470
rect 13440 2290 13500 2300
rect 13720 2460 13780 2470
rect 13720 2290 13780 2300
rect 14020 2460 14080 2470
rect 14020 2290 14080 2300
rect 14320 2460 14380 2470
rect 14320 2290 14380 2300
rect 14620 2460 14680 2470
rect 14620 2290 14680 2300
rect 14900 2460 14960 2470
rect 14900 2290 14960 2300
rect 15200 2460 15260 2470
rect 15200 2290 15260 2300
rect 15500 2460 15560 2470
rect 15500 2290 15560 2300
rect 15800 2460 15860 2470
rect 15800 2290 15860 2300
rect 16100 2460 16160 2470
rect 16100 2290 16160 2300
rect 13280 1940 13340 1950
rect 13280 1770 13340 1780
rect 13560 1940 13620 1950
rect 13560 1770 13620 1780
rect 13880 1940 13940 1950
rect 13880 1770 13940 1780
rect 14160 1940 14220 1950
rect 14160 1770 14220 1780
rect 14460 1940 14520 1950
rect 14460 1770 14520 1780
rect 14760 1940 14820 1950
rect 14760 1770 14820 1780
rect 15060 1940 15120 1950
rect 15060 1770 15120 1780
rect 15340 1940 15400 1950
rect 15340 1770 15400 1780
rect 15640 1940 15700 1950
rect 15640 1770 15700 1780
rect 15940 1940 16000 1950
rect 15940 1770 16000 1780
rect 16240 1940 16300 1950
rect 16240 1770 16300 1780
rect 16400 1940 16800 2560
rect 16400 1780 16420 1940
rect 16780 1780 16800 1940
rect 13330 1630 16230 1640
rect 3050 1570 3450 1630
rect 6350 1570 6740 1630
rect 9640 1570 10030 1630
rect 12930 1570 13330 1630
rect 150 1560 3050 1570
rect 150 1330 3050 1340
rect 3180 1330 3340 1570
rect 3450 1560 6350 1570
rect 3450 1330 6350 1340
rect 6480 1330 6620 1570
rect 6740 1560 9640 1570
rect 6740 1330 9640 1340
rect 9780 1330 9920 1570
rect 10030 1560 12930 1570
rect 10030 1330 12930 1340
rect 13060 1330 13200 1570
rect 13330 1560 16230 1570
rect 16400 1520 16800 1780
rect 16780 1380 16800 1520
rect 13330 1330 16230 1340
rect 3050 1270 3450 1330
rect 6350 1270 6740 1330
rect 9640 1270 10030 1330
rect 12930 1270 13330 1330
rect 150 1260 3050 1270
rect 100 1210 160 1220
rect 100 1020 160 1030
rect 400 1210 460 1220
rect 400 1020 460 1030
rect 700 1210 760 1220
rect 700 1020 760 1030
rect 1000 1210 1060 1220
rect 1000 1020 1060 1030
rect 1280 1210 1340 1220
rect 1280 1020 1340 1030
rect 1580 1210 1640 1220
rect 1580 1020 1640 1030
rect 1880 1210 1940 1220
rect 1880 1020 1940 1030
rect 2180 1210 2240 1220
rect 2180 1020 2240 1030
rect 2480 1210 2540 1220
rect 2480 1020 2540 1030
rect 2760 1210 2820 1220
rect 2760 1020 2820 1030
rect 3060 1210 3120 1220
rect 3060 1020 3120 1030
rect 240 950 300 960
rect 240 760 300 770
rect 540 950 600 960
rect 540 760 600 770
rect 840 950 900 960
rect 840 760 900 770
rect 1140 950 1200 960
rect 1140 760 1200 770
rect 1440 950 1500 960
rect 1440 760 1500 770
rect 1740 950 1800 960
rect 1740 760 1800 770
rect 2020 950 2080 960
rect 2020 760 2080 770
rect 2320 950 2380 960
rect 2320 760 2380 770
rect 2620 950 2680 960
rect 2620 760 2680 770
rect 2920 950 2980 960
rect 2920 760 2980 770
rect 120 690 180 700
rect 120 500 180 510
rect 400 690 460 700
rect 400 500 460 510
rect 680 690 740 700
rect 680 500 740 510
rect 980 690 1040 700
rect 980 500 1040 510
rect 1300 690 1360 700
rect 1300 500 1360 510
rect 1600 690 1660 700
rect 1600 500 1660 510
rect 1880 690 1940 700
rect 1880 500 1940 510
rect 2160 690 2220 700
rect 2160 500 2220 510
rect 2480 690 2540 700
rect 2480 500 2540 510
rect 2760 690 2820 700
rect 2760 500 2820 510
rect 3060 690 3120 700
rect 3060 500 3120 510
rect 240 430 300 440
rect 240 240 300 250
rect 540 430 600 440
rect 540 240 600 250
rect 840 430 900 440
rect 840 240 900 250
rect 1140 430 1200 440
rect 1140 240 1200 250
rect 1440 430 1500 440
rect 1440 240 1500 250
rect 1740 430 1800 440
rect 1740 240 1800 250
rect 2020 430 2080 440
rect 2020 240 2080 250
rect 2340 430 2400 440
rect 2340 240 2400 250
rect 2620 430 2680 440
rect 2620 240 2680 250
rect 2920 430 2980 440
rect 2920 240 2980 250
rect 150 120 3050 130
rect 3180 120 3340 1270
rect 3450 1260 6350 1270
rect 3400 1210 3460 1220
rect 3400 1020 3460 1030
rect 3680 1210 3740 1220
rect 3680 1020 3740 1030
rect 4000 1210 4060 1220
rect 4000 1020 4060 1030
rect 4280 1210 4340 1220
rect 4280 1020 4340 1030
rect 4580 1210 4640 1220
rect 4580 1020 4640 1030
rect 4880 1210 4940 1220
rect 4880 1020 4940 1030
rect 5160 1210 5220 1220
rect 5160 1020 5220 1030
rect 5460 1210 5520 1220
rect 5460 1020 5520 1030
rect 5760 1210 5820 1220
rect 5760 1020 5820 1030
rect 6060 1210 6120 1220
rect 6060 1020 6120 1030
rect 6360 1210 6420 1220
rect 6360 1020 6420 1030
rect 3540 950 3600 960
rect 3540 760 3600 770
rect 3840 950 3900 960
rect 3840 760 3900 770
rect 4140 950 4200 960
rect 4140 760 4200 770
rect 4440 950 4500 960
rect 4440 760 4500 770
rect 4720 950 4780 960
rect 4720 760 4780 770
rect 5020 950 5080 960
rect 5020 760 5080 770
rect 5320 950 5380 960
rect 5320 760 5380 770
rect 5620 950 5680 960
rect 5620 760 5680 770
rect 5900 950 5960 960
rect 5900 760 5960 770
rect 6220 950 6280 960
rect 6220 760 6280 770
rect 3400 690 3460 700
rect 3400 500 3460 510
rect 3700 690 3760 700
rect 3700 500 3760 510
rect 4000 690 4060 700
rect 4000 500 4060 510
rect 4280 690 4340 700
rect 4280 500 4340 510
rect 4580 690 4640 700
rect 4580 500 4640 510
rect 4880 690 4940 700
rect 4880 500 4940 510
rect 5180 690 5240 700
rect 5180 500 5240 510
rect 5460 690 5520 700
rect 5460 500 5520 510
rect 5760 690 5820 700
rect 5760 500 5820 510
rect 6060 690 6120 700
rect 6060 500 6120 510
rect 6360 690 6420 700
rect 6360 500 6420 510
rect 3540 430 3600 440
rect 3540 240 3600 250
rect 3840 430 3900 440
rect 3840 240 3900 250
rect 4140 430 4200 440
rect 4140 240 4200 250
rect 4440 430 4500 440
rect 4440 240 4500 250
rect 4720 430 4780 440
rect 4720 240 4780 250
rect 5020 430 5080 440
rect 5020 240 5080 250
rect 5320 430 5380 440
rect 5320 240 5380 250
rect 5620 430 5680 440
rect 5620 240 5680 250
rect 5900 430 5960 440
rect 5900 240 5960 250
rect 6220 430 6280 440
rect 6220 240 6280 250
rect 3450 120 6350 130
rect 6480 120 6620 1270
rect 6740 1260 9640 1270
rect 6700 1210 6760 1220
rect 6700 1020 6760 1030
rect 6980 1210 7040 1220
rect 6980 1020 7040 1030
rect 7280 1210 7340 1220
rect 7280 1020 7340 1030
rect 7580 1210 7640 1220
rect 7580 1020 7640 1030
rect 7880 1210 7940 1220
rect 7880 1020 7940 1030
rect 8180 1210 8240 1220
rect 8180 1020 8240 1030
rect 8460 1210 8520 1220
rect 8460 1020 8520 1030
rect 8760 1210 8820 1220
rect 8760 1020 8820 1030
rect 9060 1210 9120 1220
rect 9060 1020 9120 1030
rect 9360 1210 9420 1220
rect 9360 1020 9420 1030
rect 9640 1210 9700 1220
rect 9640 1020 9700 1030
rect 6840 950 6900 960
rect 6840 760 6900 770
rect 7140 950 7200 960
rect 7140 760 7200 770
rect 7420 950 7480 960
rect 7420 760 7480 770
rect 7720 950 7780 960
rect 7720 760 7780 770
rect 8020 950 8080 960
rect 8020 760 8080 770
rect 8300 950 8360 960
rect 8300 760 8360 770
rect 8620 950 8680 960
rect 8620 760 8680 770
rect 8920 950 8980 960
rect 8920 760 8980 770
rect 9220 950 9280 960
rect 9220 760 9280 770
rect 9520 950 9580 960
rect 9520 760 9580 770
rect 6700 690 6760 700
rect 6700 500 6760 510
rect 7000 690 7060 700
rect 7000 500 7060 510
rect 7280 690 7340 700
rect 7280 500 7340 510
rect 7580 690 7640 700
rect 7580 500 7640 510
rect 7860 690 7920 700
rect 7860 500 7920 510
rect 8180 690 8240 700
rect 8180 500 8240 510
rect 8480 690 8540 700
rect 8480 500 8540 510
rect 8760 690 8820 700
rect 8760 500 8820 510
rect 9060 690 9120 700
rect 9060 500 9120 510
rect 9360 690 9420 700
rect 9360 500 9420 510
rect 9660 690 9720 700
rect 9660 500 9720 510
rect 6840 430 6900 440
rect 6840 240 6900 250
rect 7140 430 7200 440
rect 7140 240 7200 250
rect 7440 430 7500 440
rect 7440 240 7500 250
rect 7720 430 7780 440
rect 7720 240 7780 250
rect 8020 430 8080 440
rect 8020 240 8080 250
rect 8320 430 8380 440
rect 8320 240 8380 250
rect 8620 430 8680 440
rect 8620 240 8680 250
rect 8920 430 8980 440
rect 8920 240 8980 250
rect 9200 430 9260 440
rect 9200 240 9260 250
rect 9520 430 9580 440
rect 9520 240 9580 250
rect 6740 120 9640 130
rect 9780 120 9920 1270
rect 10030 1260 12930 1270
rect 9980 1210 10040 1220
rect 9980 1020 10040 1030
rect 10280 1210 10340 1220
rect 10280 1020 10340 1030
rect 10560 1210 10620 1220
rect 10560 1020 10620 1030
rect 10860 1210 10920 1220
rect 10860 1020 10920 1030
rect 11160 1210 11220 1220
rect 11160 1020 11220 1030
rect 11460 1210 11520 1220
rect 11460 1020 11520 1030
rect 11760 1210 11820 1220
rect 11760 1020 11820 1030
rect 12060 1210 12120 1220
rect 12060 1020 12120 1030
rect 12360 1210 12420 1220
rect 12360 1020 12420 1030
rect 12660 1210 12720 1220
rect 12660 1020 12720 1030
rect 12940 1210 13000 1220
rect 12940 1020 13000 1030
rect 10140 950 10200 960
rect 10140 760 10200 770
rect 10420 950 10480 960
rect 10420 760 10480 770
rect 10740 950 10800 960
rect 10740 760 10800 770
rect 11020 950 11080 960
rect 11020 760 11080 770
rect 11320 950 11380 960
rect 11320 760 11380 770
rect 11620 950 11680 960
rect 11620 760 11680 770
rect 11920 950 11980 960
rect 11920 760 11980 770
rect 12220 950 12280 960
rect 12220 760 12280 770
rect 12500 950 12560 960
rect 12500 760 12560 770
rect 12800 950 12860 960
rect 12800 760 12860 770
rect 10000 690 10060 700
rect 10000 500 10060 510
rect 10280 690 10340 700
rect 10280 500 10340 510
rect 10580 690 10640 700
rect 10580 500 10640 510
rect 10860 690 10920 700
rect 10860 500 10920 510
rect 11160 690 11220 700
rect 11160 500 11220 510
rect 11480 690 11540 700
rect 11480 500 11540 510
rect 11760 690 11820 700
rect 11760 500 11820 510
rect 12060 690 12120 700
rect 12060 500 12120 510
rect 12360 690 12420 700
rect 12360 500 12420 510
rect 12660 690 12720 700
rect 12660 500 12720 510
rect 12940 690 13000 700
rect 12940 500 13000 510
rect 10140 430 10200 440
rect 10140 240 10200 250
rect 10440 430 10500 440
rect 10440 240 10500 250
rect 10740 430 10800 440
rect 10740 240 10800 250
rect 11020 430 11080 440
rect 11020 240 11080 250
rect 11300 430 11360 440
rect 11300 240 11360 250
rect 11600 430 11660 440
rect 11600 240 11660 250
rect 11900 430 11960 440
rect 11900 240 11960 250
rect 12220 430 12280 440
rect 12220 240 12280 250
rect 12500 430 12560 440
rect 12500 240 12560 250
rect 12800 430 12860 440
rect 12800 240 12860 250
rect 10030 120 12930 130
rect 13060 120 13200 1270
rect 13330 1260 16230 1270
rect 13280 1210 13340 1220
rect 13280 1020 13340 1030
rect 13580 1210 13640 1220
rect 13580 1020 13640 1030
rect 13880 1210 13940 1220
rect 13880 1020 13940 1030
rect 14180 1210 14240 1220
rect 14180 1020 14240 1030
rect 14460 1210 14520 1220
rect 14460 1020 14520 1030
rect 14760 1210 14820 1220
rect 14760 1020 14820 1030
rect 15060 1210 15120 1220
rect 15060 1020 15120 1030
rect 15360 1210 15420 1220
rect 15360 1020 15420 1030
rect 15640 1210 15700 1220
rect 15640 1020 15700 1030
rect 15960 1210 16020 1220
rect 15960 1020 16020 1030
rect 16240 1210 16300 1220
rect 16240 1020 16300 1030
rect 16400 1200 16800 1380
rect 16400 1040 16420 1200
rect 16780 1040 16800 1200
rect 13420 950 13480 960
rect 13420 760 13480 770
rect 13740 950 13800 960
rect 13740 760 13800 770
rect 14020 950 14080 960
rect 14020 760 14080 770
rect 14300 950 14360 960
rect 14300 760 14360 770
rect 14620 950 14680 960
rect 14620 760 14680 770
rect 14920 950 14980 960
rect 14920 760 14980 770
rect 15200 950 15260 960
rect 15200 760 15260 770
rect 15500 950 15560 960
rect 15500 760 15560 770
rect 15780 950 15840 960
rect 15780 760 15840 770
rect 16100 950 16160 960
rect 16100 760 16160 770
rect 13280 690 13340 700
rect 13280 500 13340 510
rect 13580 690 13640 700
rect 13580 500 13640 510
rect 13880 690 13940 700
rect 13880 500 13940 510
rect 14160 690 14220 700
rect 14160 500 14220 510
rect 14460 690 14520 700
rect 14460 500 14520 510
rect 14760 690 14820 700
rect 14760 500 14820 510
rect 15060 690 15120 700
rect 15060 500 15120 510
rect 15360 690 15420 700
rect 15360 500 15420 510
rect 15640 690 15700 700
rect 15640 500 15700 510
rect 15940 690 16000 700
rect 15940 500 16000 510
rect 16240 690 16300 700
rect 16240 500 16300 510
rect 16400 680 16800 1040
rect 16400 520 16420 680
rect 16780 520 16800 680
rect 13440 430 13500 440
rect 13440 240 13500 250
rect 13740 430 13800 440
rect 13740 240 13800 250
rect 14020 430 14080 440
rect 14020 240 14080 250
rect 14320 430 14380 440
rect 14320 240 14380 250
rect 14600 430 14660 440
rect 14600 240 14660 250
rect 14900 430 14960 440
rect 14900 240 14960 250
rect 15200 430 15260 440
rect 15200 240 15260 250
rect 15500 430 15560 440
rect 15500 240 15560 250
rect 15780 430 15840 440
rect 15780 240 15840 250
rect 16100 430 16160 440
rect 16100 240 16160 250
rect 13330 120 16230 130
rect 3050 60 3450 120
rect 6350 60 6740 120
rect 9640 60 10030 120
rect 12930 60 13330 120
rect 150 50 3050 60
rect 3180 -40 3340 60
rect 3450 50 6350 60
rect 6480 -40 6620 60
rect 6740 50 9640 60
rect 9780 -40 9920 60
rect 10030 50 12930 60
rect 13060 -40 13200 60
rect 13330 50 16230 60
rect 16400 0 16800 520
rect 16900 8520 17300 8800
rect 16900 8360 16920 8520
rect 17280 8360 17300 8520
rect 16900 7020 17300 8360
rect 16900 6860 16920 7020
rect 17280 6860 17300 7020
rect 16900 5500 17300 6860
rect 16900 5340 16920 5500
rect 17280 5340 17300 5500
rect 16900 3980 17300 5340
rect 16900 3820 16920 3980
rect 17280 3820 17300 3980
rect 16900 2460 17300 3820
rect 16900 2300 16920 2460
rect 17280 2300 17300 2460
rect 16900 940 17300 2300
rect 16900 780 16920 940
rect 17280 780 17300 940
rect 16900 420 17300 780
rect 16900 260 16920 420
rect 17280 260 17300 420
rect 16900 0 17300 260
rect 17400 6760 17800 8800
rect 17400 6600 17420 6760
rect 17780 6600 17800 6760
rect 17400 5240 17800 6600
rect 17400 5080 17420 5240
rect 17780 5080 17800 5240
rect 17400 3720 17800 5080
rect 17400 3560 17420 3720
rect 17780 3560 17800 3720
rect 17400 2200 17800 3560
rect 17400 2040 17420 2200
rect 17780 2040 17800 2200
rect 17400 0 17800 2040
rect 17900 4980 18300 8800
rect 17900 4820 17920 4980
rect 18280 4820 18300 4980
rect 17900 0 18300 4820
<< via2 >>
rect 100 8610 160 8790
rect 400 8610 460 8790
rect 690 8610 750 8790
rect 990 8610 1050 8790
rect 1290 8610 1350 8790
rect 1590 8610 1650 8790
rect 1880 8610 1940 8790
rect 2170 8610 2230 8790
rect 2470 8610 2530 8790
rect 2760 8610 2820 8790
rect 3060 8610 3120 8790
rect 250 8350 310 8530
rect 550 8350 610 8530
rect 840 8350 900 8530
rect 1140 8350 1200 8530
rect 1440 8350 1500 8530
rect 1730 8350 1790 8530
rect 2030 8350 2090 8530
rect 2320 8350 2380 8530
rect 2620 8350 2680 8530
rect 2920 8350 2980 8530
rect 100 8090 160 8270
rect 400 8090 460 8270
rect 690 8090 750 8270
rect 990 8090 1050 8270
rect 1290 8090 1350 8270
rect 1590 8090 1650 8270
rect 1880 8090 1940 8270
rect 2170 8090 2230 8270
rect 2470 8090 2530 8270
rect 2770 8090 2830 8270
rect 3060 8090 3120 8270
rect 250 7830 310 8010
rect 540 7830 600 8010
rect 840 7830 900 8010
rect 1130 7830 1190 8010
rect 1430 7830 1490 8010
rect 1730 7830 1790 8010
rect 2030 7830 2090 8010
rect 2330 7830 2390 8010
rect 2620 7830 2680 8010
rect 2920 7830 2980 8010
rect 3400 8620 3460 8800
rect 3680 8620 3740 8800
rect 3980 8620 4040 8800
rect 4280 8620 4340 8800
rect 4580 8620 4640 8800
rect 4880 8620 4940 8800
rect 5160 8620 5220 8800
rect 5460 8620 5520 8800
rect 5760 8620 5820 8800
rect 6060 8620 6120 8800
rect 6340 8620 6400 8800
rect 3540 8360 3600 8520
rect 3840 8360 3900 8520
rect 4140 8360 4200 8520
rect 4440 8360 4500 8520
rect 4720 8360 4780 8520
rect 5020 8360 5080 8520
rect 5320 8360 5380 8520
rect 5600 8360 5660 8520
rect 5920 8360 5980 8520
rect 6200 8360 6260 8520
rect 3400 8100 3460 8260
rect 3700 8100 3760 8260
rect 3980 8100 4040 8260
rect 4280 8100 4340 8260
rect 4560 8100 4620 8260
rect 4880 8100 4940 8260
rect 5160 8100 5220 8260
rect 5460 8100 5520 8260
rect 5760 8100 5820 8260
rect 6060 8100 6120 8260
rect 6360 8100 6420 8260
rect 3540 7840 3600 8000
rect 3840 7840 3900 8000
rect 4140 7840 4200 8000
rect 4420 7840 4480 8000
rect 4720 7840 4780 8000
rect 5020 7840 5080 8000
rect 5320 7840 5380 8000
rect 5620 7840 5680 8000
rect 5920 7840 5980 8000
rect 6200 7840 6260 8000
rect 6680 8640 6740 8800
rect 6980 8640 7040 8800
rect 7280 8640 7340 8800
rect 7580 8640 7640 8800
rect 7880 8640 7940 8800
rect 8160 8640 8220 8800
rect 8460 8620 8520 8780
rect 8760 8620 8820 8780
rect 9040 8620 9100 8780
rect 9340 8620 9400 8780
rect 9640 8620 9700 8780
rect 6820 8360 6880 8520
rect 7120 8360 7180 8520
rect 7420 8360 7480 8520
rect 7720 8360 7780 8520
rect 8020 8360 8080 8520
rect 8320 8360 8380 8520
rect 8620 8360 8680 8520
rect 8920 8360 8980 8520
rect 9200 8360 9260 8520
rect 9500 8360 9560 8520
rect 6680 8100 6740 8260
rect 6980 8100 7040 8260
rect 7280 8100 7340 8260
rect 7580 8100 7640 8260
rect 7860 8100 7920 8260
rect 8160 8100 8220 8260
rect 8460 8100 8520 8260
rect 8760 8100 8820 8260
rect 9060 8100 9120 8260
rect 9340 8100 9400 8260
rect 9640 8100 9700 8260
rect 6840 7840 6900 8000
rect 7140 7840 7200 8000
rect 7420 7840 7480 8000
rect 7720 7840 7780 8000
rect 8020 7840 8080 8000
rect 8300 7840 8360 8000
rect 8620 7840 8680 8000
rect 8900 7840 8960 8000
rect 9200 7840 9260 8000
rect 9500 7840 9560 8000
rect 9980 8640 10040 8800
rect 10280 8640 10340 8800
rect 10580 8640 10640 8800
rect 10880 8640 10940 8800
rect 11160 8620 11220 8780
rect 11460 8620 11520 8780
rect 11760 8620 11820 8780
rect 12040 8620 12100 8780
rect 12360 8620 12420 8780
rect 12640 8620 12700 8780
rect 12940 8620 13000 8780
rect 10140 8360 10200 8520
rect 10420 8360 10480 8520
rect 10720 8360 10780 8520
rect 11020 8360 11080 8520
rect 11320 8360 11380 8520
rect 11600 8360 11660 8520
rect 11900 8360 11960 8520
rect 12200 8360 12260 8520
rect 12500 8360 12560 8520
rect 12800 8360 12860 8520
rect 9980 8100 10040 8260
rect 10280 8100 10340 8260
rect 10580 8100 10640 8260
rect 10860 8100 10920 8260
rect 11180 8100 11240 8260
rect 11460 8100 11520 8260
rect 11760 8100 11820 8260
rect 12060 8100 12120 8260
rect 12340 8100 12400 8260
rect 12640 8100 12700 8260
rect 12940 8100 13000 8260
rect 10140 7840 10200 8000
rect 10440 7840 10500 8000
rect 10720 7840 10780 8000
rect 11020 7840 11080 8000
rect 11320 7840 11380 8000
rect 11600 7840 11660 8000
rect 11900 7840 11960 8000
rect 12200 7840 12260 8000
rect 12500 7840 12560 8000
rect 12800 7840 12860 8000
rect 13280 8620 13340 8780
rect 13580 8620 13640 8780
rect 13860 8620 13920 8780
rect 14180 8620 14240 8780
rect 14460 8620 14520 8780
rect 14760 8620 14820 8780
rect 15040 8620 15100 8780
rect 15340 8620 15400 8780
rect 15640 8620 15700 8780
rect 15940 8620 16000 8780
rect 16240 8620 16300 8780
rect 16420 8620 16780 8780
rect 13420 8360 13480 8520
rect 13720 8360 13780 8520
rect 14000 8360 14060 8520
rect 14320 8360 14380 8520
rect 14600 8360 14660 8520
rect 14900 8360 14960 8520
rect 15200 8360 15260 8520
rect 15500 8360 15560 8520
rect 15780 8360 15840 8520
rect 16080 8360 16140 8520
rect 13280 8100 13340 8260
rect 13580 8100 13640 8260
rect 13860 8100 13920 8260
rect 14180 8100 14240 8260
rect 14460 8100 14520 8260
rect 14760 8100 14820 8260
rect 15060 8100 15120 8260
rect 15360 8100 15420 8260
rect 15640 8100 15700 8260
rect 15940 8100 16000 8260
rect 16240 8100 16300 8260
rect 16420 8100 16780 8260
rect 13420 7840 13480 8000
rect 13720 7840 13780 8000
rect 14020 7840 14080 8000
rect 14320 7840 14380 8000
rect 14600 7840 14660 8000
rect 14900 7840 14960 8000
rect 15200 7840 15260 8000
rect 15500 7840 15560 8000
rect 15800 7840 15860 8000
rect 16080 7840 16140 8000
rect 100 7120 160 7280
rect 400 7120 460 7280
rect 700 7120 760 7280
rect 980 7120 1040 7280
rect 1280 7120 1340 7280
rect 1580 7120 1640 7280
rect 1880 7120 1940 7280
rect 2180 7120 2240 7280
rect 2460 7120 2520 7280
rect 2780 7120 2840 7280
rect 3060 7120 3120 7280
rect 260 6860 320 7020
rect 560 6860 620 7020
rect 840 6860 900 7020
rect 1140 6860 1200 7020
rect 1420 6860 1480 7020
rect 1720 6860 1780 7020
rect 2040 6860 2100 7020
rect 2320 6860 2380 7020
rect 2620 6860 2680 7020
rect 2900 6860 2960 7020
rect 100 6340 160 6500
rect 380 6340 440 6500
rect 700 6340 760 6500
rect 1000 6340 1060 6500
rect 1280 6340 1340 6500
rect 1580 6340 1640 6500
rect 1880 6340 1940 6500
rect 2180 6340 2240 6500
rect 2480 6340 2540 6500
rect 2760 6340 2820 6500
rect 3060 6340 3120 6500
rect 3400 7120 3460 7280
rect 3680 7120 3740 7280
rect 3980 7120 4040 7280
rect 4280 7120 4340 7280
rect 4580 7120 4640 7280
rect 4880 7120 4940 7280
rect 5180 7120 5240 7280
rect 5460 7120 5520 7280
rect 5760 7120 5820 7280
rect 6060 7120 6120 7280
rect 6360 7120 6420 7280
rect 3540 6860 3600 7020
rect 3840 6860 3900 7020
rect 4120 6860 4180 7020
rect 4420 6860 4480 7020
rect 4720 6860 4780 7020
rect 5020 6860 5080 7020
rect 5320 6860 5380 7020
rect 5620 6860 5680 7020
rect 5900 6860 5960 7020
rect 6220 6860 6280 7020
rect 3400 6340 3460 6500
rect 3680 6340 3740 6500
rect 3980 6340 4040 6500
rect 4280 6340 4340 6500
rect 4580 6340 4640 6500
rect 4880 6340 4940 6500
rect 5160 6340 5220 6500
rect 5460 6340 5520 6500
rect 5760 6340 5820 6500
rect 6060 6340 6120 6500
rect 6360 6340 6420 6500
rect 6680 7120 6740 7280
rect 6980 7120 7040 7280
rect 7280 7120 7340 7280
rect 7580 7120 7640 7280
rect 7880 7120 7940 7280
rect 8160 7120 8220 7280
rect 8460 7120 8520 7280
rect 8760 7120 8820 7280
rect 9060 7120 9120 7280
rect 9340 7120 9400 7280
rect 9640 7120 9700 7280
rect 6840 6600 6900 6760
rect 7140 6600 7200 6760
rect 7420 6600 7480 6760
rect 7720 6600 7780 6760
rect 8020 6600 8080 6760
rect 8320 6600 8380 6760
rect 8620 6600 8680 6760
rect 8920 6600 8980 6760
rect 9200 6600 9260 6760
rect 9500 6600 9560 6760
rect 6680 6340 6740 6500
rect 6980 6340 7040 6500
rect 7280 6340 7340 6500
rect 7580 6340 7640 6500
rect 7880 6340 7940 6500
rect 8180 6340 8240 6500
rect 8460 6340 8520 6500
rect 8760 6340 8820 6500
rect 9060 6340 9120 6500
rect 9360 6340 9420 6500
rect 9640 6340 9700 6500
rect 9980 7120 10040 7280
rect 10280 7120 10340 7280
rect 10580 7120 10640 7280
rect 10880 7120 10940 7280
rect 11160 7120 11220 7280
rect 11460 7120 11520 7280
rect 11760 7120 11820 7280
rect 12060 7120 12120 7280
rect 12340 7120 12400 7280
rect 12660 7120 12720 7280
rect 12940 7120 13000 7280
rect 10140 6860 10200 7020
rect 10420 6860 10480 7020
rect 10720 6860 10780 7020
rect 11020 6860 11080 7020
rect 11320 6860 11380 7020
rect 11620 6860 11680 7020
rect 11920 6860 11980 7020
rect 12200 6860 12260 7020
rect 12500 6860 12560 7020
rect 12800 6860 12860 7020
rect 10000 6340 10060 6500
rect 10280 6340 10340 6500
rect 10560 6340 10620 6500
rect 10860 6340 10920 6500
rect 11160 6340 11220 6500
rect 11460 6340 11520 6500
rect 11760 6340 11820 6500
rect 12060 6340 12120 6500
rect 12340 6340 12400 6500
rect 12640 6340 12700 6500
rect 12940 6340 13000 6500
rect 13280 7120 13340 7280
rect 13560 7120 13620 7280
rect 13880 7120 13940 7280
rect 14160 7120 14220 7280
rect 14480 7120 14540 7280
rect 14760 7120 14820 7280
rect 15060 7120 15120 7280
rect 15340 7120 15400 7280
rect 15640 7120 15700 7280
rect 15940 7120 16000 7280
rect 16240 7120 16300 7280
rect 16420 7120 16780 7280
rect 13440 6860 13500 7020
rect 13720 6860 13780 7020
rect 14020 6860 14080 7020
rect 14300 6860 14360 7020
rect 14620 6860 14680 7020
rect 14920 6860 14980 7020
rect 15200 6860 15260 7020
rect 15500 6860 15560 7020
rect 15780 6860 15840 7020
rect 16080 6860 16140 7020
rect 13260 6340 13320 6500
rect 13560 6340 13620 6500
rect 13880 6340 13940 6500
rect 14160 6340 14220 6500
rect 14460 6340 14520 6500
rect 14740 6340 14800 6500
rect 15060 6340 15120 6500
rect 15340 6340 15400 6500
rect 15660 6340 15720 6500
rect 15940 6340 16000 6500
rect 16240 6340 16300 6500
rect 16420 6340 16780 6500
rect 100 5600 160 5760
rect 400 5600 460 5760
rect 680 5600 740 5760
rect 1000 5600 1060 5760
rect 1280 5600 1340 5760
rect 1580 5600 1640 5760
rect 1880 5600 1940 5760
rect 2180 5600 2240 5760
rect 2480 5600 2540 5760
rect 2760 5600 2820 5760
rect 3060 5600 3120 5760
rect 260 5340 320 5500
rect 560 5340 620 5500
rect 840 5340 900 5500
rect 1140 5340 1200 5500
rect 1440 5340 1500 5500
rect 1720 5340 1780 5500
rect 2040 5340 2100 5500
rect 2320 5340 2380 5500
rect 2620 5340 2680 5500
rect 2920 5340 2980 5500
rect 3400 5600 3460 5760
rect 3680 5600 3740 5760
rect 3980 5600 4040 5760
rect 4280 5600 4340 5760
rect 4580 5600 4640 5760
rect 4860 5600 4920 5760
rect 5160 5600 5220 5760
rect 5460 5600 5520 5760
rect 5760 5600 5820 5760
rect 6060 5600 6120 5760
rect 6360 5600 6420 5760
rect 3560 5080 3620 5240
rect 3840 5080 3900 5240
rect 4140 5080 4200 5240
rect 4420 5080 4480 5240
rect 4740 5080 4800 5240
rect 5020 5080 5080 5240
rect 5320 5080 5380 5240
rect 5620 5080 5680 5240
rect 5900 5080 5960 5240
rect 6200 5080 6260 5240
rect 3200 4820 3320 4980
rect 6680 5600 6740 5760
rect 6980 5600 7040 5760
rect 7280 5600 7340 5760
rect 7580 5600 7640 5760
rect 7880 5600 7940 5760
rect 8180 5600 8240 5760
rect 8460 5600 8520 5760
rect 8760 5600 8820 5760
rect 9060 5600 9120 5760
rect 9360 5600 9420 5760
rect 9660 5600 9720 5760
rect 6500 4820 6600 4980
rect 6840 4820 6900 4980
rect 7140 4820 7200 4980
rect 7440 4820 7500 4980
rect 7720 4820 7780 4980
rect 8020 4820 8080 4980
rect 8320 4820 8380 4980
rect 8600 4820 8660 4980
rect 8900 4820 8960 4980
rect 9200 4820 9260 4980
rect 9500 4820 9560 4980
rect 9980 5600 10040 5760
rect 10280 5600 10340 5760
rect 10580 5600 10640 5760
rect 10880 5600 10940 5760
rect 11160 5600 11220 5760
rect 11460 5600 11520 5760
rect 11760 5600 11820 5760
rect 12060 5600 12120 5760
rect 12340 5600 12400 5760
rect 12640 5600 12700 5760
rect 12940 5600 13000 5760
rect 10120 5080 10180 5240
rect 10420 5080 10480 5240
rect 10740 5080 10800 5240
rect 11020 5080 11080 5240
rect 11320 5080 11380 5240
rect 11600 5080 11660 5240
rect 11920 5080 11980 5240
rect 12200 5080 12260 5240
rect 12500 5080 12560 5240
rect 12800 5080 12860 5240
rect 9800 4820 9900 4980
rect 13280 5600 13340 5760
rect 13560 5600 13620 5760
rect 13880 5600 13940 5760
rect 14160 5600 14220 5760
rect 14460 5600 14520 5760
rect 14740 5600 14800 5760
rect 15060 5600 15120 5760
rect 15360 5600 15420 5760
rect 15640 5600 15700 5760
rect 15940 5600 16000 5760
rect 16240 5600 16300 5760
rect 16420 5600 16780 5760
rect 13440 5340 13500 5500
rect 13720 5340 13780 5500
rect 14020 5340 14080 5500
rect 14320 5340 14380 5500
rect 14600 5340 14660 5500
rect 14900 5340 14960 5500
rect 15200 5340 15260 5500
rect 15500 5340 15560 5500
rect 15800 5340 15860 5500
rect 16080 5340 16140 5500
rect 13080 4820 13180 4980
rect 100 4080 160 4240
rect 400 4080 460 4240
rect 680 4080 740 4240
rect 980 4080 1040 4240
rect 1280 4080 1340 4240
rect 1580 4080 1640 4240
rect 1880 4080 1940 4240
rect 2180 4080 2240 4240
rect 2460 4080 2520 4240
rect 2760 4080 2820 4240
rect 3060 4080 3120 4240
rect 240 3820 300 3980
rect 540 3820 600 3980
rect 840 3820 900 3980
rect 1140 3820 1200 3980
rect 1440 3820 1500 3980
rect 1740 3820 1800 3980
rect 2020 3820 2080 3980
rect 2320 3820 2380 3980
rect 2620 3820 2680 3980
rect 2900 3820 2960 3980
rect 100 3300 160 3460
rect 400 3300 460 3460
rect 680 3300 740 3460
rect 980 3300 1040 3460
rect 1280 3300 1340 3460
rect 1580 3300 1640 3460
rect 1860 3300 1920 3460
rect 2160 3300 2220 3460
rect 2480 3300 2540 3460
rect 2760 3300 2820 3460
rect 3060 3300 3120 3460
rect 3400 4080 3460 4240
rect 3680 4080 3740 4240
rect 3980 4080 4040 4240
rect 4280 4080 4340 4240
rect 4560 4080 4620 4240
rect 4860 4080 4920 4240
rect 5160 4080 5220 4240
rect 5460 4080 5520 4240
rect 5780 4080 5840 4240
rect 6060 4080 6120 4240
rect 6360 4080 6420 4240
rect 3540 3560 3600 3720
rect 3840 3560 3900 3720
rect 4140 3560 4200 3720
rect 4420 3560 4480 3720
rect 4720 3560 4780 3720
rect 5020 3560 5080 3720
rect 5320 3560 5380 3720
rect 5620 3560 5680 3720
rect 5920 3560 5980 3720
rect 6200 3560 6260 3720
rect 3400 3300 3460 3460
rect 3680 3300 3740 3460
rect 4000 3300 4060 3460
rect 4280 3300 4340 3460
rect 4580 3300 4640 3460
rect 4860 3300 4920 3460
rect 5160 3300 5220 3460
rect 5460 3300 5520 3460
rect 5760 3300 5820 3460
rect 6060 3300 6120 3460
rect 6360 3300 6420 3460
rect 6700 4080 6760 4240
rect 6980 4080 7040 4240
rect 7280 4080 7340 4240
rect 7580 4080 7640 4240
rect 7880 4080 7940 4240
rect 8160 4080 8220 4240
rect 8460 4080 8520 4240
rect 8760 4080 8820 4240
rect 9060 4080 9120 4240
rect 9340 4080 9400 4240
rect 9640 4080 9700 4240
rect 6840 3560 6900 3720
rect 7140 3560 7200 3720
rect 7440 3560 7500 3720
rect 7720 3560 7780 3720
rect 8020 3560 8080 3720
rect 8320 3560 8380 3720
rect 8620 3560 8680 3720
rect 8900 3560 8960 3720
rect 9200 3560 9260 3720
rect 9500 3560 9560 3720
rect 6680 3300 6740 3460
rect 6980 3300 7040 3460
rect 7280 3300 7340 3460
rect 7580 3300 7640 3460
rect 7880 3300 7940 3460
rect 8160 3300 8220 3460
rect 8460 3300 8520 3460
rect 8780 3300 8840 3460
rect 9060 3300 9120 3460
rect 9360 3300 9420 3460
rect 9660 3300 9720 3460
rect 9980 4080 10040 4240
rect 10280 4080 10340 4240
rect 10560 4080 10620 4240
rect 10860 4080 10920 4240
rect 11160 4080 11220 4240
rect 11460 4080 11520 4240
rect 11760 4080 11820 4240
rect 12060 4080 12120 4240
rect 12340 4080 12400 4240
rect 12640 4080 12700 4240
rect 12940 4080 13000 4240
rect 10140 3560 10200 3720
rect 10420 3560 10480 3720
rect 10720 3560 10780 3720
rect 11020 3560 11080 3720
rect 11320 3560 11380 3720
rect 11600 3560 11660 3720
rect 11900 3560 11960 3720
rect 12200 3560 12260 3720
rect 12500 3560 12560 3720
rect 12800 3560 12860 3720
rect 10000 3300 10060 3460
rect 10280 3300 10340 3460
rect 10580 3300 10640 3460
rect 10860 3300 10920 3460
rect 11180 3300 11240 3460
rect 11460 3300 11520 3460
rect 11760 3300 11820 3460
rect 12060 3300 12120 3460
rect 12360 3300 12420 3460
rect 12640 3300 12700 3460
rect 12940 3300 13000 3460
rect 13280 4080 13340 4240
rect 13560 4080 13620 4240
rect 13860 4080 13920 4240
rect 14160 4080 14220 4240
rect 14460 4080 14520 4240
rect 14760 4080 14820 4240
rect 15060 4080 15120 4240
rect 15360 4080 15420 4240
rect 15640 4080 15700 4240
rect 15940 4080 16000 4240
rect 16220 4080 16280 4240
rect 16420 4080 16780 4240
rect 13440 3820 13500 3980
rect 13720 3820 13780 3980
rect 14020 3820 14080 3980
rect 14320 3820 14380 3980
rect 14600 3820 14660 3980
rect 14900 3820 14960 3980
rect 15200 3820 15260 3980
rect 15500 3820 15560 3980
rect 15780 3820 15840 3980
rect 16080 3820 16140 3980
rect 13280 3300 13340 3460
rect 13560 3300 13620 3460
rect 13880 3300 13940 3460
rect 14180 3300 14240 3460
rect 14460 3300 14520 3460
rect 14740 3300 14800 3460
rect 15040 3300 15100 3460
rect 15360 3300 15420 3460
rect 15640 3300 15700 3460
rect 15940 3300 16000 3460
rect 16240 3300 16300 3460
rect 16420 3300 16780 3460
rect 100 2560 160 2720
rect 400 2560 460 2720
rect 680 2560 740 2720
rect 980 2560 1040 2720
rect 1300 2560 1360 2720
rect 1600 2560 1660 2720
rect 1880 2560 1940 2720
rect 2180 2560 2240 2720
rect 2460 2560 2520 2720
rect 2760 2560 2820 2720
rect 3060 2560 3120 2720
rect 260 2300 320 2460
rect 540 2300 600 2460
rect 840 2300 900 2460
rect 1140 2300 1200 2460
rect 1440 2300 1500 2460
rect 1740 2300 1800 2460
rect 2020 2300 2080 2460
rect 2320 2300 2380 2460
rect 2620 2300 2680 2460
rect 2900 2300 2960 2460
rect 100 1780 160 1940
rect 400 1780 460 1940
rect 680 1780 740 1940
rect 1000 1780 1060 1940
rect 1300 1780 1360 1940
rect 1600 1780 1660 1940
rect 1880 1780 1940 1940
rect 2180 1780 2240 1940
rect 2460 1780 2520 1940
rect 2760 1780 2820 1940
rect 3060 1780 3120 1940
rect 3400 2560 3460 2720
rect 3680 2560 3740 2720
rect 3980 2560 4040 2720
rect 4280 2560 4340 2720
rect 4580 2560 4640 2720
rect 4880 2560 4940 2720
rect 5160 2560 5220 2720
rect 5460 2560 5520 2720
rect 5760 2560 5820 2720
rect 6060 2560 6120 2720
rect 6360 2560 6420 2720
rect 3400 1780 3460 1940
rect 3680 1780 3740 1940
rect 3980 1780 4040 1940
rect 4280 1780 4340 1940
rect 4580 1780 4640 1940
rect 4880 1780 4940 1940
rect 5160 1780 5220 1940
rect 5460 1780 5520 1940
rect 5780 1780 5840 1940
rect 6060 1780 6120 1940
rect 6340 1780 6400 1940
rect 6680 2560 6740 2720
rect 6980 2560 7040 2720
rect 7280 2560 7340 2720
rect 7580 2560 7640 2720
rect 7880 2560 7940 2720
rect 8160 2560 8220 2720
rect 8460 2560 8520 2720
rect 8760 2560 8820 2720
rect 9040 2560 9100 2720
rect 9340 2560 9400 2720
rect 9640 2560 9700 2720
rect 6840 2040 6900 2200
rect 7140 2040 7200 2200
rect 7440 2040 7500 2200
rect 7720 2040 7780 2200
rect 8020 2040 8080 2200
rect 8320 2040 8380 2200
rect 8600 2040 8660 2200
rect 8900 2040 8960 2200
rect 9200 2040 9260 2200
rect 9500 2040 9560 2200
rect 6680 1780 6740 1940
rect 7000 1780 7060 1940
rect 7280 1780 7340 1940
rect 7580 1780 7640 1940
rect 7860 1780 7920 1940
rect 8180 1780 8240 1940
rect 8460 1780 8520 1940
rect 8760 1780 8820 1940
rect 9060 1780 9120 1940
rect 9340 1780 9400 1940
rect 9640 1780 9700 1940
rect 9980 2560 10040 2720
rect 10280 2560 10340 2720
rect 10560 2560 10620 2720
rect 10860 2560 10920 2720
rect 11160 2560 11220 2720
rect 11460 2560 11520 2720
rect 11760 2560 11820 2720
rect 12040 2560 12100 2720
rect 12340 2560 12400 2720
rect 12640 2560 12700 2720
rect 12940 2560 13000 2720
rect 10140 2300 10200 2460
rect 10420 2300 10480 2460
rect 10720 2300 10780 2460
rect 11020 2300 11080 2460
rect 11320 2300 11380 2460
rect 11600 2300 11660 2460
rect 11920 2300 11980 2460
rect 12200 2300 12260 2460
rect 12500 2300 12560 2460
rect 12800 2300 12860 2460
rect 10000 1780 10060 1940
rect 10280 1780 10340 1940
rect 10580 1780 10640 1940
rect 10880 1780 10940 1940
rect 11160 1780 11220 1940
rect 11460 1780 11520 1940
rect 11760 1780 11820 1940
rect 12060 1780 12120 1940
rect 12360 1780 12420 1940
rect 12640 1780 12700 1940
rect 12940 1780 13000 1940
rect 13280 2560 13340 2720
rect 13580 2560 13640 2720
rect 13860 2560 13920 2720
rect 14160 2560 14220 2720
rect 14460 2560 14520 2720
rect 14760 2560 14820 2720
rect 15060 2560 15120 2720
rect 15340 2560 15400 2720
rect 15640 2560 15700 2720
rect 15940 2560 16000 2720
rect 16240 2560 16300 2720
rect 16420 2560 16780 2720
rect 13440 2300 13500 2460
rect 13720 2300 13780 2460
rect 14020 2300 14080 2460
rect 14320 2300 14380 2460
rect 14620 2300 14680 2460
rect 14900 2300 14960 2460
rect 15200 2300 15260 2460
rect 15500 2300 15560 2460
rect 15800 2300 15860 2460
rect 16100 2300 16160 2460
rect 13280 1780 13340 1940
rect 13560 1780 13620 1940
rect 13880 1780 13940 1940
rect 14160 1780 14220 1940
rect 14460 1780 14520 1940
rect 14760 1780 14820 1940
rect 15060 1780 15120 1940
rect 15340 1780 15400 1940
rect 15640 1780 15700 1940
rect 15940 1780 16000 1940
rect 16240 1780 16300 1940
rect 16420 1780 16780 1940
rect 100 1030 160 1210
rect 400 1030 460 1210
rect 700 1030 760 1210
rect 1000 1030 1060 1210
rect 1280 1030 1340 1210
rect 1580 1030 1640 1210
rect 1880 1030 1940 1210
rect 2180 1030 2240 1210
rect 2480 1030 2540 1210
rect 2760 1030 2820 1210
rect 3060 1030 3120 1210
rect 240 770 300 950
rect 540 770 600 950
rect 840 770 900 950
rect 1140 770 1200 950
rect 1440 770 1500 950
rect 1740 770 1800 950
rect 2020 770 2080 950
rect 2320 770 2380 950
rect 2620 770 2680 950
rect 2920 770 2980 950
rect 120 510 180 690
rect 400 510 460 690
rect 680 510 740 690
rect 980 510 1040 690
rect 1300 510 1360 690
rect 1600 510 1660 690
rect 1880 510 1940 690
rect 2160 510 2220 690
rect 2480 510 2540 690
rect 2760 510 2820 690
rect 3060 510 3120 690
rect 240 250 300 430
rect 540 250 600 430
rect 840 250 900 430
rect 1140 250 1200 430
rect 1440 250 1500 430
rect 1740 250 1800 430
rect 2020 250 2080 430
rect 2340 250 2400 430
rect 2620 250 2680 430
rect 2920 250 2980 430
rect 3400 1030 3460 1210
rect 3680 1030 3740 1210
rect 4000 1030 4060 1210
rect 4280 1030 4340 1210
rect 4580 1030 4640 1210
rect 4880 1030 4940 1210
rect 5160 1030 5220 1210
rect 5460 1030 5520 1210
rect 5760 1030 5820 1210
rect 6060 1030 6120 1210
rect 6360 1030 6420 1210
rect 3540 770 3600 950
rect 3840 770 3900 950
rect 4140 770 4200 950
rect 4440 770 4500 950
rect 4720 770 4780 950
rect 5020 770 5080 950
rect 5320 770 5380 950
rect 5620 770 5680 950
rect 5900 770 5960 950
rect 6220 770 6280 950
rect 3400 510 3460 690
rect 3700 510 3760 690
rect 4000 510 4060 690
rect 4280 510 4340 690
rect 4580 510 4640 690
rect 4880 510 4940 690
rect 5180 510 5240 690
rect 5460 510 5520 690
rect 5760 510 5820 690
rect 6060 510 6120 690
rect 6360 510 6420 690
rect 3540 250 3600 430
rect 3840 250 3900 430
rect 4140 250 4200 430
rect 4440 250 4500 430
rect 4720 250 4780 430
rect 5020 250 5080 430
rect 5320 250 5380 430
rect 5620 250 5680 430
rect 5900 250 5960 430
rect 6220 250 6280 430
rect 6700 1030 6760 1210
rect 6980 1030 7040 1210
rect 7280 1030 7340 1210
rect 7580 1030 7640 1210
rect 7880 1030 7940 1210
rect 8180 1030 8240 1210
rect 8460 1030 8520 1210
rect 8760 1030 8820 1210
rect 9060 1030 9120 1210
rect 9360 1030 9420 1210
rect 9640 1030 9700 1210
rect 6840 770 6900 950
rect 7140 770 7200 950
rect 7420 770 7480 950
rect 7720 770 7780 950
rect 8020 770 8080 950
rect 8300 770 8360 950
rect 8620 770 8680 950
rect 8920 770 8980 950
rect 9220 770 9280 950
rect 9520 770 9580 950
rect 6700 510 6760 690
rect 7000 510 7060 690
rect 7280 510 7340 690
rect 7580 510 7640 690
rect 7860 510 7920 690
rect 8180 510 8240 690
rect 8480 510 8540 690
rect 8760 510 8820 690
rect 9060 510 9120 690
rect 9360 510 9420 690
rect 9660 510 9720 690
rect 6840 250 6900 430
rect 7140 250 7200 430
rect 7440 250 7500 430
rect 7720 250 7780 430
rect 8020 250 8080 430
rect 8320 250 8380 430
rect 8620 250 8680 430
rect 8920 250 8980 430
rect 9200 250 9260 430
rect 9520 250 9580 430
rect 9980 1030 10040 1210
rect 10280 1030 10340 1210
rect 10560 1030 10620 1210
rect 10860 1030 10920 1210
rect 11160 1030 11220 1210
rect 11460 1030 11520 1210
rect 11760 1030 11820 1210
rect 12060 1030 12120 1210
rect 12360 1030 12420 1210
rect 12660 1030 12720 1210
rect 12940 1030 13000 1210
rect 10140 770 10200 950
rect 10420 770 10480 950
rect 10740 770 10800 950
rect 11020 770 11080 950
rect 11320 770 11380 950
rect 11620 770 11680 950
rect 11920 770 11980 950
rect 12220 770 12280 950
rect 12500 770 12560 950
rect 12800 770 12860 950
rect 10000 510 10060 690
rect 10280 510 10340 690
rect 10580 510 10640 690
rect 10860 510 10920 690
rect 11160 510 11220 690
rect 11480 510 11540 690
rect 11760 510 11820 690
rect 12060 510 12120 690
rect 12360 510 12420 690
rect 12660 510 12720 690
rect 12940 510 13000 690
rect 10140 250 10200 430
rect 10440 250 10500 430
rect 10740 250 10800 430
rect 11020 250 11080 430
rect 11300 250 11360 430
rect 11600 250 11660 430
rect 11900 250 11960 430
rect 12220 250 12280 430
rect 12500 250 12560 430
rect 12800 250 12860 430
rect 13280 1030 13340 1210
rect 13580 1030 13640 1210
rect 13880 1030 13940 1210
rect 14180 1030 14240 1210
rect 14460 1030 14520 1210
rect 14760 1030 14820 1210
rect 15060 1030 15120 1210
rect 15360 1030 15420 1210
rect 15640 1030 15700 1210
rect 15960 1030 16020 1210
rect 16240 1030 16300 1210
rect 16420 1040 16780 1200
rect 13420 770 13480 950
rect 13740 770 13800 950
rect 14020 770 14080 950
rect 14300 770 14360 950
rect 14620 770 14680 950
rect 14920 770 14980 950
rect 15200 770 15260 950
rect 15500 770 15560 950
rect 15780 770 15840 950
rect 16100 770 16160 950
rect 13280 510 13340 690
rect 13580 510 13640 690
rect 13880 510 13940 690
rect 14160 510 14220 690
rect 14460 510 14520 690
rect 14760 510 14820 690
rect 15060 510 15120 690
rect 15360 510 15420 690
rect 15640 510 15700 690
rect 15940 510 16000 690
rect 16240 510 16300 690
rect 16420 520 16780 680
rect 13440 250 13500 430
rect 13740 250 13800 430
rect 14020 250 14080 430
rect 14320 250 14380 430
rect 14600 250 14660 430
rect 14900 250 14960 430
rect 15200 250 15260 430
rect 15500 250 15560 430
rect 15780 250 15840 430
rect 16100 250 16160 430
rect 16920 8360 17280 8520
rect 16920 6860 17280 7020
rect 16920 5340 17280 5500
rect 16920 3820 17280 3980
rect 16920 2300 17280 2460
rect 16920 780 17280 940
rect 16920 260 17280 420
rect 17420 6600 17780 6760
rect 17420 5080 17780 5240
rect 17420 3560 17780 3720
rect 17420 2040 17780 2200
rect 17920 4820 18280 4980
<< metal3 >>
rect 3390 8800 3470 8805
rect 3670 8800 3750 8805
rect 3970 8800 4050 8805
rect 4270 8800 4350 8805
rect 4570 8800 4650 8805
rect 4870 8800 4950 8805
rect 5150 8800 5230 8805
rect 5450 8800 5530 8805
rect 5750 8800 5830 8805
rect 6050 8800 6130 8805
rect 6330 8800 6410 8805
rect 6670 8800 6750 8805
rect 6970 8800 7050 8805
rect 7270 8800 7350 8805
rect 7570 8800 7650 8805
rect 7870 8800 7950 8805
rect 8150 8800 8230 8805
rect 9970 8800 10050 8805
rect 10270 8800 10350 8805
rect 10570 8800 10650 8805
rect 10870 8800 10950 8805
rect -40 8790 3400 8800
rect -40 8610 100 8790
rect 160 8610 400 8790
rect 460 8610 690 8790
rect 750 8610 990 8790
rect 1050 8610 1290 8790
rect 1350 8610 1590 8790
rect 1650 8610 1880 8790
rect 1940 8610 2170 8790
rect 2230 8610 2470 8790
rect 2530 8610 2760 8790
rect 2820 8610 3060 8790
rect 3120 8620 3400 8790
rect 3460 8620 3680 8800
rect 3740 8620 3980 8800
rect 4040 8620 4280 8800
rect 4340 8620 4580 8800
rect 4640 8620 4880 8800
rect 4940 8620 5160 8800
rect 5220 8620 5460 8800
rect 5520 8620 5760 8800
rect 5820 8620 6060 8800
rect 6120 8620 6340 8800
rect 6400 8640 6680 8800
rect 6740 8640 6980 8800
rect 7040 8640 7280 8800
rect 7340 8640 7580 8800
rect 7640 8640 7880 8800
rect 7940 8640 8160 8800
rect 8220 8780 9980 8800
rect 8220 8640 8460 8780
rect 6400 8620 8460 8640
rect 8520 8620 8760 8780
rect 8820 8620 9040 8780
rect 9100 8620 9340 8780
rect 9400 8620 9640 8780
rect 9700 8640 9980 8780
rect 10040 8640 10280 8800
rect 10340 8640 10580 8800
rect 10640 8640 10880 8800
rect 10940 8780 18300 8800
rect 10940 8640 11160 8780
rect 9700 8620 11160 8640
rect 11220 8620 11460 8780
rect 11520 8620 11760 8780
rect 11820 8620 12040 8780
rect 12100 8620 12360 8780
rect 12420 8620 12640 8780
rect 12700 8620 12940 8780
rect 13000 8620 13280 8780
rect 13340 8620 13580 8780
rect 13640 8620 13860 8780
rect 13920 8620 14180 8780
rect 14240 8620 14460 8780
rect 14520 8620 14760 8780
rect 14820 8620 15040 8780
rect 15100 8620 15340 8780
rect 15400 8620 15640 8780
rect 15700 8620 15940 8780
rect 16000 8620 16240 8780
rect 16300 8620 16420 8780
rect 16780 8620 18300 8780
rect 3120 8610 18300 8620
rect -40 8600 18300 8610
rect -40 8530 18300 8540
rect -40 8350 250 8530
rect 310 8350 550 8530
rect 610 8350 840 8530
rect 900 8350 1140 8530
rect 1200 8350 1440 8530
rect 1500 8350 1730 8530
rect 1790 8350 2030 8530
rect 2090 8350 2320 8530
rect 2380 8350 2620 8530
rect 2680 8350 2920 8530
rect 2980 8520 18300 8530
rect 2980 8360 3540 8520
rect 3600 8360 3840 8520
rect 3900 8360 4140 8520
rect 4200 8360 4440 8520
rect 4500 8360 4720 8520
rect 4780 8360 5020 8520
rect 5080 8360 5320 8520
rect 5380 8360 5600 8520
rect 5660 8360 5920 8520
rect 5980 8360 6200 8520
rect 6260 8360 6820 8520
rect 6880 8360 7120 8520
rect 7180 8360 7420 8520
rect 7480 8360 7720 8520
rect 7780 8360 8020 8520
rect 8080 8360 8320 8520
rect 8380 8360 8620 8520
rect 8680 8360 8920 8520
rect 8980 8360 9200 8520
rect 9260 8360 9500 8520
rect 9560 8360 10140 8520
rect 10200 8360 10420 8520
rect 10480 8360 10720 8520
rect 10780 8360 11020 8520
rect 11080 8360 11320 8520
rect 11380 8360 11600 8520
rect 11660 8360 11900 8520
rect 11960 8360 12200 8520
rect 12260 8360 12500 8520
rect 12560 8360 12800 8520
rect 12860 8360 13420 8520
rect 13480 8360 13720 8520
rect 13780 8360 14000 8520
rect 14060 8360 14320 8520
rect 14380 8360 14600 8520
rect 14660 8360 14900 8520
rect 14960 8360 15200 8520
rect 15260 8360 15500 8520
rect 15560 8360 15780 8520
rect 15840 8360 16080 8520
rect 16140 8360 16920 8520
rect 17280 8360 18300 8520
rect 2980 8350 18300 8360
rect -40 8340 18300 8350
rect -40 8270 18300 8280
rect -40 8090 100 8270
rect 160 8090 400 8270
rect 460 8090 690 8270
rect 750 8090 990 8270
rect 1050 8090 1290 8270
rect 1350 8090 1590 8270
rect 1650 8090 1880 8270
rect 1940 8090 2170 8270
rect 2230 8090 2470 8270
rect 2530 8090 2770 8270
rect 2830 8090 3060 8270
rect 3120 8260 18300 8270
rect 3120 8100 3400 8260
rect 3460 8100 3700 8260
rect 3760 8100 3980 8260
rect 4040 8100 4280 8260
rect 4340 8100 4560 8260
rect 4620 8100 4880 8260
rect 4940 8100 5160 8260
rect 5220 8100 5460 8260
rect 5520 8100 5760 8260
rect 5820 8100 6060 8260
rect 6120 8100 6360 8260
rect 6420 8100 6680 8260
rect 6740 8100 6980 8260
rect 7040 8100 7280 8260
rect 7340 8100 7580 8260
rect 7640 8100 7860 8260
rect 7920 8100 8160 8260
rect 8220 8100 8460 8260
rect 8520 8100 8760 8260
rect 8820 8100 9060 8260
rect 9120 8100 9340 8260
rect 9400 8100 9640 8260
rect 9700 8100 9980 8260
rect 10040 8100 10280 8260
rect 10340 8100 10580 8260
rect 10640 8100 10860 8260
rect 10920 8100 11180 8260
rect 11240 8100 11460 8260
rect 11520 8100 11760 8260
rect 11820 8100 12060 8260
rect 12120 8100 12340 8260
rect 12400 8100 12640 8260
rect 12700 8100 12940 8260
rect 13000 8100 13280 8260
rect 13340 8100 13580 8260
rect 13640 8100 13860 8260
rect 13920 8100 14180 8260
rect 14240 8100 14460 8260
rect 14520 8100 14760 8260
rect 14820 8100 15060 8260
rect 15120 8100 15360 8260
rect 15420 8100 15640 8260
rect 15700 8100 15940 8260
rect 16000 8100 16240 8260
rect 16300 8100 16420 8260
rect 16780 8100 18300 8260
rect 3120 8090 18300 8100
rect -40 8080 18300 8090
rect -40 8010 18300 8020
rect -40 7830 250 8010
rect 310 7830 540 8010
rect 600 7830 840 8010
rect 900 7830 1130 8010
rect 1190 7830 1430 8010
rect 1490 7830 1730 8010
rect 1790 7830 2030 8010
rect 2090 7830 2330 8010
rect 2390 7830 2620 8010
rect 2680 7830 2920 8010
rect 2980 8000 18300 8010
rect 2980 7840 3540 8000
rect 3600 7840 3840 8000
rect 3900 7840 4140 8000
rect 4200 7840 4420 8000
rect 4480 7840 4720 8000
rect 4780 7840 5020 8000
rect 5080 7840 5320 8000
rect 5380 7840 5620 8000
rect 5680 7840 5920 8000
rect 5980 7840 6200 8000
rect 6260 7840 6840 8000
rect 6900 7840 7140 8000
rect 7200 7840 7420 8000
rect 7480 7840 7720 8000
rect 7780 7840 8020 8000
rect 8080 7840 8300 8000
rect 8360 7840 8620 8000
rect 8680 7840 8900 8000
rect 8960 7840 9200 8000
rect 9260 7840 9500 8000
rect 9560 7840 10140 8000
rect 10200 7840 10440 8000
rect 10500 7840 10720 8000
rect 10780 7840 11020 8000
rect 11080 7840 11320 8000
rect 11380 7840 11600 8000
rect 11660 7840 11900 8000
rect 11960 7840 12200 8000
rect 12260 7840 12500 8000
rect 12560 7840 12800 8000
rect 12860 7840 13420 8000
rect 13480 7840 13720 8000
rect 13780 7840 14020 8000
rect 14080 7840 14320 8000
rect 14380 7840 14600 8000
rect 14660 7840 14900 8000
rect 14960 7840 15200 8000
rect 15260 7840 15500 8000
rect 15560 7840 15800 8000
rect 15860 7840 16080 8000
rect 16140 7840 18300 8000
rect 2980 7830 18300 7840
rect -40 7820 18300 7830
rect -40 7280 18300 7300
rect -40 7120 100 7280
rect 160 7120 400 7280
rect 460 7120 700 7280
rect 760 7120 980 7280
rect 1040 7120 1280 7280
rect 1340 7120 1580 7280
rect 1640 7120 1880 7280
rect 1940 7120 2180 7280
rect 2240 7120 2460 7280
rect 2520 7120 2780 7280
rect 2840 7120 3060 7280
rect 3120 7120 3400 7280
rect 3460 7120 3680 7280
rect 3740 7120 3980 7280
rect 4040 7120 4280 7280
rect 4340 7120 4580 7280
rect 4640 7120 4880 7280
rect 4940 7120 5180 7280
rect 5240 7120 5460 7280
rect 5520 7120 5760 7280
rect 5820 7120 6060 7280
rect 6120 7120 6360 7280
rect 6420 7120 6680 7280
rect 6740 7120 6980 7280
rect 7040 7120 7280 7280
rect 7340 7120 7580 7280
rect 7640 7120 7880 7280
rect 7940 7120 8160 7280
rect 8220 7120 8460 7280
rect 8520 7120 8760 7280
rect 8820 7120 9060 7280
rect 9120 7120 9340 7280
rect 9400 7120 9640 7280
rect 9700 7120 9980 7280
rect 10040 7120 10280 7280
rect 10340 7120 10580 7280
rect 10640 7120 10880 7280
rect 10940 7120 11160 7280
rect 11220 7120 11460 7280
rect 11520 7120 11760 7280
rect 11820 7120 12060 7280
rect 12120 7120 12340 7280
rect 12400 7120 12660 7280
rect 12720 7120 12940 7280
rect 13000 7120 13280 7280
rect 13340 7120 13560 7280
rect 13620 7120 13880 7280
rect 13940 7120 14160 7280
rect 14220 7120 14480 7280
rect 14540 7120 14760 7280
rect 14820 7120 15060 7280
rect 15120 7120 15340 7280
rect 15400 7120 15640 7280
rect 15700 7120 15940 7280
rect 16000 7120 16240 7280
rect 16300 7120 16420 7280
rect 16780 7120 18300 7280
rect -40 7100 18300 7120
rect -40 7020 18300 7040
rect -40 6860 260 7020
rect 320 6860 560 7020
rect 620 6860 840 7020
rect 900 6860 1140 7020
rect 1200 6860 1420 7020
rect 1480 6860 1720 7020
rect 1780 6860 2040 7020
rect 2100 6860 2320 7020
rect 2380 6860 2620 7020
rect 2680 6860 2900 7020
rect 2960 6860 3540 7020
rect 3600 6860 3840 7020
rect 3900 6860 4120 7020
rect 4180 6860 4420 7020
rect 4480 6860 4720 7020
rect 4780 6860 5020 7020
rect 5080 6860 5320 7020
rect 5380 6860 5620 7020
rect 5680 6860 5900 7020
rect 5960 6860 6220 7020
rect 6280 6860 10140 7020
rect 10200 6860 10420 7020
rect 10480 6860 10720 7020
rect 10780 6860 11020 7020
rect 11080 6860 11320 7020
rect 11380 6860 11620 7020
rect 11680 6860 11920 7020
rect 11980 6860 12200 7020
rect 12260 6860 12500 7020
rect 12560 6860 12800 7020
rect 12860 6860 13440 7020
rect 13500 6860 13720 7020
rect 13780 6860 14020 7020
rect 14080 6860 14300 7020
rect 14360 6860 14620 7020
rect 14680 6860 14920 7020
rect 14980 6860 15200 7020
rect 15260 6860 15500 7020
rect 15560 6860 15780 7020
rect 15840 6860 16080 7020
rect 16140 6860 16920 7020
rect 17280 6860 18300 7020
rect -40 6840 18300 6860
rect -40 6760 18300 6780
rect -40 6600 6840 6760
rect 6900 6600 7140 6760
rect 7200 6600 7420 6760
rect 7480 6600 7720 6760
rect 7780 6600 8020 6760
rect 8080 6600 8320 6760
rect 8380 6600 8620 6760
rect 8680 6600 8920 6760
rect 8980 6600 9200 6760
rect 9260 6600 9500 6760
rect 9560 6600 17420 6760
rect 17780 6600 18300 6760
rect -40 6580 18300 6600
rect -40 6500 18300 6520
rect -40 6340 100 6500
rect 160 6340 380 6500
rect 440 6340 700 6500
rect 760 6340 1000 6500
rect 1060 6340 1280 6500
rect 1340 6340 1580 6500
rect 1640 6340 1880 6500
rect 1940 6340 2180 6500
rect 2240 6340 2480 6500
rect 2540 6340 2760 6500
rect 2820 6340 3060 6500
rect 3120 6340 3400 6500
rect 3460 6340 3680 6500
rect 3740 6340 3980 6500
rect 4040 6340 4280 6500
rect 4340 6340 4580 6500
rect 4640 6340 4880 6500
rect 4940 6340 5160 6500
rect 5220 6340 5460 6500
rect 5520 6340 5760 6500
rect 5820 6340 6060 6500
rect 6120 6340 6360 6500
rect 6420 6340 6680 6500
rect 6740 6340 6980 6500
rect 7040 6340 7280 6500
rect 7340 6340 7580 6500
rect 7640 6340 7880 6500
rect 7940 6340 8180 6500
rect 8240 6340 8460 6500
rect 8520 6340 8760 6500
rect 8820 6340 9060 6500
rect 9120 6340 9360 6500
rect 9420 6340 9640 6500
rect 9700 6340 10000 6500
rect 10060 6340 10280 6500
rect 10340 6340 10560 6500
rect 10620 6340 10860 6500
rect 10920 6340 11160 6500
rect 11220 6340 11460 6500
rect 11520 6340 11760 6500
rect 11820 6340 12060 6500
rect 12120 6340 12340 6500
rect 12400 6340 12640 6500
rect 12700 6340 12940 6500
rect 13000 6340 13260 6500
rect 13320 6340 13560 6500
rect 13620 6340 13880 6500
rect 13940 6340 14160 6500
rect 14220 6340 14460 6500
rect 14520 6340 14740 6500
rect 14800 6340 15060 6500
rect 15120 6340 15340 6500
rect 15400 6340 15660 6500
rect 15720 6340 15940 6500
rect 16000 6340 16240 6500
rect 16300 6340 16420 6500
rect 16780 6340 18300 6500
rect -40 6320 18300 6340
rect -40 5760 18300 5780
rect -40 5600 100 5760
rect 160 5600 400 5760
rect 460 5600 680 5760
rect 740 5600 1000 5760
rect 1060 5600 1280 5760
rect 1340 5600 1580 5760
rect 1640 5600 1880 5760
rect 1940 5600 2180 5760
rect 2240 5600 2480 5760
rect 2540 5600 2760 5760
rect 2820 5600 3060 5760
rect 3120 5600 3400 5760
rect 3460 5600 3680 5760
rect 3740 5600 3980 5760
rect 4040 5600 4280 5760
rect 4340 5600 4580 5760
rect 4640 5600 4860 5760
rect 4920 5600 5160 5760
rect 5220 5600 5460 5760
rect 5520 5600 5760 5760
rect 5820 5600 6060 5760
rect 6120 5600 6360 5760
rect 6420 5600 6680 5760
rect 6740 5600 6980 5760
rect 7040 5600 7280 5760
rect 7340 5600 7580 5760
rect 7640 5600 7880 5760
rect 7940 5600 8180 5760
rect 8240 5600 8460 5760
rect 8520 5600 8760 5760
rect 8820 5600 9060 5760
rect 9120 5600 9360 5760
rect 9420 5600 9660 5760
rect 9720 5600 9980 5760
rect 10040 5600 10280 5760
rect 10340 5600 10580 5760
rect 10640 5600 10880 5760
rect 10940 5600 11160 5760
rect 11220 5600 11460 5760
rect 11520 5600 11760 5760
rect 11820 5600 12060 5760
rect 12120 5600 12340 5760
rect 12400 5600 12640 5760
rect 12700 5600 12940 5760
rect 13000 5600 13280 5760
rect 13340 5600 13560 5760
rect 13620 5600 13880 5760
rect 13940 5600 14160 5760
rect 14220 5600 14460 5760
rect 14520 5600 14740 5760
rect 14800 5600 15060 5760
rect 15120 5600 15360 5760
rect 15420 5600 15640 5760
rect 15700 5600 15940 5760
rect 16000 5600 16240 5760
rect 16300 5600 16420 5760
rect 16780 5600 18300 5760
rect -40 5580 18300 5600
rect -40 5500 18300 5520
rect -40 5340 260 5500
rect 320 5340 560 5500
rect 620 5340 840 5500
rect 900 5340 1140 5500
rect 1200 5340 1440 5500
rect 1500 5340 1720 5500
rect 1780 5340 2040 5500
rect 2100 5340 2320 5500
rect 2380 5340 2620 5500
rect 2680 5340 2920 5500
rect 2980 5340 13440 5500
rect 13500 5340 13720 5500
rect 13780 5340 14020 5500
rect 14080 5340 14320 5500
rect 14380 5340 14600 5500
rect 14660 5340 14900 5500
rect 14960 5340 15200 5500
rect 15260 5340 15500 5500
rect 15560 5340 15800 5500
rect 15860 5340 16080 5500
rect 16140 5340 16920 5500
rect 17280 5340 18300 5500
rect -40 5320 18300 5340
rect -40 5240 18300 5260
rect -40 5080 3560 5240
rect 3620 5080 3840 5240
rect 3900 5080 4140 5240
rect 4200 5080 4420 5240
rect 4480 5080 4740 5240
rect 4800 5080 5020 5240
rect 5080 5080 5320 5240
rect 5380 5080 5620 5240
rect 5680 5080 5900 5240
rect 5960 5080 6200 5240
rect 6260 5080 10120 5240
rect 10180 5080 10420 5240
rect 10480 5080 10740 5240
rect 10800 5080 11020 5240
rect 11080 5080 11320 5240
rect 11380 5080 11600 5240
rect 11660 5080 11920 5240
rect 11980 5080 12200 5240
rect 12260 5080 12500 5240
rect 12560 5080 12800 5240
rect 12860 5080 17420 5240
rect 17780 5080 18300 5240
rect -40 5060 18300 5080
rect -40 4980 18300 5000
rect -40 4820 3200 4980
rect 3320 4820 6500 4980
rect 6600 4820 6840 4980
rect 6900 4820 7140 4980
rect 7200 4820 7440 4980
rect 7500 4820 7720 4980
rect 7780 4820 8020 4980
rect 8080 4820 8320 4980
rect 8380 4820 8600 4980
rect 8660 4820 8900 4980
rect 8960 4820 9200 4980
rect 9260 4820 9500 4980
rect 9560 4820 9800 4980
rect 9900 4820 13080 4980
rect 13180 4820 17920 4980
rect 18280 4820 18300 4980
rect -40 4800 18300 4820
rect -40 4240 18300 4260
rect -40 4080 100 4240
rect 160 4080 400 4240
rect 460 4080 680 4240
rect 740 4080 980 4240
rect 1040 4080 1280 4240
rect 1340 4080 1580 4240
rect 1640 4080 1880 4240
rect 1940 4080 2180 4240
rect 2240 4080 2460 4240
rect 2520 4080 2760 4240
rect 2820 4080 3060 4240
rect 3120 4080 3400 4240
rect 3460 4080 3680 4240
rect 3740 4080 3980 4240
rect 4040 4080 4280 4240
rect 4340 4080 4560 4240
rect 4620 4080 4860 4240
rect 4920 4080 5160 4240
rect 5220 4080 5460 4240
rect 5520 4080 5780 4240
rect 5840 4080 6060 4240
rect 6120 4080 6360 4240
rect 6420 4080 6700 4240
rect 6760 4080 6980 4240
rect 7040 4080 7280 4240
rect 7340 4080 7580 4240
rect 7640 4080 7880 4240
rect 7940 4080 8160 4240
rect 8220 4080 8460 4240
rect 8520 4080 8760 4240
rect 8820 4080 9060 4240
rect 9120 4080 9340 4240
rect 9400 4080 9640 4240
rect 9700 4080 9980 4240
rect 10040 4080 10280 4240
rect 10340 4080 10560 4240
rect 10620 4080 10860 4240
rect 10920 4080 11160 4240
rect 11220 4080 11460 4240
rect 11520 4080 11760 4240
rect 11820 4080 12060 4240
rect 12120 4080 12340 4240
rect 12400 4080 12640 4240
rect 12700 4080 12940 4240
rect 13000 4080 13280 4240
rect 13340 4080 13560 4240
rect 13620 4080 13860 4240
rect 13920 4080 14160 4240
rect 14220 4080 14460 4240
rect 14520 4080 14760 4240
rect 14820 4080 15060 4240
rect 15120 4080 15360 4240
rect 15420 4080 15640 4240
rect 15700 4080 15940 4240
rect 16000 4080 16220 4240
rect 16280 4080 16420 4240
rect 16780 4080 18300 4240
rect -40 4060 18300 4080
rect -40 3980 18300 4000
rect -40 3820 240 3980
rect 300 3820 540 3980
rect 600 3820 840 3980
rect 900 3820 1140 3980
rect 1200 3820 1440 3980
rect 1500 3820 1740 3980
rect 1800 3820 2020 3980
rect 2080 3820 2320 3980
rect 2380 3820 2620 3980
rect 2680 3820 2900 3980
rect 2960 3820 13440 3980
rect 13500 3820 13720 3980
rect 13780 3820 14020 3980
rect 14080 3820 14320 3980
rect 14380 3820 14600 3980
rect 14660 3820 14900 3980
rect 14960 3820 15200 3980
rect 15260 3820 15500 3980
rect 15560 3820 15780 3980
rect 15840 3820 16080 3980
rect 16140 3820 16920 3980
rect 17280 3820 18300 3980
rect -40 3800 18300 3820
rect -40 3720 18300 3740
rect -40 3560 3540 3720
rect 3600 3560 3840 3720
rect 3900 3560 4140 3720
rect 4200 3560 4420 3720
rect 4480 3560 4720 3720
rect 4780 3560 5020 3720
rect 5080 3560 5320 3720
rect 5380 3560 5620 3720
rect 5680 3560 5920 3720
rect 5980 3560 6200 3720
rect 6260 3560 6840 3720
rect 6900 3560 7140 3720
rect 7200 3560 7440 3720
rect 7500 3560 7720 3720
rect 7780 3560 8020 3720
rect 8080 3560 8320 3720
rect 8380 3560 8620 3720
rect 8680 3560 8900 3720
rect 8960 3560 9200 3720
rect 9260 3560 9500 3720
rect 9560 3560 10140 3720
rect 10200 3560 10420 3720
rect 10480 3560 10720 3720
rect 10780 3560 11020 3720
rect 11080 3560 11320 3720
rect 11380 3560 11600 3720
rect 11660 3560 11900 3720
rect 11960 3560 12200 3720
rect 12260 3560 12500 3720
rect 12560 3560 12800 3720
rect 12860 3560 17420 3720
rect 17780 3560 18300 3720
rect -40 3540 18300 3560
rect -40 3460 18300 3480
rect -40 3300 100 3460
rect 160 3300 400 3460
rect 460 3300 680 3460
rect 740 3300 980 3460
rect 1040 3300 1280 3460
rect 1340 3300 1580 3460
rect 1640 3300 1860 3460
rect 1920 3300 2160 3460
rect 2220 3300 2480 3460
rect 2540 3300 2760 3460
rect 2820 3300 3060 3460
rect 3120 3300 3400 3460
rect 3460 3300 3680 3460
rect 3740 3300 4000 3460
rect 4060 3300 4280 3460
rect 4340 3300 4580 3460
rect 4640 3300 4860 3460
rect 4920 3300 5160 3460
rect 5220 3300 5460 3460
rect 5520 3300 5760 3460
rect 5820 3300 6060 3460
rect 6120 3300 6360 3460
rect 6420 3300 6680 3460
rect 6740 3300 6980 3460
rect 7040 3300 7280 3460
rect 7340 3300 7580 3460
rect 7640 3300 7880 3460
rect 7940 3300 8160 3460
rect 8220 3300 8460 3460
rect 8520 3300 8780 3460
rect 8840 3300 9060 3460
rect 9120 3300 9360 3460
rect 9420 3300 9660 3460
rect 9720 3300 10000 3460
rect 10060 3300 10280 3460
rect 10340 3300 10580 3460
rect 10640 3300 10860 3460
rect 10920 3300 11180 3460
rect 11240 3300 11460 3460
rect 11520 3300 11760 3460
rect 11820 3300 12060 3460
rect 12120 3300 12360 3460
rect 12420 3300 12640 3460
rect 12700 3300 12940 3460
rect 13000 3300 13280 3460
rect 13340 3300 13560 3460
rect 13620 3300 13880 3460
rect 13940 3300 14180 3460
rect 14240 3300 14460 3460
rect 14520 3300 14740 3460
rect 14800 3300 15040 3460
rect 15100 3300 15360 3460
rect 15420 3300 15640 3460
rect 15700 3300 15940 3460
rect 16000 3300 16240 3460
rect 16300 3300 16420 3460
rect 16780 3300 18300 3460
rect -40 3280 18300 3300
rect -40 2720 18300 2740
rect -40 2560 100 2720
rect 160 2560 400 2720
rect 460 2560 680 2720
rect 740 2560 980 2720
rect 1040 2560 1300 2720
rect 1360 2560 1600 2720
rect 1660 2560 1880 2720
rect 1940 2560 2180 2720
rect 2240 2560 2460 2720
rect 2520 2560 2760 2720
rect 2820 2560 3060 2720
rect 3120 2560 3400 2720
rect 3460 2560 3680 2720
rect 3740 2560 3980 2720
rect 4040 2560 4280 2720
rect 4340 2560 4580 2720
rect 4640 2560 4880 2720
rect 4940 2560 5160 2720
rect 5220 2560 5460 2720
rect 5520 2560 5760 2720
rect 5820 2560 6060 2720
rect 6120 2560 6360 2720
rect 6420 2560 6680 2720
rect 6740 2560 6980 2720
rect 7040 2560 7280 2720
rect 7340 2560 7580 2720
rect 7640 2560 7880 2720
rect 7940 2560 8160 2720
rect 8220 2560 8460 2720
rect 8520 2560 8760 2720
rect 8820 2560 9040 2720
rect 9100 2560 9340 2720
rect 9400 2560 9640 2720
rect 9700 2560 9980 2720
rect 10040 2560 10280 2720
rect 10340 2560 10560 2720
rect 10620 2560 10860 2720
rect 10920 2560 11160 2720
rect 11220 2560 11460 2720
rect 11520 2560 11760 2720
rect 11820 2560 12040 2720
rect 12100 2560 12340 2720
rect 12400 2560 12640 2720
rect 12700 2560 12940 2720
rect 13000 2560 13280 2720
rect 13340 2560 13580 2720
rect 13640 2560 13860 2720
rect 13920 2560 14160 2720
rect 14220 2560 14460 2720
rect 14520 2560 14760 2720
rect 14820 2560 15060 2720
rect 15120 2560 15340 2720
rect 15400 2560 15640 2720
rect 15700 2560 15940 2720
rect 16000 2560 16240 2720
rect 16300 2560 16420 2720
rect 16780 2560 18300 2720
rect -40 2540 18300 2560
rect -40 2460 18300 2480
rect -40 2300 260 2460
rect 320 2300 540 2460
rect 600 2300 840 2460
rect 900 2300 1140 2460
rect 1200 2300 1440 2460
rect 1500 2300 1740 2460
rect 1800 2300 2020 2460
rect 2080 2300 2320 2460
rect 2380 2300 2620 2460
rect 2680 2300 2900 2460
rect 2960 2300 10140 2460
rect 10200 2300 10420 2460
rect 10480 2300 10720 2460
rect 10780 2300 11020 2460
rect 11080 2300 11320 2460
rect 11380 2300 11600 2460
rect 11660 2300 11920 2460
rect 11980 2300 12200 2460
rect 12260 2300 12500 2460
rect 12560 2300 12800 2460
rect 12860 2300 13440 2460
rect 13500 2300 13720 2460
rect 13780 2300 14020 2460
rect 14080 2300 14320 2460
rect 14380 2300 14620 2460
rect 14680 2300 14900 2460
rect 14960 2300 15200 2460
rect 15260 2300 15500 2460
rect 15560 2300 15800 2460
rect 15860 2300 16100 2460
rect 16160 2300 16920 2460
rect 17280 2300 18300 2460
rect -40 2280 18300 2300
rect -40 2200 18300 2220
rect -40 2040 6840 2200
rect 6900 2040 7140 2200
rect 7200 2040 7440 2200
rect 7500 2040 7720 2200
rect 7780 2040 8020 2200
rect 8080 2040 8320 2200
rect 8380 2040 8600 2200
rect 8660 2040 8900 2200
rect 8960 2040 9200 2200
rect 9260 2040 9500 2200
rect 9560 2040 17420 2200
rect 17780 2040 18300 2200
rect -40 2020 18300 2040
rect -40 1940 18300 1960
rect -40 1780 100 1940
rect 160 1780 400 1940
rect 460 1780 680 1940
rect 740 1780 1000 1940
rect 1060 1780 1300 1940
rect 1360 1780 1600 1940
rect 1660 1780 1880 1940
rect 1940 1780 2180 1940
rect 2240 1780 2460 1940
rect 2520 1780 2760 1940
rect 2820 1780 3060 1940
rect 3120 1780 3400 1940
rect 3460 1780 3680 1940
rect 3740 1780 3980 1940
rect 4040 1780 4280 1940
rect 4340 1780 4580 1940
rect 4640 1780 4880 1940
rect 4940 1780 5160 1940
rect 5220 1780 5460 1940
rect 5520 1780 5780 1940
rect 5840 1780 6060 1940
rect 6120 1780 6340 1940
rect 6400 1780 6680 1940
rect 6740 1780 7000 1940
rect 7060 1780 7280 1940
rect 7340 1780 7580 1940
rect 7640 1780 7860 1940
rect 7920 1780 8180 1940
rect 8240 1780 8460 1940
rect 8520 1780 8760 1940
rect 8820 1780 9060 1940
rect 9120 1780 9340 1940
rect 9400 1780 9640 1940
rect 9700 1780 10000 1940
rect 10060 1780 10280 1940
rect 10340 1780 10580 1940
rect 10640 1780 10880 1940
rect 10940 1780 11160 1940
rect 11220 1780 11460 1940
rect 11520 1780 11760 1940
rect 11820 1780 12060 1940
rect 12120 1780 12360 1940
rect 12420 1780 12640 1940
rect 12700 1780 12940 1940
rect 13000 1780 13280 1940
rect 13340 1780 13560 1940
rect 13620 1780 13880 1940
rect 13940 1780 14160 1940
rect 14220 1780 14460 1940
rect 14520 1780 14760 1940
rect 14820 1780 15060 1940
rect 15120 1780 15340 1940
rect 15400 1780 15640 1940
rect 15700 1780 15940 1940
rect 16000 1780 16240 1940
rect 16300 1780 16420 1940
rect 16780 1780 18300 1940
rect -40 1760 18300 1780
rect -40 1210 18300 1220
rect -40 1030 100 1210
rect 160 1030 400 1210
rect 460 1030 700 1210
rect 760 1030 1000 1210
rect 1060 1030 1280 1210
rect 1340 1030 1580 1210
rect 1640 1030 1880 1210
rect 1940 1030 2180 1210
rect 2240 1030 2480 1210
rect 2540 1030 2760 1210
rect 2820 1030 3060 1210
rect 3120 1030 3400 1210
rect 3460 1030 3680 1210
rect 3740 1030 4000 1210
rect 4060 1030 4280 1210
rect 4340 1030 4580 1210
rect 4640 1030 4880 1210
rect 4940 1030 5160 1210
rect 5220 1030 5460 1210
rect 5520 1030 5760 1210
rect 5820 1030 6060 1210
rect 6120 1030 6360 1210
rect 6420 1030 6700 1210
rect 6760 1030 6980 1210
rect 7040 1030 7280 1210
rect 7340 1030 7580 1210
rect 7640 1030 7880 1210
rect 7940 1030 8180 1210
rect 8240 1030 8460 1210
rect 8520 1030 8760 1210
rect 8820 1030 9060 1210
rect 9120 1030 9360 1210
rect 9420 1030 9640 1210
rect 9700 1030 9980 1210
rect 10040 1030 10280 1210
rect 10340 1030 10560 1210
rect 10620 1030 10860 1210
rect 10920 1030 11160 1210
rect 11220 1030 11460 1210
rect 11520 1030 11760 1210
rect 11820 1030 12060 1210
rect 12120 1030 12360 1210
rect 12420 1030 12660 1210
rect 12720 1030 12940 1210
rect 13000 1030 13280 1210
rect 13340 1030 13580 1210
rect 13640 1030 13880 1210
rect 13940 1030 14180 1210
rect 14240 1030 14460 1210
rect 14520 1030 14760 1210
rect 14820 1030 15060 1210
rect 15120 1030 15360 1210
rect 15420 1030 15640 1210
rect 15700 1030 15960 1210
rect 16020 1030 16240 1210
rect 16300 1200 18300 1210
rect 16300 1040 16420 1200
rect 16780 1040 18300 1200
rect 16300 1030 18300 1040
rect -40 1020 18300 1030
rect -40 950 18300 960
rect -40 770 240 950
rect 300 770 540 950
rect 600 770 840 950
rect 900 770 1140 950
rect 1200 770 1440 950
rect 1500 770 1740 950
rect 1800 770 2020 950
rect 2080 770 2320 950
rect 2380 770 2620 950
rect 2680 770 2920 950
rect 2980 770 3540 950
rect 3600 770 3840 950
rect 3900 770 4140 950
rect 4200 770 4440 950
rect 4500 770 4720 950
rect 4780 770 5020 950
rect 5080 770 5320 950
rect 5380 770 5620 950
rect 5680 770 5900 950
rect 5960 770 6220 950
rect 6280 770 6840 950
rect 6900 770 7140 950
rect 7200 770 7420 950
rect 7480 770 7720 950
rect 7780 770 8020 950
rect 8080 770 8300 950
rect 8360 770 8620 950
rect 8680 770 8920 950
rect 8980 770 9220 950
rect 9280 770 9520 950
rect 9580 770 10140 950
rect 10200 770 10420 950
rect 10480 770 10740 950
rect 10800 770 11020 950
rect 11080 770 11320 950
rect 11380 770 11620 950
rect 11680 770 11920 950
rect 11980 770 12220 950
rect 12280 770 12500 950
rect 12560 770 12800 950
rect 12860 770 13420 950
rect 13480 770 13740 950
rect 13800 770 14020 950
rect 14080 770 14300 950
rect 14360 770 14620 950
rect 14680 770 14920 950
rect 14980 770 15200 950
rect 15260 770 15500 950
rect 15560 770 15780 950
rect 15840 770 16100 950
rect 16160 940 18300 950
rect 16160 780 16920 940
rect 17280 780 18300 940
rect 16160 770 18300 780
rect -40 760 18300 770
rect -40 690 18300 700
rect -40 510 120 690
rect 180 510 400 690
rect 460 510 680 690
rect 740 510 980 690
rect 1040 510 1300 690
rect 1360 510 1600 690
rect 1660 510 1880 690
rect 1940 510 2160 690
rect 2220 510 2480 690
rect 2540 510 2760 690
rect 2820 510 3060 690
rect 3120 510 3400 690
rect 3460 510 3700 690
rect 3760 510 4000 690
rect 4060 510 4280 690
rect 4340 510 4580 690
rect 4640 510 4880 690
rect 4940 510 5180 690
rect 5240 510 5460 690
rect 5520 510 5760 690
rect 5820 510 6060 690
rect 6120 510 6360 690
rect 6420 510 6700 690
rect 6760 510 7000 690
rect 7060 510 7280 690
rect 7340 510 7580 690
rect 7640 510 7860 690
rect 7920 510 8180 690
rect 8240 510 8480 690
rect 8540 510 8760 690
rect 8820 510 9060 690
rect 9120 510 9360 690
rect 9420 510 9660 690
rect 9720 510 10000 690
rect 10060 510 10280 690
rect 10340 510 10580 690
rect 10640 510 10860 690
rect 10920 510 11160 690
rect 11220 510 11480 690
rect 11540 510 11760 690
rect 11820 510 12060 690
rect 12120 510 12360 690
rect 12420 510 12660 690
rect 12720 510 12940 690
rect 13000 510 13280 690
rect 13340 510 13580 690
rect 13640 510 13880 690
rect 13940 510 14160 690
rect 14220 510 14460 690
rect 14520 510 14760 690
rect 14820 510 15060 690
rect 15120 510 15360 690
rect 15420 510 15640 690
rect 15700 510 15940 690
rect 16000 510 16240 690
rect 16300 680 18300 690
rect 16300 520 16420 680
rect 16780 520 18300 680
rect 16300 510 18300 520
rect -40 500 18300 510
rect -40 430 18300 440
rect -40 250 240 430
rect 300 250 540 430
rect 600 250 840 430
rect 900 250 1140 430
rect 1200 250 1440 430
rect 1500 250 1740 430
rect 1800 250 2020 430
rect 2080 250 2340 430
rect 2400 250 2620 430
rect 2680 250 2920 430
rect 2980 250 3540 430
rect 3600 250 3840 430
rect 3900 250 4140 430
rect 4200 250 4440 430
rect 4500 250 4720 430
rect 4780 250 5020 430
rect 5080 250 5320 430
rect 5380 250 5620 430
rect 5680 250 5900 430
rect 5960 250 6220 430
rect 6280 250 6840 430
rect 6900 250 7140 430
rect 7200 250 7440 430
rect 7500 250 7720 430
rect 7780 250 8020 430
rect 8080 250 8320 430
rect 8380 250 8620 430
rect 8680 250 8920 430
rect 8980 250 9200 430
rect 9260 250 9520 430
rect 9580 250 10140 430
rect 10200 250 10440 430
rect 10500 250 10740 430
rect 10800 250 11020 430
rect 11080 250 11300 430
rect 11360 250 11600 430
rect 11660 250 11900 430
rect 11960 250 12220 430
rect 12280 250 12500 430
rect 12560 250 12800 430
rect 12860 250 13440 430
rect 13500 250 13740 430
rect 13800 250 14020 430
rect 14080 250 14320 430
rect 14380 250 14600 430
rect 14660 250 14900 430
rect 14960 250 15200 430
rect 15260 250 15500 430
rect 15560 250 15780 430
rect 15840 250 16100 430
rect 16160 420 18300 430
rect 16160 260 16920 420
rect 17280 260 18300 420
rect 16160 250 18300 260
rect -40 240 18300 250
use sky130_fd_pr__pfet_01v8_9CZQJE  sky130_fd_pr__pfet_01v8_9CZQJE_0
array 0 4 3294 0 5 1518
timestamp 1619109957
transform 1 0 1612 0 1 694
box -1647 -759 1647 759
<< labels >>
rlabel metal2 16900 7020 17300 8360 1 iout
rlabel metal2 17900 4980 18300 8800 1 iref
rlabel metal2 16400 1940 16800 2560 1 vdd
rlabel metal2 17400 5240 17800 6600 1 idif
rlabel metal2 16400 7600 16800 8100 1 vdd
rlabel metal2 17400 6760 17800 8800 1 idif
<< end >>
