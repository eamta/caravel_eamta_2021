magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 2083 2689 2241 2748
rect 3557 2689 3715 2748
rect 5031 2689 5189 2748
rect 6505 2689 6663 2748
rect 7979 2689 8137 2748
rect 9453 2689 9611 2748
rect 10927 2689 11003 2748
rect 2021 2688 2303 2689
rect 3495 2688 3777 2689
rect 4969 2688 5251 2689
rect 6443 2688 6725 2689
rect 7917 2688 8199 2689
rect 9391 2688 9673 2689
rect 10865 2688 11003 2689
rect 2303 2655 2336 2680
rect 3777 2655 3810 2680
rect 5251 2655 5284 2680
rect 6725 2655 6758 2680
rect 8199 2655 8232 2680
rect 9673 2655 9706 2680
rect 2021 2654 2336 2655
rect 3495 2654 3810 2655
rect 4969 2654 5284 2655
rect 6443 2654 6758 2655
rect 7917 2654 8232 2655
rect 9391 2654 9706 2655
rect 10865 2654 11003 2655
rect 2028 2592 2055 2626
rect 2118 2615 2206 2626
rect 2129 2603 2195 2615
rect 2118 2593 2206 2603
rect 2269 2593 2282 2615
rect 2118 2592 2282 2593
rect 604 2524 662 2530
rect 604 2490 616 2524
rect 604 2484 662 2490
rect 1342 2418 1400 2424
rect 774 2369 808 2387
rect 1196 2369 1230 2387
rect 1342 2384 1354 2418
rect 1342 2378 1400 2384
rect 774 2333 844 2369
rect 791 2299 862 2333
rect 604 1952 662 1958
rect 604 1918 616 1952
rect 604 1912 662 1918
rect 791 1858 861 2299
rect 973 2231 1031 2237
rect 973 2197 985 2231
rect 973 2191 1031 2197
rect 973 1899 1031 1905
rect 973 1865 985 1899
rect 973 1859 1031 1865
rect 458 1850 492 1858
rect 774 1850 861 1858
rect 458 1840 861 1850
rect 1160 1840 1230 2369
rect 1953 2281 1966 2592
rect 1512 2263 1546 2281
rect 1932 2263 1966 2281
rect 1512 2227 1582 2263
rect 1529 2193 1600 2227
rect 1896 2214 1966 2263
rect 1987 2497 2020 2592
rect 2145 2586 2179 2592
rect 2129 2570 2182 2582
rect 2147 2558 2177 2570
rect 2101 2539 2177 2558
rect 2214 2539 2223 2543
rect 1987 2222 2021 2497
rect 2089 2490 2158 2539
rect 2089 2474 2140 2490
rect 2089 2459 2135 2474
rect 2189 2471 2202 2481
rect 2046 2443 2055 2447
rect 2067 2443 2080 2447
rect 2092 2443 2135 2459
rect 2183 2469 2202 2471
rect 2034 2343 2086 2443
rect 2095 2431 2135 2443
rect 2155 2443 2168 2447
rect 2155 2442 2174 2443
rect 2147 2431 2174 2442
rect 2095 2383 2174 2431
rect 2095 2371 2114 2383
rect 2101 2367 2114 2371
rect 2134 2371 2174 2383
rect 2183 2383 2206 2469
rect 2183 2371 2202 2383
rect 2134 2358 2177 2371
rect 2111 2355 2177 2358
rect 2179 2355 2180 2371
rect 2189 2367 2202 2371
rect 2214 2371 2235 2539
rect 2214 2367 2223 2371
rect 2248 2369 2282 2592
rect 2303 2369 2336 2654
rect 3502 2592 3529 2626
rect 3592 2615 3680 2626
rect 3603 2603 3669 2615
rect 3592 2593 3680 2603
rect 3743 2593 3756 2615
rect 3592 2592 3756 2593
rect 2816 2418 2874 2424
rect 2670 2369 2704 2387
rect 2816 2384 2828 2418
rect 2816 2378 2874 2384
rect 2034 2333 2080 2343
rect 2034 2222 2075 2333
rect 2111 2324 2180 2355
rect 2248 2333 2373 2369
rect 2129 2290 2202 2324
rect 2129 2274 2180 2290
rect 2165 2259 2180 2274
rect 2265 2256 2373 2333
rect 2134 2222 2168 2256
rect 2248 2222 2373 2256
rect 1987 2214 2373 2222
rect 458 1816 1230 1840
rect 1342 1846 1400 1852
rect 1342 1838 1354 1846
rect 1529 1840 1599 2193
rect 1896 2152 2373 2214
rect 2447 2231 2505 2237
rect 2447 2197 2459 2231
rect 2447 2191 2505 2197
rect 1896 2144 2335 2152
rect 1711 2125 1769 2131
rect 1711 2091 1723 2125
rect 1711 2085 1769 2091
rect 1896 2082 2336 2144
rect 1896 1858 2337 2082
rect 2447 1899 2505 1905
rect 2447 1865 2459 1899
rect 2447 1859 2505 1865
rect 1881 1842 2337 1858
rect 1881 1840 2336 1842
rect 2634 1840 2704 2369
rect 3427 2281 3440 2592
rect 2986 2263 3020 2281
rect 3406 2263 3440 2281
rect 2986 2227 3056 2263
rect 3003 2193 3074 2227
rect 3370 2214 3440 2263
rect 3461 2497 3494 2592
rect 3619 2586 3653 2592
rect 3603 2570 3656 2582
rect 3621 2558 3651 2570
rect 3575 2539 3651 2558
rect 3688 2539 3697 2543
rect 3461 2222 3495 2497
rect 3563 2490 3632 2539
rect 3563 2474 3614 2490
rect 3563 2459 3609 2474
rect 3663 2471 3676 2481
rect 3520 2443 3529 2447
rect 3541 2443 3554 2447
rect 3566 2443 3609 2459
rect 3657 2469 3676 2471
rect 3508 2343 3560 2443
rect 3569 2431 3609 2443
rect 3629 2443 3642 2447
rect 3629 2442 3648 2443
rect 3621 2431 3648 2442
rect 3569 2383 3648 2431
rect 3569 2371 3588 2383
rect 3575 2367 3588 2371
rect 3608 2371 3648 2383
rect 3657 2383 3680 2469
rect 3657 2371 3676 2383
rect 3608 2358 3651 2371
rect 3585 2355 3651 2358
rect 3653 2355 3654 2371
rect 3663 2367 3676 2371
rect 3688 2371 3709 2539
rect 3688 2367 3697 2371
rect 3722 2369 3756 2592
rect 3777 2369 3810 2654
rect 4976 2592 5003 2626
rect 5066 2615 5154 2626
rect 5077 2603 5143 2615
rect 5066 2593 5154 2603
rect 5217 2593 5230 2615
rect 5066 2592 5230 2593
rect 4290 2418 4348 2424
rect 4144 2369 4178 2387
rect 4290 2384 4302 2418
rect 4290 2378 4348 2384
rect 3508 2333 3554 2343
rect 3508 2222 3549 2333
rect 3585 2324 3654 2355
rect 3722 2333 3847 2369
rect 3603 2290 3676 2324
rect 3603 2274 3654 2290
rect 3639 2259 3654 2274
rect 3739 2256 3847 2333
rect 3608 2222 3642 2256
rect 3722 2222 3847 2256
rect 3461 2214 3847 2222
rect 791 1804 1230 1816
rect 1338 1812 1404 1838
rect 1342 1806 1400 1812
rect 1529 1804 2704 1840
rect 2816 1846 2874 1852
rect 2816 1838 2828 1846
rect 3003 1840 3073 2193
rect 3370 2152 3847 2214
rect 3921 2231 3979 2237
rect 3921 2197 3933 2231
rect 3921 2191 3979 2197
rect 3370 2144 3809 2152
rect 3185 2125 3243 2131
rect 3185 2091 3197 2125
rect 3185 2085 3243 2091
rect 3370 2082 3810 2144
rect 3370 1858 3811 2082
rect 3921 1899 3979 1905
rect 3921 1865 3933 1899
rect 3921 1859 3979 1865
rect 3355 1842 3811 1858
rect 3355 1840 3810 1842
rect 4108 1840 4178 2369
rect 4901 2281 4914 2592
rect 4460 2263 4494 2281
rect 4880 2263 4914 2281
rect 4460 2227 4530 2263
rect 4477 2193 4548 2227
rect 4844 2214 4914 2263
rect 4935 2497 4968 2592
rect 5093 2586 5127 2592
rect 5077 2570 5130 2582
rect 5095 2558 5125 2570
rect 5049 2539 5125 2558
rect 5162 2539 5171 2543
rect 4935 2222 4969 2497
rect 5037 2490 5106 2539
rect 5037 2474 5088 2490
rect 5037 2459 5083 2474
rect 5137 2471 5150 2481
rect 4994 2443 5003 2447
rect 5015 2443 5028 2447
rect 5040 2443 5083 2459
rect 5131 2469 5150 2471
rect 4982 2343 5034 2443
rect 5043 2431 5083 2443
rect 5103 2443 5116 2447
rect 5103 2442 5122 2443
rect 5095 2431 5122 2442
rect 5043 2383 5122 2431
rect 5043 2371 5062 2383
rect 5049 2367 5062 2371
rect 5082 2371 5122 2383
rect 5131 2383 5154 2469
rect 5131 2371 5150 2383
rect 5082 2358 5125 2371
rect 5059 2355 5125 2358
rect 5127 2355 5128 2371
rect 5137 2367 5150 2371
rect 5162 2371 5183 2539
rect 5162 2367 5171 2371
rect 5196 2369 5230 2592
rect 5251 2369 5284 2654
rect 6450 2592 6477 2626
rect 6540 2615 6628 2626
rect 6551 2603 6617 2615
rect 6540 2593 6628 2603
rect 6691 2593 6704 2615
rect 6540 2592 6704 2593
rect 5764 2418 5822 2424
rect 5618 2369 5652 2387
rect 5764 2384 5776 2418
rect 5764 2378 5822 2384
rect 4982 2333 5028 2343
rect 4982 2222 5023 2333
rect 5059 2324 5128 2355
rect 5196 2333 5321 2369
rect 5077 2290 5150 2324
rect 5077 2274 5128 2290
rect 5113 2259 5128 2274
rect 5213 2256 5321 2333
rect 5082 2222 5116 2256
rect 5196 2222 5321 2256
rect 4935 2214 5321 2222
rect 2812 1812 2878 1838
rect 2816 1806 2874 1812
rect 3003 1804 4178 1840
rect 4290 1846 4348 1852
rect 4290 1838 4302 1846
rect 4477 1840 4547 2193
rect 4844 2152 5321 2214
rect 5395 2231 5453 2237
rect 5395 2197 5407 2231
rect 5395 2191 5453 2197
rect 4844 2144 5283 2152
rect 4659 2125 4717 2131
rect 4659 2091 4671 2125
rect 4659 2085 4717 2091
rect 4844 2082 5284 2144
rect 4844 1858 5285 2082
rect 5395 1899 5453 1905
rect 5395 1865 5407 1899
rect 5395 1859 5453 1865
rect 4829 1842 5285 1858
rect 4829 1840 5284 1842
rect 5582 1840 5652 2369
rect 6375 2281 6388 2592
rect 5934 2263 5968 2281
rect 6354 2263 6388 2281
rect 5934 2227 6004 2263
rect 5951 2193 6022 2227
rect 6318 2214 6388 2263
rect 6409 2497 6442 2592
rect 6567 2586 6601 2592
rect 6551 2570 6604 2582
rect 6569 2558 6599 2570
rect 6523 2539 6599 2558
rect 6636 2539 6645 2543
rect 6409 2222 6443 2497
rect 6511 2490 6580 2539
rect 6511 2474 6562 2490
rect 6511 2459 6557 2474
rect 6611 2471 6624 2481
rect 6468 2443 6477 2447
rect 6489 2443 6502 2447
rect 6514 2443 6557 2459
rect 6605 2469 6624 2471
rect 6456 2343 6508 2443
rect 6517 2431 6557 2443
rect 6577 2443 6590 2447
rect 6577 2442 6596 2443
rect 6569 2431 6596 2442
rect 6517 2383 6596 2431
rect 6517 2371 6536 2383
rect 6523 2367 6536 2371
rect 6556 2371 6596 2383
rect 6605 2383 6628 2469
rect 6605 2371 6624 2383
rect 6556 2358 6599 2371
rect 6533 2355 6599 2358
rect 6601 2355 6602 2371
rect 6611 2367 6624 2371
rect 6636 2371 6657 2539
rect 6636 2367 6645 2371
rect 6670 2369 6704 2592
rect 6725 2369 6758 2654
rect 7924 2592 7951 2626
rect 8014 2615 8102 2626
rect 8025 2603 8091 2615
rect 8014 2593 8102 2603
rect 8165 2593 8178 2615
rect 8014 2592 8178 2593
rect 7238 2418 7296 2424
rect 7092 2369 7126 2387
rect 7238 2384 7250 2418
rect 7238 2378 7296 2384
rect 6456 2333 6502 2343
rect 6456 2222 6497 2333
rect 6533 2324 6602 2355
rect 6670 2333 6795 2369
rect 6551 2290 6624 2324
rect 6551 2274 6602 2290
rect 6587 2259 6602 2274
rect 6687 2256 6795 2333
rect 6556 2222 6590 2256
rect 6670 2222 6795 2256
rect 6409 2214 6795 2222
rect 4286 1812 4352 1838
rect 4290 1806 4348 1812
rect 4477 1804 5652 1840
rect 5764 1846 5822 1852
rect 5764 1838 5776 1846
rect 5951 1840 6021 2193
rect 6318 2152 6795 2214
rect 6869 2231 6927 2237
rect 6869 2197 6881 2231
rect 6869 2191 6927 2197
rect 6318 2144 6757 2152
rect 6133 2125 6191 2131
rect 6133 2091 6145 2125
rect 6133 2085 6191 2091
rect 6318 2082 6758 2144
rect 6318 1858 6759 2082
rect 6869 1899 6927 1905
rect 6869 1865 6881 1899
rect 6869 1859 6927 1865
rect 6303 1842 6759 1858
rect 6303 1840 6758 1842
rect 7056 1840 7126 2369
rect 7849 2281 7862 2592
rect 7408 2263 7442 2281
rect 7828 2263 7862 2281
rect 7408 2227 7478 2263
rect 7425 2193 7496 2227
rect 7792 2214 7862 2263
rect 7883 2497 7916 2592
rect 8041 2586 8075 2592
rect 8025 2570 8078 2582
rect 8043 2558 8073 2570
rect 7997 2539 8073 2558
rect 8110 2539 8119 2543
rect 7883 2222 7917 2497
rect 7985 2490 8054 2539
rect 7985 2474 8036 2490
rect 7985 2459 8031 2474
rect 8085 2471 8098 2481
rect 7942 2443 7951 2447
rect 7963 2443 7976 2447
rect 7988 2443 8031 2459
rect 8079 2469 8098 2471
rect 7930 2343 7982 2443
rect 7991 2431 8031 2443
rect 8051 2443 8064 2447
rect 8051 2442 8070 2443
rect 8043 2431 8070 2442
rect 7991 2383 8070 2431
rect 7991 2371 8010 2383
rect 7997 2367 8010 2371
rect 8030 2371 8070 2383
rect 8079 2383 8102 2469
rect 8079 2371 8098 2383
rect 8030 2358 8073 2371
rect 8007 2355 8073 2358
rect 8075 2355 8076 2371
rect 8085 2367 8098 2371
rect 8110 2371 8131 2539
rect 8110 2367 8119 2371
rect 8144 2369 8178 2592
rect 8199 2369 8232 2654
rect 9398 2592 9425 2626
rect 9488 2615 9576 2626
rect 9499 2603 9565 2615
rect 9488 2593 9576 2603
rect 9639 2593 9652 2615
rect 9488 2592 9652 2593
rect 8712 2418 8770 2424
rect 8566 2369 8600 2387
rect 8712 2384 8724 2418
rect 8712 2378 8770 2384
rect 7930 2333 7976 2343
rect 7930 2222 7971 2333
rect 8007 2324 8076 2355
rect 8144 2333 8269 2369
rect 8025 2290 8098 2324
rect 8025 2274 8076 2290
rect 8061 2259 8076 2274
rect 8161 2256 8269 2333
rect 8030 2222 8064 2256
rect 8144 2222 8269 2256
rect 7883 2214 8269 2222
rect 5760 1812 5826 1838
rect 5764 1806 5822 1812
rect 5951 1804 7126 1840
rect 7238 1846 7296 1852
rect 7238 1838 7250 1846
rect 7425 1840 7495 2193
rect 7792 2152 8269 2214
rect 8343 2231 8401 2237
rect 8343 2197 8355 2231
rect 8343 2191 8401 2197
rect 7792 2144 8231 2152
rect 7607 2125 7665 2131
rect 7607 2091 7619 2125
rect 7607 2085 7665 2091
rect 7792 2082 8232 2144
rect 7792 1858 8233 2082
rect 8343 1899 8401 1905
rect 8343 1865 8355 1899
rect 8343 1859 8401 1865
rect 7777 1842 8233 1858
rect 7777 1840 8232 1842
rect 8530 1840 8600 2369
rect 9323 2281 9336 2592
rect 8882 2263 8916 2281
rect 9302 2263 9336 2281
rect 8882 2227 8952 2263
rect 8899 2193 8970 2227
rect 9266 2214 9336 2263
rect 9357 2497 9390 2592
rect 9515 2586 9549 2592
rect 9499 2570 9552 2582
rect 9517 2558 9547 2570
rect 9471 2539 9547 2558
rect 9584 2539 9593 2543
rect 9357 2222 9391 2497
rect 9459 2490 9528 2539
rect 9459 2474 9510 2490
rect 9459 2459 9505 2474
rect 9559 2471 9572 2481
rect 9416 2443 9425 2447
rect 9437 2443 9450 2447
rect 9462 2443 9505 2459
rect 9553 2469 9572 2471
rect 9404 2343 9456 2443
rect 9465 2431 9505 2443
rect 9525 2443 9538 2447
rect 9525 2442 9544 2443
rect 9517 2431 9544 2442
rect 9465 2383 9544 2431
rect 9465 2371 9484 2383
rect 9471 2367 9484 2371
rect 9504 2371 9544 2383
rect 9553 2383 9576 2469
rect 9553 2371 9572 2383
rect 9504 2358 9547 2371
rect 9481 2355 9547 2358
rect 9549 2355 9550 2371
rect 9559 2367 9572 2371
rect 9584 2371 9605 2539
rect 9584 2367 9593 2371
rect 9618 2369 9652 2592
rect 9673 2369 9706 2654
rect 10989 2586 11003 2620
rect 10186 2418 10244 2424
rect 10040 2369 10074 2387
rect 10186 2384 10198 2418
rect 10186 2378 10244 2384
rect 9404 2333 9450 2343
rect 9404 2222 9445 2333
rect 9481 2324 9550 2355
rect 9618 2333 9743 2369
rect 9499 2290 9572 2324
rect 9499 2274 9550 2290
rect 9535 2259 9550 2274
rect 9635 2256 9743 2333
rect 9504 2222 9538 2256
rect 9618 2222 9743 2256
rect 9357 2214 9743 2222
rect 7234 1812 7300 1838
rect 7238 1806 7296 1812
rect 7425 1804 8600 1840
rect 8712 1846 8770 1852
rect 8712 1838 8724 1846
rect 8899 1840 8969 2193
rect 9266 2152 9743 2214
rect 9817 2231 9875 2237
rect 9817 2197 9829 2231
rect 9817 2191 9875 2197
rect 9266 2144 9705 2152
rect 9081 2125 9139 2131
rect 9081 2091 9093 2125
rect 9081 2085 9139 2091
rect 9266 2082 9706 2144
rect 9266 1858 9707 2082
rect 9817 1899 9875 1905
rect 9817 1865 9829 1899
rect 9817 1859 9875 1865
rect 9251 1842 9707 1858
rect 9251 1840 9706 1842
rect 10004 1840 10074 2369
rect 10356 2263 10390 2281
rect 10356 2227 10426 2263
rect 10373 2193 10444 2227
rect 10831 2222 10865 2232
rect 10831 2214 11003 2222
rect 8708 1812 8774 1838
rect 8712 1806 8770 1812
rect 8899 1804 10074 1840
rect 10186 1846 10244 1852
rect 10186 1838 10198 1846
rect 10182 1812 10248 1838
rect 10186 1806 10244 1812
rect 458 1782 1213 1804
rect 1304 1798 1438 1804
rect 132 1717 290 1776
rect 791 1770 1213 1782
rect 1230 1778 1438 1798
rect 1230 1770 1404 1778
rect 1529 1770 2687 1804
rect 2778 1798 2912 1804
rect 2704 1778 2912 1798
rect 2704 1770 2878 1778
rect 3003 1770 4161 1804
rect 4252 1798 4386 1804
rect 4178 1778 4386 1798
rect 4178 1770 4352 1778
rect 4477 1770 5635 1804
rect 5726 1798 5860 1804
rect 5652 1778 5860 1798
rect 5652 1770 5826 1778
rect 5951 1770 7109 1804
rect 7200 1798 7334 1804
rect 7126 1778 7334 1798
rect 7126 1770 7300 1778
rect 7425 1770 8583 1804
rect 8674 1798 8808 1804
rect 8600 1778 8808 1798
rect 8600 1770 8774 1778
rect 8899 1770 10057 1804
rect 10148 1798 10282 1804
rect 10074 1778 10282 1798
rect 10074 1770 10248 1778
rect 791 1763 1230 1770
rect 1529 1763 2704 1770
rect 3003 1763 4178 1770
rect 4477 1763 5652 1770
rect 5951 1763 7126 1770
rect 7425 1763 8600 1770
rect 8899 1763 10074 1770
rect 791 1740 1213 1763
rect 1230 1742 1404 1744
rect 1230 1740 1450 1742
rect 791 1736 1450 1740
rect 791 1727 1332 1736
rect 70 1716 352 1717
rect 1196 1710 1332 1727
rect 1370 1710 1450 1736
rect 1529 1740 2687 1763
rect 2704 1742 2878 1744
rect 2704 1740 2924 1742
rect 1529 1736 2924 1740
rect 1529 1727 2806 1736
rect 1473 1710 1510 1717
rect 70 1682 352 1683
rect 1162 1676 1190 1702
rect 1232 1676 1298 1702
rect 1507 1676 1510 1683
rect 194 1614 228 1648
rect 1529 1621 2374 1727
rect 2670 1710 2806 1727
rect 2844 1710 2924 1736
rect 3003 1740 4161 1763
rect 4178 1742 4352 1744
rect 4178 1740 4398 1742
rect 3003 1736 4398 1740
rect 3003 1727 4280 1736
rect 2947 1710 2984 1717
rect 2636 1676 2664 1702
rect 2706 1676 2772 1702
rect 2981 1676 2984 1683
rect 3003 1621 3848 1727
rect 4144 1710 4280 1727
rect 4318 1710 4398 1736
rect 4477 1740 5635 1763
rect 5652 1742 5826 1744
rect 5652 1740 5872 1742
rect 4477 1736 5872 1740
rect 4477 1727 5754 1736
rect 4421 1710 4458 1717
rect 4110 1676 4138 1702
rect 4180 1676 4246 1702
rect 4455 1676 4458 1683
rect 4477 1621 5322 1727
rect 5618 1710 5754 1727
rect 5792 1710 5872 1736
rect 5951 1740 7109 1763
rect 7126 1742 7300 1744
rect 7126 1740 7346 1742
rect 5951 1736 7346 1740
rect 5951 1727 7228 1736
rect 5895 1710 5932 1717
rect 5584 1676 5612 1702
rect 5654 1676 5720 1702
rect 5929 1676 5932 1683
rect 5951 1621 6796 1727
rect 7092 1710 7228 1727
rect 7266 1710 7346 1736
rect 7425 1740 8583 1763
rect 8600 1742 8774 1744
rect 8600 1740 8820 1742
rect 7425 1736 8820 1740
rect 7425 1727 8702 1736
rect 7369 1710 7406 1717
rect 7058 1676 7086 1702
rect 7128 1676 7194 1702
rect 7403 1676 7406 1683
rect 7425 1621 8270 1727
rect 8566 1710 8702 1727
rect 8740 1710 8820 1736
rect 8899 1740 10057 1763
rect 10074 1742 10248 1744
rect 10074 1740 10294 1742
rect 8899 1736 10294 1740
rect 8899 1727 10176 1736
rect 8843 1710 8880 1717
rect 8532 1676 8560 1702
rect 8602 1676 8668 1702
rect 8877 1676 8880 1683
rect 8899 1621 9744 1727
rect 10040 1710 10176 1727
rect 10214 1710 10294 1736
rect 10373 1710 10443 2193
rect 10795 2152 11217 2214
rect 10555 2125 10613 2131
rect 10555 2091 10567 2125
rect 10555 2085 10613 2091
rect 10957 1862 10977 1870
rect 10555 1793 10613 1799
rect 10555 1759 10567 1793
rect 10555 1753 10613 1759
rect 10006 1676 10034 1702
rect 10076 1676 10142 1702
rect 10373 1674 10426 1710
rect 1668 1614 1702 1621
rect 3142 1614 3176 1621
rect 4616 1614 4650 1621
rect 6090 1614 6124 1621
rect 7564 1614 7598 1621
rect 9038 1614 9072 1621
rect 2182 1411 2198 1433
rect 3656 1411 3672 1433
rect 5130 1411 5146 1433
rect 6604 1411 6620 1433
rect 8078 1411 8094 1433
rect 9552 1411 9568 1433
rect 2182 1383 2204 1405
rect 3656 1383 3678 1405
rect 5130 1383 5152 1405
rect 6604 1383 6626 1405
rect 8078 1383 8100 1405
rect 9552 1383 9574 1405
rect 36 1250 70 1260
rect 352 1250 386 1260
rect 36 1242 386 1250
rect 1510 1250 1544 1260
rect 1826 1250 1860 1260
rect 1510 1242 1860 1250
rect 2984 1250 3018 1260
rect 3300 1250 3334 1260
rect 2984 1242 3334 1250
rect 4458 1250 4492 1260
rect 4774 1250 4808 1260
rect 4458 1242 4808 1250
rect 5932 1250 5966 1260
rect 6248 1250 6282 1260
rect 5932 1242 6282 1250
rect 7406 1250 7440 1260
rect 7722 1250 7756 1260
rect 7406 1242 7756 1250
rect 8880 1250 8914 1260
rect 9196 1250 9230 1260
rect 8880 1242 9230 1250
rect 0 1180 422 1242
rect 1474 1180 1896 1242
rect 2948 1180 3370 1242
rect 4422 1180 4844 1242
rect 5896 1180 6318 1242
rect 7370 1180 7792 1242
rect 8844 1180 9266 1242
rect 668 928 675 1033
rect 696 956 703 1020
rect 2142 1005 2149 1033
rect 2170 1005 2177 1020
rect 3616 1005 3623 1033
rect 3644 1005 3651 1020
rect 5090 1005 5097 1033
rect 5118 1005 5125 1020
rect 6564 1005 6571 1033
rect 6592 1005 6599 1020
rect 8038 1005 8045 1033
rect 8066 1005 8073 1020
rect 9512 1005 9519 1033
rect 9540 1005 9547 1020
rect 162 890 182 898
rect 1636 890 1656 898
rect 3110 890 3130 898
rect 4584 890 4604 898
rect 6058 890 6078 898
rect 7532 890 7552 898
rect 9006 890 9026 898
rect 2098 808 2204 810
rect 3572 808 3678 810
rect 5046 808 5152 810
rect 6520 808 6626 810
rect 7994 808 8100 810
rect 9468 808 9574 810
rect 2088 805 2204 808
rect 3562 805 3678 808
rect 5036 805 5152 808
rect 6510 805 6626 808
rect 7984 805 8100 808
rect 9458 805 9574 808
rect 2126 780 2192 782
rect 3600 780 3666 782
rect 5074 780 5140 782
rect 6548 780 6614 782
rect 8022 780 8088 782
rect 9496 780 9562 782
rect 2116 777 2232 780
rect 3590 777 3706 780
rect 5064 777 5180 780
rect 6538 777 6654 780
rect 8012 777 8128 780
rect 9486 777 9602 780
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
use mux_2to1_logic  x1
timestamp 1624053917
transform 1 0 475 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x2
timestamp 1624053917
transform 1 0 1949 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x3
timestamp 1624053917
transform 1 0 3423 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x5
timestamp 1624053917
transform 1 0 4897 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x6
timestamp 1624053917
transform 1 0 6371 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x7
timestamp 1624053917
transform 1 0 7845 0 1 1233
box -475 -2400 1898 1551
use mux_2to1_logic  x8
timestamp 1624053917
transform 1 0 9319 0 1 1233
box -475 -2400 1898 1551
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd1p8
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 avss1p8
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 mux_i7
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 mux_i6
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 mux_i5
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 out_mux
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 mux_i4
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 mux_i3
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 reg0
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 mux_i2
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 mux_i1
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 {}
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 mux_i0
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 reg1
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 reg2
port 15 nsew
<< end >>
