magic
tech sky130A
magscale 1 2
timestamp 1623255091
<< error_p >>
rect -1823 -1511 -1761 -1505
rect -1695 -1511 -1633 -1505
rect -1567 -1511 -1505 -1505
rect -1439 -1511 -1377 -1505
rect -1311 -1511 -1249 -1505
rect -1183 -1511 -1121 -1505
rect -1055 -1511 -993 -1505
rect -927 -1511 -865 -1505
rect -799 -1511 -737 -1505
rect -671 -1511 -609 -1505
rect -543 -1511 -481 -1505
rect -415 -1511 -353 -1505
rect -287 -1511 -225 -1505
rect -159 -1511 -97 -1505
rect -31 -1511 31 -1505
rect 97 -1511 159 -1505
rect 225 -1511 287 -1505
rect 353 -1511 415 -1505
rect 481 -1511 543 -1505
rect 609 -1511 671 -1505
rect 737 -1511 799 -1505
rect 865 -1511 927 -1505
rect 993 -1511 1055 -1505
rect 1121 -1511 1183 -1505
rect 1249 -1511 1311 -1505
rect 1377 -1511 1439 -1505
rect 1505 -1511 1567 -1505
rect 1633 -1511 1695 -1505
rect 1761 -1511 1823 -1505
rect -1823 -1545 -1811 -1511
rect -1695 -1545 -1683 -1511
rect -1567 -1545 -1555 -1511
rect -1439 -1545 -1427 -1511
rect -1311 -1545 -1299 -1511
rect -1183 -1545 -1171 -1511
rect -1055 -1545 -1043 -1511
rect -927 -1545 -915 -1511
rect -799 -1545 -787 -1511
rect -671 -1545 -659 -1511
rect -543 -1545 -531 -1511
rect -415 -1545 -403 -1511
rect -287 -1545 -275 -1511
rect -159 -1545 -147 -1511
rect -31 -1545 -19 -1511
rect 97 -1545 109 -1511
rect 225 -1545 237 -1511
rect 353 -1545 365 -1511
rect 481 -1545 493 -1511
rect 609 -1545 621 -1511
rect 737 -1545 749 -1511
rect 865 -1545 877 -1511
rect 993 -1545 1005 -1511
rect 1121 -1545 1133 -1511
rect 1249 -1545 1261 -1511
rect 1377 -1545 1389 -1511
rect 1505 -1545 1517 -1511
rect 1633 -1545 1645 -1511
rect 1761 -1545 1773 -1511
rect -1823 -1551 -1761 -1545
rect -1695 -1551 -1633 -1545
rect -1567 -1551 -1505 -1545
rect -1439 -1551 -1377 -1545
rect -1311 -1551 -1249 -1545
rect -1183 -1551 -1121 -1545
rect -1055 -1551 -993 -1545
rect -927 -1551 -865 -1545
rect -799 -1551 -737 -1545
rect -671 -1551 -609 -1545
rect -543 -1551 -481 -1545
rect -415 -1551 -353 -1545
rect -287 -1551 -225 -1545
rect -159 -1551 -97 -1545
rect -31 -1551 31 -1545
rect 97 -1551 159 -1545
rect 225 -1551 287 -1545
rect 353 -1551 415 -1545
rect 481 -1551 543 -1545
rect 609 -1551 671 -1545
rect 737 -1551 799 -1545
rect 865 -1551 927 -1545
rect 993 -1551 1055 -1545
rect 1121 -1551 1183 -1545
rect 1249 -1551 1311 -1545
rect 1377 -1551 1439 -1545
rect 1505 -1551 1567 -1545
rect 1633 -1551 1695 -1545
rect 1761 -1551 1823 -1545
<< nwell >>
rect -2023 -1684 2023 1684
<< pmoslvt >>
rect -1827 -1464 -1757 1536
rect -1699 -1464 -1629 1536
rect -1571 -1464 -1501 1536
rect -1443 -1464 -1373 1536
rect -1315 -1464 -1245 1536
rect -1187 -1464 -1117 1536
rect -1059 -1464 -989 1536
rect -931 -1464 -861 1536
rect -803 -1464 -733 1536
rect -675 -1464 -605 1536
rect -547 -1464 -477 1536
rect -419 -1464 -349 1536
rect -291 -1464 -221 1536
rect -163 -1464 -93 1536
rect -35 -1464 35 1536
rect 93 -1464 163 1536
rect 221 -1464 291 1536
rect 349 -1464 419 1536
rect 477 -1464 547 1536
rect 605 -1464 675 1536
rect 733 -1464 803 1536
rect 861 -1464 931 1536
rect 989 -1464 1059 1536
rect 1117 -1464 1187 1536
rect 1245 -1464 1315 1536
rect 1373 -1464 1443 1536
rect 1501 -1464 1571 1536
rect 1629 -1464 1699 1536
rect 1757 -1464 1827 1536
<< pdiff >>
rect -1885 1524 -1827 1536
rect -1885 -1452 -1873 1524
rect -1839 -1452 -1827 1524
rect -1885 -1464 -1827 -1452
rect -1757 1524 -1699 1536
rect -1757 -1452 -1745 1524
rect -1711 -1452 -1699 1524
rect -1757 -1464 -1699 -1452
rect -1629 1524 -1571 1536
rect -1629 -1452 -1617 1524
rect -1583 -1452 -1571 1524
rect -1629 -1464 -1571 -1452
rect -1501 1524 -1443 1536
rect -1501 -1452 -1489 1524
rect -1455 -1452 -1443 1524
rect -1501 -1464 -1443 -1452
rect -1373 1524 -1315 1536
rect -1373 -1452 -1361 1524
rect -1327 -1452 -1315 1524
rect -1373 -1464 -1315 -1452
rect -1245 1524 -1187 1536
rect -1245 -1452 -1233 1524
rect -1199 -1452 -1187 1524
rect -1245 -1464 -1187 -1452
rect -1117 1524 -1059 1536
rect -1117 -1452 -1105 1524
rect -1071 -1452 -1059 1524
rect -1117 -1464 -1059 -1452
rect -989 1524 -931 1536
rect -989 -1452 -977 1524
rect -943 -1452 -931 1524
rect -989 -1464 -931 -1452
rect -861 1524 -803 1536
rect -861 -1452 -849 1524
rect -815 -1452 -803 1524
rect -861 -1464 -803 -1452
rect -733 1524 -675 1536
rect -733 -1452 -721 1524
rect -687 -1452 -675 1524
rect -733 -1464 -675 -1452
rect -605 1524 -547 1536
rect -605 -1452 -593 1524
rect -559 -1452 -547 1524
rect -605 -1464 -547 -1452
rect -477 1524 -419 1536
rect -477 -1452 -465 1524
rect -431 -1452 -419 1524
rect -477 -1464 -419 -1452
rect -349 1524 -291 1536
rect -349 -1452 -337 1524
rect -303 -1452 -291 1524
rect -349 -1464 -291 -1452
rect -221 1524 -163 1536
rect -221 -1452 -209 1524
rect -175 -1452 -163 1524
rect -221 -1464 -163 -1452
rect -93 1524 -35 1536
rect -93 -1452 -81 1524
rect -47 -1452 -35 1524
rect -93 -1464 -35 -1452
rect 35 1524 93 1536
rect 35 -1452 47 1524
rect 81 -1452 93 1524
rect 35 -1464 93 -1452
rect 163 1524 221 1536
rect 163 -1452 175 1524
rect 209 -1452 221 1524
rect 163 -1464 221 -1452
rect 291 1524 349 1536
rect 291 -1452 303 1524
rect 337 -1452 349 1524
rect 291 -1464 349 -1452
rect 419 1524 477 1536
rect 419 -1452 431 1524
rect 465 -1452 477 1524
rect 419 -1464 477 -1452
rect 547 1524 605 1536
rect 547 -1452 559 1524
rect 593 -1452 605 1524
rect 547 -1464 605 -1452
rect 675 1524 733 1536
rect 675 -1452 687 1524
rect 721 -1452 733 1524
rect 675 -1464 733 -1452
rect 803 1524 861 1536
rect 803 -1452 815 1524
rect 849 -1452 861 1524
rect 803 -1464 861 -1452
rect 931 1524 989 1536
rect 931 -1452 943 1524
rect 977 -1452 989 1524
rect 931 -1464 989 -1452
rect 1059 1524 1117 1536
rect 1059 -1452 1071 1524
rect 1105 -1452 1117 1524
rect 1059 -1464 1117 -1452
rect 1187 1524 1245 1536
rect 1187 -1452 1199 1524
rect 1233 -1452 1245 1524
rect 1187 -1464 1245 -1452
rect 1315 1524 1373 1536
rect 1315 -1452 1327 1524
rect 1361 -1452 1373 1524
rect 1315 -1464 1373 -1452
rect 1443 1524 1501 1536
rect 1443 -1452 1455 1524
rect 1489 -1452 1501 1524
rect 1443 -1464 1501 -1452
rect 1571 1524 1629 1536
rect 1571 -1452 1583 1524
rect 1617 -1452 1629 1524
rect 1571 -1464 1629 -1452
rect 1699 1524 1757 1536
rect 1699 -1452 1711 1524
rect 1745 -1452 1757 1524
rect 1699 -1464 1757 -1452
rect 1827 1524 1885 1536
rect 1827 -1452 1839 1524
rect 1873 -1452 1885 1524
rect 1827 -1464 1885 -1452
<< pdiffc >>
rect -1873 -1452 -1839 1524
rect -1745 -1452 -1711 1524
rect -1617 -1452 -1583 1524
rect -1489 -1452 -1455 1524
rect -1361 -1452 -1327 1524
rect -1233 -1452 -1199 1524
rect -1105 -1452 -1071 1524
rect -977 -1452 -943 1524
rect -849 -1452 -815 1524
rect -721 -1452 -687 1524
rect -593 -1452 -559 1524
rect -465 -1452 -431 1524
rect -337 -1452 -303 1524
rect -209 -1452 -175 1524
rect -81 -1452 -47 1524
rect 47 -1452 81 1524
rect 175 -1452 209 1524
rect 303 -1452 337 1524
rect 431 -1452 465 1524
rect 559 -1452 593 1524
rect 687 -1452 721 1524
rect 815 -1452 849 1524
rect 943 -1452 977 1524
rect 1071 -1452 1105 1524
rect 1199 -1452 1233 1524
rect 1327 -1452 1361 1524
rect 1455 -1452 1489 1524
rect 1583 -1452 1617 1524
rect 1711 -1452 1745 1524
rect 1839 -1452 1873 1524
<< nsubdiff >>
rect -1987 1614 -1891 1648
rect 1891 1614 1987 1648
rect -1987 1551 -1953 1614
rect 1953 1551 1987 1614
rect -1987 -1614 -1953 -1551
rect 1953 -1614 1987 -1551
rect -1987 -1648 -1891 -1614
rect 1891 -1648 1987 -1614
<< nsubdiffcont >>
rect -1891 1614 1891 1648
rect -1987 -1551 -1953 1551
rect 1953 -1551 1987 1551
rect -1891 -1648 1891 -1614
<< poly >>
rect -1827 1536 -1757 1562
rect -1699 1536 -1629 1562
rect -1571 1536 -1501 1562
rect -1443 1536 -1373 1562
rect -1315 1536 -1245 1562
rect -1187 1536 -1117 1562
rect -1059 1536 -989 1562
rect -931 1536 -861 1562
rect -803 1536 -733 1562
rect -675 1536 -605 1562
rect -547 1536 -477 1562
rect -419 1536 -349 1562
rect -291 1536 -221 1562
rect -163 1536 -93 1562
rect -35 1536 35 1562
rect 93 1536 163 1562
rect 221 1536 291 1562
rect 349 1536 419 1562
rect 477 1536 547 1562
rect 605 1536 675 1562
rect 733 1536 803 1562
rect 861 1536 931 1562
rect 989 1536 1059 1562
rect 1117 1536 1187 1562
rect 1245 1536 1315 1562
rect 1373 1536 1443 1562
rect 1501 1536 1571 1562
rect 1629 1536 1699 1562
rect 1757 1536 1827 1562
rect -1827 -1511 -1757 -1464
rect -1827 -1545 -1811 -1511
rect -1773 -1545 -1757 -1511
rect -1827 -1561 -1757 -1545
rect -1699 -1511 -1629 -1464
rect -1699 -1545 -1683 -1511
rect -1645 -1545 -1629 -1511
rect -1699 -1561 -1629 -1545
rect -1571 -1511 -1501 -1464
rect -1571 -1545 -1555 -1511
rect -1517 -1545 -1501 -1511
rect -1571 -1561 -1501 -1545
rect -1443 -1511 -1373 -1464
rect -1443 -1545 -1427 -1511
rect -1389 -1545 -1373 -1511
rect -1443 -1561 -1373 -1545
rect -1315 -1511 -1245 -1464
rect -1315 -1545 -1299 -1511
rect -1261 -1545 -1245 -1511
rect -1315 -1561 -1245 -1545
rect -1187 -1511 -1117 -1464
rect -1187 -1545 -1171 -1511
rect -1133 -1545 -1117 -1511
rect -1187 -1561 -1117 -1545
rect -1059 -1511 -989 -1464
rect -1059 -1545 -1043 -1511
rect -1005 -1545 -989 -1511
rect -1059 -1561 -989 -1545
rect -931 -1511 -861 -1464
rect -931 -1545 -915 -1511
rect -877 -1545 -861 -1511
rect -931 -1561 -861 -1545
rect -803 -1511 -733 -1464
rect -803 -1545 -787 -1511
rect -749 -1545 -733 -1511
rect -803 -1561 -733 -1545
rect -675 -1511 -605 -1464
rect -675 -1545 -659 -1511
rect -621 -1545 -605 -1511
rect -675 -1561 -605 -1545
rect -547 -1511 -477 -1464
rect -547 -1545 -531 -1511
rect -493 -1545 -477 -1511
rect -547 -1561 -477 -1545
rect -419 -1511 -349 -1464
rect -419 -1545 -403 -1511
rect -365 -1545 -349 -1511
rect -419 -1561 -349 -1545
rect -291 -1511 -221 -1464
rect -291 -1545 -275 -1511
rect -237 -1545 -221 -1511
rect -291 -1561 -221 -1545
rect -163 -1511 -93 -1464
rect -163 -1545 -147 -1511
rect -109 -1545 -93 -1511
rect -163 -1561 -93 -1545
rect -35 -1511 35 -1464
rect -35 -1545 -19 -1511
rect 19 -1545 35 -1511
rect -35 -1561 35 -1545
rect 93 -1511 163 -1464
rect 93 -1545 109 -1511
rect 147 -1545 163 -1511
rect 93 -1561 163 -1545
rect 221 -1511 291 -1464
rect 221 -1545 237 -1511
rect 275 -1545 291 -1511
rect 221 -1561 291 -1545
rect 349 -1511 419 -1464
rect 349 -1545 365 -1511
rect 403 -1545 419 -1511
rect 349 -1561 419 -1545
rect 477 -1511 547 -1464
rect 477 -1545 493 -1511
rect 531 -1545 547 -1511
rect 477 -1561 547 -1545
rect 605 -1511 675 -1464
rect 605 -1545 621 -1511
rect 659 -1545 675 -1511
rect 605 -1561 675 -1545
rect 733 -1511 803 -1464
rect 733 -1545 749 -1511
rect 787 -1545 803 -1511
rect 733 -1561 803 -1545
rect 861 -1511 931 -1464
rect 861 -1545 877 -1511
rect 915 -1545 931 -1511
rect 861 -1561 931 -1545
rect 989 -1511 1059 -1464
rect 989 -1545 1005 -1511
rect 1043 -1545 1059 -1511
rect 989 -1561 1059 -1545
rect 1117 -1511 1187 -1464
rect 1117 -1545 1133 -1511
rect 1171 -1545 1187 -1511
rect 1117 -1561 1187 -1545
rect 1245 -1511 1315 -1464
rect 1245 -1545 1261 -1511
rect 1299 -1545 1315 -1511
rect 1245 -1561 1315 -1545
rect 1373 -1511 1443 -1464
rect 1373 -1545 1389 -1511
rect 1427 -1545 1443 -1511
rect 1373 -1561 1443 -1545
rect 1501 -1511 1571 -1464
rect 1501 -1545 1517 -1511
rect 1555 -1545 1571 -1511
rect 1501 -1561 1571 -1545
rect 1629 -1511 1699 -1464
rect 1629 -1545 1645 -1511
rect 1683 -1545 1699 -1511
rect 1629 -1561 1699 -1545
rect 1757 -1511 1827 -1464
rect 1757 -1545 1773 -1511
rect 1811 -1545 1827 -1511
rect 1757 -1561 1827 -1545
<< polycont >>
rect -1811 -1545 -1773 -1511
rect -1683 -1545 -1645 -1511
rect -1555 -1545 -1517 -1511
rect -1427 -1545 -1389 -1511
rect -1299 -1545 -1261 -1511
rect -1171 -1545 -1133 -1511
rect -1043 -1545 -1005 -1511
rect -915 -1545 -877 -1511
rect -787 -1545 -749 -1511
rect -659 -1545 -621 -1511
rect -531 -1545 -493 -1511
rect -403 -1545 -365 -1511
rect -275 -1545 -237 -1511
rect -147 -1545 -109 -1511
rect -19 -1545 19 -1511
rect 109 -1545 147 -1511
rect 237 -1545 275 -1511
rect 365 -1545 403 -1511
rect 493 -1545 531 -1511
rect 621 -1545 659 -1511
rect 749 -1545 787 -1511
rect 877 -1545 915 -1511
rect 1005 -1545 1043 -1511
rect 1133 -1545 1171 -1511
rect 1261 -1545 1299 -1511
rect 1389 -1545 1427 -1511
rect 1517 -1545 1555 -1511
rect 1645 -1545 1683 -1511
rect 1773 -1545 1811 -1511
<< locali >>
rect -1987 1614 -1891 1648
rect 1891 1614 1987 1648
rect -1987 1551 -1953 1614
rect 1953 1551 1987 1614
rect -1873 1524 -1839 1540
rect -1873 -1468 -1839 -1452
rect -1745 1524 -1711 1540
rect -1745 -1468 -1711 -1452
rect -1617 1524 -1583 1540
rect -1617 -1468 -1583 -1452
rect -1489 1524 -1455 1540
rect -1489 -1468 -1455 -1452
rect -1361 1524 -1327 1540
rect -1361 -1468 -1327 -1452
rect -1233 1524 -1199 1540
rect -1233 -1468 -1199 -1452
rect -1105 1524 -1071 1540
rect -1105 -1468 -1071 -1452
rect -977 1524 -943 1540
rect -977 -1468 -943 -1452
rect -849 1524 -815 1540
rect -849 -1468 -815 -1452
rect -721 1524 -687 1540
rect -721 -1468 -687 -1452
rect -593 1524 -559 1540
rect -593 -1468 -559 -1452
rect -465 1524 -431 1540
rect -465 -1468 -431 -1452
rect -337 1524 -303 1540
rect -337 -1468 -303 -1452
rect -209 1524 -175 1540
rect -209 -1468 -175 -1452
rect -81 1524 -47 1540
rect -81 -1468 -47 -1452
rect 47 1524 81 1540
rect 47 -1468 81 -1452
rect 175 1524 209 1540
rect 175 -1468 209 -1452
rect 303 1524 337 1540
rect 303 -1468 337 -1452
rect 431 1524 465 1540
rect 431 -1468 465 -1452
rect 559 1524 593 1540
rect 559 -1468 593 -1452
rect 687 1524 721 1540
rect 687 -1468 721 -1452
rect 815 1524 849 1540
rect 815 -1468 849 -1452
rect 943 1524 977 1540
rect 943 -1468 977 -1452
rect 1071 1524 1105 1540
rect 1071 -1468 1105 -1452
rect 1199 1524 1233 1540
rect 1199 -1468 1233 -1452
rect 1327 1524 1361 1540
rect 1327 -1468 1361 -1452
rect 1455 1524 1489 1540
rect 1455 -1468 1489 -1452
rect 1583 1524 1617 1540
rect 1583 -1468 1617 -1452
rect 1711 1524 1745 1540
rect 1711 -1468 1745 -1452
rect 1839 1524 1873 1540
rect 1839 -1468 1873 -1452
rect -1827 -1545 -1811 -1511
rect -1773 -1545 -1757 -1511
rect -1699 -1545 -1683 -1511
rect -1645 -1545 -1629 -1511
rect -1571 -1545 -1555 -1511
rect -1517 -1545 -1501 -1511
rect -1443 -1545 -1427 -1511
rect -1389 -1545 -1373 -1511
rect -1315 -1545 -1299 -1511
rect -1261 -1545 -1245 -1511
rect -1187 -1545 -1171 -1511
rect -1133 -1545 -1117 -1511
rect -1059 -1545 -1043 -1511
rect -1005 -1545 -989 -1511
rect -931 -1545 -915 -1511
rect -877 -1545 -861 -1511
rect -803 -1545 -787 -1511
rect -749 -1545 -733 -1511
rect -675 -1545 -659 -1511
rect -621 -1545 -605 -1511
rect -547 -1545 -531 -1511
rect -493 -1545 -477 -1511
rect -419 -1545 -403 -1511
rect -365 -1545 -349 -1511
rect -291 -1545 -275 -1511
rect -237 -1545 -221 -1511
rect -163 -1545 -147 -1511
rect -109 -1545 -93 -1511
rect -35 -1545 -19 -1511
rect 19 -1545 35 -1511
rect 93 -1545 109 -1511
rect 147 -1545 163 -1511
rect 221 -1545 237 -1511
rect 275 -1545 291 -1511
rect 349 -1545 365 -1511
rect 403 -1545 419 -1511
rect 477 -1545 493 -1511
rect 531 -1545 547 -1511
rect 605 -1545 621 -1511
rect 659 -1545 675 -1511
rect 733 -1545 749 -1511
rect 787 -1545 803 -1511
rect 861 -1545 877 -1511
rect 915 -1545 931 -1511
rect 989 -1545 1005 -1511
rect 1043 -1545 1059 -1511
rect 1117 -1545 1133 -1511
rect 1171 -1545 1187 -1511
rect 1245 -1545 1261 -1511
rect 1299 -1545 1315 -1511
rect 1373 -1545 1389 -1511
rect 1427 -1545 1443 -1511
rect 1501 -1545 1517 -1511
rect 1555 -1545 1571 -1511
rect 1629 -1545 1645 -1511
rect 1683 -1545 1699 -1511
rect 1757 -1545 1773 -1511
rect 1811 -1545 1827 -1511
rect -1987 -1614 -1953 -1551
rect 1953 -1614 1987 -1551
rect -1987 -1648 -1891 -1614
rect 1891 -1648 1987 -1614
<< viali >>
rect -1873 -1452 -1839 1524
rect -1745 -1452 -1711 1524
rect -1617 -1452 -1583 1524
rect -1489 -1452 -1455 1524
rect -1361 -1452 -1327 1524
rect -1233 -1452 -1199 1524
rect -1105 -1452 -1071 1524
rect -977 -1452 -943 1524
rect -849 -1452 -815 1524
rect -721 -1452 -687 1524
rect -593 -1452 -559 1524
rect -465 -1452 -431 1524
rect -337 -1452 -303 1524
rect -209 -1452 -175 1524
rect -81 -1452 -47 1524
rect 47 -1452 81 1524
rect 175 -1452 209 1524
rect 303 -1452 337 1524
rect 431 -1452 465 1524
rect 559 -1452 593 1524
rect 687 -1452 721 1524
rect 815 -1452 849 1524
rect 943 -1452 977 1524
rect 1071 -1452 1105 1524
rect 1199 -1452 1233 1524
rect 1327 -1452 1361 1524
rect 1455 -1452 1489 1524
rect 1583 -1452 1617 1524
rect 1711 -1452 1745 1524
rect 1839 -1452 1873 1524
rect -1811 -1545 -1773 -1511
rect -1683 -1545 -1645 -1511
rect -1555 -1545 -1517 -1511
rect -1427 -1545 -1389 -1511
rect -1299 -1545 -1261 -1511
rect -1171 -1545 -1133 -1511
rect -1043 -1545 -1005 -1511
rect -915 -1545 -877 -1511
rect -787 -1545 -749 -1511
rect -659 -1545 -621 -1511
rect -531 -1545 -493 -1511
rect -403 -1545 -365 -1511
rect -275 -1545 -237 -1511
rect -147 -1545 -109 -1511
rect -19 -1545 19 -1511
rect 109 -1545 147 -1511
rect 237 -1545 275 -1511
rect 365 -1545 403 -1511
rect 493 -1545 531 -1511
rect 621 -1545 659 -1511
rect 749 -1545 787 -1511
rect 877 -1545 915 -1511
rect 1005 -1545 1043 -1511
rect 1133 -1545 1171 -1511
rect 1261 -1545 1299 -1511
rect 1389 -1545 1427 -1511
rect 1517 -1545 1555 -1511
rect 1645 -1545 1683 -1511
rect 1773 -1545 1811 -1511
<< metal1 >>
rect -1879 1524 -1833 1536
rect -1879 -1452 -1873 1524
rect -1839 -1452 -1833 1524
rect -1879 -1464 -1833 -1452
rect -1751 1524 -1705 1536
rect -1751 -1452 -1745 1524
rect -1711 -1452 -1705 1524
rect -1751 -1464 -1705 -1452
rect -1623 1524 -1577 1536
rect -1623 -1452 -1617 1524
rect -1583 -1452 -1577 1524
rect -1623 -1464 -1577 -1452
rect -1495 1524 -1449 1536
rect -1495 -1452 -1489 1524
rect -1455 -1452 -1449 1524
rect -1495 -1464 -1449 -1452
rect -1367 1524 -1321 1536
rect -1367 -1452 -1361 1524
rect -1327 -1452 -1321 1524
rect -1367 -1464 -1321 -1452
rect -1239 1524 -1193 1536
rect -1239 -1452 -1233 1524
rect -1199 -1452 -1193 1524
rect -1239 -1464 -1193 -1452
rect -1111 1524 -1065 1536
rect -1111 -1452 -1105 1524
rect -1071 -1452 -1065 1524
rect -1111 -1464 -1065 -1452
rect -983 1524 -937 1536
rect -983 -1452 -977 1524
rect -943 -1452 -937 1524
rect -983 -1464 -937 -1452
rect -855 1524 -809 1536
rect -855 -1452 -849 1524
rect -815 -1452 -809 1524
rect -855 -1464 -809 -1452
rect -727 1524 -681 1536
rect -727 -1452 -721 1524
rect -687 -1452 -681 1524
rect -727 -1464 -681 -1452
rect -599 1524 -553 1536
rect -599 -1452 -593 1524
rect -559 -1452 -553 1524
rect -599 -1464 -553 -1452
rect -471 1524 -425 1536
rect -471 -1452 -465 1524
rect -431 -1452 -425 1524
rect -471 -1464 -425 -1452
rect -343 1524 -297 1536
rect -343 -1452 -337 1524
rect -303 -1452 -297 1524
rect -343 -1464 -297 -1452
rect -215 1524 -169 1536
rect -215 -1452 -209 1524
rect -175 -1452 -169 1524
rect -215 -1464 -169 -1452
rect -87 1524 -41 1536
rect -87 -1452 -81 1524
rect -47 -1452 -41 1524
rect -87 -1464 -41 -1452
rect 41 1524 87 1536
rect 41 -1452 47 1524
rect 81 -1452 87 1524
rect 41 -1464 87 -1452
rect 169 1524 215 1536
rect 169 -1452 175 1524
rect 209 -1452 215 1524
rect 169 -1464 215 -1452
rect 297 1524 343 1536
rect 297 -1452 303 1524
rect 337 -1452 343 1524
rect 297 -1464 343 -1452
rect 425 1524 471 1536
rect 425 -1452 431 1524
rect 465 -1452 471 1524
rect 425 -1464 471 -1452
rect 553 1524 599 1536
rect 553 -1452 559 1524
rect 593 -1452 599 1524
rect 553 -1464 599 -1452
rect 681 1524 727 1536
rect 681 -1452 687 1524
rect 721 -1452 727 1524
rect 681 -1464 727 -1452
rect 809 1524 855 1536
rect 809 -1452 815 1524
rect 849 -1452 855 1524
rect 809 -1464 855 -1452
rect 937 1524 983 1536
rect 937 -1452 943 1524
rect 977 -1452 983 1524
rect 937 -1464 983 -1452
rect 1065 1524 1111 1536
rect 1065 -1452 1071 1524
rect 1105 -1452 1111 1524
rect 1065 -1464 1111 -1452
rect 1193 1524 1239 1536
rect 1193 -1452 1199 1524
rect 1233 -1452 1239 1524
rect 1193 -1464 1239 -1452
rect 1321 1524 1367 1536
rect 1321 -1452 1327 1524
rect 1361 -1452 1367 1524
rect 1321 -1464 1367 -1452
rect 1449 1524 1495 1536
rect 1449 -1452 1455 1524
rect 1489 -1452 1495 1524
rect 1449 -1464 1495 -1452
rect 1577 1524 1623 1536
rect 1577 -1452 1583 1524
rect 1617 -1452 1623 1524
rect 1577 -1464 1623 -1452
rect 1705 1524 1751 1536
rect 1705 -1452 1711 1524
rect 1745 -1452 1751 1524
rect 1705 -1464 1751 -1452
rect 1833 1524 1879 1536
rect 1833 -1452 1839 1524
rect 1873 -1452 1879 1524
rect 1833 -1464 1879 -1452
rect -1823 -1511 -1761 -1505
rect -1823 -1545 -1811 -1511
rect -1773 -1545 -1761 -1511
rect -1823 -1551 -1761 -1545
rect -1695 -1511 -1633 -1505
rect -1695 -1545 -1683 -1511
rect -1645 -1545 -1633 -1511
rect -1695 -1551 -1633 -1545
rect -1567 -1511 -1505 -1505
rect -1567 -1545 -1555 -1511
rect -1517 -1545 -1505 -1511
rect -1567 -1551 -1505 -1545
rect -1439 -1511 -1377 -1505
rect -1439 -1545 -1427 -1511
rect -1389 -1545 -1377 -1511
rect -1439 -1551 -1377 -1545
rect -1311 -1511 -1249 -1505
rect -1311 -1545 -1299 -1511
rect -1261 -1545 -1249 -1511
rect -1311 -1551 -1249 -1545
rect -1183 -1511 -1121 -1505
rect -1183 -1545 -1171 -1511
rect -1133 -1545 -1121 -1511
rect -1183 -1551 -1121 -1545
rect -1055 -1511 -993 -1505
rect -1055 -1545 -1043 -1511
rect -1005 -1545 -993 -1511
rect -1055 -1551 -993 -1545
rect -927 -1511 -865 -1505
rect -927 -1545 -915 -1511
rect -877 -1545 -865 -1511
rect -927 -1551 -865 -1545
rect -799 -1511 -737 -1505
rect -799 -1545 -787 -1511
rect -749 -1545 -737 -1511
rect -799 -1551 -737 -1545
rect -671 -1511 -609 -1505
rect -671 -1545 -659 -1511
rect -621 -1545 -609 -1511
rect -671 -1551 -609 -1545
rect -543 -1511 -481 -1505
rect -543 -1545 -531 -1511
rect -493 -1545 -481 -1511
rect -543 -1551 -481 -1545
rect -415 -1511 -353 -1505
rect -415 -1545 -403 -1511
rect -365 -1545 -353 -1511
rect -415 -1551 -353 -1545
rect -287 -1511 -225 -1505
rect -287 -1545 -275 -1511
rect -237 -1545 -225 -1511
rect -287 -1551 -225 -1545
rect -159 -1511 -97 -1505
rect -159 -1545 -147 -1511
rect -109 -1545 -97 -1511
rect -159 -1551 -97 -1545
rect -31 -1511 31 -1505
rect -31 -1545 -19 -1511
rect 19 -1545 31 -1511
rect -31 -1551 31 -1545
rect 97 -1511 159 -1505
rect 97 -1545 109 -1511
rect 147 -1545 159 -1511
rect 97 -1551 159 -1545
rect 225 -1511 287 -1505
rect 225 -1545 237 -1511
rect 275 -1545 287 -1511
rect 225 -1551 287 -1545
rect 353 -1511 415 -1505
rect 353 -1545 365 -1511
rect 403 -1545 415 -1511
rect 353 -1551 415 -1545
rect 481 -1511 543 -1505
rect 481 -1545 493 -1511
rect 531 -1545 543 -1511
rect 481 -1551 543 -1545
rect 609 -1511 671 -1505
rect 609 -1545 621 -1511
rect 659 -1545 671 -1511
rect 609 -1551 671 -1545
rect 737 -1511 799 -1505
rect 737 -1545 749 -1511
rect 787 -1545 799 -1511
rect 737 -1551 799 -1545
rect 865 -1511 927 -1505
rect 865 -1545 877 -1511
rect 915 -1545 927 -1511
rect 865 -1551 927 -1545
rect 993 -1511 1055 -1505
rect 993 -1545 1005 -1511
rect 1043 -1545 1055 -1511
rect 993 -1551 1055 -1545
rect 1121 -1511 1183 -1505
rect 1121 -1545 1133 -1511
rect 1171 -1545 1183 -1511
rect 1121 -1551 1183 -1545
rect 1249 -1511 1311 -1505
rect 1249 -1545 1261 -1511
rect 1299 -1545 1311 -1511
rect 1249 -1551 1311 -1545
rect 1377 -1511 1439 -1505
rect 1377 -1545 1389 -1511
rect 1427 -1545 1439 -1511
rect 1377 -1551 1439 -1545
rect 1505 -1511 1567 -1505
rect 1505 -1545 1517 -1511
rect 1555 -1545 1567 -1511
rect 1505 -1551 1567 -1545
rect 1633 -1511 1695 -1505
rect 1633 -1545 1645 -1511
rect 1683 -1545 1695 -1511
rect 1633 -1551 1695 -1545
rect 1761 -1511 1823 -1505
rect 1761 -1545 1773 -1511
rect 1811 -1545 1823 -1511
rect 1761 -1551 1823 -1545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -1970 -1631 1970 1631
string parameters w 15 l 0.35 m 1 nf 29 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
