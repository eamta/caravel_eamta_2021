magic
tech sky130A
magscale 1 2
timestamp 1619113446
<< error_p >>
rect -1901 1787 -1843 1793
rect -1709 1787 -1651 1793
rect -1517 1787 -1459 1793
rect -1325 1787 -1267 1793
rect -1133 1787 -1075 1793
rect -941 1787 -883 1793
rect -749 1787 -691 1793
rect -557 1787 -499 1793
rect -365 1787 -307 1793
rect -173 1787 -115 1793
rect 19 1787 77 1793
rect 211 1787 269 1793
rect 403 1787 461 1793
rect 595 1787 653 1793
rect 787 1787 845 1793
rect 979 1787 1037 1793
rect 1171 1787 1229 1793
rect 1363 1787 1421 1793
rect 1555 1787 1613 1793
rect 1747 1787 1805 1793
rect -1901 1753 -1889 1787
rect -1709 1753 -1697 1787
rect -1517 1753 -1505 1787
rect -1325 1753 -1313 1787
rect -1133 1753 -1121 1787
rect -941 1753 -929 1787
rect -749 1753 -737 1787
rect -557 1753 -545 1787
rect -365 1753 -353 1787
rect -173 1753 -161 1787
rect 19 1753 31 1787
rect 211 1753 223 1787
rect 403 1753 415 1787
rect 595 1753 607 1787
rect 787 1753 799 1787
rect 979 1753 991 1787
rect 1171 1753 1183 1787
rect 1363 1753 1375 1787
rect 1555 1753 1567 1787
rect 1747 1753 1759 1787
rect -1901 1747 -1843 1753
rect -1709 1747 -1651 1753
rect -1517 1747 -1459 1753
rect -1325 1747 -1267 1753
rect -1133 1747 -1075 1753
rect -941 1747 -883 1753
rect -749 1747 -691 1753
rect -557 1747 -499 1753
rect -365 1747 -307 1753
rect -173 1747 -115 1753
rect 19 1747 77 1753
rect 211 1747 269 1753
rect 403 1747 461 1753
rect 595 1747 653 1753
rect 787 1747 845 1753
rect 979 1747 1037 1753
rect 1171 1747 1229 1753
rect 1363 1747 1421 1753
rect 1555 1747 1613 1753
rect 1747 1747 1805 1753
rect -1805 1287 -1747 1293
rect -1613 1287 -1555 1293
rect -1421 1287 -1363 1293
rect -1229 1287 -1171 1293
rect -1037 1287 -979 1293
rect -845 1287 -787 1293
rect -653 1287 -595 1293
rect -461 1287 -403 1293
rect -269 1287 -211 1293
rect -77 1287 -19 1293
rect 115 1287 173 1293
rect 307 1287 365 1293
rect 499 1287 557 1293
rect 691 1287 749 1293
rect 883 1287 941 1293
rect 1075 1287 1133 1293
rect 1267 1287 1325 1293
rect 1459 1287 1517 1293
rect 1651 1287 1709 1293
rect 1843 1287 1901 1293
rect -1805 1253 -1793 1287
rect -1613 1253 -1601 1287
rect -1421 1253 -1409 1287
rect -1229 1253 -1217 1287
rect -1037 1253 -1025 1287
rect -845 1253 -833 1287
rect -653 1253 -641 1287
rect -461 1253 -449 1287
rect -269 1253 -257 1287
rect -77 1253 -65 1287
rect 115 1253 127 1287
rect 307 1253 319 1287
rect 499 1253 511 1287
rect 691 1253 703 1287
rect 883 1253 895 1287
rect 1075 1253 1087 1287
rect 1267 1253 1279 1287
rect 1459 1253 1471 1287
rect 1651 1253 1663 1287
rect 1843 1253 1855 1287
rect -1805 1247 -1747 1253
rect -1613 1247 -1555 1253
rect -1421 1247 -1363 1253
rect -1229 1247 -1171 1253
rect -1037 1247 -979 1253
rect -845 1247 -787 1253
rect -653 1247 -595 1253
rect -461 1247 -403 1253
rect -269 1247 -211 1253
rect -77 1247 -19 1253
rect 115 1247 173 1253
rect 307 1247 365 1253
rect 499 1247 557 1253
rect 691 1247 749 1253
rect 883 1247 941 1253
rect 1075 1247 1133 1253
rect 1267 1247 1325 1253
rect 1459 1247 1517 1253
rect 1651 1247 1709 1253
rect 1843 1247 1901 1253
rect -1805 1179 -1747 1185
rect -1613 1179 -1555 1185
rect -1421 1179 -1363 1185
rect -1229 1179 -1171 1185
rect -1037 1179 -979 1185
rect -845 1179 -787 1185
rect -653 1179 -595 1185
rect -461 1179 -403 1185
rect -269 1179 -211 1185
rect -77 1179 -19 1185
rect 115 1179 173 1185
rect 307 1179 365 1185
rect 499 1179 557 1185
rect 691 1179 749 1185
rect 883 1179 941 1185
rect 1075 1179 1133 1185
rect 1267 1179 1325 1185
rect 1459 1179 1517 1185
rect 1651 1179 1709 1185
rect 1843 1179 1901 1185
rect -1805 1145 -1793 1179
rect -1613 1145 -1601 1179
rect -1421 1145 -1409 1179
rect -1229 1145 -1217 1179
rect -1037 1145 -1025 1179
rect -845 1145 -833 1179
rect -653 1145 -641 1179
rect -461 1145 -449 1179
rect -269 1145 -257 1179
rect -77 1145 -65 1179
rect 115 1145 127 1179
rect 307 1145 319 1179
rect 499 1145 511 1179
rect 691 1145 703 1179
rect 883 1145 895 1179
rect 1075 1145 1087 1179
rect 1267 1145 1279 1179
rect 1459 1145 1471 1179
rect 1651 1145 1663 1179
rect 1843 1145 1855 1179
rect -1805 1139 -1747 1145
rect -1613 1139 -1555 1145
rect -1421 1139 -1363 1145
rect -1229 1139 -1171 1145
rect -1037 1139 -979 1145
rect -845 1139 -787 1145
rect -653 1139 -595 1145
rect -461 1139 -403 1145
rect -269 1139 -211 1145
rect -77 1139 -19 1145
rect 115 1139 173 1145
rect 307 1139 365 1145
rect 499 1139 557 1145
rect 691 1139 749 1145
rect 883 1139 941 1145
rect 1075 1139 1133 1145
rect 1267 1139 1325 1145
rect 1459 1139 1517 1145
rect 1651 1139 1709 1145
rect 1843 1139 1901 1145
rect -1901 679 -1843 685
rect -1709 679 -1651 685
rect -1517 679 -1459 685
rect -1325 679 -1267 685
rect -1133 679 -1075 685
rect -941 679 -883 685
rect -749 679 -691 685
rect -557 679 -499 685
rect -365 679 -307 685
rect -173 679 -115 685
rect 19 679 77 685
rect 211 679 269 685
rect 403 679 461 685
rect 595 679 653 685
rect 787 679 845 685
rect 979 679 1037 685
rect 1171 679 1229 685
rect 1363 679 1421 685
rect 1555 679 1613 685
rect 1747 679 1805 685
rect -1901 645 -1889 679
rect -1709 645 -1697 679
rect -1517 645 -1505 679
rect -1325 645 -1313 679
rect -1133 645 -1121 679
rect -941 645 -929 679
rect -749 645 -737 679
rect -557 645 -545 679
rect -365 645 -353 679
rect -173 645 -161 679
rect 19 645 31 679
rect 211 645 223 679
rect 403 645 415 679
rect 595 645 607 679
rect 787 645 799 679
rect 979 645 991 679
rect 1171 645 1183 679
rect 1363 645 1375 679
rect 1555 645 1567 679
rect 1747 645 1759 679
rect -1901 639 -1843 645
rect -1709 639 -1651 645
rect -1517 639 -1459 645
rect -1325 639 -1267 645
rect -1133 639 -1075 645
rect -941 639 -883 645
rect -749 639 -691 645
rect -557 639 -499 645
rect -365 639 -307 645
rect -173 639 -115 645
rect 19 639 77 645
rect 211 639 269 645
rect 403 639 461 645
rect 595 639 653 645
rect 787 639 845 645
rect 979 639 1037 645
rect 1171 639 1229 645
rect 1363 639 1421 645
rect 1555 639 1613 645
rect 1747 639 1805 645
rect -1901 571 -1843 577
rect -1709 571 -1651 577
rect -1517 571 -1459 577
rect -1325 571 -1267 577
rect -1133 571 -1075 577
rect -941 571 -883 577
rect -749 571 -691 577
rect -557 571 -499 577
rect -365 571 -307 577
rect -173 571 -115 577
rect 19 571 77 577
rect 211 571 269 577
rect 403 571 461 577
rect 595 571 653 577
rect 787 571 845 577
rect 979 571 1037 577
rect 1171 571 1229 577
rect 1363 571 1421 577
rect 1555 571 1613 577
rect 1747 571 1805 577
rect -1901 537 -1889 571
rect -1709 537 -1697 571
rect -1517 537 -1505 571
rect -1325 537 -1313 571
rect -1133 537 -1121 571
rect -941 537 -929 571
rect -749 537 -737 571
rect -557 537 -545 571
rect -365 537 -353 571
rect -173 537 -161 571
rect 19 537 31 571
rect 211 537 223 571
rect 403 537 415 571
rect 595 537 607 571
rect 787 537 799 571
rect 979 537 991 571
rect 1171 537 1183 571
rect 1363 537 1375 571
rect 1555 537 1567 571
rect 1747 537 1759 571
rect -1901 531 -1843 537
rect -1709 531 -1651 537
rect -1517 531 -1459 537
rect -1325 531 -1267 537
rect -1133 531 -1075 537
rect -941 531 -883 537
rect -749 531 -691 537
rect -557 531 -499 537
rect -365 531 -307 537
rect -173 531 -115 537
rect 19 531 77 537
rect 211 531 269 537
rect 403 531 461 537
rect 595 531 653 537
rect 787 531 845 537
rect 979 531 1037 537
rect 1171 531 1229 537
rect 1363 531 1421 537
rect 1555 531 1613 537
rect 1747 531 1805 537
rect -1805 71 -1747 77
rect -1613 71 -1555 77
rect -1421 71 -1363 77
rect -1229 71 -1171 77
rect -1037 71 -979 77
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect 1075 71 1133 77
rect 1267 71 1325 77
rect 1459 71 1517 77
rect 1651 71 1709 77
rect 1843 71 1901 77
rect -1805 37 -1793 71
rect -1613 37 -1601 71
rect -1421 37 -1409 71
rect -1229 37 -1217 71
rect -1037 37 -1025 71
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect 1075 37 1087 71
rect 1267 37 1279 71
rect 1459 37 1471 71
rect 1651 37 1663 71
rect 1843 37 1855 71
rect -1805 31 -1747 37
rect -1613 31 -1555 37
rect -1421 31 -1363 37
rect -1229 31 -1171 37
rect -1037 31 -979 37
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect 1075 31 1133 37
rect 1267 31 1325 37
rect 1459 31 1517 37
rect 1651 31 1709 37
rect 1843 31 1901 37
rect -1805 -37 -1747 -31
rect -1613 -37 -1555 -31
rect -1421 -37 -1363 -31
rect -1229 -37 -1171 -31
rect -1037 -37 -979 -31
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect 1075 -37 1133 -31
rect 1267 -37 1325 -31
rect 1459 -37 1517 -31
rect 1651 -37 1709 -31
rect 1843 -37 1901 -31
rect -1805 -71 -1793 -37
rect -1613 -71 -1601 -37
rect -1421 -71 -1409 -37
rect -1229 -71 -1217 -37
rect -1037 -71 -1025 -37
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect 1075 -71 1087 -37
rect 1267 -71 1279 -37
rect 1459 -71 1471 -37
rect 1651 -71 1663 -37
rect 1843 -71 1855 -37
rect -1805 -77 -1747 -71
rect -1613 -77 -1555 -71
rect -1421 -77 -1363 -71
rect -1229 -77 -1171 -71
rect -1037 -77 -979 -71
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect 1075 -77 1133 -71
rect 1267 -77 1325 -71
rect 1459 -77 1517 -71
rect 1651 -77 1709 -71
rect 1843 -77 1901 -71
rect -1901 -537 -1843 -531
rect -1709 -537 -1651 -531
rect -1517 -537 -1459 -531
rect -1325 -537 -1267 -531
rect -1133 -537 -1075 -531
rect -941 -537 -883 -531
rect -749 -537 -691 -531
rect -557 -537 -499 -531
rect -365 -537 -307 -531
rect -173 -537 -115 -531
rect 19 -537 77 -531
rect 211 -537 269 -531
rect 403 -537 461 -531
rect 595 -537 653 -531
rect 787 -537 845 -531
rect 979 -537 1037 -531
rect 1171 -537 1229 -531
rect 1363 -537 1421 -531
rect 1555 -537 1613 -531
rect 1747 -537 1805 -531
rect -1901 -571 -1889 -537
rect -1709 -571 -1697 -537
rect -1517 -571 -1505 -537
rect -1325 -571 -1313 -537
rect -1133 -571 -1121 -537
rect -941 -571 -929 -537
rect -749 -571 -737 -537
rect -557 -571 -545 -537
rect -365 -571 -353 -537
rect -173 -571 -161 -537
rect 19 -571 31 -537
rect 211 -571 223 -537
rect 403 -571 415 -537
rect 595 -571 607 -537
rect 787 -571 799 -537
rect 979 -571 991 -537
rect 1171 -571 1183 -537
rect 1363 -571 1375 -537
rect 1555 -571 1567 -537
rect 1747 -571 1759 -537
rect -1901 -577 -1843 -571
rect -1709 -577 -1651 -571
rect -1517 -577 -1459 -571
rect -1325 -577 -1267 -571
rect -1133 -577 -1075 -571
rect -941 -577 -883 -571
rect -749 -577 -691 -571
rect -557 -577 -499 -571
rect -365 -577 -307 -571
rect -173 -577 -115 -571
rect 19 -577 77 -571
rect 211 -577 269 -571
rect 403 -577 461 -571
rect 595 -577 653 -571
rect 787 -577 845 -571
rect 979 -577 1037 -571
rect 1171 -577 1229 -571
rect 1363 -577 1421 -571
rect 1555 -577 1613 -571
rect 1747 -577 1805 -571
rect -1901 -645 -1843 -639
rect -1709 -645 -1651 -639
rect -1517 -645 -1459 -639
rect -1325 -645 -1267 -639
rect -1133 -645 -1075 -639
rect -941 -645 -883 -639
rect -749 -645 -691 -639
rect -557 -645 -499 -639
rect -365 -645 -307 -639
rect -173 -645 -115 -639
rect 19 -645 77 -639
rect 211 -645 269 -639
rect 403 -645 461 -639
rect 595 -645 653 -639
rect 787 -645 845 -639
rect 979 -645 1037 -639
rect 1171 -645 1229 -639
rect 1363 -645 1421 -639
rect 1555 -645 1613 -639
rect 1747 -645 1805 -639
rect -1901 -679 -1889 -645
rect -1709 -679 -1697 -645
rect -1517 -679 -1505 -645
rect -1325 -679 -1313 -645
rect -1133 -679 -1121 -645
rect -941 -679 -929 -645
rect -749 -679 -737 -645
rect -557 -679 -545 -645
rect -365 -679 -353 -645
rect -173 -679 -161 -645
rect 19 -679 31 -645
rect 211 -679 223 -645
rect 403 -679 415 -645
rect 595 -679 607 -645
rect 787 -679 799 -645
rect 979 -679 991 -645
rect 1171 -679 1183 -645
rect 1363 -679 1375 -645
rect 1555 -679 1567 -645
rect 1747 -679 1759 -645
rect -1901 -685 -1843 -679
rect -1709 -685 -1651 -679
rect -1517 -685 -1459 -679
rect -1325 -685 -1267 -679
rect -1133 -685 -1075 -679
rect -941 -685 -883 -679
rect -749 -685 -691 -679
rect -557 -685 -499 -679
rect -365 -685 -307 -679
rect -173 -685 -115 -679
rect 19 -685 77 -679
rect 211 -685 269 -679
rect 403 -685 461 -679
rect 595 -685 653 -679
rect 787 -685 845 -679
rect 979 -685 1037 -679
rect 1171 -685 1229 -679
rect 1363 -685 1421 -679
rect 1555 -685 1613 -679
rect 1747 -685 1805 -679
rect -1805 -1145 -1747 -1139
rect -1613 -1145 -1555 -1139
rect -1421 -1145 -1363 -1139
rect -1229 -1145 -1171 -1139
rect -1037 -1145 -979 -1139
rect -845 -1145 -787 -1139
rect -653 -1145 -595 -1139
rect -461 -1145 -403 -1139
rect -269 -1145 -211 -1139
rect -77 -1145 -19 -1139
rect 115 -1145 173 -1139
rect 307 -1145 365 -1139
rect 499 -1145 557 -1139
rect 691 -1145 749 -1139
rect 883 -1145 941 -1139
rect 1075 -1145 1133 -1139
rect 1267 -1145 1325 -1139
rect 1459 -1145 1517 -1139
rect 1651 -1145 1709 -1139
rect 1843 -1145 1901 -1139
rect -1805 -1179 -1793 -1145
rect -1613 -1179 -1601 -1145
rect -1421 -1179 -1409 -1145
rect -1229 -1179 -1217 -1145
rect -1037 -1179 -1025 -1145
rect -845 -1179 -833 -1145
rect -653 -1179 -641 -1145
rect -461 -1179 -449 -1145
rect -269 -1179 -257 -1145
rect -77 -1179 -65 -1145
rect 115 -1179 127 -1145
rect 307 -1179 319 -1145
rect 499 -1179 511 -1145
rect 691 -1179 703 -1145
rect 883 -1179 895 -1145
rect 1075 -1179 1087 -1145
rect 1267 -1179 1279 -1145
rect 1459 -1179 1471 -1145
rect 1651 -1179 1663 -1145
rect 1843 -1179 1855 -1145
rect -1805 -1185 -1747 -1179
rect -1613 -1185 -1555 -1179
rect -1421 -1185 -1363 -1179
rect -1229 -1185 -1171 -1179
rect -1037 -1185 -979 -1179
rect -845 -1185 -787 -1179
rect -653 -1185 -595 -1179
rect -461 -1185 -403 -1179
rect -269 -1185 -211 -1179
rect -77 -1185 -19 -1179
rect 115 -1185 173 -1179
rect 307 -1185 365 -1179
rect 499 -1185 557 -1179
rect 691 -1185 749 -1179
rect 883 -1185 941 -1179
rect 1075 -1185 1133 -1179
rect 1267 -1185 1325 -1179
rect 1459 -1185 1517 -1179
rect 1651 -1185 1709 -1179
rect 1843 -1185 1901 -1179
rect -1805 -1253 -1747 -1247
rect -1613 -1253 -1555 -1247
rect -1421 -1253 -1363 -1247
rect -1229 -1253 -1171 -1247
rect -1037 -1253 -979 -1247
rect -845 -1253 -787 -1247
rect -653 -1253 -595 -1247
rect -461 -1253 -403 -1247
rect -269 -1253 -211 -1247
rect -77 -1253 -19 -1247
rect 115 -1253 173 -1247
rect 307 -1253 365 -1247
rect 499 -1253 557 -1247
rect 691 -1253 749 -1247
rect 883 -1253 941 -1247
rect 1075 -1253 1133 -1247
rect 1267 -1253 1325 -1247
rect 1459 -1253 1517 -1247
rect 1651 -1253 1709 -1247
rect 1843 -1253 1901 -1247
rect -1805 -1287 -1793 -1253
rect -1613 -1287 -1601 -1253
rect -1421 -1287 -1409 -1253
rect -1229 -1287 -1217 -1253
rect -1037 -1287 -1025 -1253
rect -845 -1287 -833 -1253
rect -653 -1287 -641 -1253
rect -461 -1287 -449 -1253
rect -269 -1287 -257 -1253
rect -77 -1287 -65 -1253
rect 115 -1287 127 -1253
rect 307 -1287 319 -1253
rect 499 -1287 511 -1253
rect 691 -1287 703 -1253
rect 883 -1287 895 -1253
rect 1075 -1287 1087 -1253
rect 1267 -1287 1279 -1253
rect 1459 -1287 1471 -1253
rect 1651 -1287 1663 -1253
rect 1843 -1287 1855 -1253
rect -1805 -1293 -1747 -1287
rect -1613 -1293 -1555 -1287
rect -1421 -1293 -1363 -1287
rect -1229 -1293 -1171 -1287
rect -1037 -1293 -979 -1287
rect -845 -1293 -787 -1287
rect -653 -1293 -595 -1287
rect -461 -1293 -403 -1287
rect -269 -1293 -211 -1287
rect -77 -1293 -19 -1287
rect 115 -1293 173 -1287
rect 307 -1293 365 -1287
rect 499 -1293 557 -1287
rect 691 -1293 749 -1287
rect 883 -1293 941 -1287
rect 1075 -1293 1133 -1287
rect 1267 -1293 1325 -1287
rect 1459 -1293 1517 -1287
rect 1651 -1293 1709 -1287
rect 1843 -1293 1901 -1287
rect -1901 -1753 -1843 -1747
rect -1709 -1753 -1651 -1747
rect -1517 -1753 -1459 -1747
rect -1325 -1753 -1267 -1747
rect -1133 -1753 -1075 -1747
rect -941 -1753 -883 -1747
rect -749 -1753 -691 -1747
rect -557 -1753 -499 -1747
rect -365 -1753 -307 -1747
rect -173 -1753 -115 -1747
rect 19 -1753 77 -1747
rect 211 -1753 269 -1747
rect 403 -1753 461 -1747
rect 595 -1753 653 -1747
rect 787 -1753 845 -1747
rect 979 -1753 1037 -1747
rect 1171 -1753 1229 -1747
rect 1363 -1753 1421 -1747
rect 1555 -1753 1613 -1747
rect 1747 -1753 1805 -1747
rect -1901 -1787 -1889 -1753
rect -1709 -1787 -1697 -1753
rect -1517 -1787 -1505 -1753
rect -1325 -1787 -1313 -1753
rect -1133 -1787 -1121 -1753
rect -941 -1787 -929 -1753
rect -749 -1787 -737 -1753
rect -557 -1787 -545 -1753
rect -365 -1787 -353 -1753
rect -173 -1787 -161 -1753
rect 19 -1787 31 -1753
rect 211 -1787 223 -1753
rect 403 -1787 415 -1753
rect 595 -1787 607 -1753
rect 787 -1787 799 -1753
rect 979 -1787 991 -1753
rect 1171 -1787 1183 -1753
rect 1363 -1787 1375 -1753
rect 1555 -1787 1567 -1753
rect 1747 -1787 1759 -1753
rect -1901 -1793 -1843 -1787
rect -1709 -1793 -1651 -1787
rect -1517 -1793 -1459 -1787
rect -1325 -1793 -1267 -1787
rect -1133 -1793 -1075 -1787
rect -941 -1793 -883 -1787
rect -749 -1793 -691 -1787
rect -557 -1793 -499 -1787
rect -365 -1793 -307 -1787
rect -173 -1793 -115 -1787
rect 19 -1793 77 -1787
rect 211 -1793 269 -1787
rect 403 -1793 461 -1787
rect 595 -1793 653 -1787
rect 787 -1793 845 -1787
rect 979 -1793 1037 -1787
rect 1171 -1793 1229 -1787
rect 1363 -1793 1421 -1787
rect 1555 -1793 1613 -1787
rect 1747 -1793 1805 -1787
<< pwell >>
rect -2087 -1925 2087 1925
<< nmos >>
rect -1887 1325 -1857 1715
rect -1791 1325 -1761 1715
rect -1695 1325 -1665 1715
rect -1599 1325 -1569 1715
rect -1503 1325 -1473 1715
rect -1407 1325 -1377 1715
rect -1311 1325 -1281 1715
rect -1215 1325 -1185 1715
rect -1119 1325 -1089 1715
rect -1023 1325 -993 1715
rect -927 1325 -897 1715
rect -831 1325 -801 1715
rect -735 1325 -705 1715
rect -639 1325 -609 1715
rect -543 1325 -513 1715
rect -447 1325 -417 1715
rect -351 1325 -321 1715
rect -255 1325 -225 1715
rect -159 1325 -129 1715
rect -63 1325 -33 1715
rect 33 1325 63 1715
rect 129 1325 159 1715
rect 225 1325 255 1715
rect 321 1325 351 1715
rect 417 1325 447 1715
rect 513 1325 543 1715
rect 609 1325 639 1715
rect 705 1325 735 1715
rect 801 1325 831 1715
rect 897 1325 927 1715
rect 993 1325 1023 1715
rect 1089 1325 1119 1715
rect 1185 1325 1215 1715
rect 1281 1325 1311 1715
rect 1377 1325 1407 1715
rect 1473 1325 1503 1715
rect 1569 1325 1599 1715
rect 1665 1325 1695 1715
rect 1761 1325 1791 1715
rect 1857 1325 1887 1715
rect -1887 717 -1857 1107
rect -1791 717 -1761 1107
rect -1695 717 -1665 1107
rect -1599 717 -1569 1107
rect -1503 717 -1473 1107
rect -1407 717 -1377 1107
rect -1311 717 -1281 1107
rect -1215 717 -1185 1107
rect -1119 717 -1089 1107
rect -1023 717 -993 1107
rect -927 717 -897 1107
rect -831 717 -801 1107
rect -735 717 -705 1107
rect -639 717 -609 1107
rect -543 717 -513 1107
rect -447 717 -417 1107
rect -351 717 -321 1107
rect -255 717 -225 1107
rect -159 717 -129 1107
rect -63 717 -33 1107
rect 33 717 63 1107
rect 129 717 159 1107
rect 225 717 255 1107
rect 321 717 351 1107
rect 417 717 447 1107
rect 513 717 543 1107
rect 609 717 639 1107
rect 705 717 735 1107
rect 801 717 831 1107
rect 897 717 927 1107
rect 993 717 1023 1107
rect 1089 717 1119 1107
rect 1185 717 1215 1107
rect 1281 717 1311 1107
rect 1377 717 1407 1107
rect 1473 717 1503 1107
rect 1569 717 1599 1107
rect 1665 717 1695 1107
rect 1761 717 1791 1107
rect 1857 717 1887 1107
rect -1887 109 -1857 499
rect -1791 109 -1761 499
rect -1695 109 -1665 499
rect -1599 109 -1569 499
rect -1503 109 -1473 499
rect -1407 109 -1377 499
rect -1311 109 -1281 499
rect -1215 109 -1185 499
rect -1119 109 -1089 499
rect -1023 109 -993 499
rect -927 109 -897 499
rect -831 109 -801 499
rect -735 109 -705 499
rect -639 109 -609 499
rect -543 109 -513 499
rect -447 109 -417 499
rect -351 109 -321 499
rect -255 109 -225 499
rect -159 109 -129 499
rect -63 109 -33 499
rect 33 109 63 499
rect 129 109 159 499
rect 225 109 255 499
rect 321 109 351 499
rect 417 109 447 499
rect 513 109 543 499
rect 609 109 639 499
rect 705 109 735 499
rect 801 109 831 499
rect 897 109 927 499
rect 993 109 1023 499
rect 1089 109 1119 499
rect 1185 109 1215 499
rect 1281 109 1311 499
rect 1377 109 1407 499
rect 1473 109 1503 499
rect 1569 109 1599 499
rect 1665 109 1695 499
rect 1761 109 1791 499
rect 1857 109 1887 499
rect -1887 -499 -1857 -109
rect -1791 -499 -1761 -109
rect -1695 -499 -1665 -109
rect -1599 -499 -1569 -109
rect -1503 -499 -1473 -109
rect -1407 -499 -1377 -109
rect -1311 -499 -1281 -109
rect -1215 -499 -1185 -109
rect -1119 -499 -1089 -109
rect -1023 -499 -993 -109
rect -927 -499 -897 -109
rect -831 -499 -801 -109
rect -735 -499 -705 -109
rect -639 -499 -609 -109
rect -543 -499 -513 -109
rect -447 -499 -417 -109
rect -351 -499 -321 -109
rect -255 -499 -225 -109
rect -159 -499 -129 -109
rect -63 -499 -33 -109
rect 33 -499 63 -109
rect 129 -499 159 -109
rect 225 -499 255 -109
rect 321 -499 351 -109
rect 417 -499 447 -109
rect 513 -499 543 -109
rect 609 -499 639 -109
rect 705 -499 735 -109
rect 801 -499 831 -109
rect 897 -499 927 -109
rect 993 -499 1023 -109
rect 1089 -499 1119 -109
rect 1185 -499 1215 -109
rect 1281 -499 1311 -109
rect 1377 -499 1407 -109
rect 1473 -499 1503 -109
rect 1569 -499 1599 -109
rect 1665 -499 1695 -109
rect 1761 -499 1791 -109
rect 1857 -499 1887 -109
rect -1887 -1107 -1857 -717
rect -1791 -1107 -1761 -717
rect -1695 -1107 -1665 -717
rect -1599 -1107 -1569 -717
rect -1503 -1107 -1473 -717
rect -1407 -1107 -1377 -717
rect -1311 -1107 -1281 -717
rect -1215 -1107 -1185 -717
rect -1119 -1107 -1089 -717
rect -1023 -1107 -993 -717
rect -927 -1107 -897 -717
rect -831 -1107 -801 -717
rect -735 -1107 -705 -717
rect -639 -1107 -609 -717
rect -543 -1107 -513 -717
rect -447 -1107 -417 -717
rect -351 -1107 -321 -717
rect -255 -1107 -225 -717
rect -159 -1107 -129 -717
rect -63 -1107 -33 -717
rect 33 -1107 63 -717
rect 129 -1107 159 -717
rect 225 -1107 255 -717
rect 321 -1107 351 -717
rect 417 -1107 447 -717
rect 513 -1107 543 -717
rect 609 -1107 639 -717
rect 705 -1107 735 -717
rect 801 -1107 831 -717
rect 897 -1107 927 -717
rect 993 -1107 1023 -717
rect 1089 -1107 1119 -717
rect 1185 -1107 1215 -717
rect 1281 -1107 1311 -717
rect 1377 -1107 1407 -717
rect 1473 -1107 1503 -717
rect 1569 -1107 1599 -717
rect 1665 -1107 1695 -717
rect 1761 -1107 1791 -717
rect 1857 -1107 1887 -717
rect -1887 -1715 -1857 -1325
rect -1791 -1715 -1761 -1325
rect -1695 -1715 -1665 -1325
rect -1599 -1715 -1569 -1325
rect -1503 -1715 -1473 -1325
rect -1407 -1715 -1377 -1325
rect -1311 -1715 -1281 -1325
rect -1215 -1715 -1185 -1325
rect -1119 -1715 -1089 -1325
rect -1023 -1715 -993 -1325
rect -927 -1715 -897 -1325
rect -831 -1715 -801 -1325
rect -735 -1715 -705 -1325
rect -639 -1715 -609 -1325
rect -543 -1715 -513 -1325
rect -447 -1715 -417 -1325
rect -351 -1715 -321 -1325
rect -255 -1715 -225 -1325
rect -159 -1715 -129 -1325
rect -63 -1715 -33 -1325
rect 33 -1715 63 -1325
rect 129 -1715 159 -1325
rect 225 -1715 255 -1325
rect 321 -1715 351 -1325
rect 417 -1715 447 -1325
rect 513 -1715 543 -1325
rect 609 -1715 639 -1325
rect 705 -1715 735 -1325
rect 801 -1715 831 -1325
rect 897 -1715 927 -1325
rect 993 -1715 1023 -1325
rect 1089 -1715 1119 -1325
rect 1185 -1715 1215 -1325
rect 1281 -1715 1311 -1325
rect 1377 -1715 1407 -1325
rect 1473 -1715 1503 -1325
rect 1569 -1715 1599 -1325
rect 1665 -1715 1695 -1325
rect 1761 -1715 1791 -1325
rect 1857 -1715 1887 -1325
<< ndiff >>
rect -1949 1703 -1887 1715
rect -1949 1337 -1937 1703
rect -1903 1337 -1887 1703
rect -1949 1325 -1887 1337
rect -1857 1703 -1791 1715
rect -1857 1337 -1841 1703
rect -1807 1337 -1791 1703
rect -1857 1325 -1791 1337
rect -1761 1703 -1695 1715
rect -1761 1337 -1745 1703
rect -1711 1337 -1695 1703
rect -1761 1325 -1695 1337
rect -1665 1703 -1599 1715
rect -1665 1337 -1649 1703
rect -1615 1337 -1599 1703
rect -1665 1325 -1599 1337
rect -1569 1703 -1503 1715
rect -1569 1337 -1553 1703
rect -1519 1337 -1503 1703
rect -1569 1325 -1503 1337
rect -1473 1703 -1407 1715
rect -1473 1337 -1457 1703
rect -1423 1337 -1407 1703
rect -1473 1325 -1407 1337
rect -1377 1703 -1311 1715
rect -1377 1337 -1361 1703
rect -1327 1337 -1311 1703
rect -1377 1325 -1311 1337
rect -1281 1703 -1215 1715
rect -1281 1337 -1265 1703
rect -1231 1337 -1215 1703
rect -1281 1325 -1215 1337
rect -1185 1703 -1119 1715
rect -1185 1337 -1169 1703
rect -1135 1337 -1119 1703
rect -1185 1325 -1119 1337
rect -1089 1703 -1023 1715
rect -1089 1337 -1073 1703
rect -1039 1337 -1023 1703
rect -1089 1325 -1023 1337
rect -993 1703 -927 1715
rect -993 1337 -977 1703
rect -943 1337 -927 1703
rect -993 1325 -927 1337
rect -897 1703 -831 1715
rect -897 1337 -881 1703
rect -847 1337 -831 1703
rect -897 1325 -831 1337
rect -801 1703 -735 1715
rect -801 1337 -785 1703
rect -751 1337 -735 1703
rect -801 1325 -735 1337
rect -705 1703 -639 1715
rect -705 1337 -689 1703
rect -655 1337 -639 1703
rect -705 1325 -639 1337
rect -609 1703 -543 1715
rect -609 1337 -593 1703
rect -559 1337 -543 1703
rect -609 1325 -543 1337
rect -513 1703 -447 1715
rect -513 1337 -497 1703
rect -463 1337 -447 1703
rect -513 1325 -447 1337
rect -417 1703 -351 1715
rect -417 1337 -401 1703
rect -367 1337 -351 1703
rect -417 1325 -351 1337
rect -321 1703 -255 1715
rect -321 1337 -305 1703
rect -271 1337 -255 1703
rect -321 1325 -255 1337
rect -225 1703 -159 1715
rect -225 1337 -209 1703
rect -175 1337 -159 1703
rect -225 1325 -159 1337
rect -129 1703 -63 1715
rect -129 1337 -113 1703
rect -79 1337 -63 1703
rect -129 1325 -63 1337
rect -33 1703 33 1715
rect -33 1337 -17 1703
rect 17 1337 33 1703
rect -33 1325 33 1337
rect 63 1703 129 1715
rect 63 1337 79 1703
rect 113 1337 129 1703
rect 63 1325 129 1337
rect 159 1703 225 1715
rect 159 1337 175 1703
rect 209 1337 225 1703
rect 159 1325 225 1337
rect 255 1703 321 1715
rect 255 1337 271 1703
rect 305 1337 321 1703
rect 255 1325 321 1337
rect 351 1703 417 1715
rect 351 1337 367 1703
rect 401 1337 417 1703
rect 351 1325 417 1337
rect 447 1703 513 1715
rect 447 1337 463 1703
rect 497 1337 513 1703
rect 447 1325 513 1337
rect 543 1703 609 1715
rect 543 1337 559 1703
rect 593 1337 609 1703
rect 543 1325 609 1337
rect 639 1703 705 1715
rect 639 1337 655 1703
rect 689 1337 705 1703
rect 639 1325 705 1337
rect 735 1703 801 1715
rect 735 1337 751 1703
rect 785 1337 801 1703
rect 735 1325 801 1337
rect 831 1703 897 1715
rect 831 1337 847 1703
rect 881 1337 897 1703
rect 831 1325 897 1337
rect 927 1703 993 1715
rect 927 1337 943 1703
rect 977 1337 993 1703
rect 927 1325 993 1337
rect 1023 1703 1089 1715
rect 1023 1337 1039 1703
rect 1073 1337 1089 1703
rect 1023 1325 1089 1337
rect 1119 1703 1185 1715
rect 1119 1337 1135 1703
rect 1169 1337 1185 1703
rect 1119 1325 1185 1337
rect 1215 1703 1281 1715
rect 1215 1337 1231 1703
rect 1265 1337 1281 1703
rect 1215 1325 1281 1337
rect 1311 1703 1377 1715
rect 1311 1337 1327 1703
rect 1361 1337 1377 1703
rect 1311 1325 1377 1337
rect 1407 1703 1473 1715
rect 1407 1337 1423 1703
rect 1457 1337 1473 1703
rect 1407 1325 1473 1337
rect 1503 1703 1569 1715
rect 1503 1337 1519 1703
rect 1553 1337 1569 1703
rect 1503 1325 1569 1337
rect 1599 1703 1665 1715
rect 1599 1337 1615 1703
rect 1649 1337 1665 1703
rect 1599 1325 1665 1337
rect 1695 1703 1761 1715
rect 1695 1337 1711 1703
rect 1745 1337 1761 1703
rect 1695 1325 1761 1337
rect 1791 1703 1857 1715
rect 1791 1337 1807 1703
rect 1841 1337 1857 1703
rect 1791 1325 1857 1337
rect 1887 1703 1949 1715
rect 1887 1337 1903 1703
rect 1937 1337 1949 1703
rect 1887 1325 1949 1337
rect -1949 1095 -1887 1107
rect -1949 729 -1937 1095
rect -1903 729 -1887 1095
rect -1949 717 -1887 729
rect -1857 1095 -1791 1107
rect -1857 729 -1841 1095
rect -1807 729 -1791 1095
rect -1857 717 -1791 729
rect -1761 1095 -1695 1107
rect -1761 729 -1745 1095
rect -1711 729 -1695 1095
rect -1761 717 -1695 729
rect -1665 1095 -1599 1107
rect -1665 729 -1649 1095
rect -1615 729 -1599 1095
rect -1665 717 -1599 729
rect -1569 1095 -1503 1107
rect -1569 729 -1553 1095
rect -1519 729 -1503 1095
rect -1569 717 -1503 729
rect -1473 1095 -1407 1107
rect -1473 729 -1457 1095
rect -1423 729 -1407 1095
rect -1473 717 -1407 729
rect -1377 1095 -1311 1107
rect -1377 729 -1361 1095
rect -1327 729 -1311 1095
rect -1377 717 -1311 729
rect -1281 1095 -1215 1107
rect -1281 729 -1265 1095
rect -1231 729 -1215 1095
rect -1281 717 -1215 729
rect -1185 1095 -1119 1107
rect -1185 729 -1169 1095
rect -1135 729 -1119 1095
rect -1185 717 -1119 729
rect -1089 1095 -1023 1107
rect -1089 729 -1073 1095
rect -1039 729 -1023 1095
rect -1089 717 -1023 729
rect -993 1095 -927 1107
rect -993 729 -977 1095
rect -943 729 -927 1095
rect -993 717 -927 729
rect -897 1095 -831 1107
rect -897 729 -881 1095
rect -847 729 -831 1095
rect -897 717 -831 729
rect -801 1095 -735 1107
rect -801 729 -785 1095
rect -751 729 -735 1095
rect -801 717 -735 729
rect -705 1095 -639 1107
rect -705 729 -689 1095
rect -655 729 -639 1095
rect -705 717 -639 729
rect -609 1095 -543 1107
rect -609 729 -593 1095
rect -559 729 -543 1095
rect -609 717 -543 729
rect -513 1095 -447 1107
rect -513 729 -497 1095
rect -463 729 -447 1095
rect -513 717 -447 729
rect -417 1095 -351 1107
rect -417 729 -401 1095
rect -367 729 -351 1095
rect -417 717 -351 729
rect -321 1095 -255 1107
rect -321 729 -305 1095
rect -271 729 -255 1095
rect -321 717 -255 729
rect -225 1095 -159 1107
rect -225 729 -209 1095
rect -175 729 -159 1095
rect -225 717 -159 729
rect -129 1095 -63 1107
rect -129 729 -113 1095
rect -79 729 -63 1095
rect -129 717 -63 729
rect -33 1095 33 1107
rect -33 729 -17 1095
rect 17 729 33 1095
rect -33 717 33 729
rect 63 1095 129 1107
rect 63 729 79 1095
rect 113 729 129 1095
rect 63 717 129 729
rect 159 1095 225 1107
rect 159 729 175 1095
rect 209 729 225 1095
rect 159 717 225 729
rect 255 1095 321 1107
rect 255 729 271 1095
rect 305 729 321 1095
rect 255 717 321 729
rect 351 1095 417 1107
rect 351 729 367 1095
rect 401 729 417 1095
rect 351 717 417 729
rect 447 1095 513 1107
rect 447 729 463 1095
rect 497 729 513 1095
rect 447 717 513 729
rect 543 1095 609 1107
rect 543 729 559 1095
rect 593 729 609 1095
rect 543 717 609 729
rect 639 1095 705 1107
rect 639 729 655 1095
rect 689 729 705 1095
rect 639 717 705 729
rect 735 1095 801 1107
rect 735 729 751 1095
rect 785 729 801 1095
rect 735 717 801 729
rect 831 1095 897 1107
rect 831 729 847 1095
rect 881 729 897 1095
rect 831 717 897 729
rect 927 1095 993 1107
rect 927 729 943 1095
rect 977 729 993 1095
rect 927 717 993 729
rect 1023 1095 1089 1107
rect 1023 729 1039 1095
rect 1073 729 1089 1095
rect 1023 717 1089 729
rect 1119 1095 1185 1107
rect 1119 729 1135 1095
rect 1169 729 1185 1095
rect 1119 717 1185 729
rect 1215 1095 1281 1107
rect 1215 729 1231 1095
rect 1265 729 1281 1095
rect 1215 717 1281 729
rect 1311 1095 1377 1107
rect 1311 729 1327 1095
rect 1361 729 1377 1095
rect 1311 717 1377 729
rect 1407 1095 1473 1107
rect 1407 729 1423 1095
rect 1457 729 1473 1095
rect 1407 717 1473 729
rect 1503 1095 1569 1107
rect 1503 729 1519 1095
rect 1553 729 1569 1095
rect 1503 717 1569 729
rect 1599 1095 1665 1107
rect 1599 729 1615 1095
rect 1649 729 1665 1095
rect 1599 717 1665 729
rect 1695 1095 1761 1107
rect 1695 729 1711 1095
rect 1745 729 1761 1095
rect 1695 717 1761 729
rect 1791 1095 1857 1107
rect 1791 729 1807 1095
rect 1841 729 1857 1095
rect 1791 717 1857 729
rect 1887 1095 1949 1107
rect 1887 729 1903 1095
rect 1937 729 1949 1095
rect 1887 717 1949 729
rect -1949 487 -1887 499
rect -1949 121 -1937 487
rect -1903 121 -1887 487
rect -1949 109 -1887 121
rect -1857 487 -1791 499
rect -1857 121 -1841 487
rect -1807 121 -1791 487
rect -1857 109 -1791 121
rect -1761 487 -1695 499
rect -1761 121 -1745 487
rect -1711 121 -1695 487
rect -1761 109 -1695 121
rect -1665 487 -1599 499
rect -1665 121 -1649 487
rect -1615 121 -1599 487
rect -1665 109 -1599 121
rect -1569 487 -1503 499
rect -1569 121 -1553 487
rect -1519 121 -1503 487
rect -1569 109 -1503 121
rect -1473 487 -1407 499
rect -1473 121 -1457 487
rect -1423 121 -1407 487
rect -1473 109 -1407 121
rect -1377 487 -1311 499
rect -1377 121 -1361 487
rect -1327 121 -1311 487
rect -1377 109 -1311 121
rect -1281 487 -1215 499
rect -1281 121 -1265 487
rect -1231 121 -1215 487
rect -1281 109 -1215 121
rect -1185 487 -1119 499
rect -1185 121 -1169 487
rect -1135 121 -1119 487
rect -1185 109 -1119 121
rect -1089 487 -1023 499
rect -1089 121 -1073 487
rect -1039 121 -1023 487
rect -1089 109 -1023 121
rect -993 487 -927 499
rect -993 121 -977 487
rect -943 121 -927 487
rect -993 109 -927 121
rect -897 487 -831 499
rect -897 121 -881 487
rect -847 121 -831 487
rect -897 109 -831 121
rect -801 487 -735 499
rect -801 121 -785 487
rect -751 121 -735 487
rect -801 109 -735 121
rect -705 487 -639 499
rect -705 121 -689 487
rect -655 121 -639 487
rect -705 109 -639 121
rect -609 487 -543 499
rect -609 121 -593 487
rect -559 121 -543 487
rect -609 109 -543 121
rect -513 487 -447 499
rect -513 121 -497 487
rect -463 121 -447 487
rect -513 109 -447 121
rect -417 487 -351 499
rect -417 121 -401 487
rect -367 121 -351 487
rect -417 109 -351 121
rect -321 487 -255 499
rect -321 121 -305 487
rect -271 121 -255 487
rect -321 109 -255 121
rect -225 487 -159 499
rect -225 121 -209 487
rect -175 121 -159 487
rect -225 109 -159 121
rect -129 487 -63 499
rect -129 121 -113 487
rect -79 121 -63 487
rect -129 109 -63 121
rect -33 487 33 499
rect -33 121 -17 487
rect 17 121 33 487
rect -33 109 33 121
rect 63 487 129 499
rect 63 121 79 487
rect 113 121 129 487
rect 63 109 129 121
rect 159 487 225 499
rect 159 121 175 487
rect 209 121 225 487
rect 159 109 225 121
rect 255 487 321 499
rect 255 121 271 487
rect 305 121 321 487
rect 255 109 321 121
rect 351 487 417 499
rect 351 121 367 487
rect 401 121 417 487
rect 351 109 417 121
rect 447 487 513 499
rect 447 121 463 487
rect 497 121 513 487
rect 447 109 513 121
rect 543 487 609 499
rect 543 121 559 487
rect 593 121 609 487
rect 543 109 609 121
rect 639 487 705 499
rect 639 121 655 487
rect 689 121 705 487
rect 639 109 705 121
rect 735 487 801 499
rect 735 121 751 487
rect 785 121 801 487
rect 735 109 801 121
rect 831 487 897 499
rect 831 121 847 487
rect 881 121 897 487
rect 831 109 897 121
rect 927 487 993 499
rect 927 121 943 487
rect 977 121 993 487
rect 927 109 993 121
rect 1023 487 1089 499
rect 1023 121 1039 487
rect 1073 121 1089 487
rect 1023 109 1089 121
rect 1119 487 1185 499
rect 1119 121 1135 487
rect 1169 121 1185 487
rect 1119 109 1185 121
rect 1215 487 1281 499
rect 1215 121 1231 487
rect 1265 121 1281 487
rect 1215 109 1281 121
rect 1311 487 1377 499
rect 1311 121 1327 487
rect 1361 121 1377 487
rect 1311 109 1377 121
rect 1407 487 1473 499
rect 1407 121 1423 487
rect 1457 121 1473 487
rect 1407 109 1473 121
rect 1503 487 1569 499
rect 1503 121 1519 487
rect 1553 121 1569 487
rect 1503 109 1569 121
rect 1599 487 1665 499
rect 1599 121 1615 487
rect 1649 121 1665 487
rect 1599 109 1665 121
rect 1695 487 1761 499
rect 1695 121 1711 487
rect 1745 121 1761 487
rect 1695 109 1761 121
rect 1791 487 1857 499
rect 1791 121 1807 487
rect 1841 121 1857 487
rect 1791 109 1857 121
rect 1887 487 1949 499
rect 1887 121 1903 487
rect 1937 121 1949 487
rect 1887 109 1949 121
rect -1949 -121 -1887 -109
rect -1949 -487 -1937 -121
rect -1903 -487 -1887 -121
rect -1949 -499 -1887 -487
rect -1857 -121 -1791 -109
rect -1857 -487 -1841 -121
rect -1807 -487 -1791 -121
rect -1857 -499 -1791 -487
rect -1761 -121 -1695 -109
rect -1761 -487 -1745 -121
rect -1711 -487 -1695 -121
rect -1761 -499 -1695 -487
rect -1665 -121 -1599 -109
rect -1665 -487 -1649 -121
rect -1615 -487 -1599 -121
rect -1665 -499 -1599 -487
rect -1569 -121 -1503 -109
rect -1569 -487 -1553 -121
rect -1519 -487 -1503 -121
rect -1569 -499 -1503 -487
rect -1473 -121 -1407 -109
rect -1473 -487 -1457 -121
rect -1423 -487 -1407 -121
rect -1473 -499 -1407 -487
rect -1377 -121 -1311 -109
rect -1377 -487 -1361 -121
rect -1327 -487 -1311 -121
rect -1377 -499 -1311 -487
rect -1281 -121 -1215 -109
rect -1281 -487 -1265 -121
rect -1231 -487 -1215 -121
rect -1281 -499 -1215 -487
rect -1185 -121 -1119 -109
rect -1185 -487 -1169 -121
rect -1135 -487 -1119 -121
rect -1185 -499 -1119 -487
rect -1089 -121 -1023 -109
rect -1089 -487 -1073 -121
rect -1039 -487 -1023 -121
rect -1089 -499 -1023 -487
rect -993 -121 -927 -109
rect -993 -487 -977 -121
rect -943 -487 -927 -121
rect -993 -499 -927 -487
rect -897 -121 -831 -109
rect -897 -487 -881 -121
rect -847 -487 -831 -121
rect -897 -499 -831 -487
rect -801 -121 -735 -109
rect -801 -487 -785 -121
rect -751 -487 -735 -121
rect -801 -499 -735 -487
rect -705 -121 -639 -109
rect -705 -487 -689 -121
rect -655 -487 -639 -121
rect -705 -499 -639 -487
rect -609 -121 -543 -109
rect -609 -487 -593 -121
rect -559 -487 -543 -121
rect -609 -499 -543 -487
rect -513 -121 -447 -109
rect -513 -487 -497 -121
rect -463 -487 -447 -121
rect -513 -499 -447 -487
rect -417 -121 -351 -109
rect -417 -487 -401 -121
rect -367 -487 -351 -121
rect -417 -499 -351 -487
rect -321 -121 -255 -109
rect -321 -487 -305 -121
rect -271 -487 -255 -121
rect -321 -499 -255 -487
rect -225 -121 -159 -109
rect -225 -487 -209 -121
rect -175 -487 -159 -121
rect -225 -499 -159 -487
rect -129 -121 -63 -109
rect -129 -487 -113 -121
rect -79 -487 -63 -121
rect -129 -499 -63 -487
rect -33 -121 33 -109
rect -33 -487 -17 -121
rect 17 -487 33 -121
rect -33 -499 33 -487
rect 63 -121 129 -109
rect 63 -487 79 -121
rect 113 -487 129 -121
rect 63 -499 129 -487
rect 159 -121 225 -109
rect 159 -487 175 -121
rect 209 -487 225 -121
rect 159 -499 225 -487
rect 255 -121 321 -109
rect 255 -487 271 -121
rect 305 -487 321 -121
rect 255 -499 321 -487
rect 351 -121 417 -109
rect 351 -487 367 -121
rect 401 -487 417 -121
rect 351 -499 417 -487
rect 447 -121 513 -109
rect 447 -487 463 -121
rect 497 -487 513 -121
rect 447 -499 513 -487
rect 543 -121 609 -109
rect 543 -487 559 -121
rect 593 -487 609 -121
rect 543 -499 609 -487
rect 639 -121 705 -109
rect 639 -487 655 -121
rect 689 -487 705 -121
rect 639 -499 705 -487
rect 735 -121 801 -109
rect 735 -487 751 -121
rect 785 -487 801 -121
rect 735 -499 801 -487
rect 831 -121 897 -109
rect 831 -487 847 -121
rect 881 -487 897 -121
rect 831 -499 897 -487
rect 927 -121 993 -109
rect 927 -487 943 -121
rect 977 -487 993 -121
rect 927 -499 993 -487
rect 1023 -121 1089 -109
rect 1023 -487 1039 -121
rect 1073 -487 1089 -121
rect 1023 -499 1089 -487
rect 1119 -121 1185 -109
rect 1119 -487 1135 -121
rect 1169 -487 1185 -121
rect 1119 -499 1185 -487
rect 1215 -121 1281 -109
rect 1215 -487 1231 -121
rect 1265 -487 1281 -121
rect 1215 -499 1281 -487
rect 1311 -121 1377 -109
rect 1311 -487 1327 -121
rect 1361 -487 1377 -121
rect 1311 -499 1377 -487
rect 1407 -121 1473 -109
rect 1407 -487 1423 -121
rect 1457 -487 1473 -121
rect 1407 -499 1473 -487
rect 1503 -121 1569 -109
rect 1503 -487 1519 -121
rect 1553 -487 1569 -121
rect 1503 -499 1569 -487
rect 1599 -121 1665 -109
rect 1599 -487 1615 -121
rect 1649 -487 1665 -121
rect 1599 -499 1665 -487
rect 1695 -121 1761 -109
rect 1695 -487 1711 -121
rect 1745 -487 1761 -121
rect 1695 -499 1761 -487
rect 1791 -121 1857 -109
rect 1791 -487 1807 -121
rect 1841 -487 1857 -121
rect 1791 -499 1857 -487
rect 1887 -121 1949 -109
rect 1887 -487 1903 -121
rect 1937 -487 1949 -121
rect 1887 -499 1949 -487
rect -1949 -729 -1887 -717
rect -1949 -1095 -1937 -729
rect -1903 -1095 -1887 -729
rect -1949 -1107 -1887 -1095
rect -1857 -729 -1791 -717
rect -1857 -1095 -1841 -729
rect -1807 -1095 -1791 -729
rect -1857 -1107 -1791 -1095
rect -1761 -729 -1695 -717
rect -1761 -1095 -1745 -729
rect -1711 -1095 -1695 -729
rect -1761 -1107 -1695 -1095
rect -1665 -729 -1599 -717
rect -1665 -1095 -1649 -729
rect -1615 -1095 -1599 -729
rect -1665 -1107 -1599 -1095
rect -1569 -729 -1503 -717
rect -1569 -1095 -1553 -729
rect -1519 -1095 -1503 -729
rect -1569 -1107 -1503 -1095
rect -1473 -729 -1407 -717
rect -1473 -1095 -1457 -729
rect -1423 -1095 -1407 -729
rect -1473 -1107 -1407 -1095
rect -1377 -729 -1311 -717
rect -1377 -1095 -1361 -729
rect -1327 -1095 -1311 -729
rect -1377 -1107 -1311 -1095
rect -1281 -729 -1215 -717
rect -1281 -1095 -1265 -729
rect -1231 -1095 -1215 -729
rect -1281 -1107 -1215 -1095
rect -1185 -729 -1119 -717
rect -1185 -1095 -1169 -729
rect -1135 -1095 -1119 -729
rect -1185 -1107 -1119 -1095
rect -1089 -729 -1023 -717
rect -1089 -1095 -1073 -729
rect -1039 -1095 -1023 -729
rect -1089 -1107 -1023 -1095
rect -993 -729 -927 -717
rect -993 -1095 -977 -729
rect -943 -1095 -927 -729
rect -993 -1107 -927 -1095
rect -897 -729 -831 -717
rect -897 -1095 -881 -729
rect -847 -1095 -831 -729
rect -897 -1107 -831 -1095
rect -801 -729 -735 -717
rect -801 -1095 -785 -729
rect -751 -1095 -735 -729
rect -801 -1107 -735 -1095
rect -705 -729 -639 -717
rect -705 -1095 -689 -729
rect -655 -1095 -639 -729
rect -705 -1107 -639 -1095
rect -609 -729 -543 -717
rect -609 -1095 -593 -729
rect -559 -1095 -543 -729
rect -609 -1107 -543 -1095
rect -513 -729 -447 -717
rect -513 -1095 -497 -729
rect -463 -1095 -447 -729
rect -513 -1107 -447 -1095
rect -417 -729 -351 -717
rect -417 -1095 -401 -729
rect -367 -1095 -351 -729
rect -417 -1107 -351 -1095
rect -321 -729 -255 -717
rect -321 -1095 -305 -729
rect -271 -1095 -255 -729
rect -321 -1107 -255 -1095
rect -225 -729 -159 -717
rect -225 -1095 -209 -729
rect -175 -1095 -159 -729
rect -225 -1107 -159 -1095
rect -129 -729 -63 -717
rect -129 -1095 -113 -729
rect -79 -1095 -63 -729
rect -129 -1107 -63 -1095
rect -33 -729 33 -717
rect -33 -1095 -17 -729
rect 17 -1095 33 -729
rect -33 -1107 33 -1095
rect 63 -729 129 -717
rect 63 -1095 79 -729
rect 113 -1095 129 -729
rect 63 -1107 129 -1095
rect 159 -729 225 -717
rect 159 -1095 175 -729
rect 209 -1095 225 -729
rect 159 -1107 225 -1095
rect 255 -729 321 -717
rect 255 -1095 271 -729
rect 305 -1095 321 -729
rect 255 -1107 321 -1095
rect 351 -729 417 -717
rect 351 -1095 367 -729
rect 401 -1095 417 -729
rect 351 -1107 417 -1095
rect 447 -729 513 -717
rect 447 -1095 463 -729
rect 497 -1095 513 -729
rect 447 -1107 513 -1095
rect 543 -729 609 -717
rect 543 -1095 559 -729
rect 593 -1095 609 -729
rect 543 -1107 609 -1095
rect 639 -729 705 -717
rect 639 -1095 655 -729
rect 689 -1095 705 -729
rect 639 -1107 705 -1095
rect 735 -729 801 -717
rect 735 -1095 751 -729
rect 785 -1095 801 -729
rect 735 -1107 801 -1095
rect 831 -729 897 -717
rect 831 -1095 847 -729
rect 881 -1095 897 -729
rect 831 -1107 897 -1095
rect 927 -729 993 -717
rect 927 -1095 943 -729
rect 977 -1095 993 -729
rect 927 -1107 993 -1095
rect 1023 -729 1089 -717
rect 1023 -1095 1039 -729
rect 1073 -1095 1089 -729
rect 1023 -1107 1089 -1095
rect 1119 -729 1185 -717
rect 1119 -1095 1135 -729
rect 1169 -1095 1185 -729
rect 1119 -1107 1185 -1095
rect 1215 -729 1281 -717
rect 1215 -1095 1231 -729
rect 1265 -1095 1281 -729
rect 1215 -1107 1281 -1095
rect 1311 -729 1377 -717
rect 1311 -1095 1327 -729
rect 1361 -1095 1377 -729
rect 1311 -1107 1377 -1095
rect 1407 -729 1473 -717
rect 1407 -1095 1423 -729
rect 1457 -1095 1473 -729
rect 1407 -1107 1473 -1095
rect 1503 -729 1569 -717
rect 1503 -1095 1519 -729
rect 1553 -1095 1569 -729
rect 1503 -1107 1569 -1095
rect 1599 -729 1665 -717
rect 1599 -1095 1615 -729
rect 1649 -1095 1665 -729
rect 1599 -1107 1665 -1095
rect 1695 -729 1761 -717
rect 1695 -1095 1711 -729
rect 1745 -1095 1761 -729
rect 1695 -1107 1761 -1095
rect 1791 -729 1857 -717
rect 1791 -1095 1807 -729
rect 1841 -1095 1857 -729
rect 1791 -1107 1857 -1095
rect 1887 -729 1949 -717
rect 1887 -1095 1903 -729
rect 1937 -1095 1949 -729
rect 1887 -1107 1949 -1095
rect -1949 -1337 -1887 -1325
rect -1949 -1703 -1937 -1337
rect -1903 -1703 -1887 -1337
rect -1949 -1715 -1887 -1703
rect -1857 -1337 -1791 -1325
rect -1857 -1703 -1841 -1337
rect -1807 -1703 -1791 -1337
rect -1857 -1715 -1791 -1703
rect -1761 -1337 -1695 -1325
rect -1761 -1703 -1745 -1337
rect -1711 -1703 -1695 -1337
rect -1761 -1715 -1695 -1703
rect -1665 -1337 -1599 -1325
rect -1665 -1703 -1649 -1337
rect -1615 -1703 -1599 -1337
rect -1665 -1715 -1599 -1703
rect -1569 -1337 -1503 -1325
rect -1569 -1703 -1553 -1337
rect -1519 -1703 -1503 -1337
rect -1569 -1715 -1503 -1703
rect -1473 -1337 -1407 -1325
rect -1473 -1703 -1457 -1337
rect -1423 -1703 -1407 -1337
rect -1473 -1715 -1407 -1703
rect -1377 -1337 -1311 -1325
rect -1377 -1703 -1361 -1337
rect -1327 -1703 -1311 -1337
rect -1377 -1715 -1311 -1703
rect -1281 -1337 -1215 -1325
rect -1281 -1703 -1265 -1337
rect -1231 -1703 -1215 -1337
rect -1281 -1715 -1215 -1703
rect -1185 -1337 -1119 -1325
rect -1185 -1703 -1169 -1337
rect -1135 -1703 -1119 -1337
rect -1185 -1715 -1119 -1703
rect -1089 -1337 -1023 -1325
rect -1089 -1703 -1073 -1337
rect -1039 -1703 -1023 -1337
rect -1089 -1715 -1023 -1703
rect -993 -1337 -927 -1325
rect -993 -1703 -977 -1337
rect -943 -1703 -927 -1337
rect -993 -1715 -927 -1703
rect -897 -1337 -831 -1325
rect -897 -1703 -881 -1337
rect -847 -1703 -831 -1337
rect -897 -1715 -831 -1703
rect -801 -1337 -735 -1325
rect -801 -1703 -785 -1337
rect -751 -1703 -735 -1337
rect -801 -1715 -735 -1703
rect -705 -1337 -639 -1325
rect -705 -1703 -689 -1337
rect -655 -1703 -639 -1337
rect -705 -1715 -639 -1703
rect -609 -1337 -543 -1325
rect -609 -1703 -593 -1337
rect -559 -1703 -543 -1337
rect -609 -1715 -543 -1703
rect -513 -1337 -447 -1325
rect -513 -1703 -497 -1337
rect -463 -1703 -447 -1337
rect -513 -1715 -447 -1703
rect -417 -1337 -351 -1325
rect -417 -1703 -401 -1337
rect -367 -1703 -351 -1337
rect -417 -1715 -351 -1703
rect -321 -1337 -255 -1325
rect -321 -1703 -305 -1337
rect -271 -1703 -255 -1337
rect -321 -1715 -255 -1703
rect -225 -1337 -159 -1325
rect -225 -1703 -209 -1337
rect -175 -1703 -159 -1337
rect -225 -1715 -159 -1703
rect -129 -1337 -63 -1325
rect -129 -1703 -113 -1337
rect -79 -1703 -63 -1337
rect -129 -1715 -63 -1703
rect -33 -1337 33 -1325
rect -33 -1703 -17 -1337
rect 17 -1703 33 -1337
rect -33 -1715 33 -1703
rect 63 -1337 129 -1325
rect 63 -1703 79 -1337
rect 113 -1703 129 -1337
rect 63 -1715 129 -1703
rect 159 -1337 225 -1325
rect 159 -1703 175 -1337
rect 209 -1703 225 -1337
rect 159 -1715 225 -1703
rect 255 -1337 321 -1325
rect 255 -1703 271 -1337
rect 305 -1703 321 -1337
rect 255 -1715 321 -1703
rect 351 -1337 417 -1325
rect 351 -1703 367 -1337
rect 401 -1703 417 -1337
rect 351 -1715 417 -1703
rect 447 -1337 513 -1325
rect 447 -1703 463 -1337
rect 497 -1703 513 -1337
rect 447 -1715 513 -1703
rect 543 -1337 609 -1325
rect 543 -1703 559 -1337
rect 593 -1703 609 -1337
rect 543 -1715 609 -1703
rect 639 -1337 705 -1325
rect 639 -1703 655 -1337
rect 689 -1703 705 -1337
rect 639 -1715 705 -1703
rect 735 -1337 801 -1325
rect 735 -1703 751 -1337
rect 785 -1703 801 -1337
rect 735 -1715 801 -1703
rect 831 -1337 897 -1325
rect 831 -1703 847 -1337
rect 881 -1703 897 -1337
rect 831 -1715 897 -1703
rect 927 -1337 993 -1325
rect 927 -1703 943 -1337
rect 977 -1703 993 -1337
rect 927 -1715 993 -1703
rect 1023 -1337 1089 -1325
rect 1023 -1703 1039 -1337
rect 1073 -1703 1089 -1337
rect 1023 -1715 1089 -1703
rect 1119 -1337 1185 -1325
rect 1119 -1703 1135 -1337
rect 1169 -1703 1185 -1337
rect 1119 -1715 1185 -1703
rect 1215 -1337 1281 -1325
rect 1215 -1703 1231 -1337
rect 1265 -1703 1281 -1337
rect 1215 -1715 1281 -1703
rect 1311 -1337 1377 -1325
rect 1311 -1703 1327 -1337
rect 1361 -1703 1377 -1337
rect 1311 -1715 1377 -1703
rect 1407 -1337 1473 -1325
rect 1407 -1703 1423 -1337
rect 1457 -1703 1473 -1337
rect 1407 -1715 1473 -1703
rect 1503 -1337 1569 -1325
rect 1503 -1703 1519 -1337
rect 1553 -1703 1569 -1337
rect 1503 -1715 1569 -1703
rect 1599 -1337 1665 -1325
rect 1599 -1703 1615 -1337
rect 1649 -1703 1665 -1337
rect 1599 -1715 1665 -1703
rect 1695 -1337 1761 -1325
rect 1695 -1703 1711 -1337
rect 1745 -1703 1761 -1337
rect 1695 -1715 1761 -1703
rect 1791 -1337 1857 -1325
rect 1791 -1703 1807 -1337
rect 1841 -1703 1857 -1337
rect 1791 -1715 1857 -1703
rect 1887 -1337 1949 -1325
rect 1887 -1703 1903 -1337
rect 1937 -1703 1949 -1337
rect 1887 -1715 1949 -1703
<< ndiffc >>
rect -1937 1337 -1903 1703
rect -1841 1337 -1807 1703
rect -1745 1337 -1711 1703
rect -1649 1337 -1615 1703
rect -1553 1337 -1519 1703
rect -1457 1337 -1423 1703
rect -1361 1337 -1327 1703
rect -1265 1337 -1231 1703
rect -1169 1337 -1135 1703
rect -1073 1337 -1039 1703
rect -977 1337 -943 1703
rect -881 1337 -847 1703
rect -785 1337 -751 1703
rect -689 1337 -655 1703
rect -593 1337 -559 1703
rect -497 1337 -463 1703
rect -401 1337 -367 1703
rect -305 1337 -271 1703
rect -209 1337 -175 1703
rect -113 1337 -79 1703
rect -17 1337 17 1703
rect 79 1337 113 1703
rect 175 1337 209 1703
rect 271 1337 305 1703
rect 367 1337 401 1703
rect 463 1337 497 1703
rect 559 1337 593 1703
rect 655 1337 689 1703
rect 751 1337 785 1703
rect 847 1337 881 1703
rect 943 1337 977 1703
rect 1039 1337 1073 1703
rect 1135 1337 1169 1703
rect 1231 1337 1265 1703
rect 1327 1337 1361 1703
rect 1423 1337 1457 1703
rect 1519 1337 1553 1703
rect 1615 1337 1649 1703
rect 1711 1337 1745 1703
rect 1807 1337 1841 1703
rect 1903 1337 1937 1703
rect -1937 729 -1903 1095
rect -1841 729 -1807 1095
rect -1745 729 -1711 1095
rect -1649 729 -1615 1095
rect -1553 729 -1519 1095
rect -1457 729 -1423 1095
rect -1361 729 -1327 1095
rect -1265 729 -1231 1095
rect -1169 729 -1135 1095
rect -1073 729 -1039 1095
rect -977 729 -943 1095
rect -881 729 -847 1095
rect -785 729 -751 1095
rect -689 729 -655 1095
rect -593 729 -559 1095
rect -497 729 -463 1095
rect -401 729 -367 1095
rect -305 729 -271 1095
rect -209 729 -175 1095
rect -113 729 -79 1095
rect -17 729 17 1095
rect 79 729 113 1095
rect 175 729 209 1095
rect 271 729 305 1095
rect 367 729 401 1095
rect 463 729 497 1095
rect 559 729 593 1095
rect 655 729 689 1095
rect 751 729 785 1095
rect 847 729 881 1095
rect 943 729 977 1095
rect 1039 729 1073 1095
rect 1135 729 1169 1095
rect 1231 729 1265 1095
rect 1327 729 1361 1095
rect 1423 729 1457 1095
rect 1519 729 1553 1095
rect 1615 729 1649 1095
rect 1711 729 1745 1095
rect 1807 729 1841 1095
rect 1903 729 1937 1095
rect -1937 121 -1903 487
rect -1841 121 -1807 487
rect -1745 121 -1711 487
rect -1649 121 -1615 487
rect -1553 121 -1519 487
rect -1457 121 -1423 487
rect -1361 121 -1327 487
rect -1265 121 -1231 487
rect -1169 121 -1135 487
rect -1073 121 -1039 487
rect -977 121 -943 487
rect -881 121 -847 487
rect -785 121 -751 487
rect -689 121 -655 487
rect -593 121 -559 487
rect -497 121 -463 487
rect -401 121 -367 487
rect -305 121 -271 487
rect -209 121 -175 487
rect -113 121 -79 487
rect -17 121 17 487
rect 79 121 113 487
rect 175 121 209 487
rect 271 121 305 487
rect 367 121 401 487
rect 463 121 497 487
rect 559 121 593 487
rect 655 121 689 487
rect 751 121 785 487
rect 847 121 881 487
rect 943 121 977 487
rect 1039 121 1073 487
rect 1135 121 1169 487
rect 1231 121 1265 487
rect 1327 121 1361 487
rect 1423 121 1457 487
rect 1519 121 1553 487
rect 1615 121 1649 487
rect 1711 121 1745 487
rect 1807 121 1841 487
rect 1903 121 1937 487
rect -1937 -487 -1903 -121
rect -1841 -487 -1807 -121
rect -1745 -487 -1711 -121
rect -1649 -487 -1615 -121
rect -1553 -487 -1519 -121
rect -1457 -487 -1423 -121
rect -1361 -487 -1327 -121
rect -1265 -487 -1231 -121
rect -1169 -487 -1135 -121
rect -1073 -487 -1039 -121
rect -977 -487 -943 -121
rect -881 -487 -847 -121
rect -785 -487 -751 -121
rect -689 -487 -655 -121
rect -593 -487 -559 -121
rect -497 -487 -463 -121
rect -401 -487 -367 -121
rect -305 -487 -271 -121
rect -209 -487 -175 -121
rect -113 -487 -79 -121
rect -17 -487 17 -121
rect 79 -487 113 -121
rect 175 -487 209 -121
rect 271 -487 305 -121
rect 367 -487 401 -121
rect 463 -487 497 -121
rect 559 -487 593 -121
rect 655 -487 689 -121
rect 751 -487 785 -121
rect 847 -487 881 -121
rect 943 -487 977 -121
rect 1039 -487 1073 -121
rect 1135 -487 1169 -121
rect 1231 -487 1265 -121
rect 1327 -487 1361 -121
rect 1423 -487 1457 -121
rect 1519 -487 1553 -121
rect 1615 -487 1649 -121
rect 1711 -487 1745 -121
rect 1807 -487 1841 -121
rect 1903 -487 1937 -121
rect -1937 -1095 -1903 -729
rect -1841 -1095 -1807 -729
rect -1745 -1095 -1711 -729
rect -1649 -1095 -1615 -729
rect -1553 -1095 -1519 -729
rect -1457 -1095 -1423 -729
rect -1361 -1095 -1327 -729
rect -1265 -1095 -1231 -729
rect -1169 -1095 -1135 -729
rect -1073 -1095 -1039 -729
rect -977 -1095 -943 -729
rect -881 -1095 -847 -729
rect -785 -1095 -751 -729
rect -689 -1095 -655 -729
rect -593 -1095 -559 -729
rect -497 -1095 -463 -729
rect -401 -1095 -367 -729
rect -305 -1095 -271 -729
rect -209 -1095 -175 -729
rect -113 -1095 -79 -729
rect -17 -1095 17 -729
rect 79 -1095 113 -729
rect 175 -1095 209 -729
rect 271 -1095 305 -729
rect 367 -1095 401 -729
rect 463 -1095 497 -729
rect 559 -1095 593 -729
rect 655 -1095 689 -729
rect 751 -1095 785 -729
rect 847 -1095 881 -729
rect 943 -1095 977 -729
rect 1039 -1095 1073 -729
rect 1135 -1095 1169 -729
rect 1231 -1095 1265 -729
rect 1327 -1095 1361 -729
rect 1423 -1095 1457 -729
rect 1519 -1095 1553 -729
rect 1615 -1095 1649 -729
rect 1711 -1095 1745 -729
rect 1807 -1095 1841 -729
rect 1903 -1095 1937 -729
rect -1937 -1703 -1903 -1337
rect -1841 -1703 -1807 -1337
rect -1745 -1703 -1711 -1337
rect -1649 -1703 -1615 -1337
rect -1553 -1703 -1519 -1337
rect -1457 -1703 -1423 -1337
rect -1361 -1703 -1327 -1337
rect -1265 -1703 -1231 -1337
rect -1169 -1703 -1135 -1337
rect -1073 -1703 -1039 -1337
rect -977 -1703 -943 -1337
rect -881 -1703 -847 -1337
rect -785 -1703 -751 -1337
rect -689 -1703 -655 -1337
rect -593 -1703 -559 -1337
rect -497 -1703 -463 -1337
rect -401 -1703 -367 -1337
rect -305 -1703 -271 -1337
rect -209 -1703 -175 -1337
rect -113 -1703 -79 -1337
rect -17 -1703 17 -1337
rect 79 -1703 113 -1337
rect 175 -1703 209 -1337
rect 271 -1703 305 -1337
rect 367 -1703 401 -1337
rect 463 -1703 497 -1337
rect 559 -1703 593 -1337
rect 655 -1703 689 -1337
rect 751 -1703 785 -1337
rect 847 -1703 881 -1337
rect 943 -1703 977 -1337
rect 1039 -1703 1073 -1337
rect 1135 -1703 1169 -1337
rect 1231 -1703 1265 -1337
rect 1327 -1703 1361 -1337
rect 1423 -1703 1457 -1337
rect 1519 -1703 1553 -1337
rect 1615 -1703 1649 -1337
rect 1711 -1703 1745 -1337
rect 1807 -1703 1841 -1337
rect 1903 -1703 1937 -1337
<< psubdiff >>
rect -2051 1855 -1955 1889
rect 1955 1855 2051 1889
rect -2051 1793 -2017 1855
rect 2017 1793 2051 1855
rect -2051 -1855 -2017 -1793
rect 2017 -1855 2051 -1793
rect -2051 -1889 -1955 -1855
rect 1955 -1889 2051 -1855
<< psubdiffcont >>
rect -1955 1855 1955 1889
rect -2051 -1793 -2017 1793
rect 2017 -1793 2051 1793
rect -1955 -1889 1955 -1855
<< poly >>
rect -1905 1787 -1839 1803
rect -1905 1753 -1889 1787
rect -1855 1753 -1839 1787
rect -1905 1737 -1839 1753
rect -1713 1787 -1647 1803
rect -1713 1753 -1697 1787
rect -1663 1753 -1647 1787
rect -1887 1715 -1857 1737
rect -1791 1715 -1761 1741
rect -1713 1737 -1647 1753
rect -1521 1787 -1455 1803
rect -1521 1753 -1505 1787
rect -1471 1753 -1455 1787
rect -1695 1715 -1665 1737
rect -1599 1715 -1569 1741
rect -1521 1737 -1455 1753
rect -1329 1787 -1263 1803
rect -1329 1753 -1313 1787
rect -1279 1753 -1263 1787
rect -1503 1715 -1473 1737
rect -1407 1715 -1377 1741
rect -1329 1737 -1263 1753
rect -1137 1787 -1071 1803
rect -1137 1753 -1121 1787
rect -1087 1753 -1071 1787
rect -1311 1715 -1281 1737
rect -1215 1715 -1185 1741
rect -1137 1737 -1071 1753
rect -945 1787 -879 1803
rect -945 1753 -929 1787
rect -895 1753 -879 1787
rect -1119 1715 -1089 1737
rect -1023 1715 -993 1741
rect -945 1737 -879 1753
rect -753 1787 -687 1803
rect -753 1753 -737 1787
rect -703 1753 -687 1787
rect -927 1715 -897 1737
rect -831 1715 -801 1741
rect -753 1737 -687 1753
rect -561 1787 -495 1803
rect -561 1753 -545 1787
rect -511 1753 -495 1787
rect -735 1715 -705 1737
rect -639 1715 -609 1741
rect -561 1737 -495 1753
rect -369 1787 -303 1803
rect -369 1753 -353 1787
rect -319 1753 -303 1787
rect -543 1715 -513 1737
rect -447 1715 -417 1741
rect -369 1737 -303 1753
rect -177 1787 -111 1803
rect -177 1753 -161 1787
rect -127 1753 -111 1787
rect -351 1715 -321 1737
rect -255 1715 -225 1741
rect -177 1737 -111 1753
rect 15 1787 81 1803
rect 15 1753 31 1787
rect 65 1753 81 1787
rect -159 1715 -129 1737
rect -63 1715 -33 1741
rect 15 1737 81 1753
rect 207 1787 273 1803
rect 207 1753 223 1787
rect 257 1753 273 1787
rect 33 1715 63 1737
rect 129 1715 159 1741
rect 207 1737 273 1753
rect 399 1787 465 1803
rect 399 1753 415 1787
rect 449 1753 465 1787
rect 225 1715 255 1737
rect 321 1715 351 1741
rect 399 1737 465 1753
rect 591 1787 657 1803
rect 591 1753 607 1787
rect 641 1753 657 1787
rect 417 1715 447 1737
rect 513 1715 543 1741
rect 591 1737 657 1753
rect 783 1787 849 1803
rect 783 1753 799 1787
rect 833 1753 849 1787
rect 609 1715 639 1737
rect 705 1715 735 1741
rect 783 1737 849 1753
rect 975 1787 1041 1803
rect 975 1753 991 1787
rect 1025 1753 1041 1787
rect 801 1715 831 1737
rect 897 1715 927 1741
rect 975 1737 1041 1753
rect 1167 1787 1233 1803
rect 1167 1753 1183 1787
rect 1217 1753 1233 1787
rect 993 1715 1023 1737
rect 1089 1715 1119 1741
rect 1167 1737 1233 1753
rect 1359 1787 1425 1803
rect 1359 1753 1375 1787
rect 1409 1753 1425 1787
rect 1185 1715 1215 1737
rect 1281 1715 1311 1741
rect 1359 1737 1425 1753
rect 1551 1787 1617 1803
rect 1551 1753 1567 1787
rect 1601 1753 1617 1787
rect 1377 1715 1407 1737
rect 1473 1715 1503 1741
rect 1551 1737 1617 1753
rect 1743 1787 1809 1803
rect 1743 1753 1759 1787
rect 1793 1753 1809 1787
rect 1569 1715 1599 1737
rect 1665 1715 1695 1741
rect 1743 1737 1809 1753
rect 1761 1715 1791 1737
rect 1857 1715 1887 1741
rect -1887 1299 -1857 1325
rect -1791 1303 -1761 1325
rect -1809 1287 -1743 1303
rect -1695 1299 -1665 1325
rect -1599 1303 -1569 1325
rect -1809 1253 -1793 1287
rect -1759 1253 -1743 1287
rect -1809 1237 -1743 1253
rect -1617 1287 -1551 1303
rect -1503 1299 -1473 1325
rect -1407 1303 -1377 1325
rect -1617 1253 -1601 1287
rect -1567 1253 -1551 1287
rect -1617 1237 -1551 1253
rect -1425 1287 -1359 1303
rect -1311 1299 -1281 1325
rect -1215 1303 -1185 1325
rect -1425 1253 -1409 1287
rect -1375 1253 -1359 1287
rect -1425 1237 -1359 1253
rect -1233 1287 -1167 1303
rect -1119 1299 -1089 1325
rect -1023 1303 -993 1325
rect -1233 1253 -1217 1287
rect -1183 1253 -1167 1287
rect -1233 1237 -1167 1253
rect -1041 1287 -975 1303
rect -927 1299 -897 1325
rect -831 1303 -801 1325
rect -1041 1253 -1025 1287
rect -991 1253 -975 1287
rect -1041 1237 -975 1253
rect -849 1287 -783 1303
rect -735 1299 -705 1325
rect -639 1303 -609 1325
rect -849 1253 -833 1287
rect -799 1253 -783 1287
rect -849 1237 -783 1253
rect -657 1287 -591 1303
rect -543 1299 -513 1325
rect -447 1303 -417 1325
rect -657 1253 -641 1287
rect -607 1253 -591 1287
rect -657 1237 -591 1253
rect -465 1287 -399 1303
rect -351 1299 -321 1325
rect -255 1303 -225 1325
rect -465 1253 -449 1287
rect -415 1253 -399 1287
rect -465 1237 -399 1253
rect -273 1287 -207 1303
rect -159 1299 -129 1325
rect -63 1303 -33 1325
rect -273 1253 -257 1287
rect -223 1253 -207 1287
rect -273 1237 -207 1253
rect -81 1287 -15 1303
rect 33 1299 63 1325
rect 129 1303 159 1325
rect -81 1253 -65 1287
rect -31 1253 -15 1287
rect -81 1237 -15 1253
rect 111 1287 177 1303
rect 225 1299 255 1325
rect 321 1303 351 1325
rect 111 1253 127 1287
rect 161 1253 177 1287
rect 111 1237 177 1253
rect 303 1287 369 1303
rect 417 1299 447 1325
rect 513 1303 543 1325
rect 303 1253 319 1287
rect 353 1253 369 1287
rect 303 1237 369 1253
rect 495 1287 561 1303
rect 609 1299 639 1325
rect 705 1303 735 1325
rect 495 1253 511 1287
rect 545 1253 561 1287
rect 495 1237 561 1253
rect 687 1287 753 1303
rect 801 1299 831 1325
rect 897 1303 927 1325
rect 687 1253 703 1287
rect 737 1253 753 1287
rect 687 1237 753 1253
rect 879 1287 945 1303
rect 993 1299 1023 1325
rect 1089 1303 1119 1325
rect 879 1253 895 1287
rect 929 1253 945 1287
rect 879 1237 945 1253
rect 1071 1287 1137 1303
rect 1185 1299 1215 1325
rect 1281 1303 1311 1325
rect 1071 1253 1087 1287
rect 1121 1253 1137 1287
rect 1071 1237 1137 1253
rect 1263 1287 1329 1303
rect 1377 1299 1407 1325
rect 1473 1303 1503 1325
rect 1263 1253 1279 1287
rect 1313 1253 1329 1287
rect 1263 1237 1329 1253
rect 1455 1287 1521 1303
rect 1569 1299 1599 1325
rect 1665 1303 1695 1325
rect 1455 1253 1471 1287
rect 1505 1253 1521 1287
rect 1455 1237 1521 1253
rect 1647 1287 1713 1303
rect 1761 1299 1791 1325
rect 1857 1303 1887 1325
rect 1647 1253 1663 1287
rect 1697 1253 1713 1287
rect 1647 1237 1713 1253
rect 1839 1287 1905 1303
rect 1839 1253 1855 1287
rect 1889 1253 1905 1287
rect 1839 1237 1905 1253
rect -1809 1179 -1743 1195
rect -1809 1145 -1793 1179
rect -1759 1145 -1743 1179
rect -1887 1107 -1857 1133
rect -1809 1129 -1743 1145
rect -1617 1179 -1551 1195
rect -1617 1145 -1601 1179
rect -1567 1145 -1551 1179
rect -1791 1107 -1761 1129
rect -1695 1107 -1665 1133
rect -1617 1129 -1551 1145
rect -1425 1179 -1359 1195
rect -1425 1145 -1409 1179
rect -1375 1145 -1359 1179
rect -1599 1107 -1569 1129
rect -1503 1107 -1473 1133
rect -1425 1129 -1359 1145
rect -1233 1179 -1167 1195
rect -1233 1145 -1217 1179
rect -1183 1145 -1167 1179
rect -1407 1107 -1377 1129
rect -1311 1107 -1281 1133
rect -1233 1129 -1167 1145
rect -1041 1179 -975 1195
rect -1041 1145 -1025 1179
rect -991 1145 -975 1179
rect -1215 1107 -1185 1129
rect -1119 1107 -1089 1133
rect -1041 1129 -975 1145
rect -849 1179 -783 1195
rect -849 1145 -833 1179
rect -799 1145 -783 1179
rect -1023 1107 -993 1129
rect -927 1107 -897 1133
rect -849 1129 -783 1145
rect -657 1179 -591 1195
rect -657 1145 -641 1179
rect -607 1145 -591 1179
rect -831 1107 -801 1129
rect -735 1107 -705 1133
rect -657 1129 -591 1145
rect -465 1179 -399 1195
rect -465 1145 -449 1179
rect -415 1145 -399 1179
rect -639 1107 -609 1129
rect -543 1107 -513 1133
rect -465 1129 -399 1145
rect -273 1179 -207 1195
rect -273 1145 -257 1179
rect -223 1145 -207 1179
rect -447 1107 -417 1129
rect -351 1107 -321 1133
rect -273 1129 -207 1145
rect -81 1179 -15 1195
rect -81 1145 -65 1179
rect -31 1145 -15 1179
rect -255 1107 -225 1129
rect -159 1107 -129 1133
rect -81 1129 -15 1145
rect 111 1179 177 1195
rect 111 1145 127 1179
rect 161 1145 177 1179
rect -63 1107 -33 1129
rect 33 1107 63 1133
rect 111 1129 177 1145
rect 303 1179 369 1195
rect 303 1145 319 1179
rect 353 1145 369 1179
rect 129 1107 159 1129
rect 225 1107 255 1133
rect 303 1129 369 1145
rect 495 1179 561 1195
rect 495 1145 511 1179
rect 545 1145 561 1179
rect 321 1107 351 1129
rect 417 1107 447 1133
rect 495 1129 561 1145
rect 687 1179 753 1195
rect 687 1145 703 1179
rect 737 1145 753 1179
rect 513 1107 543 1129
rect 609 1107 639 1133
rect 687 1129 753 1145
rect 879 1179 945 1195
rect 879 1145 895 1179
rect 929 1145 945 1179
rect 705 1107 735 1129
rect 801 1107 831 1133
rect 879 1129 945 1145
rect 1071 1179 1137 1195
rect 1071 1145 1087 1179
rect 1121 1145 1137 1179
rect 897 1107 927 1129
rect 993 1107 1023 1133
rect 1071 1129 1137 1145
rect 1263 1179 1329 1195
rect 1263 1145 1279 1179
rect 1313 1145 1329 1179
rect 1089 1107 1119 1129
rect 1185 1107 1215 1133
rect 1263 1129 1329 1145
rect 1455 1179 1521 1195
rect 1455 1145 1471 1179
rect 1505 1145 1521 1179
rect 1281 1107 1311 1129
rect 1377 1107 1407 1133
rect 1455 1129 1521 1145
rect 1647 1179 1713 1195
rect 1647 1145 1663 1179
rect 1697 1145 1713 1179
rect 1473 1107 1503 1129
rect 1569 1107 1599 1133
rect 1647 1129 1713 1145
rect 1839 1179 1905 1195
rect 1839 1145 1855 1179
rect 1889 1145 1905 1179
rect 1665 1107 1695 1129
rect 1761 1107 1791 1133
rect 1839 1129 1905 1145
rect 1857 1107 1887 1129
rect -1887 695 -1857 717
rect -1905 679 -1839 695
rect -1791 691 -1761 717
rect -1695 695 -1665 717
rect -1905 645 -1889 679
rect -1855 645 -1839 679
rect -1905 629 -1839 645
rect -1713 679 -1647 695
rect -1599 691 -1569 717
rect -1503 695 -1473 717
rect -1713 645 -1697 679
rect -1663 645 -1647 679
rect -1713 629 -1647 645
rect -1521 679 -1455 695
rect -1407 691 -1377 717
rect -1311 695 -1281 717
rect -1521 645 -1505 679
rect -1471 645 -1455 679
rect -1521 629 -1455 645
rect -1329 679 -1263 695
rect -1215 691 -1185 717
rect -1119 695 -1089 717
rect -1329 645 -1313 679
rect -1279 645 -1263 679
rect -1329 629 -1263 645
rect -1137 679 -1071 695
rect -1023 691 -993 717
rect -927 695 -897 717
rect -1137 645 -1121 679
rect -1087 645 -1071 679
rect -1137 629 -1071 645
rect -945 679 -879 695
rect -831 691 -801 717
rect -735 695 -705 717
rect -945 645 -929 679
rect -895 645 -879 679
rect -945 629 -879 645
rect -753 679 -687 695
rect -639 691 -609 717
rect -543 695 -513 717
rect -753 645 -737 679
rect -703 645 -687 679
rect -753 629 -687 645
rect -561 679 -495 695
rect -447 691 -417 717
rect -351 695 -321 717
rect -561 645 -545 679
rect -511 645 -495 679
rect -561 629 -495 645
rect -369 679 -303 695
rect -255 691 -225 717
rect -159 695 -129 717
rect -369 645 -353 679
rect -319 645 -303 679
rect -369 629 -303 645
rect -177 679 -111 695
rect -63 691 -33 717
rect 33 695 63 717
rect -177 645 -161 679
rect -127 645 -111 679
rect -177 629 -111 645
rect 15 679 81 695
rect 129 691 159 717
rect 225 695 255 717
rect 15 645 31 679
rect 65 645 81 679
rect 15 629 81 645
rect 207 679 273 695
rect 321 691 351 717
rect 417 695 447 717
rect 207 645 223 679
rect 257 645 273 679
rect 207 629 273 645
rect 399 679 465 695
rect 513 691 543 717
rect 609 695 639 717
rect 399 645 415 679
rect 449 645 465 679
rect 399 629 465 645
rect 591 679 657 695
rect 705 691 735 717
rect 801 695 831 717
rect 591 645 607 679
rect 641 645 657 679
rect 591 629 657 645
rect 783 679 849 695
rect 897 691 927 717
rect 993 695 1023 717
rect 783 645 799 679
rect 833 645 849 679
rect 783 629 849 645
rect 975 679 1041 695
rect 1089 691 1119 717
rect 1185 695 1215 717
rect 975 645 991 679
rect 1025 645 1041 679
rect 975 629 1041 645
rect 1167 679 1233 695
rect 1281 691 1311 717
rect 1377 695 1407 717
rect 1167 645 1183 679
rect 1217 645 1233 679
rect 1167 629 1233 645
rect 1359 679 1425 695
rect 1473 691 1503 717
rect 1569 695 1599 717
rect 1359 645 1375 679
rect 1409 645 1425 679
rect 1359 629 1425 645
rect 1551 679 1617 695
rect 1665 691 1695 717
rect 1761 695 1791 717
rect 1551 645 1567 679
rect 1601 645 1617 679
rect 1551 629 1617 645
rect 1743 679 1809 695
rect 1857 691 1887 717
rect 1743 645 1759 679
rect 1793 645 1809 679
rect 1743 629 1809 645
rect -1905 571 -1839 587
rect -1905 537 -1889 571
rect -1855 537 -1839 571
rect -1905 521 -1839 537
rect -1713 571 -1647 587
rect -1713 537 -1697 571
rect -1663 537 -1647 571
rect -1887 499 -1857 521
rect -1791 499 -1761 525
rect -1713 521 -1647 537
rect -1521 571 -1455 587
rect -1521 537 -1505 571
rect -1471 537 -1455 571
rect -1695 499 -1665 521
rect -1599 499 -1569 525
rect -1521 521 -1455 537
rect -1329 571 -1263 587
rect -1329 537 -1313 571
rect -1279 537 -1263 571
rect -1503 499 -1473 521
rect -1407 499 -1377 525
rect -1329 521 -1263 537
rect -1137 571 -1071 587
rect -1137 537 -1121 571
rect -1087 537 -1071 571
rect -1311 499 -1281 521
rect -1215 499 -1185 525
rect -1137 521 -1071 537
rect -945 571 -879 587
rect -945 537 -929 571
rect -895 537 -879 571
rect -1119 499 -1089 521
rect -1023 499 -993 525
rect -945 521 -879 537
rect -753 571 -687 587
rect -753 537 -737 571
rect -703 537 -687 571
rect -927 499 -897 521
rect -831 499 -801 525
rect -753 521 -687 537
rect -561 571 -495 587
rect -561 537 -545 571
rect -511 537 -495 571
rect -735 499 -705 521
rect -639 499 -609 525
rect -561 521 -495 537
rect -369 571 -303 587
rect -369 537 -353 571
rect -319 537 -303 571
rect -543 499 -513 521
rect -447 499 -417 525
rect -369 521 -303 537
rect -177 571 -111 587
rect -177 537 -161 571
rect -127 537 -111 571
rect -351 499 -321 521
rect -255 499 -225 525
rect -177 521 -111 537
rect 15 571 81 587
rect 15 537 31 571
rect 65 537 81 571
rect -159 499 -129 521
rect -63 499 -33 525
rect 15 521 81 537
rect 207 571 273 587
rect 207 537 223 571
rect 257 537 273 571
rect 33 499 63 521
rect 129 499 159 525
rect 207 521 273 537
rect 399 571 465 587
rect 399 537 415 571
rect 449 537 465 571
rect 225 499 255 521
rect 321 499 351 525
rect 399 521 465 537
rect 591 571 657 587
rect 591 537 607 571
rect 641 537 657 571
rect 417 499 447 521
rect 513 499 543 525
rect 591 521 657 537
rect 783 571 849 587
rect 783 537 799 571
rect 833 537 849 571
rect 609 499 639 521
rect 705 499 735 525
rect 783 521 849 537
rect 975 571 1041 587
rect 975 537 991 571
rect 1025 537 1041 571
rect 801 499 831 521
rect 897 499 927 525
rect 975 521 1041 537
rect 1167 571 1233 587
rect 1167 537 1183 571
rect 1217 537 1233 571
rect 993 499 1023 521
rect 1089 499 1119 525
rect 1167 521 1233 537
rect 1359 571 1425 587
rect 1359 537 1375 571
rect 1409 537 1425 571
rect 1185 499 1215 521
rect 1281 499 1311 525
rect 1359 521 1425 537
rect 1551 571 1617 587
rect 1551 537 1567 571
rect 1601 537 1617 571
rect 1377 499 1407 521
rect 1473 499 1503 525
rect 1551 521 1617 537
rect 1743 571 1809 587
rect 1743 537 1759 571
rect 1793 537 1809 571
rect 1569 499 1599 521
rect 1665 499 1695 525
rect 1743 521 1809 537
rect 1761 499 1791 521
rect 1857 499 1887 525
rect -1887 83 -1857 109
rect -1791 87 -1761 109
rect -1809 71 -1743 87
rect -1695 83 -1665 109
rect -1599 87 -1569 109
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1809 21 -1743 37
rect -1617 71 -1551 87
rect -1503 83 -1473 109
rect -1407 87 -1377 109
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1617 21 -1551 37
rect -1425 71 -1359 87
rect -1311 83 -1281 109
rect -1215 87 -1185 109
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1425 21 -1359 37
rect -1233 71 -1167 87
rect -1119 83 -1089 109
rect -1023 87 -993 109
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1233 21 -1167 37
rect -1041 71 -975 87
rect -927 83 -897 109
rect -831 87 -801 109
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -1041 21 -975 37
rect -849 71 -783 87
rect -735 83 -705 109
rect -639 87 -609 109
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -543 83 -513 109
rect -447 87 -417 109
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -351 83 -321 109
rect -255 87 -225 109
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -159 83 -129 109
rect -63 87 -33 109
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect 33 83 63 109
rect 129 87 159 109
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 225 83 255 109
rect 321 87 351 109
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 417 83 447 109
rect 513 87 543 109
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 609 83 639 109
rect 705 87 735 109
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 801 83 831 109
rect 897 87 927 109
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 993 83 1023 109
rect 1089 87 1119 109
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect 1071 71 1137 87
rect 1185 83 1215 109
rect 1281 87 1311 109
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1071 21 1137 37
rect 1263 71 1329 87
rect 1377 83 1407 109
rect 1473 87 1503 109
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1263 21 1329 37
rect 1455 71 1521 87
rect 1569 83 1599 109
rect 1665 87 1695 109
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1455 21 1521 37
rect 1647 71 1713 87
rect 1761 83 1791 109
rect 1857 87 1887 109
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1647 21 1713 37
rect 1839 71 1905 87
rect 1839 37 1855 71
rect 1889 37 1905 71
rect 1839 21 1905 37
rect -1809 -37 -1743 -21
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1887 -109 -1857 -83
rect -1809 -87 -1743 -71
rect -1617 -37 -1551 -21
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1791 -109 -1761 -87
rect -1695 -109 -1665 -83
rect -1617 -87 -1551 -71
rect -1425 -37 -1359 -21
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1599 -109 -1569 -87
rect -1503 -109 -1473 -83
rect -1425 -87 -1359 -71
rect -1233 -37 -1167 -21
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1407 -109 -1377 -87
rect -1311 -109 -1281 -83
rect -1233 -87 -1167 -71
rect -1041 -37 -975 -21
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -1215 -109 -1185 -87
rect -1119 -109 -1089 -83
rect -1041 -87 -975 -71
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -1023 -109 -993 -87
rect -927 -109 -897 -83
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -831 -109 -801 -87
rect -735 -109 -705 -83
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -639 -109 -609 -87
rect -543 -109 -513 -83
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -447 -109 -417 -87
rect -351 -109 -321 -83
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -255 -109 -225 -87
rect -159 -109 -129 -83
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect -63 -109 -33 -87
rect 33 -109 63 -83
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 129 -109 159 -87
rect 225 -109 255 -83
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 321 -109 351 -87
rect 417 -109 447 -83
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 513 -109 543 -87
rect 609 -109 639 -83
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 705 -109 735 -87
rect 801 -109 831 -83
rect 879 -87 945 -71
rect 1071 -37 1137 -21
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 897 -109 927 -87
rect 993 -109 1023 -83
rect 1071 -87 1137 -71
rect 1263 -37 1329 -21
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1089 -109 1119 -87
rect 1185 -109 1215 -83
rect 1263 -87 1329 -71
rect 1455 -37 1521 -21
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1281 -109 1311 -87
rect 1377 -109 1407 -83
rect 1455 -87 1521 -71
rect 1647 -37 1713 -21
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1473 -109 1503 -87
rect 1569 -109 1599 -83
rect 1647 -87 1713 -71
rect 1839 -37 1905 -21
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect 1665 -109 1695 -87
rect 1761 -109 1791 -83
rect 1839 -87 1905 -71
rect 1857 -109 1887 -87
rect -1887 -521 -1857 -499
rect -1905 -537 -1839 -521
rect -1791 -525 -1761 -499
rect -1695 -521 -1665 -499
rect -1905 -571 -1889 -537
rect -1855 -571 -1839 -537
rect -1905 -587 -1839 -571
rect -1713 -537 -1647 -521
rect -1599 -525 -1569 -499
rect -1503 -521 -1473 -499
rect -1713 -571 -1697 -537
rect -1663 -571 -1647 -537
rect -1713 -587 -1647 -571
rect -1521 -537 -1455 -521
rect -1407 -525 -1377 -499
rect -1311 -521 -1281 -499
rect -1521 -571 -1505 -537
rect -1471 -571 -1455 -537
rect -1521 -587 -1455 -571
rect -1329 -537 -1263 -521
rect -1215 -525 -1185 -499
rect -1119 -521 -1089 -499
rect -1329 -571 -1313 -537
rect -1279 -571 -1263 -537
rect -1329 -587 -1263 -571
rect -1137 -537 -1071 -521
rect -1023 -525 -993 -499
rect -927 -521 -897 -499
rect -1137 -571 -1121 -537
rect -1087 -571 -1071 -537
rect -1137 -587 -1071 -571
rect -945 -537 -879 -521
rect -831 -525 -801 -499
rect -735 -521 -705 -499
rect -945 -571 -929 -537
rect -895 -571 -879 -537
rect -945 -587 -879 -571
rect -753 -537 -687 -521
rect -639 -525 -609 -499
rect -543 -521 -513 -499
rect -753 -571 -737 -537
rect -703 -571 -687 -537
rect -753 -587 -687 -571
rect -561 -537 -495 -521
rect -447 -525 -417 -499
rect -351 -521 -321 -499
rect -561 -571 -545 -537
rect -511 -571 -495 -537
rect -561 -587 -495 -571
rect -369 -537 -303 -521
rect -255 -525 -225 -499
rect -159 -521 -129 -499
rect -369 -571 -353 -537
rect -319 -571 -303 -537
rect -369 -587 -303 -571
rect -177 -537 -111 -521
rect -63 -525 -33 -499
rect 33 -521 63 -499
rect -177 -571 -161 -537
rect -127 -571 -111 -537
rect -177 -587 -111 -571
rect 15 -537 81 -521
rect 129 -525 159 -499
rect 225 -521 255 -499
rect 15 -571 31 -537
rect 65 -571 81 -537
rect 15 -587 81 -571
rect 207 -537 273 -521
rect 321 -525 351 -499
rect 417 -521 447 -499
rect 207 -571 223 -537
rect 257 -571 273 -537
rect 207 -587 273 -571
rect 399 -537 465 -521
rect 513 -525 543 -499
rect 609 -521 639 -499
rect 399 -571 415 -537
rect 449 -571 465 -537
rect 399 -587 465 -571
rect 591 -537 657 -521
rect 705 -525 735 -499
rect 801 -521 831 -499
rect 591 -571 607 -537
rect 641 -571 657 -537
rect 591 -587 657 -571
rect 783 -537 849 -521
rect 897 -525 927 -499
rect 993 -521 1023 -499
rect 783 -571 799 -537
rect 833 -571 849 -537
rect 783 -587 849 -571
rect 975 -537 1041 -521
rect 1089 -525 1119 -499
rect 1185 -521 1215 -499
rect 975 -571 991 -537
rect 1025 -571 1041 -537
rect 975 -587 1041 -571
rect 1167 -537 1233 -521
rect 1281 -525 1311 -499
rect 1377 -521 1407 -499
rect 1167 -571 1183 -537
rect 1217 -571 1233 -537
rect 1167 -587 1233 -571
rect 1359 -537 1425 -521
rect 1473 -525 1503 -499
rect 1569 -521 1599 -499
rect 1359 -571 1375 -537
rect 1409 -571 1425 -537
rect 1359 -587 1425 -571
rect 1551 -537 1617 -521
rect 1665 -525 1695 -499
rect 1761 -521 1791 -499
rect 1551 -571 1567 -537
rect 1601 -571 1617 -537
rect 1551 -587 1617 -571
rect 1743 -537 1809 -521
rect 1857 -525 1887 -499
rect 1743 -571 1759 -537
rect 1793 -571 1809 -537
rect 1743 -587 1809 -571
rect -1905 -645 -1839 -629
rect -1905 -679 -1889 -645
rect -1855 -679 -1839 -645
rect -1905 -695 -1839 -679
rect -1713 -645 -1647 -629
rect -1713 -679 -1697 -645
rect -1663 -679 -1647 -645
rect -1887 -717 -1857 -695
rect -1791 -717 -1761 -691
rect -1713 -695 -1647 -679
rect -1521 -645 -1455 -629
rect -1521 -679 -1505 -645
rect -1471 -679 -1455 -645
rect -1695 -717 -1665 -695
rect -1599 -717 -1569 -691
rect -1521 -695 -1455 -679
rect -1329 -645 -1263 -629
rect -1329 -679 -1313 -645
rect -1279 -679 -1263 -645
rect -1503 -717 -1473 -695
rect -1407 -717 -1377 -691
rect -1329 -695 -1263 -679
rect -1137 -645 -1071 -629
rect -1137 -679 -1121 -645
rect -1087 -679 -1071 -645
rect -1311 -717 -1281 -695
rect -1215 -717 -1185 -691
rect -1137 -695 -1071 -679
rect -945 -645 -879 -629
rect -945 -679 -929 -645
rect -895 -679 -879 -645
rect -1119 -717 -1089 -695
rect -1023 -717 -993 -691
rect -945 -695 -879 -679
rect -753 -645 -687 -629
rect -753 -679 -737 -645
rect -703 -679 -687 -645
rect -927 -717 -897 -695
rect -831 -717 -801 -691
rect -753 -695 -687 -679
rect -561 -645 -495 -629
rect -561 -679 -545 -645
rect -511 -679 -495 -645
rect -735 -717 -705 -695
rect -639 -717 -609 -691
rect -561 -695 -495 -679
rect -369 -645 -303 -629
rect -369 -679 -353 -645
rect -319 -679 -303 -645
rect -543 -717 -513 -695
rect -447 -717 -417 -691
rect -369 -695 -303 -679
rect -177 -645 -111 -629
rect -177 -679 -161 -645
rect -127 -679 -111 -645
rect -351 -717 -321 -695
rect -255 -717 -225 -691
rect -177 -695 -111 -679
rect 15 -645 81 -629
rect 15 -679 31 -645
rect 65 -679 81 -645
rect -159 -717 -129 -695
rect -63 -717 -33 -691
rect 15 -695 81 -679
rect 207 -645 273 -629
rect 207 -679 223 -645
rect 257 -679 273 -645
rect 33 -717 63 -695
rect 129 -717 159 -691
rect 207 -695 273 -679
rect 399 -645 465 -629
rect 399 -679 415 -645
rect 449 -679 465 -645
rect 225 -717 255 -695
rect 321 -717 351 -691
rect 399 -695 465 -679
rect 591 -645 657 -629
rect 591 -679 607 -645
rect 641 -679 657 -645
rect 417 -717 447 -695
rect 513 -717 543 -691
rect 591 -695 657 -679
rect 783 -645 849 -629
rect 783 -679 799 -645
rect 833 -679 849 -645
rect 609 -717 639 -695
rect 705 -717 735 -691
rect 783 -695 849 -679
rect 975 -645 1041 -629
rect 975 -679 991 -645
rect 1025 -679 1041 -645
rect 801 -717 831 -695
rect 897 -717 927 -691
rect 975 -695 1041 -679
rect 1167 -645 1233 -629
rect 1167 -679 1183 -645
rect 1217 -679 1233 -645
rect 993 -717 1023 -695
rect 1089 -717 1119 -691
rect 1167 -695 1233 -679
rect 1359 -645 1425 -629
rect 1359 -679 1375 -645
rect 1409 -679 1425 -645
rect 1185 -717 1215 -695
rect 1281 -717 1311 -691
rect 1359 -695 1425 -679
rect 1551 -645 1617 -629
rect 1551 -679 1567 -645
rect 1601 -679 1617 -645
rect 1377 -717 1407 -695
rect 1473 -717 1503 -691
rect 1551 -695 1617 -679
rect 1743 -645 1809 -629
rect 1743 -679 1759 -645
rect 1793 -679 1809 -645
rect 1569 -717 1599 -695
rect 1665 -717 1695 -691
rect 1743 -695 1809 -679
rect 1761 -717 1791 -695
rect 1857 -717 1887 -691
rect -1887 -1133 -1857 -1107
rect -1791 -1129 -1761 -1107
rect -1809 -1145 -1743 -1129
rect -1695 -1133 -1665 -1107
rect -1599 -1129 -1569 -1107
rect -1809 -1179 -1793 -1145
rect -1759 -1179 -1743 -1145
rect -1809 -1195 -1743 -1179
rect -1617 -1145 -1551 -1129
rect -1503 -1133 -1473 -1107
rect -1407 -1129 -1377 -1107
rect -1617 -1179 -1601 -1145
rect -1567 -1179 -1551 -1145
rect -1617 -1195 -1551 -1179
rect -1425 -1145 -1359 -1129
rect -1311 -1133 -1281 -1107
rect -1215 -1129 -1185 -1107
rect -1425 -1179 -1409 -1145
rect -1375 -1179 -1359 -1145
rect -1425 -1195 -1359 -1179
rect -1233 -1145 -1167 -1129
rect -1119 -1133 -1089 -1107
rect -1023 -1129 -993 -1107
rect -1233 -1179 -1217 -1145
rect -1183 -1179 -1167 -1145
rect -1233 -1195 -1167 -1179
rect -1041 -1145 -975 -1129
rect -927 -1133 -897 -1107
rect -831 -1129 -801 -1107
rect -1041 -1179 -1025 -1145
rect -991 -1179 -975 -1145
rect -1041 -1195 -975 -1179
rect -849 -1145 -783 -1129
rect -735 -1133 -705 -1107
rect -639 -1129 -609 -1107
rect -849 -1179 -833 -1145
rect -799 -1179 -783 -1145
rect -849 -1195 -783 -1179
rect -657 -1145 -591 -1129
rect -543 -1133 -513 -1107
rect -447 -1129 -417 -1107
rect -657 -1179 -641 -1145
rect -607 -1179 -591 -1145
rect -657 -1195 -591 -1179
rect -465 -1145 -399 -1129
rect -351 -1133 -321 -1107
rect -255 -1129 -225 -1107
rect -465 -1179 -449 -1145
rect -415 -1179 -399 -1145
rect -465 -1195 -399 -1179
rect -273 -1145 -207 -1129
rect -159 -1133 -129 -1107
rect -63 -1129 -33 -1107
rect -273 -1179 -257 -1145
rect -223 -1179 -207 -1145
rect -273 -1195 -207 -1179
rect -81 -1145 -15 -1129
rect 33 -1133 63 -1107
rect 129 -1129 159 -1107
rect -81 -1179 -65 -1145
rect -31 -1179 -15 -1145
rect -81 -1195 -15 -1179
rect 111 -1145 177 -1129
rect 225 -1133 255 -1107
rect 321 -1129 351 -1107
rect 111 -1179 127 -1145
rect 161 -1179 177 -1145
rect 111 -1195 177 -1179
rect 303 -1145 369 -1129
rect 417 -1133 447 -1107
rect 513 -1129 543 -1107
rect 303 -1179 319 -1145
rect 353 -1179 369 -1145
rect 303 -1195 369 -1179
rect 495 -1145 561 -1129
rect 609 -1133 639 -1107
rect 705 -1129 735 -1107
rect 495 -1179 511 -1145
rect 545 -1179 561 -1145
rect 495 -1195 561 -1179
rect 687 -1145 753 -1129
rect 801 -1133 831 -1107
rect 897 -1129 927 -1107
rect 687 -1179 703 -1145
rect 737 -1179 753 -1145
rect 687 -1195 753 -1179
rect 879 -1145 945 -1129
rect 993 -1133 1023 -1107
rect 1089 -1129 1119 -1107
rect 879 -1179 895 -1145
rect 929 -1179 945 -1145
rect 879 -1195 945 -1179
rect 1071 -1145 1137 -1129
rect 1185 -1133 1215 -1107
rect 1281 -1129 1311 -1107
rect 1071 -1179 1087 -1145
rect 1121 -1179 1137 -1145
rect 1071 -1195 1137 -1179
rect 1263 -1145 1329 -1129
rect 1377 -1133 1407 -1107
rect 1473 -1129 1503 -1107
rect 1263 -1179 1279 -1145
rect 1313 -1179 1329 -1145
rect 1263 -1195 1329 -1179
rect 1455 -1145 1521 -1129
rect 1569 -1133 1599 -1107
rect 1665 -1129 1695 -1107
rect 1455 -1179 1471 -1145
rect 1505 -1179 1521 -1145
rect 1455 -1195 1521 -1179
rect 1647 -1145 1713 -1129
rect 1761 -1133 1791 -1107
rect 1857 -1129 1887 -1107
rect 1647 -1179 1663 -1145
rect 1697 -1179 1713 -1145
rect 1647 -1195 1713 -1179
rect 1839 -1145 1905 -1129
rect 1839 -1179 1855 -1145
rect 1889 -1179 1905 -1145
rect 1839 -1195 1905 -1179
rect -1809 -1253 -1743 -1237
rect -1809 -1287 -1793 -1253
rect -1759 -1287 -1743 -1253
rect -1887 -1325 -1857 -1299
rect -1809 -1303 -1743 -1287
rect -1617 -1253 -1551 -1237
rect -1617 -1287 -1601 -1253
rect -1567 -1287 -1551 -1253
rect -1791 -1325 -1761 -1303
rect -1695 -1325 -1665 -1299
rect -1617 -1303 -1551 -1287
rect -1425 -1253 -1359 -1237
rect -1425 -1287 -1409 -1253
rect -1375 -1287 -1359 -1253
rect -1599 -1325 -1569 -1303
rect -1503 -1325 -1473 -1299
rect -1425 -1303 -1359 -1287
rect -1233 -1253 -1167 -1237
rect -1233 -1287 -1217 -1253
rect -1183 -1287 -1167 -1253
rect -1407 -1325 -1377 -1303
rect -1311 -1325 -1281 -1299
rect -1233 -1303 -1167 -1287
rect -1041 -1253 -975 -1237
rect -1041 -1287 -1025 -1253
rect -991 -1287 -975 -1253
rect -1215 -1325 -1185 -1303
rect -1119 -1325 -1089 -1299
rect -1041 -1303 -975 -1287
rect -849 -1253 -783 -1237
rect -849 -1287 -833 -1253
rect -799 -1287 -783 -1253
rect -1023 -1325 -993 -1303
rect -927 -1325 -897 -1299
rect -849 -1303 -783 -1287
rect -657 -1253 -591 -1237
rect -657 -1287 -641 -1253
rect -607 -1287 -591 -1253
rect -831 -1325 -801 -1303
rect -735 -1325 -705 -1299
rect -657 -1303 -591 -1287
rect -465 -1253 -399 -1237
rect -465 -1287 -449 -1253
rect -415 -1287 -399 -1253
rect -639 -1325 -609 -1303
rect -543 -1325 -513 -1299
rect -465 -1303 -399 -1287
rect -273 -1253 -207 -1237
rect -273 -1287 -257 -1253
rect -223 -1287 -207 -1253
rect -447 -1325 -417 -1303
rect -351 -1325 -321 -1299
rect -273 -1303 -207 -1287
rect -81 -1253 -15 -1237
rect -81 -1287 -65 -1253
rect -31 -1287 -15 -1253
rect -255 -1325 -225 -1303
rect -159 -1325 -129 -1299
rect -81 -1303 -15 -1287
rect 111 -1253 177 -1237
rect 111 -1287 127 -1253
rect 161 -1287 177 -1253
rect -63 -1325 -33 -1303
rect 33 -1325 63 -1299
rect 111 -1303 177 -1287
rect 303 -1253 369 -1237
rect 303 -1287 319 -1253
rect 353 -1287 369 -1253
rect 129 -1325 159 -1303
rect 225 -1325 255 -1299
rect 303 -1303 369 -1287
rect 495 -1253 561 -1237
rect 495 -1287 511 -1253
rect 545 -1287 561 -1253
rect 321 -1325 351 -1303
rect 417 -1325 447 -1299
rect 495 -1303 561 -1287
rect 687 -1253 753 -1237
rect 687 -1287 703 -1253
rect 737 -1287 753 -1253
rect 513 -1325 543 -1303
rect 609 -1325 639 -1299
rect 687 -1303 753 -1287
rect 879 -1253 945 -1237
rect 879 -1287 895 -1253
rect 929 -1287 945 -1253
rect 705 -1325 735 -1303
rect 801 -1325 831 -1299
rect 879 -1303 945 -1287
rect 1071 -1253 1137 -1237
rect 1071 -1287 1087 -1253
rect 1121 -1287 1137 -1253
rect 897 -1325 927 -1303
rect 993 -1325 1023 -1299
rect 1071 -1303 1137 -1287
rect 1263 -1253 1329 -1237
rect 1263 -1287 1279 -1253
rect 1313 -1287 1329 -1253
rect 1089 -1325 1119 -1303
rect 1185 -1325 1215 -1299
rect 1263 -1303 1329 -1287
rect 1455 -1253 1521 -1237
rect 1455 -1287 1471 -1253
rect 1505 -1287 1521 -1253
rect 1281 -1325 1311 -1303
rect 1377 -1325 1407 -1299
rect 1455 -1303 1521 -1287
rect 1647 -1253 1713 -1237
rect 1647 -1287 1663 -1253
rect 1697 -1287 1713 -1253
rect 1473 -1325 1503 -1303
rect 1569 -1325 1599 -1299
rect 1647 -1303 1713 -1287
rect 1839 -1253 1905 -1237
rect 1839 -1287 1855 -1253
rect 1889 -1287 1905 -1253
rect 1665 -1325 1695 -1303
rect 1761 -1325 1791 -1299
rect 1839 -1303 1905 -1287
rect 1857 -1325 1887 -1303
rect -1887 -1737 -1857 -1715
rect -1905 -1753 -1839 -1737
rect -1791 -1741 -1761 -1715
rect -1695 -1737 -1665 -1715
rect -1905 -1787 -1889 -1753
rect -1855 -1787 -1839 -1753
rect -1905 -1803 -1839 -1787
rect -1713 -1753 -1647 -1737
rect -1599 -1741 -1569 -1715
rect -1503 -1737 -1473 -1715
rect -1713 -1787 -1697 -1753
rect -1663 -1787 -1647 -1753
rect -1713 -1803 -1647 -1787
rect -1521 -1753 -1455 -1737
rect -1407 -1741 -1377 -1715
rect -1311 -1737 -1281 -1715
rect -1521 -1787 -1505 -1753
rect -1471 -1787 -1455 -1753
rect -1521 -1803 -1455 -1787
rect -1329 -1753 -1263 -1737
rect -1215 -1741 -1185 -1715
rect -1119 -1737 -1089 -1715
rect -1329 -1787 -1313 -1753
rect -1279 -1787 -1263 -1753
rect -1329 -1803 -1263 -1787
rect -1137 -1753 -1071 -1737
rect -1023 -1741 -993 -1715
rect -927 -1737 -897 -1715
rect -1137 -1787 -1121 -1753
rect -1087 -1787 -1071 -1753
rect -1137 -1803 -1071 -1787
rect -945 -1753 -879 -1737
rect -831 -1741 -801 -1715
rect -735 -1737 -705 -1715
rect -945 -1787 -929 -1753
rect -895 -1787 -879 -1753
rect -945 -1803 -879 -1787
rect -753 -1753 -687 -1737
rect -639 -1741 -609 -1715
rect -543 -1737 -513 -1715
rect -753 -1787 -737 -1753
rect -703 -1787 -687 -1753
rect -753 -1803 -687 -1787
rect -561 -1753 -495 -1737
rect -447 -1741 -417 -1715
rect -351 -1737 -321 -1715
rect -561 -1787 -545 -1753
rect -511 -1787 -495 -1753
rect -561 -1803 -495 -1787
rect -369 -1753 -303 -1737
rect -255 -1741 -225 -1715
rect -159 -1737 -129 -1715
rect -369 -1787 -353 -1753
rect -319 -1787 -303 -1753
rect -369 -1803 -303 -1787
rect -177 -1753 -111 -1737
rect -63 -1741 -33 -1715
rect 33 -1737 63 -1715
rect -177 -1787 -161 -1753
rect -127 -1787 -111 -1753
rect -177 -1803 -111 -1787
rect 15 -1753 81 -1737
rect 129 -1741 159 -1715
rect 225 -1737 255 -1715
rect 15 -1787 31 -1753
rect 65 -1787 81 -1753
rect 15 -1803 81 -1787
rect 207 -1753 273 -1737
rect 321 -1741 351 -1715
rect 417 -1737 447 -1715
rect 207 -1787 223 -1753
rect 257 -1787 273 -1753
rect 207 -1803 273 -1787
rect 399 -1753 465 -1737
rect 513 -1741 543 -1715
rect 609 -1737 639 -1715
rect 399 -1787 415 -1753
rect 449 -1787 465 -1753
rect 399 -1803 465 -1787
rect 591 -1753 657 -1737
rect 705 -1741 735 -1715
rect 801 -1737 831 -1715
rect 591 -1787 607 -1753
rect 641 -1787 657 -1753
rect 591 -1803 657 -1787
rect 783 -1753 849 -1737
rect 897 -1741 927 -1715
rect 993 -1737 1023 -1715
rect 783 -1787 799 -1753
rect 833 -1787 849 -1753
rect 783 -1803 849 -1787
rect 975 -1753 1041 -1737
rect 1089 -1741 1119 -1715
rect 1185 -1737 1215 -1715
rect 975 -1787 991 -1753
rect 1025 -1787 1041 -1753
rect 975 -1803 1041 -1787
rect 1167 -1753 1233 -1737
rect 1281 -1741 1311 -1715
rect 1377 -1737 1407 -1715
rect 1167 -1787 1183 -1753
rect 1217 -1787 1233 -1753
rect 1167 -1803 1233 -1787
rect 1359 -1753 1425 -1737
rect 1473 -1741 1503 -1715
rect 1569 -1737 1599 -1715
rect 1359 -1787 1375 -1753
rect 1409 -1787 1425 -1753
rect 1359 -1803 1425 -1787
rect 1551 -1753 1617 -1737
rect 1665 -1741 1695 -1715
rect 1761 -1737 1791 -1715
rect 1551 -1787 1567 -1753
rect 1601 -1787 1617 -1753
rect 1551 -1803 1617 -1787
rect 1743 -1753 1809 -1737
rect 1857 -1741 1887 -1715
rect 1743 -1787 1759 -1753
rect 1793 -1787 1809 -1753
rect 1743 -1803 1809 -1787
<< polycont >>
rect -1889 1753 -1855 1787
rect -1697 1753 -1663 1787
rect -1505 1753 -1471 1787
rect -1313 1753 -1279 1787
rect -1121 1753 -1087 1787
rect -929 1753 -895 1787
rect -737 1753 -703 1787
rect -545 1753 -511 1787
rect -353 1753 -319 1787
rect -161 1753 -127 1787
rect 31 1753 65 1787
rect 223 1753 257 1787
rect 415 1753 449 1787
rect 607 1753 641 1787
rect 799 1753 833 1787
rect 991 1753 1025 1787
rect 1183 1753 1217 1787
rect 1375 1753 1409 1787
rect 1567 1753 1601 1787
rect 1759 1753 1793 1787
rect -1793 1253 -1759 1287
rect -1601 1253 -1567 1287
rect -1409 1253 -1375 1287
rect -1217 1253 -1183 1287
rect -1025 1253 -991 1287
rect -833 1253 -799 1287
rect -641 1253 -607 1287
rect -449 1253 -415 1287
rect -257 1253 -223 1287
rect -65 1253 -31 1287
rect 127 1253 161 1287
rect 319 1253 353 1287
rect 511 1253 545 1287
rect 703 1253 737 1287
rect 895 1253 929 1287
rect 1087 1253 1121 1287
rect 1279 1253 1313 1287
rect 1471 1253 1505 1287
rect 1663 1253 1697 1287
rect 1855 1253 1889 1287
rect -1793 1145 -1759 1179
rect -1601 1145 -1567 1179
rect -1409 1145 -1375 1179
rect -1217 1145 -1183 1179
rect -1025 1145 -991 1179
rect -833 1145 -799 1179
rect -641 1145 -607 1179
rect -449 1145 -415 1179
rect -257 1145 -223 1179
rect -65 1145 -31 1179
rect 127 1145 161 1179
rect 319 1145 353 1179
rect 511 1145 545 1179
rect 703 1145 737 1179
rect 895 1145 929 1179
rect 1087 1145 1121 1179
rect 1279 1145 1313 1179
rect 1471 1145 1505 1179
rect 1663 1145 1697 1179
rect 1855 1145 1889 1179
rect -1889 645 -1855 679
rect -1697 645 -1663 679
rect -1505 645 -1471 679
rect -1313 645 -1279 679
rect -1121 645 -1087 679
rect -929 645 -895 679
rect -737 645 -703 679
rect -545 645 -511 679
rect -353 645 -319 679
rect -161 645 -127 679
rect 31 645 65 679
rect 223 645 257 679
rect 415 645 449 679
rect 607 645 641 679
rect 799 645 833 679
rect 991 645 1025 679
rect 1183 645 1217 679
rect 1375 645 1409 679
rect 1567 645 1601 679
rect 1759 645 1793 679
rect -1889 537 -1855 571
rect -1697 537 -1663 571
rect -1505 537 -1471 571
rect -1313 537 -1279 571
rect -1121 537 -1087 571
rect -929 537 -895 571
rect -737 537 -703 571
rect -545 537 -511 571
rect -353 537 -319 571
rect -161 537 -127 571
rect 31 537 65 571
rect 223 537 257 571
rect 415 537 449 571
rect 607 537 641 571
rect 799 537 833 571
rect 991 537 1025 571
rect 1183 537 1217 571
rect 1375 537 1409 571
rect 1567 537 1601 571
rect 1759 537 1793 571
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect -1889 -571 -1855 -537
rect -1697 -571 -1663 -537
rect -1505 -571 -1471 -537
rect -1313 -571 -1279 -537
rect -1121 -571 -1087 -537
rect -929 -571 -895 -537
rect -737 -571 -703 -537
rect -545 -571 -511 -537
rect -353 -571 -319 -537
rect -161 -571 -127 -537
rect 31 -571 65 -537
rect 223 -571 257 -537
rect 415 -571 449 -537
rect 607 -571 641 -537
rect 799 -571 833 -537
rect 991 -571 1025 -537
rect 1183 -571 1217 -537
rect 1375 -571 1409 -537
rect 1567 -571 1601 -537
rect 1759 -571 1793 -537
rect -1889 -679 -1855 -645
rect -1697 -679 -1663 -645
rect -1505 -679 -1471 -645
rect -1313 -679 -1279 -645
rect -1121 -679 -1087 -645
rect -929 -679 -895 -645
rect -737 -679 -703 -645
rect -545 -679 -511 -645
rect -353 -679 -319 -645
rect -161 -679 -127 -645
rect 31 -679 65 -645
rect 223 -679 257 -645
rect 415 -679 449 -645
rect 607 -679 641 -645
rect 799 -679 833 -645
rect 991 -679 1025 -645
rect 1183 -679 1217 -645
rect 1375 -679 1409 -645
rect 1567 -679 1601 -645
rect 1759 -679 1793 -645
rect -1793 -1179 -1759 -1145
rect -1601 -1179 -1567 -1145
rect -1409 -1179 -1375 -1145
rect -1217 -1179 -1183 -1145
rect -1025 -1179 -991 -1145
rect -833 -1179 -799 -1145
rect -641 -1179 -607 -1145
rect -449 -1179 -415 -1145
rect -257 -1179 -223 -1145
rect -65 -1179 -31 -1145
rect 127 -1179 161 -1145
rect 319 -1179 353 -1145
rect 511 -1179 545 -1145
rect 703 -1179 737 -1145
rect 895 -1179 929 -1145
rect 1087 -1179 1121 -1145
rect 1279 -1179 1313 -1145
rect 1471 -1179 1505 -1145
rect 1663 -1179 1697 -1145
rect 1855 -1179 1889 -1145
rect -1793 -1287 -1759 -1253
rect -1601 -1287 -1567 -1253
rect -1409 -1287 -1375 -1253
rect -1217 -1287 -1183 -1253
rect -1025 -1287 -991 -1253
rect -833 -1287 -799 -1253
rect -641 -1287 -607 -1253
rect -449 -1287 -415 -1253
rect -257 -1287 -223 -1253
rect -65 -1287 -31 -1253
rect 127 -1287 161 -1253
rect 319 -1287 353 -1253
rect 511 -1287 545 -1253
rect 703 -1287 737 -1253
rect 895 -1287 929 -1253
rect 1087 -1287 1121 -1253
rect 1279 -1287 1313 -1253
rect 1471 -1287 1505 -1253
rect 1663 -1287 1697 -1253
rect 1855 -1287 1889 -1253
rect -1889 -1787 -1855 -1753
rect -1697 -1787 -1663 -1753
rect -1505 -1787 -1471 -1753
rect -1313 -1787 -1279 -1753
rect -1121 -1787 -1087 -1753
rect -929 -1787 -895 -1753
rect -737 -1787 -703 -1753
rect -545 -1787 -511 -1753
rect -353 -1787 -319 -1753
rect -161 -1787 -127 -1753
rect 31 -1787 65 -1753
rect 223 -1787 257 -1753
rect 415 -1787 449 -1753
rect 607 -1787 641 -1753
rect 799 -1787 833 -1753
rect 991 -1787 1025 -1753
rect 1183 -1787 1217 -1753
rect 1375 -1787 1409 -1753
rect 1567 -1787 1601 -1753
rect 1759 -1787 1793 -1753
<< locali >>
rect -2051 1855 -1955 1889
rect 1955 1855 2051 1889
rect -2051 1793 -2017 1855
rect 2017 1793 2051 1855
rect -1905 1753 -1889 1787
rect -1855 1753 -1839 1787
rect -1713 1753 -1697 1787
rect -1663 1753 -1647 1787
rect -1521 1753 -1505 1787
rect -1471 1753 -1455 1787
rect -1329 1753 -1313 1787
rect -1279 1753 -1263 1787
rect -1137 1753 -1121 1787
rect -1087 1753 -1071 1787
rect -945 1753 -929 1787
rect -895 1753 -879 1787
rect -753 1753 -737 1787
rect -703 1753 -687 1787
rect -561 1753 -545 1787
rect -511 1753 -495 1787
rect -369 1753 -353 1787
rect -319 1753 -303 1787
rect -177 1753 -161 1787
rect -127 1753 -111 1787
rect 15 1753 31 1787
rect 65 1753 81 1787
rect 207 1753 223 1787
rect 257 1753 273 1787
rect 399 1753 415 1787
rect 449 1753 465 1787
rect 591 1753 607 1787
rect 641 1753 657 1787
rect 783 1753 799 1787
rect 833 1753 849 1787
rect 975 1753 991 1787
rect 1025 1753 1041 1787
rect 1167 1753 1183 1787
rect 1217 1753 1233 1787
rect 1359 1753 1375 1787
rect 1409 1753 1425 1787
rect 1551 1753 1567 1787
rect 1601 1753 1617 1787
rect 1743 1753 1759 1787
rect 1793 1753 1809 1787
rect -1937 1703 -1903 1719
rect -1937 1321 -1903 1337
rect -1841 1703 -1807 1719
rect -1841 1321 -1807 1337
rect -1745 1703 -1711 1719
rect -1745 1321 -1711 1337
rect -1649 1703 -1615 1719
rect -1649 1321 -1615 1337
rect -1553 1703 -1519 1719
rect -1553 1321 -1519 1337
rect -1457 1703 -1423 1719
rect -1457 1321 -1423 1337
rect -1361 1703 -1327 1719
rect -1361 1321 -1327 1337
rect -1265 1703 -1231 1719
rect -1265 1321 -1231 1337
rect -1169 1703 -1135 1719
rect -1169 1321 -1135 1337
rect -1073 1703 -1039 1719
rect -1073 1321 -1039 1337
rect -977 1703 -943 1719
rect -977 1321 -943 1337
rect -881 1703 -847 1719
rect -881 1321 -847 1337
rect -785 1703 -751 1719
rect -785 1321 -751 1337
rect -689 1703 -655 1719
rect -689 1321 -655 1337
rect -593 1703 -559 1719
rect -593 1321 -559 1337
rect -497 1703 -463 1719
rect -497 1321 -463 1337
rect -401 1703 -367 1719
rect -401 1321 -367 1337
rect -305 1703 -271 1719
rect -305 1321 -271 1337
rect -209 1703 -175 1719
rect -209 1321 -175 1337
rect -113 1703 -79 1719
rect -113 1321 -79 1337
rect -17 1703 17 1719
rect -17 1321 17 1337
rect 79 1703 113 1719
rect 79 1321 113 1337
rect 175 1703 209 1719
rect 175 1321 209 1337
rect 271 1703 305 1719
rect 271 1321 305 1337
rect 367 1703 401 1719
rect 367 1321 401 1337
rect 463 1703 497 1719
rect 463 1321 497 1337
rect 559 1703 593 1719
rect 559 1321 593 1337
rect 655 1703 689 1719
rect 655 1321 689 1337
rect 751 1703 785 1719
rect 751 1321 785 1337
rect 847 1703 881 1719
rect 847 1321 881 1337
rect 943 1703 977 1719
rect 943 1321 977 1337
rect 1039 1703 1073 1719
rect 1039 1321 1073 1337
rect 1135 1703 1169 1719
rect 1135 1321 1169 1337
rect 1231 1703 1265 1719
rect 1231 1321 1265 1337
rect 1327 1703 1361 1719
rect 1327 1321 1361 1337
rect 1423 1703 1457 1719
rect 1423 1321 1457 1337
rect 1519 1703 1553 1719
rect 1519 1321 1553 1337
rect 1615 1703 1649 1719
rect 1615 1321 1649 1337
rect 1711 1703 1745 1719
rect 1711 1321 1745 1337
rect 1807 1703 1841 1719
rect 1807 1321 1841 1337
rect 1903 1703 1937 1719
rect 1903 1321 1937 1337
rect -1809 1253 -1793 1287
rect -1759 1253 -1743 1287
rect -1617 1253 -1601 1287
rect -1567 1253 -1551 1287
rect -1425 1253 -1409 1287
rect -1375 1253 -1359 1287
rect -1233 1253 -1217 1287
rect -1183 1253 -1167 1287
rect -1041 1253 -1025 1287
rect -991 1253 -975 1287
rect -849 1253 -833 1287
rect -799 1253 -783 1287
rect -657 1253 -641 1287
rect -607 1253 -591 1287
rect -465 1253 -449 1287
rect -415 1253 -399 1287
rect -273 1253 -257 1287
rect -223 1253 -207 1287
rect -81 1253 -65 1287
rect -31 1253 -15 1287
rect 111 1253 127 1287
rect 161 1253 177 1287
rect 303 1253 319 1287
rect 353 1253 369 1287
rect 495 1253 511 1287
rect 545 1253 561 1287
rect 687 1253 703 1287
rect 737 1253 753 1287
rect 879 1253 895 1287
rect 929 1253 945 1287
rect 1071 1253 1087 1287
rect 1121 1253 1137 1287
rect 1263 1253 1279 1287
rect 1313 1253 1329 1287
rect 1455 1253 1471 1287
rect 1505 1253 1521 1287
rect 1647 1253 1663 1287
rect 1697 1253 1713 1287
rect 1839 1253 1855 1287
rect 1889 1253 1905 1287
rect -1809 1145 -1793 1179
rect -1759 1145 -1743 1179
rect -1617 1145 -1601 1179
rect -1567 1145 -1551 1179
rect -1425 1145 -1409 1179
rect -1375 1145 -1359 1179
rect -1233 1145 -1217 1179
rect -1183 1145 -1167 1179
rect -1041 1145 -1025 1179
rect -991 1145 -975 1179
rect -849 1145 -833 1179
rect -799 1145 -783 1179
rect -657 1145 -641 1179
rect -607 1145 -591 1179
rect -465 1145 -449 1179
rect -415 1145 -399 1179
rect -273 1145 -257 1179
rect -223 1145 -207 1179
rect -81 1145 -65 1179
rect -31 1145 -15 1179
rect 111 1145 127 1179
rect 161 1145 177 1179
rect 303 1145 319 1179
rect 353 1145 369 1179
rect 495 1145 511 1179
rect 545 1145 561 1179
rect 687 1145 703 1179
rect 737 1145 753 1179
rect 879 1145 895 1179
rect 929 1145 945 1179
rect 1071 1145 1087 1179
rect 1121 1145 1137 1179
rect 1263 1145 1279 1179
rect 1313 1145 1329 1179
rect 1455 1145 1471 1179
rect 1505 1145 1521 1179
rect 1647 1145 1663 1179
rect 1697 1145 1713 1179
rect 1839 1145 1855 1179
rect 1889 1145 1905 1179
rect -1937 1095 -1903 1111
rect -1937 713 -1903 729
rect -1841 1095 -1807 1111
rect -1841 713 -1807 729
rect -1745 1095 -1711 1111
rect -1745 713 -1711 729
rect -1649 1095 -1615 1111
rect -1649 713 -1615 729
rect -1553 1095 -1519 1111
rect -1553 713 -1519 729
rect -1457 1095 -1423 1111
rect -1457 713 -1423 729
rect -1361 1095 -1327 1111
rect -1361 713 -1327 729
rect -1265 1095 -1231 1111
rect -1265 713 -1231 729
rect -1169 1095 -1135 1111
rect -1169 713 -1135 729
rect -1073 1095 -1039 1111
rect -1073 713 -1039 729
rect -977 1095 -943 1111
rect -977 713 -943 729
rect -881 1095 -847 1111
rect -881 713 -847 729
rect -785 1095 -751 1111
rect -785 713 -751 729
rect -689 1095 -655 1111
rect -689 713 -655 729
rect -593 1095 -559 1111
rect -593 713 -559 729
rect -497 1095 -463 1111
rect -497 713 -463 729
rect -401 1095 -367 1111
rect -401 713 -367 729
rect -305 1095 -271 1111
rect -305 713 -271 729
rect -209 1095 -175 1111
rect -209 713 -175 729
rect -113 1095 -79 1111
rect -113 713 -79 729
rect -17 1095 17 1111
rect -17 713 17 729
rect 79 1095 113 1111
rect 79 713 113 729
rect 175 1095 209 1111
rect 175 713 209 729
rect 271 1095 305 1111
rect 271 713 305 729
rect 367 1095 401 1111
rect 367 713 401 729
rect 463 1095 497 1111
rect 463 713 497 729
rect 559 1095 593 1111
rect 559 713 593 729
rect 655 1095 689 1111
rect 655 713 689 729
rect 751 1095 785 1111
rect 751 713 785 729
rect 847 1095 881 1111
rect 847 713 881 729
rect 943 1095 977 1111
rect 943 713 977 729
rect 1039 1095 1073 1111
rect 1039 713 1073 729
rect 1135 1095 1169 1111
rect 1135 713 1169 729
rect 1231 1095 1265 1111
rect 1231 713 1265 729
rect 1327 1095 1361 1111
rect 1327 713 1361 729
rect 1423 1095 1457 1111
rect 1423 713 1457 729
rect 1519 1095 1553 1111
rect 1519 713 1553 729
rect 1615 1095 1649 1111
rect 1615 713 1649 729
rect 1711 1095 1745 1111
rect 1711 713 1745 729
rect 1807 1095 1841 1111
rect 1807 713 1841 729
rect 1903 1095 1937 1111
rect 1903 713 1937 729
rect -1905 645 -1889 679
rect -1855 645 -1839 679
rect -1713 645 -1697 679
rect -1663 645 -1647 679
rect -1521 645 -1505 679
rect -1471 645 -1455 679
rect -1329 645 -1313 679
rect -1279 645 -1263 679
rect -1137 645 -1121 679
rect -1087 645 -1071 679
rect -945 645 -929 679
rect -895 645 -879 679
rect -753 645 -737 679
rect -703 645 -687 679
rect -561 645 -545 679
rect -511 645 -495 679
rect -369 645 -353 679
rect -319 645 -303 679
rect -177 645 -161 679
rect -127 645 -111 679
rect 15 645 31 679
rect 65 645 81 679
rect 207 645 223 679
rect 257 645 273 679
rect 399 645 415 679
rect 449 645 465 679
rect 591 645 607 679
rect 641 645 657 679
rect 783 645 799 679
rect 833 645 849 679
rect 975 645 991 679
rect 1025 645 1041 679
rect 1167 645 1183 679
rect 1217 645 1233 679
rect 1359 645 1375 679
rect 1409 645 1425 679
rect 1551 645 1567 679
rect 1601 645 1617 679
rect 1743 645 1759 679
rect 1793 645 1809 679
rect -1905 537 -1889 571
rect -1855 537 -1839 571
rect -1713 537 -1697 571
rect -1663 537 -1647 571
rect -1521 537 -1505 571
rect -1471 537 -1455 571
rect -1329 537 -1313 571
rect -1279 537 -1263 571
rect -1137 537 -1121 571
rect -1087 537 -1071 571
rect -945 537 -929 571
rect -895 537 -879 571
rect -753 537 -737 571
rect -703 537 -687 571
rect -561 537 -545 571
rect -511 537 -495 571
rect -369 537 -353 571
rect -319 537 -303 571
rect -177 537 -161 571
rect -127 537 -111 571
rect 15 537 31 571
rect 65 537 81 571
rect 207 537 223 571
rect 257 537 273 571
rect 399 537 415 571
rect 449 537 465 571
rect 591 537 607 571
rect 641 537 657 571
rect 783 537 799 571
rect 833 537 849 571
rect 975 537 991 571
rect 1025 537 1041 571
rect 1167 537 1183 571
rect 1217 537 1233 571
rect 1359 537 1375 571
rect 1409 537 1425 571
rect 1551 537 1567 571
rect 1601 537 1617 571
rect 1743 537 1759 571
rect 1793 537 1809 571
rect -1937 487 -1903 503
rect -1937 105 -1903 121
rect -1841 487 -1807 503
rect -1841 105 -1807 121
rect -1745 487 -1711 503
rect -1745 105 -1711 121
rect -1649 487 -1615 503
rect -1649 105 -1615 121
rect -1553 487 -1519 503
rect -1553 105 -1519 121
rect -1457 487 -1423 503
rect -1457 105 -1423 121
rect -1361 487 -1327 503
rect -1361 105 -1327 121
rect -1265 487 -1231 503
rect -1265 105 -1231 121
rect -1169 487 -1135 503
rect -1169 105 -1135 121
rect -1073 487 -1039 503
rect -1073 105 -1039 121
rect -977 487 -943 503
rect -977 105 -943 121
rect -881 487 -847 503
rect -881 105 -847 121
rect -785 487 -751 503
rect -785 105 -751 121
rect -689 487 -655 503
rect -689 105 -655 121
rect -593 487 -559 503
rect -593 105 -559 121
rect -497 487 -463 503
rect -497 105 -463 121
rect -401 487 -367 503
rect -401 105 -367 121
rect -305 487 -271 503
rect -305 105 -271 121
rect -209 487 -175 503
rect -209 105 -175 121
rect -113 487 -79 503
rect -113 105 -79 121
rect -17 487 17 503
rect -17 105 17 121
rect 79 487 113 503
rect 79 105 113 121
rect 175 487 209 503
rect 175 105 209 121
rect 271 487 305 503
rect 271 105 305 121
rect 367 487 401 503
rect 367 105 401 121
rect 463 487 497 503
rect 463 105 497 121
rect 559 487 593 503
rect 559 105 593 121
rect 655 487 689 503
rect 655 105 689 121
rect 751 487 785 503
rect 751 105 785 121
rect 847 487 881 503
rect 847 105 881 121
rect 943 487 977 503
rect 943 105 977 121
rect 1039 487 1073 503
rect 1039 105 1073 121
rect 1135 487 1169 503
rect 1135 105 1169 121
rect 1231 487 1265 503
rect 1231 105 1265 121
rect 1327 487 1361 503
rect 1327 105 1361 121
rect 1423 487 1457 503
rect 1423 105 1457 121
rect 1519 487 1553 503
rect 1519 105 1553 121
rect 1615 487 1649 503
rect 1615 105 1649 121
rect 1711 487 1745 503
rect 1711 105 1745 121
rect 1807 487 1841 503
rect 1807 105 1841 121
rect 1903 487 1937 503
rect 1903 105 1937 121
rect -1809 37 -1793 71
rect -1759 37 -1743 71
rect -1617 37 -1601 71
rect -1567 37 -1551 71
rect -1425 37 -1409 71
rect -1375 37 -1359 71
rect -1233 37 -1217 71
rect -1183 37 -1167 71
rect -1041 37 -1025 71
rect -991 37 -975 71
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect 1071 37 1087 71
rect 1121 37 1137 71
rect 1263 37 1279 71
rect 1313 37 1329 71
rect 1455 37 1471 71
rect 1505 37 1521 71
rect 1647 37 1663 71
rect 1697 37 1713 71
rect 1839 37 1855 71
rect 1889 37 1905 71
rect -1809 -71 -1793 -37
rect -1759 -71 -1743 -37
rect -1617 -71 -1601 -37
rect -1567 -71 -1551 -37
rect -1425 -71 -1409 -37
rect -1375 -71 -1359 -37
rect -1233 -71 -1217 -37
rect -1183 -71 -1167 -37
rect -1041 -71 -1025 -37
rect -991 -71 -975 -37
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 1071 -71 1087 -37
rect 1121 -71 1137 -37
rect 1263 -71 1279 -37
rect 1313 -71 1329 -37
rect 1455 -71 1471 -37
rect 1505 -71 1521 -37
rect 1647 -71 1663 -37
rect 1697 -71 1713 -37
rect 1839 -71 1855 -37
rect 1889 -71 1905 -37
rect -1937 -121 -1903 -105
rect -1937 -503 -1903 -487
rect -1841 -121 -1807 -105
rect -1841 -503 -1807 -487
rect -1745 -121 -1711 -105
rect -1745 -503 -1711 -487
rect -1649 -121 -1615 -105
rect -1649 -503 -1615 -487
rect -1553 -121 -1519 -105
rect -1553 -503 -1519 -487
rect -1457 -121 -1423 -105
rect -1457 -503 -1423 -487
rect -1361 -121 -1327 -105
rect -1361 -503 -1327 -487
rect -1265 -121 -1231 -105
rect -1265 -503 -1231 -487
rect -1169 -121 -1135 -105
rect -1169 -503 -1135 -487
rect -1073 -121 -1039 -105
rect -1073 -503 -1039 -487
rect -977 -121 -943 -105
rect -977 -503 -943 -487
rect -881 -121 -847 -105
rect -881 -503 -847 -487
rect -785 -121 -751 -105
rect -785 -503 -751 -487
rect -689 -121 -655 -105
rect -689 -503 -655 -487
rect -593 -121 -559 -105
rect -593 -503 -559 -487
rect -497 -121 -463 -105
rect -497 -503 -463 -487
rect -401 -121 -367 -105
rect -401 -503 -367 -487
rect -305 -121 -271 -105
rect -305 -503 -271 -487
rect -209 -121 -175 -105
rect -209 -503 -175 -487
rect -113 -121 -79 -105
rect -113 -503 -79 -487
rect -17 -121 17 -105
rect -17 -503 17 -487
rect 79 -121 113 -105
rect 79 -503 113 -487
rect 175 -121 209 -105
rect 175 -503 209 -487
rect 271 -121 305 -105
rect 271 -503 305 -487
rect 367 -121 401 -105
rect 367 -503 401 -487
rect 463 -121 497 -105
rect 463 -503 497 -487
rect 559 -121 593 -105
rect 559 -503 593 -487
rect 655 -121 689 -105
rect 655 -503 689 -487
rect 751 -121 785 -105
rect 751 -503 785 -487
rect 847 -121 881 -105
rect 847 -503 881 -487
rect 943 -121 977 -105
rect 943 -503 977 -487
rect 1039 -121 1073 -105
rect 1039 -503 1073 -487
rect 1135 -121 1169 -105
rect 1135 -503 1169 -487
rect 1231 -121 1265 -105
rect 1231 -503 1265 -487
rect 1327 -121 1361 -105
rect 1327 -503 1361 -487
rect 1423 -121 1457 -105
rect 1423 -503 1457 -487
rect 1519 -121 1553 -105
rect 1519 -503 1553 -487
rect 1615 -121 1649 -105
rect 1615 -503 1649 -487
rect 1711 -121 1745 -105
rect 1711 -503 1745 -487
rect 1807 -121 1841 -105
rect 1807 -503 1841 -487
rect 1903 -121 1937 -105
rect 1903 -503 1937 -487
rect -1905 -571 -1889 -537
rect -1855 -571 -1839 -537
rect -1713 -571 -1697 -537
rect -1663 -571 -1647 -537
rect -1521 -571 -1505 -537
rect -1471 -571 -1455 -537
rect -1329 -571 -1313 -537
rect -1279 -571 -1263 -537
rect -1137 -571 -1121 -537
rect -1087 -571 -1071 -537
rect -945 -571 -929 -537
rect -895 -571 -879 -537
rect -753 -571 -737 -537
rect -703 -571 -687 -537
rect -561 -571 -545 -537
rect -511 -571 -495 -537
rect -369 -571 -353 -537
rect -319 -571 -303 -537
rect -177 -571 -161 -537
rect -127 -571 -111 -537
rect 15 -571 31 -537
rect 65 -571 81 -537
rect 207 -571 223 -537
rect 257 -571 273 -537
rect 399 -571 415 -537
rect 449 -571 465 -537
rect 591 -571 607 -537
rect 641 -571 657 -537
rect 783 -571 799 -537
rect 833 -571 849 -537
rect 975 -571 991 -537
rect 1025 -571 1041 -537
rect 1167 -571 1183 -537
rect 1217 -571 1233 -537
rect 1359 -571 1375 -537
rect 1409 -571 1425 -537
rect 1551 -571 1567 -537
rect 1601 -571 1617 -537
rect 1743 -571 1759 -537
rect 1793 -571 1809 -537
rect -1905 -679 -1889 -645
rect -1855 -679 -1839 -645
rect -1713 -679 -1697 -645
rect -1663 -679 -1647 -645
rect -1521 -679 -1505 -645
rect -1471 -679 -1455 -645
rect -1329 -679 -1313 -645
rect -1279 -679 -1263 -645
rect -1137 -679 -1121 -645
rect -1087 -679 -1071 -645
rect -945 -679 -929 -645
rect -895 -679 -879 -645
rect -753 -679 -737 -645
rect -703 -679 -687 -645
rect -561 -679 -545 -645
rect -511 -679 -495 -645
rect -369 -679 -353 -645
rect -319 -679 -303 -645
rect -177 -679 -161 -645
rect -127 -679 -111 -645
rect 15 -679 31 -645
rect 65 -679 81 -645
rect 207 -679 223 -645
rect 257 -679 273 -645
rect 399 -679 415 -645
rect 449 -679 465 -645
rect 591 -679 607 -645
rect 641 -679 657 -645
rect 783 -679 799 -645
rect 833 -679 849 -645
rect 975 -679 991 -645
rect 1025 -679 1041 -645
rect 1167 -679 1183 -645
rect 1217 -679 1233 -645
rect 1359 -679 1375 -645
rect 1409 -679 1425 -645
rect 1551 -679 1567 -645
rect 1601 -679 1617 -645
rect 1743 -679 1759 -645
rect 1793 -679 1809 -645
rect -1937 -729 -1903 -713
rect -1937 -1111 -1903 -1095
rect -1841 -729 -1807 -713
rect -1841 -1111 -1807 -1095
rect -1745 -729 -1711 -713
rect -1745 -1111 -1711 -1095
rect -1649 -729 -1615 -713
rect -1649 -1111 -1615 -1095
rect -1553 -729 -1519 -713
rect -1553 -1111 -1519 -1095
rect -1457 -729 -1423 -713
rect -1457 -1111 -1423 -1095
rect -1361 -729 -1327 -713
rect -1361 -1111 -1327 -1095
rect -1265 -729 -1231 -713
rect -1265 -1111 -1231 -1095
rect -1169 -729 -1135 -713
rect -1169 -1111 -1135 -1095
rect -1073 -729 -1039 -713
rect -1073 -1111 -1039 -1095
rect -977 -729 -943 -713
rect -977 -1111 -943 -1095
rect -881 -729 -847 -713
rect -881 -1111 -847 -1095
rect -785 -729 -751 -713
rect -785 -1111 -751 -1095
rect -689 -729 -655 -713
rect -689 -1111 -655 -1095
rect -593 -729 -559 -713
rect -593 -1111 -559 -1095
rect -497 -729 -463 -713
rect -497 -1111 -463 -1095
rect -401 -729 -367 -713
rect -401 -1111 -367 -1095
rect -305 -729 -271 -713
rect -305 -1111 -271 -1095
rect -209 -729 -175 -713
rect -209 -1111 -175 -1095
rect -113 -729 -79 -713
rect -113 -1111 -79 -1095
rect -17 -729 17 -713
rect -17 -1111 17 -1095
rect 79 -729 113 -713
rect 79 -1111 113 -1095
rect 175 -729 209 -713
rect 175 -1111 209 -1095
rect 271 -729 305 -713
rect 271 -1111 305 -1095
rect 367 -729 401 -713
rect 367 -1111 401 -1095
rect 463 -729 497 -713
rect 463 -1111 497 -1095
rect 559 -729 593 -713
rect 559 -1111 593 -1095
rect 655 -729 689 -713
rect 655 -1111 689 -1095
rect 751 -729 785 -713
rect 751 -1111 785 -1095
rect 847 -729 881 -713
rect 847 -1111 881 -1095
rect 943 -729 977 -713
rect 943 -1111 977 -1095
rect 1039 -729 1073 -713
rect 1039 -1111 1073 -1095
rect 1135 -729 1169 -713
rect 1135 -1111 1169 -1095
rect 1231 -729 1265 -713
rect 1231 -1111 1265 -1095
rect 1327 -729 1361 -713
rect 1327 -1111 1361 -1095
rect 1423 -729 1457 -713
rect 1423 -1111 1457 -1095
rect 1519 -729 1553 -713
rect 1519 -1111 1553 -1095
rect 1615 -729 1649 -713
rect 1615 -1111 1649 -1095
rect 1711 -729 1745 -713
rect 1711 -1111 1745 -1095
rect 1807 -729 1841 -713
rect 1807 -1111 1841 -1095
rect 1903 -729 1937 -713
rect 1903 -1111 1937 -1095
rect -1809 -1179 -1793 -1145
rect -1759 -1179 -1743 -1145
rect -1617 -1179 -1601 -1145
rect -1567 -1179 -1551 -1145
rect -1425 -1179 -1409 -1145
rect -1375 -1179 -1359 -1145
rect -1233 -1179 -1217 -1145
rect -1183 -1179 -1167 -1145
rect -1041 -1179 -1025 -1145
rect -991 -1179 -975 -1145
rect -849 -1179 -833 -1145
rect -799 -1179 -783 -1145
rect -657 -1179 -641 -1145
rect -607 -1179 -591 -1145
rect -465 -1179 -449 -1145
rect -415 -1179 -399 -1145
rect -273 -1179 -257 -1145
rect -223 -1179 -207 -1145
rect -81 -1179 -65 -1145
rect -31 -1179 -15 -1145
rect 111 -1179 127 -1145
rect 161 -1179 177 -1145
rect 303 -1179 319 -1145
rect 353 -1179 369 -1145
rect 495 -1179 511 -1145
rect 545 -1179 561 -1145
rect 687 -1179 703 -1145
rect 737 -1179 753 -1145
rect 879 -1179 895 -1145
rect 929 -1179 945 -1145
rect 1071 -1179 1087 -1145
rect 1121 -1179 1137 -1145
rect 1263 -1179 1279 -1145
rect 1313 -1179 1329 -1145
rect 1455 -1179 1471 -1145
rect 1505 -1179 1521 -1145
rect 1647 -1179 1663 -1145
rect 1697 -1179 1713 -1145
rect 1839 -1179 1855 -1145
rect 1889 -1179 1905 -1145
rect -1809 -1287 -1793 -1253
rect -1759 -1287 -1743 -1253
rect -1617 -1287 -1601 -1253
rect -1567 -1287 -1551 -1253
rect -1425 -1287 -1409 -1253
rect -1375 -1287 -1359 -1253
rect -1233 -1287 -1217 -1253
rect -1183 -1287 -1167 -1253
rect -1041 -1287 -1025 -1253
rect -991 -1287 -975 -1253
rect -849 -1287 -833 -1253
rect -799 -1287 -783 -1253
rect -657 -1287 -641 -1253
rect -607 -1287 -591 -1253
rect -465 -1287 -449 -1253
rect -415 -1287 -399 -1253
rect -273 -1287 -257 -1253
rect -223 -1287 -207 -1253
rect -81 -1287 -65 -1253
rect -31 -1287 -15 -1253
rect 111 -1287 127 -1253
rect 161 -1287 177 -1253
rect 303 -1287 319 -1253
rect 353 -1287 369 -1253
rect 495 -1287 511 -1253
rect 545 -1287 561 -1253
rect 687 -1287 703 -1253
rect 737 -1287 753 -1253
rect 879 -1287 895 -1253
rect 929 -1287 945 -1253
rect 1071 -1287 1087 -1253
rect 1121 -1287 1137 -1253
rect 1263 -1287 1279 -1253
rect 1313 -1287 1329 -1253
rect 1455 -1287 1471 -1253
rect 1505 -1287 1521 -1253
rect 1647 -1287 1663 -1253
rect 1697 -1287 1713 -1253
rect 1839 -1287 1855 -1253
rect 1889 -1287 1905 -1253
rect -1937 -1337 -1903 -1321
rect -1937 -1719 -1903 -1703
rect -1841 -1337 -1807 -1321
rect -1841 -1719 -1807 -1703
rect -1745 -1337 -1711 -1321
rect -1745 -1719 -1711 -1703
rect -1649 -1337 -1615 -1321
rect -1649 -1719 -1615 -1703
rect -1553 -1337 -1519 -1321
rect -1553 -1719 -1519 -1703
rect -1457 -1337 -1423 -1321
rect -1457 -1719 -1423 -1703
rect -1361 -1337 -1327 -1321
rect -1361 -1719 -1327 -1703
rect -1265 -1337 -1231 -1321
rect -1265 -1719 -1231 -1703
rect -1169 -1337 -1135 -1321
rect -1169 -1719 -1135 -1703
rect -1073 -1337 -1039 -1321
rect -1073 -1719 -1039 -1703
rect -977 -1337 -943 -1321
rect -977 -1719 -943 -1703
rect -881 -1337 -847 -1321
rect -881 -1719 -847 -1703
rect -785 -1337 -751 -1321
rect -785 -1719 -751 -1703
rect -689 -1337 -655 -1321
rect -689 -1719 -655 -1703
rect -593 -1337 -559 -1321
rect -593 -1719 -559 -1703
rect -497 -1337 -463 -1321
rect -497 -1719 -463 -1703
rect -401 -1337 -367 -1321
rect -401 -1719 -367 -1703
rect -305 -1337 -271 -1321
rect -305 -1719 -271 -1703
rect -209 -1337 -175 -1321
rect -209 -1719 -175 -1703
rect -113 -1337 -79 -1321
rect -113 -1719 -79 -1703
rect -17 -1337 17 -1321
rect -17 -1719 17 -1703
rect 79 -1337 113 -1321
rect 79 -1719 113 -1703
rect 175 -1337 209 -1321
rect 175 -1719 209 -1703
rect 271 -1337 305 -1321
rect 271 -1719 305 -1703
rect 367 -1337 401 -1321
rect 367 -1719 401 -1703
rect 463 -1337 497 -1321
rect 463 -1719 497 -1703
rect 559 -1337 593 -1321
rect 559 -1719 593 -1703
rect 655 -1337 689 -1321
rect 655 -1719 689 -1703
rect 751 -1337 785 -1321
rect 751 -1719 785 -1703
rect 847 -1337 881 -1321
rect 847 -1719 881 -1703
rect 943 -1337 977 -1321
rect 943 -1719 977 -1703
rect 1039 -1337 1073 -1321
rect 1039 -1719 1073 -1703
rect 1135 -1337 1169 -1321
rect 1135 -1719 1169 -1703
rect 1231 -1337 1265 -1321
rect 1231 -1719 1265 -1703
rect 1327 -1337 1361 -1321
rect 1327 -1719 1361 -1703
rect 1423 -1337 1457 -1321
rect 1423 -1719 1457 -1703
rect 1519 -1337 1553 -1321
rect 1519 -1719 1553 -1703
rect 1615 -1337 1649 -1321
rect 1615 -1719 1649 -1703
rect 1711 -1337 1745 -1321
rect 1711 -1719 1745 -1703
rect 1807 -1337 1841 -1321
rect 1807 -1719 1841 -1703
rect 1903 -1337 1937 -1321
rect 1903 -1719 1937 -1703
rect -1905 -1787 -1889 -1753
rect -1855 -1787 -1839 -1753
rect -1713 -1787 -1697 -1753
rect -1663 -1787 -1647 -1753
rect -1521 -1787 -1505 -1753
rect -1471 -1787 -1455 -1753
rect -1329 -1787 -1313 -1753
rect -1279 -1787 -1263 -1753
rect -1137 -1787 -1121 -1753
rect -1087 -1787 -1071 -1753
rect -945 -1787 -929 -1753
rect -895 -1787 -879 -1753
rect -753 -1787 -737 -1753
rect -703 -1787 -687 -1753
rect -561 -1787 -545 -1753
rect -511 -1787 -495 -1753
rect -369 -1787 -353 -1753
rect -319 -1787 -303 -1753
rect -177 -1787 -161 -1753
rect -127 -1787 -111 -1753
rect 15 -1787 31 -1753
rect 65 -1787 81 -1753
rect 207 -1787 223 -1753
rect 257 -1787 273 -1753
rect 399 -1787 415 -1753
rect 449 -1787 465 -1753
rect 591 -1787 607 -1753
rect 641 -1787 657 -1753
rect 783 -1787 799 -1753
rect 833 -1787 849 -1753
rect 975 -1787 991 -1753
rect 1025 -1787 1041 -1753
rect 1167 -1787 1183 -1753
rect 1217 -1787 1233 -1753
rect 1359 -1787 1375 -1753
rect 1409 -1787 1425 -1753
rect 1551 -1787 1567 -1753
rect 1601 -1787 1617 -1753
rect 1743 -1787 1759 -1753
rect 1793 -1787 1809 -1753
rect -2051 -1855 -2017 -1793
rect 2017 -1855 2051 -1793
rect -2051 -1889 -1955 -1855
rect 1955 -1889 2051 -1855
<< viali >>
rect -1889 1753 -1855 1787
rect -1697 1753 -1663 1787
rect -1505 1753 -1471 1787
rect -1313 1753 -1279 1787
rect -1121 1753 -1087 1787
rect -929 1753 -895 1787
rect -737 1753 -703 1787
rect -545 1753 -511 1787
rect -353 1753 -319 1787
rect -161 1753 -127 1787
rect 31 1753 65 1787
rect 223 1753 257 1787
rect 415 1753 449 1787
rect 607 1753 641 1787
rect 799 1753 833 1787
rect 991 1753 1025 1787
rect 1183 1753 1217 1787
rect 1375 1753 1409 1787
rect 1567 1753 1601 1787
rect 1759 1753 1793 1787
rect -1937 1337 -1903 1703
rect -1841 1337 -1807 1703
rect -1745 1337 -1711 1703
rect -1649 1337 -1615 1703
rect -1553 1337 -1519 1703
rect -1457 1337 -1423 1703
rect -1361 1337 -1327 1703
rect -1265 1337 -1231 1703
rect -1169 1337 -1135 1703
rect -1073 1337 -1039 1703
rect -977 1337 -943 1703
rect -881 1337 -847 1703
rect -785 1337 -751 1703
rect -689 1337 -655 1703
rect -593 1337 -559 1703
rect -497 1337 -463 1703
rect -401 1337 -367 1703
rect -305 1337 -271 1703
rect -209 1337 -175 1703
rect -113 1337 -79 1703
rect -17 1337 17 1703
rect 79 1337 113 1703
rect 175 1337 209 1703
rect 271 1337 305 1703
rect 367 1337 401 1703
rect 463 1337 497 1703
rect 559 1337 593 1703
rect 655 1337 689 1703
rect 751 1337 785 1703
rect 847 1337 881 1703
rect 943 1337 977 1703
rect 1039 1337 1073 1703
rect 1135 1337 1169 1703
rect 1231 1337 1265 1703
rect 1327 1337 1361 1703
rect 1423 1337 1457 1703
rect 1519 1337 1553 1703
rect 1615 1337 1649 1703
rect 1711 1337 1745 1703
rect 1807 1337 1841 1703
rect 1903 1337 1937 1703
rect -1793 1253 -1759 1287
rect -1601 1253 -1567 1287
rect -1409 1253 -1375 1287
rect -1217 1253 -1183 1287
rect -1025 1253 -991 1287
rect -833 1253 -799 1287
rect -641 1253 -607 1287
rect -449 1253 -415 1287
rect -257 1253 -223 1287
rect -65 1253 -31 1287
rect 127 1253 161 1287
rect 319 1253 353 1287
rect 511 1253 545 1287
rect 703 1253 737 1287
rect 895 1253 929 1287
rect 1087 1253 1121 1287
rect 1279 1253 1313 1287
rect 1471 1253 1505 1287
rect 1663 1253 1697 1287
rect 1855 1253 1889 1287
rect -1793 1145 -1759 1179
rect -1601 1145 -1567 1179
rect -1409 1145 -1375 1179
rect -1217 1145 -1183 1179
rect -1025 1145 -991 1179
rect -833 1145 -799 1179
rect -641 1145 -607 1179
rect -449 1145 -415 1179
rect -257 1145 -223 1179
rect -65 1145 -31 1179
rect 127 1145 161 1179
rect 319 1145 353 1179
rect 511 1145 545 1179
rect 703 1145 737 1179
rect 895 1145 929 1179
rect 1087 1145 1121 1179
rect 1279 1145 1313 1179
rect 1471 1145 1505 1179
rect 1663 1145 1697 1179
rect 1855 1145 1889 1179
rect -1937 729 -1903 1095
rect -1841 729 -1807 1095
rect -1745 729 -1711 1095
rect -1649 729 -1615 1095
rect -1553 729 -1519 1095
rect -1457 729 -1423 1095
rect -1361 729 -1327 1095
rect -1265 729 -1231 1095
rect -1169 729 -1135 1095
rect -1073 729 -1039 1095
rect -977 729 -943 1095
rect -881 729 -847 1095
rect -785 729 -751 1095
rect -689 729 -655 1095
rect -593 729 -559 1095
rect -497 729 -463 1095
rect -401 729 -367 1095
rect -305 729 -271 1095
rect -209 729 -175 1095
rect -113 729 -79 1095
rect -17 729 17 1095
rect 79 729 113 1095
rect 175 729 209 1095
rect 271 729 305 1095
rect 367 729 401 1095
rect 463 729 497 1095
rect 559 729 593 1095
rect 655 729 689 1095
rect 751 729 785 1095
rect 847 729 881 1095
rect 943 729 977 1095
rect 1039 729 1073 1095
rect 1135 729 1169 1095
rect 1231 729 1265 1095
rect 1327 729 1361 1095
rect 1423 729 1457 1095
rect 1519 729 1553 1095
rect 1615 729 1649 1095
rect 1711 729 1745 1095
rect 1807 729 1841 1095
rect 1903 729 1937 1095
rect -1889 645 -1855 679
rect -1697 645 -1663 679
rect -1505 645 -1471 679
rect -1313 645 -1279 679
rect -1121 645 -1087 679
rect -929 645 -895 679
rect -737 645 -703 679
rect -545 645 -511 679
rect -353 645 -319 679
rect -161 645 -127 679
rect 31 645 65 679
rect 223 645 257 679
rect 415 645 449 679
rect 607 645 641 679
rect 799 645 833 679
rect 991 645 1025 679
rect 1183 645 1217 679
rect 1375 645 1409 679
rect 1567 645 1601 679
rect 1759 645 1793 679
rect -1889 537 -1855 571
rect -1697 537 -1663 571
rect -1505 537 -1471 571
rect -1313 537 -1279 571
rect -1121 537 -1087 571
rect -929 537 -895 571
rect -737 537 -703 571
rect -545 537 -511 571
rect -353 537 -319 571
rect -161 537 -127 571
rect 31 537 65 571
rect 223 537 257 571
rect 415 537 449 571
rect 607 537 641 571
rect 799 537 833 571
rect 991 537 1025 571
rect 1183 537 1217 571
rect 1375 537 1409 571
rect 1567 537 1601 571
rect 1759 537 1793 571
rect -1937 121 -1903 487
rect -1841 121 -1807 487
rect -1745 121 -1711 487
rect -1649 121 -1615 487
rect -1553 121 -1519 487
rect -1457 121 -1423 487
rect -1361 121 -1327 487
rect -1265 121 -1231 487
rect -1169 121 -1135 487
rect -1073 121 -1039 487
rect -977 121 -943 487
rect -881 121 -847 487
rect -785 121 -751 487
rect -689 121 -655 487
rect -593 121 -559 487
rect -497 121 -463 487
rect -401 121 -367 487
rect -305 121 -271 487
rect -209 121 -175 487
rect -113 121 -79 487
rect -17 121 17 487
rect 79 121 113 487
rect 175 121 209 487
rect 271 121 305 487
rect 367 121 401 487
rect 463 121 497 487
rect 559 121 593 487
rect 655 121 689 487
rect 751 121 785 487
rect 847 121 881 487
rect 943 121 977 487
rect 1039 121 1073 487
rect 1135 121 1169 487
rect 1231 121 1265 487
rect 1327 121 1361 487
rect 1423 121 1457 487
rect 1519 121 1553 487
rect 1615 121 1649 487
rect 1711 121 1745 487
rect 1807 121 1841 487
rect 1903 121 1937 487
rect -1793 37 -1759 71
rect -1601 37 -1567 71
rect -1409 37 -1375 71
rect -1217 37 -1183 71
rect -1025 37 -991 71
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect 1087 37 1121 71
rect 1279 37 1313 71
rect 1471 37 1505 71
rect 1663 37 1697 71
rect 1855 37 1889 71
rect -1793 -71 -1759 -37
rect -1601 -71 -1567 -37
rect -1409 -71 -1375 -37
rect -1217 -71 -1183 -37
rect -1025 -71 -991 -37
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect 1087 -71 1121 -37
rect 1279 -71 1313 -37
rect 1471 -71 1505 -37
rect 1663 -71 1697 -37
rect 1855 -71 1889 -37
rect -1937 -487 -1903 -121
rect -1841 -487 -1807 -121
rect -1745 -487 -1711 -121
rect -1649 -487 -1615 -121
rect -1553 -487 -1519 -121
rect -1457 -487 -1423 -121
rect -1361 -487 -1327 -121
rect -1265 -487 -1231 -121
rect -1169 -487 -1135 -121
rect -1073 -487 -1039 -121
rect -977 -487 -943 -121
rect -881 -487 -847 -121
rect -785 -487 -751 -121
rect -689 -487 -655 -121
rect -593 -487 -559 -121
rect -497 -487 -463 -121
rect -401 -487 -367 -121
rect -305 -487 -271 -121
rect -209 -487 -175 -121
rect -113 -487 -79 -121
rect -17 -487 17 -121
rect 79 -487 113 -121
rect 175 -487 209 -121
rect 271 -487 305 -121
rect 367 -487 401 -121
rect 463 -487 497 -121
rect 559 -487 593 -121
rect 655 -487 689 -121
rect 751 -487 785 -121
rect 847 -487 881 -121
rect 943 -487 977 -121
rect 1039 -487 1073 -121
rect 1135 -487 1169 -121
rect 1231 -487 1265 -121
rect 1327 -487 1361 -121
rect 1423 -487 1457 -121
rect 1519 -487 1553 -121
rect 1615 -487 1649 -121
rect 1711 -487 1745 -121
rect 1807 -487 1841 -121
rect 1903 -487 1937 -121
rect -1889 -571 -1855 -537
rect -1697 -571 -1663 -537
rect -1505 -571 -1471 -537
rect -1313 -571 -1279 -537
rect -1121 -571 -1087 -537
rect -929 -571 -895 -537
rect -737 -571 -703 -537
rect -545 -571 -511 -537
rect -353 -571 -319 -537
rect -161 -571 -127 -537
rect 31 -571 65 -537
rect 223 -571 257 -537
rect 415 -571 449 -537
rect 607 -571 641 -537
rect 799 -571 833 -537
rect 991 -571 1025 -537
rect 1183 -571 1217 -537
rect 1375 -571 1409 -537
rect 1567 -571 1601 -537
rect 1759 -571 1793 -537
rect -1889 -679 -1855 -645
rect -1697 -679 -1663 -645
rect -1505 -679 -1471 -645
rect -1313 -679 -1279 -645
rect -1121 -679 -1087 -645
rect -929 -679 -895 -645
rect -737 -679 -703 -645
rect -545 -679 -511 -645
rect -353 -679 -319 -645
rect -161 -679 -127 -645
rect 31 -679 65 -645
rect 223 -679 257 -645
rect 415 -679 449 -645
rect 607 -679 641 -645
rect 799 -679 833 -645
rect 991 -679 1025 -645
rect 1183 -679 1217 -645
rect 1375 -679 1409 -645
rect 1567 -679 1601 -645
rect 1759 -679 1793 -645
rect -1937 -1095 -1903 -729
rect -1841 -1095 -1807 -729
rect -1745 -1095 -1711 -729
rect -1649 -1095 -1615 -729
rect -1553 -1095 -1519 -729
rect -1457 -1095 -1423 -729
rect -1361 -1095 -1327 -729
rect -1265 -1095 -1231 -729
rect -1169 -1095 -1135 -729
rect -1073 -1095 -1039 -729
rect -977 -1095 -943 -729
rect -881 -1095 -847 -729
rect -785 -1095 -751 -729
rect -689 -1095 -655 -729
rect -593 -1095 -559 -729
rect -497 -1095 -463 -729
rect -401 -1095 -367 -729
rect -305 -1095 -271 -729
rect -209 -1095 -175 -729
rect -113 -1095 -79 -729
rect -17 -1095 17 -729
rect 79 -1095 113 -729
rect 175 -1095 209 -729
rect 271 -1095 305 -729
rect 367 -1095 401 -729
rect 463 -1095 497 -729
rect 559 -1095 593 -729
rect 655 -1095 689 -729
rect 751 -1095 785 -729
rect 847 -1095 881 -729
rect 943 -1095 977 -729
rect 1039 -1095 1073 -729
rect 1135 -1095 1169 -729
rect 1231 -1095 1265 -729
rect 1327 -1095 1361 -729
rect 1423 -1095 1457 -729
rect 1519 -1095 1553 -729
rect 1615 -1095 1649 -729
rect 1711 -1095 1745 -729
rect 1807 -1095 1841 -729
rect 1903 -1095 1937 -729
rect -1793 -1179 -1759 -1145
rect -1601 -1179 -1567 -1145
rect -1409 -1179 -1375 -1145
rect -1217 -1179 -1183 -1145
rect -1025 -1179 -991 -1145
rect -833 -1179 -799 -1145
rect -641 -1179 -607 -1145
rect -449 -1179 -415 -1145
rect -257 -1179 -223 -1145
rect -65 -1179 -31 -1145
rect 127 -1179 161 -1145
rect 319 -1179 353 -1145
rect 511 -1179 545 -1145
rect 703 -1179 737 -1145
rect 895 -1179 929 -1145
rect 1087 -1179 1121 -1145
rect 1279 -1179 1313 -1145
rect 1471 -1179 1505 -1145
rect 1663 -1179 1697 -1145
rect 1855 -1179 1889 -1145
rect -1793 -1287 -1759 -1253
rect -1601 -1287 -1567 -1253
rect -1409 -1287 -1375 -1253
rect -1217 -1287 -1183 -1253
rect -1025 -1287 -991 -1253
rect -833 -1287 -799 -1253
rect -641 -1287 -607 -1253
rect -449 -1287 -415 -1253
rect -257 -1287 -223 -1253
rect -65 -1287 -31 -1253
rect 127 -1287 161 -1253
rect 319 -1287 353 -1253
rect 511 -1287 545 -1253
rect 703 -1287 737 -1253
rect 895 -1287 929 -1253
rect 1087 -1287 1121 -1253
rect 1279 -1287 1313 -1253
rect 1471 -1287 1505 -1253
rect 1663 -1287 1697 -1253
rect 1855 -1287 1889 -1253
rect -1937 -1703 -1903 -1337
rect -1841 -1703 -1807 -1337
rect -1745 -1703 -1711 -1337
rect -1649 -1703 -1615 -1337
rect -1553 -1703 -1519 -1337
rect -1457 -1703 -1423 -1337
rect -1361 -1703 -1327 -1337
rect -1265 -1703 -1231 -1337
rect -1169 -1703 -1135 -1337
rect -1073 -1703 -1039 -1337
rect -977 -1703 -943 -1337
rect -881 -1703 -847 -1337
rect -785 -1703 -751 -1337
rect -689 -1703 -655 -1337
rect -593 -1703 -559 -1337
rect -497 -1703 -463 -1337
rect -401 -1703 -367 -1337
rect -305 -1703 -271 -1337
rect -209 -1703 -175 -1337
rect -113 -1703 -79 -1337
rect -17 -1703 17 -1337
rect 79 -1703 113 -1337
rect 175 -1703 209 -1337
rect 271 -1703 305 -1337
rect 367 -1703 401 -1337
rect 463 -1703 497 -1337
rect 559 -1703 593 -1337
rect 655 -1703 689 -1337
rect 751 -1703 785 -1337
rect 847 -1703 881 -1337
rect 943 -1703 977 -1337
rect 1039 -1703 1073 -1337
rect 1135 -1703 1169 -1337
rect 1231 -1703 1265 -1337
rect 1327 -1703 1361 -1337
rect 1423 -1703 1457 -1337
rect 1519 -1703 1553 -1337
rect 1615 -1703 1649 -1337
rect 1711 -1703 1745 -1337
rect 1807 -1703 1841 -1337
rect 1903 -1703 1937 -1337
rect -1889 -1787 -1855 -1753
rect -1697 -1787 -1663 -1753
rect -1505 -1787 -1471 -1753
rect -1313 -1787 -1279 -1753
rect -1121 -1787 -1087 -1753
rect -929 -1787 -895 -1753
rect -737 -1787 -703 -1753
rect -545 -1787 -511 -1753
rect -353 -1787 -319 -1753
rect -161 -1787 -127 -1753
rect 31 -1787 65 -1753
rect 223 -1787 257 -1753
rect 415 -1787 449 -1753
rect 607 -1787 641 -1753
rect 799 -1787 833 -1753
rect 991 -1787 1025 -1753
rect 1183 -1787 1217 -1753
rect 1375 -1787 1409 -1753
rect 1567 -1787 1601 -1753
rect 1759 -1787 1793 -1753
<< metal1 >>
rect -1901 1787 -1843 1793
rect -1901 1753 -1889 1787
rect -1855 1753 -1843 1787
rect -1901 1747 -1843 1753
rect -1709 1787 -1651 1793
rect -1709 1753 -1697 1787
rect -1663 1753 -1651 1787
rect -1709 1747 -1651 1753
rect -1517 1787 -1459 1793
rect -1517 1753 -1505 1787
rect -1471 1753 -1459 1787
rect -1517 1747 -1459 1753
rect -1325 1787 -1267 1793
rect -1325 1753 -1313 1787
rect -1279 1753 -1267 1787
rect -1325 1747 -1267 1753
rect -1133 1787 -1075 1793
rect -1133 1753 -1121 1787
rect -1087 1753 -1075 1787
rect -1133 1747 -1075 1753
rect -941 1787 -883 1793
rect -941 1753 -929 1787
rect -895 1753 -883 1787
rect -941 1747 -883 1753
rect -749 1787 -691 1793
rect -749 1753 -737 1787
rect -703 1753 -691 1787
rect -749 1747 -691 1753
rect -557 1787 -499 1793
rect -557 1753 -545 1787
rect -511 1753 -499 1787
rect -557 1747 -499 1753
rect -365 1787 -307 1793
rect -365 1753 -353 1787
rect -319 1753 -307 1787
rect -365 1747 -307 1753
rect -173 1787 -115 1793
rect -173 1753 -161 1787
rect -127 1753 -115 1787
rect -173 1747 -115 1753
rect 19 1787 77 1793
rect 19 1753 31 1787
rect 65 1753 77 1787
rect 19 1747 77 1753
rect 211 1787 269 1793
rect 211 1753 223 1787
rect 257 1753 269 1787
rect 211 1747 269 1753
rect 403 1787 461 1793
rect 403 1753 415 1787
rect 449 1753 461 1787
rect 403 1747 461 1753
rect 595 1787 653 1793
rect 595 1753 607 1787
rect 641 1753 653 1787
rect 595 1747 653 1753
rect 787 1787 845 1793
rect 787 1753 799 1787
rect 833 1753 845 1787
rect 787 1747 845 1753
rect 979 1787 1037 1793
rect 979 1753 991 1787
rect 1025 1753 1037 1787
rect 979 1747 1037 1753
rect 1171 1787 1229 1793
rect 1171 1753 1183 1787
rect 1217 1753 1229 1787
rect 1171 1747 1229 1753
rect 1363 1787 1421 1793
rect 1363 1753 1375 1787
rect 1409 1753 1421 1787
rect 1363 1747 1421 1753
rect 1555 1787 1613 1793
rect 1555 1753 1567 1787
rect 1601 1753 1613 1787
rect 1555 1747 1613 1753
rect 1747 1787 1805 1793
rect 1747 1753 1759 1787
rect 1793 1753 1805 1787
rect 1747 1747 1805 1753
rect -1943 1703 -1897 1715
rect -1943 1337 -1937 1703
rect -1903 1337 -1897 1703
rect -1943 1325 -1897 1337
rect -1847 1703 -1801 1715
rect -1847 1337 -1841 1703
rect -1807 1337 -1801 1703
rect -1847 1325 -1801 1337
rect -1751 1703 -1705 1715
rect -1751 1337 -1745 1703
rect -1711 1337 -1705 1703
rect -1751 1325 -1705 1337
rect -1655 1703 -1609 1715
rect -1655 1337 -1649 1703
rect -1615 1337 -1609 1703
rect -1655 1325 -1609 1337
rect -1559 1703 -1513 1715
rect -1559 1337 -1553 1703
rect -1519 1337 -1513 1703
rect -1559 1325 -1513 1337
rect -1463 1703 -1417 1715
rect -1463 1337 -1457 1703
rect -1423 1337 -1417 1703
rect -1463 1325 -1417 1337
rect -1367 1703 -1321 1715
rect -1367 1337 -1361 1703
rect -1327 1337 -1321 1703
rect -1367 1325 -1321 1337
rect -1271 1703 -1225 1715
rect -1271 1337 -1265 1703
rect -1231 1337 -1225 1703
rect -1271 1325 -1225 1337
rect -1175 1703 -1129 1715
rect -1175 1337 -1169 1703
rect -1135 1337 -1129 1703
rect -1175 1325 -1129 1337
rect -1079 1703 -1033 1715
rect -1079 1337 -1073 1703
rect -1039 1337 -1033 1703
rect -1079 1325 -1033 1337
rect -983 1703 -937 1715
rect -983 1337 -977 1703
rect -943 1337 -937 1703
rect -983 1325 -937 1337
rect -887 1703 -841 1715
rect -887 1337 -881 1703
rect -847 1337 -841 1703
rect -887 1325 -841 1337
rect -791 1703 -745 1715
rect -791 1337 -785 1703
rect -751 1337 -745 1703
rect -791 1325 -745 1337
rect -695 1703 -649 1715
rect -695 1337 -689 1703
rect -655 1337 -649 1703
rect -695 1325 -649 1337
rect -599 1703 -553 1715
rect -599 1337 -593 1703
rect -559 1337 -553 1703
rect -599 1325 -553 1337
rect -503 1703 -457 1715
rect -503 1337 -497 1703
rect -463 1337 -457 1703
rect -503 1325 -457 1337
rect -407 1703 -361 1715
rect -407 1337 -401 1703
rect -367 1337 -361 1703
rect -407 1325 -361 1337
rect -311 1703 -265 1715
rect -311 1337 -305 1703
rect -271 1337 -265 1703
rect -311 1325 -265 1337
rect -215 1703 -169 1715
rect -215 1337 -209 1703
rect -175 1337 -169 1703
rect -215 1325 -169 1337
rect -119 1703 -73 1715
rect -119 1337 -113 1703
rect -79 1337 -73 1703
rect -119 1325 -73 1337
rect -23 1703 23 1715
rect -23 1337 -17 1703
rect 17 1337 23 1703
rect -23 1325 23 1337
rect 73 1703 119 1715
rect 73 1337 79 1703
rect 113 1337 119 1703
rect 73 1325 119 1337
rect 169 1703 215 1715
rect 169 1337 175 1703
rect 209 1337 215 1703
rect 169 1325 215 1337
rect 265 1703 311 1715
rect 265 1337 271 1703
rect 305 1337 311 1703
rect 265 1325 311 1337
rect 361 1703 407 1715
rect 361 1337 367 1703
rect 401 1337 407 1703
rect 361 1325 407 1337
rect 457 1703 503 1715
rect 457 1337 463 1703
rect 497 1337 503 1703
rect 457 1325 503 1337
rect 553 1703 599 1715
rect 553 1337 559 1703
rect 593 1337 599 1703
rect 553 1325 599 1337
rect 649 1703 695 1715
rect 649 1337 655 1703
rect 689 1337 695 1703
rect 649 1325 695 1337
rect 745 1703 791 1715
rect 745 1337 751 1703
rect 785 1337 791 1703
rect 745 1325 791 1337
rect 841 1703 887 1715
rect 841 1337 847 1703
rect 881 1337 887 1703
rect 841 1325 887 1337
rect 937 1703 983 1715
rect 937 1337 943 1703
rect 977 1337 983 1703
rect 937 1325 983 1337
rect 1033 1703 1079 1715
rect 1033 1337 1039 1703
rect 1073 1337 1079 1703
rect 1033 1325 1079 1337
rect 1129 1703 1175 1715
rect 1129 1337 1135 1703
rect 1169 1337 1175 1703
rect 1129 1325 1175 1337
rect 1225 1703 1271 1715
rect 1225 1337 1231 1703
rect 1265 1337 1271 1703
rect 1225 1325 1271 1337
rect 1321 1703 1367 1715
rect 1321 1337 1327 1703
rect 1361 1337 1367 1703
rect 1321 1325 1367 1337
rect 1417 1703 1463 1715
rect 1417 1337 1423 1703
rect 1457 1337 1463 1703
rect 1417 1325 1463 1337
rect 1513 1703 1559 1715
rect 1513 1337 1519 1703
rect 1553 1337 1559 1703
rect 1513 1325 1559 1337
rect 1609 1703 1655 1715
rect 1609 1337 1615 1703
rect 1649 1337 1655 1703
rect 1609 1325 1655 1337
rect 1705 1703 1751 1715
rect 1705 1337 1711 1703
rect 1745 1337 1751 1703
rect 1705 1325 1751 1337
rect 1801 1703 1847 1715
rect 1801 1337 1807 1703
rect 1841 1337 1847 1703
rect 1801 1325 1847 1337
rect 1897 1703 1943 1715
rect 1897 1337 1903 1703
rect 1937 1337 1943 1703
rect 1897 1325 1943 1337
rect -1805 1287 -1747 1293
rect -1805 1253 -1793 1287
rect -1759 1253 -1747 1287
rect -1805 1247 -1747 1253
rect -1613 1287 -1555 1293
rect -1613 1253 -1601 1287
rect -1567 1253 -1555 1287
rect -1613 1247 -1555 1253
rect -1421 1287 -1363 1293
rect -1421 1253 -1409 1287
rect -1375 1253 -1363 1287
rect -1421 1247 -1363 1253
rect -1229 1287 -1171 1293
rect -1229 1253 -1217 1287
rect -1183 1253 -1171 1287
rect -1229 1247 -1171 1253
rect -1037 1287 -979 1293
rect -1037 1253 -1025 1287
rect -991 1253 -979 1287
rect -1037 1247 -979 1253
rect -845 1287 -787 1293
rect -845 1253 -833 1287
rect -799 1253 -787 1287
rect -845 1247 -787 1253
rect -653 1287 -595 1293
rect -653 1253 -641 1287
rect -607 1253 -595 1287
rect -653 1247 -595 1253
rect -461 1287 -403 1293
rect -461 1253 -449 1287
rect -415 1253 -403 1287
rect -461 1247 -403 1253
rect -269 1287 -211 1293
rect -269 1253 -257 1287
rect -223 1253 -211 1287
rect -269 1247 -211 1253
rect -77 1287 -19 1293
rect -77 1253 -65 1287
rect -31 1253 -19 1287
rect -77 1247 -19 1253
rect 115 1287 173 1293
rect 115 1253 127 1287
rect 161 1253 173 1287
rect 115 1247 173 1253
rect 307 1287 365 1293
rect 307 1253 319 1287
rect 353 1253 365 1287
rect 307 1247 365 1253
rect 499 1287 557 1293
rect 499 1253 511 1287
rect 545 1253 557 1287
rect 499 1247 557 1253
rect 691 1287 749 1293
rect 691 1253 703 1287
rect 737 1253 749 1287
rect 691 1247 749 1253
rect 883 1287 941 1293
rect 883 1253 895 1287
rect 929 1253 941 1287
rect 883 1247 941 1253
rect 1075 1287 1133 1293
rect 1075 1253 1087 1287
rect 1121 1253 1133 1287
rect 1075 1247 1133 1253
rect 1267 1287 1325 1293
rect 1267 1253 1279 1287
rect 1313 1253 1325 1287
rect 1267 1247 1325 1253
rect 1459 1287 1517 1293
rect 1459 1253 1471 1287
rect 1505 1253 1517 1287
rect 1459 1247 1517 1253
rect 1651 1287 1709 1293
rect 1651 1253 1663 1287
rect 1697 1253 1709 1287
rect 1651 1247 1709 1253
rect 1843 1287 1901 1293
rect 1843 1253 1855 1287
rect 1889 1253 1901 1287
rect 1843 1247 1901 1253
rect -1805 1179 -1747 1185
rect -1805 1145 -1793 1179
rect -1759 1145 -1747 1179
rect -1805 1139 -1747 1145
rect -1613 1179 -1555 1185
rect -1613 1145 -1601 1179
rect -1567 1145 -1555 1179
rect -1613 1139 -1555 1145
rect -1421 1179 -1363 1185
rect -1421 1145 -1409 1179
rect -1375 1145 -1363 1179
rect -1421 1139 -1363 1145
rect -1229 1179 -1171 1185
rect -1229 1145 -1217 1179
rect -1183 1145 -1171 1179
rect -1229 1139 -1171 1145
rect -1037 1179 -979 1185
rect -1037 1145 -1025 1179
rect -991 1145 -979 1179
rect -1037 1139 -979 1145
rect -845 1179 -787 1185
rect -845 1145 -833 1179
rect -799 1145 -787 1179
rect -845 1139 -787 1145
rect -653 1179 -595 1185
rect -653 1145 -641 1179
rect -607 1145 -595 1179
rect -653 1139 -595 1145
rect -461 1179 -403 1185
rect -461 1145 -449 1179
rect -415 1145 -403 1179
rect -461 1139 -403 1145
rect -269 1179 -211 1185
rect -269 1145 -257 1179
rect -223 1145 -211 1179
rect -269 1139 -211 1145
rect -77 1179 -19 1185
rect -77 1145 -65 1179
rect -31 1145 -19 1179
rect -77 1139 -19 1145
rect 115 1179 173 1185
rect 115 1145 127 1179
rect 161 1145 173 1179
rect 115 1139 173 1145
rect 307 1179 365 1185
rect 307 1145 319 1179
rect 353 1145 365 1179
rect 307 1139 365 1145
rect 499 1179 557 1185
rect 499 1145 511 1179
rect 545 1145 557 1179
rect 499 1139 557 1145
rect 691 1179 749 1185
rect 691 1145 703 1179
rect 737 1145 749 1179
rect 691 1139 749 1145
rect 883 1179 941 1185
rect 883 1145 895 1179
rect 929 1145 941 1179
rect 883 1139 941 1145
rect 1075 1179 1133 1185
rect 1075 1145 1087 1179
rect 1121 1145 1133 1179
rect 1075 1139 1133 1145
rect 1267 1179 1325 1185
rect 1267 1145 1279 1179
rect 1313 1145 1325 1179
rect 1267 1139 1325 1145
rect 1459 1179 1517 1185
rect 1459 1145 1471 1179
rect 1505 1145 1517 1179
rect 1459 1139 1517 1145
rect 1651 1179 1709 1185
rect 1651 1145 1663 1179
rect 1697 1145 1709 1179
rect 1651 1139 1709 1145
rect 1843 1179 1901 1185
rect 1843 1145 1855 1179
rect 1889 1145 1901 1179
rect 1843 1139 1901 1145
rect -1943 1095 -1897 1107
rect -1943 729 -1937 1095
rect -1903 729 -1897 1095
rect -1943 717 -1897 729
rect -1847 1095 -1801 1107
rect -1847 729 -1841 1095
rect -1807 729 -1801 1095
rect -1847 717 -1801 729
rect -1751 1095 -1705 1107
rect -1751 729 -1745 1095
rect -1711 729 -1705 1095
rect -1751 717 -1705 729
rect -1655 1095 -1609 1107
rect -1655 729 -1649 1095
rect -1615 729 -1609 1095
rect -1655 717 -1609 729
rect -1559 1095 -1513 1107
rect -1559 729 -1553 1095
rect -1519 729 -1513 1095
rect -1559 717 -1513 729
rect -1463 1095 -1417 1107
rect -1463 729 -1457 1095
rect -1423 729 -1417 1095
rect -1463 717 -1417 729
rect -1367 1095 -1321 1107
rect -1367 729 -1361 1095
rect -1327 729 -1321 1095
rect -1367 717 -1321 729
rect -1271 1095 -1225 1107
rect -1271 729 -1265 1095
rect -1231 729 -1225 1095
rect -1271 717 -1225 729
rect -1175 1095 -1129 1107
rect -1175 729 -1169 1095
rect -1135 729 -1129 1095
rect -1175 717 -1129 729
rect -1079 1095 -1033 1107
rect -1079 729 -1073 1095
rect -1039 729 -1033 1095
rect -1079 717 -1033 729
rect -983 1095 -937 1107
rect -983 729 -977 1095
rect -943 729 -937 1095
rect -983 717 -937 729
rect -887 1095 -841 1107
rect -887 729 -881 1095
rect -847 729 -841 1095
rect -887 717 -841 729
rect -791 1095 -745 1107
rect -791 729 -785 1095
rect -751 729 -745 1095
rect -791 717 -745 729
rect -695 1095 -649 1107
rect -695 729 -689 1095
rect -655 729 -649 1095
rect -695 717 -649 729
rect -599 1095 -553 1107
rect -599 729 -593 1095
rect -559 729 -553 1095
rect -599 717 -553 729
rect -503 1095 -457 1107
rect -503 729 -497 1095
rect -463 729 -457 1095
rect -503 717 -457 729
rect -407 1095 -361 1107
rect -407 729 -401 1095
rect -367 729 -361 1095
rect -407 717 -361 729
rect -311 1095 -265 1107
rect -311 729 -305 1095
rect -271 729 -265 1095
rect -311 717 -265 729
rect -215 1095 -169 1107
rect -215 729 -209 1095
rect -175 729 -169 1095
rect -215 717 -169 729
rect -119 1095 -73 1107
rect -119 729 -113 1095
rect -79 729 -73 1095
rect -119 717 -73 729
rect -23 1095 23 1107
rect -23 729 -17 1095
rect 17 729 23 1095
rect -23 717 23 729
rect 73 1095 119 1107
rect 73 729 79 1095
rect 113 729 119 1095
rect 73 717 119 729
rect 169 1095 215 1107
rect 169 729 175 1095
rect 209 729 215 1095
rect 169 717 215 729
rect 265 1095 311 1107
rect 265 729 271 1095
rect 305 729 311 1095
rect 265 717 311 729
rect 361 1095 407 1107
rect 361 729 367 1095
rect 401 729 407 1095
rect 361 717 407 729
rect 457 1095 503 1107
rect 457 729 463 1095
rect 497 729 503 1095
rect 457 717 503 729
rect 553 1095 599 1107
rect 553 729 559 1095
rect 593 729 599 1095
rect 553 717 599 729
rect 649 1095 695 1107
rect 649 729 655 1095
rect 689 729 695 1095
rect 649 717 695 729
rect 745 1095 791 1107
rect 745 729 751 1095
rect 785 729 791 1095
rect 745 717 791 729
rect 841 1095 887 1107
rect 841 729 847 1095
rect 881 729 887 1095
rect 841 717 887 729
rect 937 1095 983 1107
rect 937 729 943 1095
rect 977 729 983 1095
rect 937 717 983 729
rect 1033 1095 1079 1107
rect 1033 729 1039 1095
rect 1073 729 1079 1095
rect 1033 717 1079 729
rect 1129 1095 1175 1107
rect 1129 729 1135 1095
rect 1169 729 1175 1095
rect 1129 717 1175 729
rect 1225 1095 1271 1107
rect 1225 729 1231 1095
rect 1265 729 1271 1095
rect 1225 717 1271 729
rect 1321 1095 1367 1107
rect 1321 729 1327 1095
rect 1361 729 1367 1095
rect 1321 717 1367 729
rect 1417 1095 1463 1107
rect 1417 729 1423 1095
rect 1457 729 1463 1095
rect 1417 717 1463 729
rect 1513 1095 1559 1107
rect 1513 729 1519 1095
rect 1553 729 1559 1095
rect 1513 717 1559 729
rect 1609 1095 1655 1107
rect 1609 729 1615 1095
rect 1649 729 1655 1095
rect 1609 717 1655 729
rect 1705 1095 1751 1107
rect 1705 729 1711 1095
rect 1745 729 1751 1095
rect 1705 717 1751 729
rect 1801 1095 1847 1107
rect 1801 729 1807 1095
rect 1841 729 1847 1095
rect 1801 717 1847 729
rect 1897 1095 1943 1107
rect 1897 729 1903 1095
rect 1937 729 1943 1095
rect 1897 717 1943 729
rect -1901 679 -1843 685
rect -1901 645 -1889 679
rect -1855 645 -1843 679
rect -1901 639 -1843 645
rect -1709 679 -1651 685
rect -1709 645 -1697 679
rect -1663 645 -1651 679
rect -1709 639 -1651 645
rect -1517 679 -1459 685
rect -1517 645 -1505 679
rect -1471 645 -1459 679
rect -1517 639 -1459 645
rect -1325 679 -1267 685
rect -1325 645 -1313 679
rect -1279 645 -1267 679
rect -1325 639 -1267 645
rect -1133 679 -1075 685
rect -1133 645 -1121 679
rect -1087 645 -1075 679
rect -1133 639 -1075 645
rect -941 679 -883 685
rect -941 645 -929 679
rect -895 645 -883 679
rect -941 639 -883 645
rect -749 679 -691 685
rect -749 645 -737 679
rect -703 645 -691 679
rect -749 639 -691 645
rect -557 679 -499 685
rect -557 645 -545 679
rect -511 645 -499 679
rect -557 639 -499 645
rect -365 679 -307 685
rect -365 645 -353 679
rect -319 645 -307 679
rect -365 639 -307 645
rect -173 679 -115 685
rect -173 645 -161 679
rect -127 645 -115 679
rect -173 639 -115 645
rect 19 679 77 685
rect 19 645 31 679
rect 65 645 77 679
rect 19 639 77 645
rect 211 679 269 685
rect 211 645 223 679
rect 257 645 269 679
rect 211 639 269 645
rect 403 679 461 685
rect 403 645 415 679
rect 449 645 461 679
rect 403 639 461 645
rect 595 679 653 685
rect 595 645 607 679
rect 641 645 653 679
rect 595 639 653 645
rect 787 679 845 685
rect 787 645 799 679
rect 833 645 845 679
rect 787 639 845 645
rect 979 679 1037 685
rect 979 645 991 679
rect 1025 645 1037 679
rect 979 639 1037 645
rect 1171 679 1229 685
rect 1171 645 1183 679
rect 1217 645 1229 679
rect 1171 639 1229 645
rect 1363 679 1421 685
rect 1363 645 1375 679
rect 1409 645 1421 679
rect 1363 639 1421 645
rect 1555 679 1613 685
rect 1555 645 1567 679
rect 1601 645 1613 679
rect 1555 639 1613 645
rect 1747 679 1805 685
rect 1747 645 1759 679
rect 1793 645 1805 679
rect 1747 639 1805 645
rect -1901 571 -1843 577
rect -1901 537 -1889 571
rect -1855 537 -1843 571
rect -1901 531 -1843 537
rect -1709 571 -1651 577
rect -1709 537 -1697 571
rect -1663 537 -1651 571
rect -1709 531 -1651 537
rect -1517 571 -1459 577
rect -1517 537 -1505 571
rect -1471 537 -1459 571
rect -1517 531 -1459 537
rect -1325 571 -1267 577
rect -1325 537 -1313 571
rect -1279 537 -1267 571
rect -1325 531 -1267 537
rect -1133 571 -1075 577
rect -1133 537 -1121 571
rect -1087 537 -1075 571
rect -1133 531 -1075 537
rect -941 571 -883 577
rect -941 537 -929 571
rect -895 537 -883 571
rect -941 531 -883 537
rect -749 571 -691 577
rect -749 537 -737 571
rect -703 537 -691 571
rect -749 531 -691 537
rect -557 571 -499 577
rect -557 537 -545 571
rect -511 537 -499 571
rect -557 531 -499 537
rect -365 571 -307 577
rect -365 537 -353 571
rect -319 537 -307 571
rect -365 531 -307 537
rect -173 571 -115 577
rect -173 537 -161 571
rect -127 537 -115 571
rect -173 531 -115 537
rect 19 571 77 577
rect 19 537 31 571
rect 65 537 77 571
rect 19 531 77 537
rect 211 571 269 577
rect 211 537 223 571
rect 257 537 269 571
rect 211 531 269 537
rect 403 571 461 577
rect 403 537 415 571
rect 449 537 461 571
rect 403 531 461 537
rect 595 571 653 577
rect 595 537 607 571
rect 641 537 653 571
rect 595 531 653 537
rect 787 571 845 577
rect 787 537 799 571
rect 833 537 845 571
rect 787 531 845 537
rect 979 571 1037 577
rect 979 537 991 571
rect 1025 537 1037 571
rect 979 531 1037 537
rect 1171 571 1229 577
rect 1171 537 1183 571
rect 1217 537 1229 571
rect 1171 531 1229 537
rect 1363 571 1421 577
rect 1363 537 1375 571
rect 1409 537 1421 571
rect 1363 531 1421 537
rect 1555 571 1613 577
rect 1555 537 1567 571
rect 1601 537 1613 571
rect 1555 531 1613 537
rect 1747 571 1805 577
rect 1747 537 1759 571
rect 1793 537 1805 571
rect 1747 531 1805 537
rect -1943 487 -1897 499
rect -1943 121 -1937 487
rect -1903 121 -1897 487
rect -1943 109 -1897 121
rect -1847 487 -1801 499
rect -1847 121 -1841 487
rect -1807 121 -1801 487
rect -1847 109 -1801 121
rect -1751 487 -1705 499
rect -1751 121 -1745 487
rect -1711 121 -1705 487
rect -1751 109 -1705 121
rect -1655 487 -1609 499
rect -1655 121 -1649 487
rect -1615 121 -1609 487
rect -1655 109 -1609 121
rect -1559 487 -1513 499
rect -1559 121 -1553 487
rect -1519 121 -1513 487
rect -1559 109 -1513 121
rect -1463 487 -1417 499
rect -1463 121 -1457 487
rect -1423 121 -1417 487
rect -1463 109 -1417 121
rect -1367 487 -1321 499
rect -1367 121 -1361 487
rect -1327 121 -1321 487
rect -1367 109 -1321 121
rect -1271 487 -1225 499
rect -1271 121 -1265 487
rect -1231 121 -1225 487
rect -1271 109 -1225 121
rect -1175 487 -1129 499
rect -1175 121 -1169 487
rect -1135 121 -1129 487
rect -1175 109 -1129 121
rect -1079 487 -1033 499
rect -1079 121 -1073 487
rect -1039 121 -1033 487
rect -1079 109 -1033 121
rect -983 487 -937 499
rect -983 121 -977 487
rect -943 121 -937 487
rect -983 109 -937 121
rect -887 487 -841 499
rect -887 121 -881 487
rect -847 121 -841 487
rect -887 109 -841 121
rect -791 487 -745 499
rect -791 121 -785 487
rect -751 121 -745 487
rect -791 109 -745 121
rect -695 487 -649 499
rect -695 121 -689 487
rect -655 121 -649 487
rect -695 109 -649 121
rect -599 487 -553 499
rect -599 121 -593 487
rect -559 121 -553 487
rect -599 109 -553 121
rect -503 487 -457 499
rect -503 121 -497 487
rect -463 121 -457 487
rect -503 109 -457 121
rect -407 487 -361 499
rect -407 121 -401 487
rect -367 121 -361 487
rect -407 109 -361 121
rect -311 487 -265 499
rect -311 121 -305 487
rect -271 121 -265 487
rect -311 109 -265 121
rect -215 487 -169 499
rect -215 121 -209 487
rect -175 121 -169 487
rect -215 109 -169 121
rect -119 487 -73 499
rect -119 121 -113 487
rect -79 121 -73 487
rect -119 109 -73 121
rect -23 487 23 499
rect -23 121 -17 487
rect 17 121 23 487
rect -23 109 23 121
rect 73 487 119 499
rect 73 121 79 487
rect 113 121 119 487
rect 73 109 119 121
rect 169 487 215 499
rect 169 121 175 487
rect 209 121 215 487
rect 169 109 215 121
rect 265 487 311 499
rect 265 121 271 487
rect 305 121 311 487
rect 265 109 311 121
rect 361 487 407 499
rect 361 121 367 487
rect 401 121 407 487
rect 361 109 407 121
rect 457 487 503 499
rect 457 121 463 487
rect 497 121 503 487
rect 457 109 503 121
rect 553 487 599 499
rect 553 121 559 487
rect 593 121 599 487
rect 553 109 599 121
rect 649 487 695 499
rect 649 121 655 487
rect 689 121 695 487
rect 649 109 695 121
rect 745 487 791 499
rect 745 121 751 487
rect 785 121 791 487
rect 745 109 791 121
rect 841 487 887 499
rect 841 121 847 487
rect 881 121 887 487
rect 841 109 887 121
rect 937 487 983 499
rect 937 121 943 487
rect 977 121 983 487
rect 937 109 983 121
rect 1033 487 1079 499
rect 1033 121 1039 487
rect 1073 121 1079 487
rect 1033 109 1079 121
rect 1129 487 1175 499
rect 1129 121 1135 487
rect 1169 121 1175 487
rect 1129 109 1175 121
rect 1225 487 1271 499
rect 1225 121 1231 487
rect 1265 121 1271 487
rect 1225 109 1271 121
rect 1321 487 1367 499
rect 1321 121 1327 487
rect 1361 121 1367 487
rect 1321 109 1367 121
rect 1417 487 1463 499
rect 1417 121 1423 487
rect 1457 121 1463 487
rect 1417 109 1463 121
rect 1513 487 1559 499
rect 1513 121 1519 487
rect 1553 121 1559 487
rect 1513 109 1559 121
rect 1609 487 1655 499
rect 1609 121 1615 487
rect 1649 121 1655 487
rect 1609 109 1655 121
rect 1705 487 1751 499
rect 1705 121 1711 487
rect 1745 121 1751 487
rect 1705 109 1751 121
rect 1801 487 1847 499
rect 1801 121 1807 487
rect 1841 121 1847 487
rect 1801 109 1847 121
rect 1897 487 1943 499
rect 1897 121 1903 487
rect 1937 121 1943 487
rect 1897 109 1943 121
rect -1805 71 -1747 77
rect -1805 37 -1793 71
rect -1759 37 -1747 71
rect -1805 31 -1747 37
rect -1613 71 -1555 77
rect -1613 37 -1601 71
rect -1567 37 -1555 71
rect -1613 31 -1555 37
rect -1421 71 -1363 77
rect -1421 37 -1409 71
rect -1375 37 -1363 71
rect -1421 31 -1363 37
rect -1229 71 -1171 77
rect -1229 37 -1217 71
rect -1183 37 -1171 71
rect -1229 31 -1171 37
rect -1037 71 -979 77
rect -1037 37 -1025 71
rect -991 37 -979 71
rect -1037 31 -979 37
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect 1075 71 1133 77
rect 1075 37 1087 71
rect 1121 37 1133 71
rect 1075 31 1133 37
rect 1267 71 1325 77
rect 1267 37 1279 71
rect 1313 37 1325 71
rect 1267 31 1325 37
rect 1459 71 1517 77
rect 1459 37 1471 71
rect 1505 37 1517 71
rect 1459 31 1517 37
rect 1651 71 1709 77
rect 1651 37 1663 71
rect 1697 37 1709 71
rect 1651 31 1709 37
rect 1843 71 1901 77
rect 1843 37 1855 71
rect 1889 37 1901 71
rect 1843 31 1901 37
rect -1805 -37 -1747 -31
rect -1805 -71 -1793 -37
rect -1759 -71 -1747 -37
rect -1805 -77 -1747 -71
rect -1613 -37 -1555 -31
rect -1613 -71 -1601 -37
rect -1567 -71 -1555 -37
rect -1613 -77 -1555 -71
rect -1421 -37 -1363 -31
rect -1421 -71 -1409 -37
rect -1375 -71 -1363 -37
rect -1421 -77 -1363 -71
rect -1229 -37 -1171 -31
rect -1229 -71 -1217 -37
rect -1183 -71 -1171 -37
rect -1229 -77 -1171 -71
rect -1037 -37 -979 -31
rect -1037 -71 -1025 -37
rect -991 -71 -979 -37
rect -1037 -77 -979 -71
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect 1075 -37 1133 -31
rect 1075 -71 1087 -37
rect 1121 -71 1133 -37
rect 1075 -77 1133 -71
rect 1267 -37 1325 -31
rect 1267 -71 1279 -37
rect 1313 -71 1325 -37
rect 1267 -77 1325 -71
rect 1459 -37 1517 -31
rect 1459 -71 1471 -37
rect 1505 -71 1517 -37
rect 1459 -77 1517 -71
rect 1651 -37 1709 -31
rect 1651 -71 1663 -37
rect 1697 -71 1709 -37
rect 1651 -77 1709 -71
rect 1843 -37 1901 -31
rect 1843 -71 1855 -37
rect 1889 -71 1901 -37
rect 1843 -77 1901 -71
rect -1943 -121 -1897 -109
rect -1943 -487 -1937 -121
rect -1903 -487 -1897 -121
rect -1943 -499 -1897 -487
rect -1847 -121 -1801 -109
rect -1847 -487 -1841 -121
rect -1807 -487 -1801 -121
rect -1847 -499 -1801 -487
rect -1751 -121 -1705 -109
rect -1751 -487 -1745 -121
rect -1711 -487 -1705 -121
rect -1751 -499 -1705 -487
rect -1655 -121 -1609 -109
rect -1655 -487 -1649 -121
rect -1615 -487 -1609 -121
rect -1655 -499 -1609 -487
rect -1559 -121 -1513 -109
rect -1559 -487 -1553 -121
rect -1519 -487 -1513 -121
rect -1559 -499 -1513 -487
rect -1463 -121 -1417 -109
rect -1463 -487 -1457 -121
rect -1423 -487 -1417 -121
rect -1463 -499 -1417 -487
rect -1367 -121 -1321 -109
rect -1367 -487 -1361 -121
rect -1327 -487 -1321 -121
rect -1367 -499 -1321 -487
rect -1271 -121 -1225 -109
rect -1271 -487 -1265 -121
rect -1231 -487 -1225 -121
rect -1271 -499 -1225 -487
rect -1175 -121 -1129 -109
rect -1175 -487 -1169 -121
rect -1135 -487 -1129 -121
rect -1175 -499 -1129 -487
rect -1079 -121 -1033 -109
rect -1079 -487 -1073 -121
rect -1039 -487 -1033 -121
rect -1079 -499 -1033 -487
rect -983 -121 -937 -109
rect -983 -487 -977 -121
rect -943 -487 -937 -121
rect -983 -499 -937 -487
rect -887 -121 -841 -109
rect -887 -487 -881 -121
rect -847 -487 -841 -121
rect -887 -499 -841 -487
rect -791 -121 -745 -109
rect -791 -487 -785 -121
rect -751 -487 -745 -121
rect -791 -499 -745 -487
rect -695 -121 -649 -109
rect -695 -487 -689 -121
rect -655 -487 -649 -121
rect -695 -499 -649 -487
rect -599 -121 -553 -109
rect -599 -487 -593 -121
rect -559 -487 -553 -121
rect -599 -499 -553 -487
rect -503 -121 -457 -109
rect -503 -487 -497 -121
rect -463 -487 -457 -121
rect -503 -499 -457 -487
rect -407 -121 -361 -109
rect -407 -487 -401 -121
rect -367 -487 -361 -121
rect -407 -499 -361 -487
rect -311 -121 -265 -109
rect -311 -487 -305 -121
rect -271 -487 -265 -121
rect -311 -499 -265 -487
rect -215 -121 -169 -109
rect -215 -487 -209 -121
rect -175 -487 -169 -121
rect -215 -499 -169 -487
rect -119 -121 -73 -109
rect -119 -487 -113 -121
rect -79 -487 -73 -121
rect -119 -499 -73 -487
rect -23 -121 23 -109
rect -23 -487 -17 -121
rect 17 -487 23 -121
rect -23 -499 23 -487
rect 73 -121 119 -109
rect 73 -487 79 -121
rect 113 -487 119 -121
rect 73 -499 119 -487
rect 169 -121 215 -109
rect 169 -487 175 -121
rect 209 -487 215 -121
rect 169 -499 215 -487
rect 265 -121 311 -109
rect 265 -487 271 -121
rect 305 -487 311 -121
rect 265 -499 311 -487
rect 361 -121 407 -109
rect 361 -487 367 -121
rect 401 -487 407 -121
rect 361 -499 407 -487
rect 457 -121 503 -109
rect 457 -487 463 -121
rect 497 -487 503 -121
rect 457 -499 503 -487
rect 553 -121 599 -109
rect 553 -487 559 -121
rect 593 -487 599 -121
rect 553 -499 599 -487
rect 649 -121 695 -109
rect 649 -487 655 -121
rect 689 -487 695 -121
rect 649 -499 695 -487
rect 745 -121 791 -109
rect 745 -487 751 -121
rect 785 -487 791 -121
rect 745 -499 791 -487
rect 841 -121 887 -109
rect 841 -487 847 -121
rect 881 -487 887 -121
rect 841 -499 887 -487
rect 937 -121 983 -109
rect 937 -487 943 -121
rect 977 -487 983 -121
rect 937 -499 983 -487
rect 1033 -121 1079 -109
rect 1033 -487 1039 -121
rect 1073 -487 1079 -121
rect 1033 -499 1079 -487
rect 1129 -121 1175 -109
rect 1129 -487 1135 -121
rect 1169 -487 1175 -121
rect 1129 -499 1175 -487
rect 1225 -121 1271 -109
rect 1225 -487 1231 -121
rect 1265 -487 1271 -121
rect 1225 -499 1271 -487
rect 1321 -121 1367 -109
rect 1321 -487 1327 -121
rect 1361 -487 1367 -121
rect 1321 -499 1367 -487
rect 1417 -121 1463 -109
rect 1417 -487 1423 -121
rect 1457 -487 1463 -121
rect 1417 -499 1463 -487
rect 1513 -121 1559 -109
rect 1513 -487 1519 -121
rect 1553 -487 1559 -121
rect 1513 -499 1559 -487
rect 1609 -121 1655 -109
rect 1609 -487 1615 -121
rect 1649 -487 1655 -121
rect 1609 -499 1655 -487
rect 1705 -121 1751 -109
rect 1705 -487 1711 -121
rect 1745 -487 1751 -121
rect 1705 -499 1751 -487
rect 1801 -121 1847 -109
rect 1801 -487 1807 -121
rect 1841 -487 1847 -121
rect 1801 -499 1847 -487
rect 1897 -121 1943 -109
rect 1897 -487 1903 -121
rect 1937 -487 1943 -121
rect 1897 -499 1943 -487
rect -1901 -537 -1843 -531
rect -1901 -571 -1889 -537
rect -1855 -571 -1843 -537
rect -1901 -577 -1843 -571
rect -1709 -537 -1651 -531
rect -1709 -571 -1697 -537
rect -1663 -571 -1651 -537
rect -1709 -577 -1651 -571
rect -1517 -537 -1459 -531
rect -1517 -571 -1505 -537
rect -1471 -571 -1459 -537
rect -1517 -577 -1459 -571
rect -1325 -537 -1267 -531
rect -1325 -571 -1313 -537
rect -1279 -571 -1267 -537
rect -1325 -577 -1267 -571
rect -1133 -537 -1075 -531
rect -1133 -571 -1121 -537
rect -1087 -571 -1075 -537
rect -1133 -577 -1075 -571
rect -941 -537 -883 -531
rect -941 -571 -929 -537
rect -895 -571 -883 -537
rect -941 -577 -883 -571
rect -749 -537 -691 -531
rect -749 -571 -737 -537
rect -703 -571 -691 -537
rect -749 -577 -691 -571
rect -557 -537 -499 -531
rect -557 -571 -545 -537
rect -511 -571 -499 -537
rect -557 -577 -499 -571
rect -365 -537 -307 -531
rect -365 -571 -353 -537
rect -319 -571 -307 -537
rect -365 -577 -307 -571
rect -173 -537 -115 -531
rect -173 -571 -161 -537
rect -127 -571 -115 -537
rect -173 -577 -115 -571
rect 19 -537 77 -531
rect 19 -571 31 -537
rect 65 -571 77 -537
rect 19 -577 77 -571
rect 211 -537 269 -531
rect 211 -571 223 -537
rect 257 -571 269 -537
rect 211 -577 269 -571
rect 403 -537 461 -531
rect 403 -571 415 -537
rect 449 -571 461 -537
rect 403 -577 461 -571
rect 595 -537 653 -531
rect 595 -571 607 -537
rect 641 -571 653 -537
rect 595 -577 653 -571
rect 787 -537 845 -531
rect 787 -571 799 -537
rect 833 -571 845 -537
rect 787 -577 845 -571
rect 979 -537 1037 -531
rect 979 -571 991 -537
rect 1025 -571 1037 -537
rect 979 -577 1037 -571
rect 1171 -537 1229 -531
rect 1171 -571 1183 -537
rect 1217 -571 1229 -537
rect 1171 -577 1229 -571
rect 1363 -537 1421 -531
rect 1363 -571 1375 -537
rect 1409 -571 1421 -537
rect 1363 -577 1421 -571
rect 1555 -537 1613 -531
rect 1555 -571 1567 -537
rect 1601 -571 1613 -537
rect 1555 -577 1613 -571
rect 1747 -537 1805 -531
rect 1747 -571 1759 -537
rect 1793 -571 1805 -537
rect 1747 -577 1805 -571
rect -1901 -645 -1843 -639
rect -1901 -679 -1889 -645
rect -1855 -679 -1843 -645
rect -1901 -685 -1843 -679
rect -1709 -645 -1651 -639
rect -1709 -679 -1697 -645
rect -1663 -679 -1651 -645
rect -1709 -685 -1651 -679
rect -1517 -645 -1459 -639
rect -1517 -679 -1505 -645
rect -1471 -679 -1459 -645
rect -1517 -685 -1459 -679
rect -1325 -645 -1267 -639
rect -1325 -679 -1313 -645
rect -1279 -679 -1267 -645
rect -1325 -685 -1267 -679
rect -1133 -645 -1075 -639
rect -1133 -679 -1121 -645
rect -1087 -679 -1075 -645
rect -1133 -685 -1075 -679
rect -941 -645 -883 -639
rect -941 -679 -929 -645
rect -895 -679 -883 -645
rect -941 -685 -883 -679
rect -749 -645 -691 -639
rect -749 -679 -737 -645
rect -703 -679 -691 -645
rect -749 -685 -691 -679
rect -557 -645 -499 -639
rect -557 -679 -545 -645
rect -511 -679 -499 -645
rect -557 -685 -499 -679
rect -365 -645 -307 -639
rect -365 -679 -353 -645
rect -319 -679 -307 -645
rect -365 -685 -307 -679
rect -173 -645 -115 -639
rect -173 -679 -161 -645
rect -127 -679 -115 -645
rect -173 -685 -115 -679
rect 19 -645 77 -639
rect 19 -679 31 -645
rect 65 -679 77 -645
rect 19 -685 77 -679
rect 211 -645 269 -639
rect 211 -679 223 -645
rect 257 -679 269 -645
rect 211 -685 269 -679
rect 403 -645 461 -639
rect 403 -679 415 -645
rect 449 -679 461 -645
rect 403 -685 461 -679
rect 595 -645 653 -639
rect 595 -679 607 -645
rect 641 -679 653 -645
rect 595 -685 653 -679
rect 787 -645 845 -639
rect 787 -679 799 -645
rect 833 -679 845 -645
rect 787 -685 845 -679
rect 979 -645 1037 -639
rect 979 -679 991 -645
rect 1025 -679 1037 -645
rect 979 -685 1037 -679
rect 1171 -645 1229 -639
rect 1171 -679 1183 -645
rect 1217 -679 1229 -645
rect 1171 -685 1229 -679
rect 1363 -645 1421 -639
rect 1363 -679 1375 -645
rect 1409 -679 1421 -645
rect 1363 -685 1421 -679
rect 1555 -645 1613 -639
rect 1555 -679 1567 -645
rect 1601 -679 1613 -645
rect 1555 -685 1613 -679
rect 1747 -645 1805 -639
rect 1747 -679 1759 -645
rect 1793 -679 1805 -645
rect 1747 -685 1805 -679
rect -1943 -729 -1897 -717
rect -1943 -1095 -1937 -729
rect -1903 -1095 -1897 -729
rect -1943 -1107 -1897 -1095
rect -1847 -729 -1801 -717
rect -1847 -1095 -1841 -729
rect -1807 -1095 -1801 -729
rect -1847 -1107 -1801 -1095
rect -1751 -729 -1705 -717
rect -1751 -1095 -1745 -729
rect -1711 -1095 -1705 -729
rect -1751 -1107 -1705 -1095
rect -1655 -729 -1609 -717
rect -1655 -1095 -1649 -729
rect -1615 -1095 -1609 -729
rect -1655 -1107 -1609 -1095
rect -1559 -729 -1513 -717
rect -1559 -1095 -1553 -729
rect -1519 -1095 -1513 -729
rect -1559 -1107 -1513 -1095
rect -1463 -729 -1417 -717
rect -1463 -1095 -1457 -729
rect -1423 -1095 -1417 -729
rect -1463 -1107 -1417 -1095
rect -1367 -729 -1321 -717
rect -1367 -1095 -1361 -729
rect -1327 -1095 -1321 -729
rect -1367 -1107 -1321 -1095
rect -1271 -729 -1225 -717
rect -1271 -1095 -1265 -729
rect -1231 -1095 -1225 -729
rect -1271 -1107 -1225 -1095
rect -1175 -729 -1129 -717
rect -1175 -1095 -1169 -729
rect -1135 -1095 -1129 -729
rect -1175 -1107 -1129 -1095
rect -1079 -729 -1033 -717
rect -1079 -1095 -1073 -729
rect -1039 -1095 -1033 -729
rect -1079 -1107 -1033 -1095
rect -983 -729 -937 -717
rect -983 -1095 -977 -729
rect -943 -1095 -937 -729
rect -983 -1107 -937 -1095
rect -887 -729 -841 -717
rect -887 -1095 -881 -729
rect -847 -1095 -841 -729
rect -887 -1107 -841 -1095
rect -791 -729 -745 -717
rect -791 -1095 -785 -729
rect -751 -1095 -745 -729
rect -791 -1107 -745 -1095
rect -695 -729 -649 -717
rect -695 -1095 -689 -729
rect -655 -1095 -649 -729
rect -695 -1107 -649 -1095
rect -599 -729 -553 -717
rect -599 -1095 -593 -729
rect -559 -1095 -553 -729
rect -599 -1107 -553 -1095
rect -503 -729 -457 -717
rect -503 -1095 -497 -729
rect -463 -1095 -457 -729
rect -503 -1107 -457 -1095
rect -407 -729 -361 -717
rect -407 -1095 -401 -729
rect -367 -1095 -361 -729
rect -407 -1107 -361 -1095
rect -311 -729 -265 -717
rect -311 -1095 -305 -729
rect -271 -1095 -265 -729
rect -311 -1107 -265 -1095
rect -215 -729 -169 -717
rect -215 -1095 -209 -729
rect -175 -1095 -169 -729
rect -215 -1107 -169 -1095
rect -119 -729 -73 -717
rect -119 -1095 -113 -729
rect -79 -1095 -73 -729
rect -119 -1107 -73 -1095
rect -23 -729 23 -717
rect -23 -1095 -17 -729
rect 17 -1095 23 -729
rect -23 -1107 23 -1095
rect 73 -729 119 -717
rect 73 -1095 79 -729
rect 113 -1095 119 -729
rect 73 -1107 119 -1095
rect 169 -729 215 -717
rect 169 -1095 175 -729
rect 209 -1095 215 -729
rect 169 -1107 215 -1095
rect 265 -729 311 -717
rect 265 -1095 271 -729
rect 305 -1095 311 -729
rect 265 -1107 311 -1095
rect 361 -729 407 -717
rect 361 -1095 367 -729
rect 401 -1095 407 -729
rect 361 -1107 407 -1095
rect 457 -729 503 -717
rect 457 -1095 463 -729
rect 497 -1095 503 -729
rect 457 -1107 503 -1095
rect 553 -729 599 -717
rect 553 -1095 559 -729
rect 593 -1095 599 -729
rect 553 -1107 599 -1095
rect 649 -729 695 -717
rect 649 -1095 655 -729
rect 689 -1095 695 -729
rect 649 -1107 695 -1095
rect 745 -729 791 -717
rect 745 -1095 751 -729
rect 785 -1095 791 -729
rect 745 -1107 791 -1095
rect 841 -729 887 -717
rect 841 -1095 847 -729
rect 881 -1095 887 -729
rect 841 -1107 887 -1095
rect 937 -729 983 -717
rect 937 -1095 943 -729
rect 977 -1095 983 -729
rect 937 -1107 983 -1095
rect 1033 -729 1079 -717
rect 1033 -1095 1039 -729
rect 1073 -1095 1079 -729
rect 1033 -1107 1079 -1095
rect 1129 -729 1175 -717
rect 1129 -1095 1135 -729
rect 1169 -1095 1175 -729
rect 1129 -1107 1175 -1095
rect 1225 -729 1271 -717
rect 1225 -1095 1231 -729
rect 1265 -1095 1271 -729
rect 1225 -1107 1271 -1095
rect 1321 -729 1367 -717
rect 1321 -1095 1327 -729
rect 1361 -1095 1367 -729
rect 1321 -1107 1367 -1095
rect 1417 -729 1463 -717
rect 1417 -1095 1423 -729
rect 1457 -1095 1463 -729
rect 1417 -1107 1463 -1095
rect 1513 -729 1559 -717
rect 1513 -1095 1519 -729
rect 1553 -1095 1559 -729
rect 1513 -1107 1559 -1095
rect 1609 -729 1655 -717
rect 1609 -1095 1615 -729
rect 1649 -1095 1655 -729
rect 1609 -1107 1655 -1095
rect 1705 -729 1751 -717
rect 1705 -1095 1711 -729
rect 1745 -1095 1751 -729
rect 1705 -1107 1751 -1095
rect 1801 -729 1847 -717
rect 1801 -1095 1807 -729
rect 1841 -1095 1847 -729
rect 1801 -1107 1847 -1095
rect 1897 -729 1943 -717
rect 1897 -1095 1903 -729
rect 1937 -1095 1943 -729
rect 1897 -1107 1943 -1095
rect -1805 -1145 -1747 -1139
rect -1805 -1179 -1793 -1145
rect -1759 -1179 -1747 -1145
rect -1805 -1185 -1747 -1179
rect -1613 -1145 -1555 -1139
rect -1613 -1179 -1601 -1145
rect -1567 -1179 -1555 -1145
rect -1613 -1185 -1555 -1179
rect -1421 -1145 -1363 -1139
rect -1421 -1179 -1409 -1145
rect -1375 -1179 -1363 -1145
rect -1421 -1185 -1363 -1179
rect -1229 -1145 -1171 -1139
rect -1229 -1179 -1217 -1145
rect -1183 -1179 -1171 -1145
rect -1229 -1185 -1171 -1179
rect -1037 -1145 -979 -1139
rect -1037 -1179 -1025 -1145
rect -991 -1179 -979 -1145
rect -1037 -1185 -979 -1179
rect -845 -1145 -787 -1139
rect -845 -1179 -833 -1145
rect -799 -1179 -787 -1145
rect -845 -1185 -787 -1179
rect -653 -1145 -595 -1139
rect -653 -1179 -641 -1145
rect -607 -1179 -595 -1145
rect -653 -1185 -595 -1179
rect -461 -1145 -403 -1139
rect -461 -1179 -449 -1145
rect -415 -1179 -403 -1145
rect -461 -1185 -403 -1179
rect -269 -1145 -211 -1139
rect -269 -1179 -257 -1145
rect -223 -1179 -211 -1145
rect -269 -1185 -211 -1179
rect -77 -1145 -19 -1139
rect -77 -1179 -65 -1145
rect -31 -1179 -19 -1145
rect -77 -1185 -19 -1179
rect 115 -1145 173 -1139
rect 115 -1179 127 -1145
rect 161 -1179 173 -1145
rect 115 -1185 173 -1179
rect 307 -1145 365 -1139
rect 307 -1179 319 -1145
rect 353 -1179 365 -1145
rect 307 -1185 365 -1179
rect 499 -1145 557 -1139
rect 499 -1179 511 -1145
rect 545 -1179 557 -1145
rect 499 -1185 557 -1179
rect 691 -1145 749 -1139
rect 691 -1179 703 -1145
rect 737 -1179 749 -1145
rect 691 -1185 749 -1179
rect 883 -1145 941 -1139
rect 883 -1179 895 -1145
rect 929 -1179 941 -1145
rect 883 -1185 941 -1179
rect 1075 -1145 1133 -1139
rect 1075 -1179 1087 -1145
rect 1121 -1179 1133 -1145
rect 1075 -1185 1133 -1179
rect 1267 -1145 1325 -1139
rect 1267 -1179 1279 -1145
rect 1313 -1179 1325 -1145
rect 1267 -1185 1325 -1179
rect 1459 -1145 1517 -1139
rect 1459 -1179 1471 -1145
rect 1505 -1179 1517 -1145
rect 1459 -1185 1517 -1179
rect 1651 -1145 1709 -1139
rect 1651 -1179 1663 -1145
rect 1697 -1179 1709 -1145
rect 1651 -1185 1709 -1179
rect 1843 -1145 1901 -1139
rect 1843 -1179 1855 -1145
rect 1889 -1179 1901 -1145
rect 1843 -1185 1901 -1179
rect -1805 -1253 -1747 -1247
rect -1805 -1287 -1793 -1253
rect -1759 -1287 -1747 -1253
rect -1805 -1293 -1747 -1287
rect -1613 -1253 -1555 -1247
rect -1613 -1287 -1601 -1253
rect -1567 -1287 -1555 -1253
rect -1613 -1293 -1555 -1287
rect -1421 -1253 -1363 -1247
rect -1421 -1287 -1409 -1253
rect -1375 -1287 -1363 -1253
rect -1421 -1293 -1363 -1287
rect -1229 -1253 -1171 -1247
rect -1229 -1287 -1217 -1253
rect -1183 -1287 -1171 -1253
rect -1229 -1293 -1171 -1287
rect -1037 -1253 -979 -1247
rect -1037 -1287 -1025 -1253
rect -991 -1287 -979 -1253
rect -1037 -1293 -979 -1287
rect -845 -1253 -787 -1247
rect -845 -1287 -833 -1253
rect -799 -1287 -787 -1253
rect -845 -1293 -787 -1287
rect -653 -1253 -595 -1247
rect -653 -1287 -641 -1253
rect -607 -1287 -595 -1253
rect -653 -1293 -595 -1287
rect -461 -1253 -403 -1247
rect -461 -1287 -449 -1253
rect -415 -1287 -403 -1253
rect -461 -1293 -403 -1287
rect -269 -1253 -211 -1247
rect -269 -1287 -257 -1253
rect -223 -1287 -211 -1253
rect -269 -1293 -211 -1287
rect -77 -1253 -19 -1247
rect -77 -1287 -65 -1253
rect -31 -1287 -19 -1253
rect -77 -1293 -19 -1287
rect 115 -1253 173 -1247
rect 115 -1287 127 -1253
rect 161 -1287 173 -1253
rect 115 -1293 173 -1287
rect 307 -1253 365 -1247
rect 307 -1287 319 -1253
rect 353 -1287 365 -1253
rect 307 -1293 365 -1287
rect 499 -1253 557 -1247
rect 499 -1287 511 -1253
rect 545 -1287 557 -1253
rect 499 -1293 557 -1287
rect 691 -1253 749 -1247
rect 691 -1287 703 -1253
rect 737 -1287 749 -1253
rect 691 -1293 749 -1287
rect 883 -1253 941 -1247
rect 883 -1287 895 -1253
rect 929 -1287 941 -1253
rect 883 -1293 941 -1287
rect 1075 -1253 1133 -1247
rect 1075 -1287 1087 -1253
rect 1121 -1287 1133 -1253
rect 1075 -1293 1133 -1287
rect 1267 -1253 1325 -1247
rect 1267 -1287 1279 -1253
rect 1313 -1287 1325 -1253
rect 1267 -1293 1325 -1287
rect 1459 -1253 1517 -1247
rect 1459 -1287 1471 -1253
rect 1505 -1287 1517 -1253
rect 1459 -1293 1517 -1287
rect 1651 -1253 1709 -1247
rect 1651 -1287 1663 -1253
rect 1697 -1287 1709 -1253
rect 1651 -1293 1709 -1287
rect 1843 -1253 1901 -1247
rect 1843 -1287 1855 -1253
rect 1889 -1287 1901 -1253
rect 1843 -1293 1901 -1287
rect -1943 -1337 -1897 -1325
rect -1943 -1703 -1937 -1337
rect -1903 -1703 -1897 -1337
rect -1943 -1715 -1897 -1703
rect -1847 -1337 -1801 -1325
rect -1847 -1703 -1841 -1337
rect -1807 -1703 -1801 -1337
rect -1847 -1715 -1801 -1703
rect -1751 -1337 -1705 -1325
rect -1751 -1703 -1745 -1337
rect -1711 -1703 -1705 -1337
rect -1751 -1715 -1705 -1703
rect -1655 -1337 -1609 -1325
rect -1655 -1703 -1649 -1337
rect -1615 -1703 -1609 -1337
rect -1655 -1715 -1609 -1703
rect -1559 -1337 -1513 -1325
rect -1559 -1703 -1553 -1337
rect -1519 -1703 -1513 -1337
rect -1559 -1715 -1513 -1703
rect -1463 -1337 -1417 -1325
rect -1463 -1703 -1457 -1337
rect -1423 -1703 -1417 -1337
rect -1463 -1715 -1417 -1703
rect -1367 -1337 -1321 -1325
rect -1367 -1703 -1361 -1337
rect -1327 -1703 -1321 -1337
rect -1367 -1715 -1321 -1703
rect -1271 -1337 -1225 -1325
rect -1271 -1703 -1265 -1337
rect -1231 -1703 -1225 -1337
rect -1271 -1715 -1225 -1703
rect -1175 -1337 -1129 -1325
rect -1175 -1703 -1169 -1337
rect -1135 -1703 -1129 -1337
rect -1175 -1715 -1129 -1703
rect -1079 -1337 -1033 -1325
rect -1079 -1703 -1073 -1337
rect -1039 -1703 -1033 -1337
rect -1079 -1715 -1033 -1703
rect -983 -1337 -937 -1325
rect -983 -1703 -977 -1337
rect -943 -1703 -937 -1337
rect -983 -1715 -937 -1703
rect -887 -1337 -841 -1325
rect -887 -1703 -881 -1337
rect -847 -1703 -841 -1337
rect -887 -1715 -841 -1703
rect -791 -1337 -745 -1325
rect -791 -1703 -785 -1337
rect -751 -1703 -745 -1337
rect -791 -1715 -745 -1703
rect -695 -1337 -649 -1325
rect -695 -1703 -689 -1337
rect -655 -1703 -649 -1337
rect -695 -1715 -649 -1703
rect -599 -1337 -553 -1325
rect -599 -1703 -593 -1337
rect -559 -1703 -553 -1337
rect -599 -1715 -553 -1703
rect -503 -1337 -457 -1325
rect -503 -1703 -497 -1337
rect -463 -1703 -457 -1337
rect -503 -1715 -457 -1703
rect -407 -1337 -361 -1325
rect -407 -1703 -401 -1337
rect -367 -1703 -361 -1337
rect -407 -1715 -361 -1703
rect -311 -1337 -265 -1325
rect -311 -1703 -305 -1337
rect -271 -1703 -265 -1337
rect -311 -1715 -265 -1703
rect -215 -1337 -169 -1325
rect -215 -1703 -209 -1337
rect -175 -1703 -169 -1337
rect -215 -1715 -169 -1703
rect -119 -1337 -73 -1325
rect -119 -1703 -113 -1337
rect -79 -1703 -73 -1337
rect -119 -1715 -73 -1703
rect -23 -1337 23 -1325
rect -23 -1703 -17 -1337
rect 17 -1703 23 -1337
rect -23 -1715 23 -1703
rect 73 -1337 119 -1325
rect 73 -1703 79 -1337
rect 113 -1703 119 -1337
rect 73 -1715 119 -1703
rect 169 -1337 215 -1325
rect 169 -1703 175 -1337
rect 209 -1703 215 -1337
rect 169 -1715 215 -1703
rect 265 -1337 311 -1325
rect 265 -1703 271 -1337
rect 305 -1703 311 -1337
rect 265 -1715 311 -1703
rect 361 -1337 407 -1325
rect 361 -1703 367 -1337
rect 401 -1703 407 -1337
rect 361 -1715 407 -1703
rect 457 -1337 503 -1325
rect 457 -1703 463 -1337
rect 497 -1703 503 -1337
rect 457 -1715 503 -1703
rect 553 -1337 599 -1325
rect 553 -1703 559 -1337
rect 593 -1703 599 -1337
rect 553 -1715 599 -1703
rect 649 -1337 695 -1325
rect 649 -1703 655 -1337
rect 689 -1703 695 -1337
rect 649 -1715 695 -1703
rect 745 -1337 791 -1325
rect 745 -1703 751 -1337
rect 785 -1703 791 -1337
rect 745 -1715 791 -1703
rect 841 -1337 887 -1325
rect 841 -1703 847 -1337
rect 881 -1703 887 -1337
rect 841 -1715 887 -1703
rect 937 -1337 983 -1325
rect 937 -1703 943 -1337
rect 977 -1703 983 -1337
rect 937 -1715 983 -1703
rect 1033 -1337 1079 -1325
rect 1033 -1703 1039 -1337
rect 1073 -1703 1079 -1337
rect 1033 -1715 1079 -1703
rect 1129 -1337 1175 -1325
rect 1129 -1703 1135 -1337
rect 1169 -1703 1175 -1337
rect 1129 -1715 1175 -1703
rect 1225 -1337 1271 -1325
rect 1225 -1703 1231 -1337
rect 1265 -1703 1271 -1337
rect 1225 -1715 1271 -1703
rect 1321 -1337 1367 -1325
rect 1321 -1703 1327 -1337
rect 1361 -1703 1367 -1337
rect 1321 -1715 1367 -1703
rect 1417 -1337 1463 -1325
rect 1417 -1703 1423 -1337
rect 1457 -1703 1463 -1337
rect 1417 -1715 1463 -1703
rect 1513 -1337 1559 -1325
rect 1513 -1703 1519 -1337
rect 1553 -1703 1559 -1337
rect 1513 -1715 1559 -1703
rect 1609 -1337 1655 -1325
rect 1609 -1703 1615 -1337
rect 1649 -1703 1655 -1337
rect 1609 -1715 1655 -1703
rect 1705 -1337 1751 -1325
rect 1705 -1703 1711 -1337
rect 1745 -1703 1751 -1337
rect 1705 -1715 1751 -1703
rect 1801 -1337 1847 -1325
rect 1801 -1703 1807 -1337
rect 1841 -1703 1847 -1337
rect 1801 -1715 1847 -1703
rect 1897 -1337 1943 -1325
rect 1897 -1703 1903 -1337
rect 1937 -1703 1943 -1337
rect 1897 -1715 1943 -1703
rect -1901 -1753 -1843 -1747
rect -1901 -1787 -1889 -1753
rect -1855 -1787 -1843 -1753
rect -1901 -1793 -1843 -1787
rect -1709 -1753 -1651 -1747
rect -1709 -1787 -1697 -1753
rect -1663 -1787 -1651 -1753
rect -1709 -1793 -1651 -1787
rect -1517 -1753 -1459 -1747
rect -1517 -1787 -1505 -1753
rect -1471 -1787 -1459 -1753
rect -1517 -1793 -1459 -1787
rect -1325 -1753 -1267 -1747
rect -1325 -1787 -1313 -1753
rect -1279 -1787 -1267 -1753
rect -1325 -1793 -1267 -1787
rect -1133 -1753 -1075 -1747
rect -1133 -1787 -1121 -1753
rect -1087 -1787 -1075 -1753
rect -1133 -1793 -1075 -1787
rect -941 -1753 -883 -1747
rect -941 -1787 -929 -1753
rect -895 -1787 -883 -1753
rect -941 -1793 -883 -1787
rect -749 -1753 -691 -1747
rect -749 -1787 -737 -1753
rect -703 -1787 -691 -1753
rect -749 -1793 -691 -1787
rect -557 -1753 -499 -1747
rect -557 -1787 -545 -1753
rect -511 -1787 -499 -1753
rect -557 -1793 -499 -1787
rect -365 -1753 -307 -1747
rect -365 -1787 -353 -1753
rect -319 -1787 -307 -1753
rect -365 -1793 -307 -1787
rect -173 -1753 -115 -1747
rect -173 -1787 -161 -1753
rect -127 -1787 -115 -1753
rect -173 -1793 -115 -1787
rect 19 -1753 77 -1747
rect 19 -1787 31 -1753
rect 65 -1787 77 -1753
rect 19 -1793 77 -1787
rect 211 -1753 269 -1747
rect 211 -1787 223 -1753
rect 257 -1787 269 -1753
rect 211 -1793 269 -1787
rect 403 -1753 461 -1747
rect 403 -1787 415 -1753
rect 449 -1787 461 -1753
rect 403 -1793 461 -1787
rect 595 -1753 653 -1747
rect 595 -1787 607 -1753
rect 641 -1787 653 -1753
rect 595 -1793 653 -1787
rect 787 -1753 845 -1747
rect 787 -1787 799 -1753
rect 833 -1787 845 -1753
rect 787 -1793 845 -1787
rect 979 -1753 1037 -1747
rect 979 -1787 991 -1753
rect 1025 -1787 1037 -1753
rect 979 -1793 1037 -1787
rect 1171 -1753 1229 -1747
rect 1171 -1787 1183 -1753
rect 1217 -1787 1229 -1753
rect 1171 -1793 1229 -1787
rect 1363 -1753 1421 -1747
rect 1363 -1787 1375 -1753
rect 1409 -1787 1421 -1753
rect 1363 -1793 1421 -1787
rect 1555 -1753 1613 -1747
rect 1555 -1787 1567 -1753
rect 1601 -1787 1613 -1753
rect 1555 -1793 1613 -1787
rect 1747 -1753 1805 -1747
rect 1747 -1787 1759 -1753
rect 1793 -1787 1805 -1753
rect 1747 -1793 1805 -1787
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -2034 -1872 2034 1872
string parameters w 1.95 l 0.150 m 6 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
