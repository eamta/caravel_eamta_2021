magic
tech sky130A
magscale 1 2
timestamp 1623262251
<< nwell >>
rect -54 3270 3993 3545
<< nsubdiff >>
rect 54 3337 78 3509
rect 3860 3337 3884 3509
<< nsubdiffcont >>
rect 78 3337 3860 3509
<< locali >>
rect 62 3337 78 3509
rect 3860 3337 3876 3509
<< viali >>
rect 78 3337 3860 3509
rect 78 3245 3860 3279
rect -18 80 16 3182
rect 3922 80 3956 3182
rect 78 -377 2068 -343
rect -18 -3542 16 -440
rect 2130 -3542 2164 -440
<< metal1 >>
rect -24 3509 3962 3515
rect -24 3337 78 3509
rect 3860 3337 3962 3509
rect -24 3279 3962 3337
rect -24 3245 78 3279
rect 3860 3245 3962 3279
rect -24 3239 3962 3245
rect -24 3182 22 3239
rect -24 80 -18 3182
rect 16 80 22 3182
rect 218 3154 264 3239
rect 474 3164 520 3239
rect 730 3165 776 3239
rect 986 3163 1032 3239
rect 1242 3163 1288 3239
rect 1498 3162 1544 3239
rect 1754 3164 1800 3239
rect 2010 3163 2056 3239
rect 2266 3163 2312 3239
rect 2522 3163 2568 3239
rect 2778 3164 2824 3239
rect 3034 3162 3080 3239
rect 3290 3163 3336 3239
rect 3546 3162 3592 3239
rect 3802 3164 3848 3239
rect 3916 3182 3962 3239
rect -24 68 22 80
rect 90 126 136 212
rect 346 126 392 240
rect 602 126 648 243
rect 858 126 904 245
rect 1114 126 1160 245
rect 1370 126 1416 246
rect 1626 126 1672 241
rect 1882 126 1928 244
rect 2137 126 2184 187
rect 2393 126 2440 186
rect 2649 126 2696 195
rect 2905 126 2952 190
rect 3162 126 3209 191
rect 3418 126 3465 194
rect 3674 126 3721 193
rect 90 -120 3796 126
rect 3916 80 3922 3182
rect 3956 80 3962 3182
rect 3916 68 3962 80
rect 90 -239 3222 -120
rect -24 -343 3222 -239
rect -24 -377 78 -343
rect 2068 -377 3222 -343
rect -24 -383 3222 -377
rect -24 -440 22 -383
rect -24 -3542 -18 -440
rect 16 -3542 22 -440
rect 90 -413 3222 -383
rect 3796 -413 3806 -120
rect 90 -494 136 -413
rect 346 -466 392 -413
rect 602 -463 648 -413
rect 858 -461 904 -413
rect 1114 -461 1160 -413
rect 1370 -460 1416 -413
rect 1626 -465 1672 -413
rect 1882 -462 1928 -413
rect 2124 -440 2170 -413
rect 218 -3495 264 -3450
rect 474 -3495 520 -3449
rect 730 -3495 776 -3452
rect 986 -3495 1032 -3452
rect 1242 -3495 1288 -3450
rect 1498 -3495 1544 -3450
rect 1754 -3495 1800 -3450
rect 2010 -3495 2056 -3451
rect -24 -3554 22 -3542
rect 142 -3682 2056 -3495
rect 2124 -3542 2130 -440
rect 2164 -3542 2170 -440
rect 2124 -3554 2170 -3542
rect 2344 -3682 2354 -3254
rect 142 -3948 2354 -3682
rect 2686 -3948 2696 -3254
<< via1 >>
rect 3222 -413 3796 -120
rect 2354 -3948 2686 -3254
<< metal2 >>
rect 3222 -120 3796 -110
rect 3222 -423 3796 -413
rect 2354 -3254 2686 -3244
rect 2354 -3958 2686 -3948
use sky130_fd_pr__pfet_01v8_lvt_NRCKZ4  M7
timestamp 1623256316
transform 1 0 1073 0 1 -1991
box -1127 -1684 1127 1684
use sky130_fd_pr__pfet_01v8_lvt_NRU274  M8
timestamp 1623255091
transform 1 0 1969 0 1 1631
box -2023 -1684 2023 1684
<< labels >>
rlabel via1 2354 -3948 2686 -3254 1 ibias
rlabel via1 3222 -413 3796 -120 1 vbias_1
rlabel nwell 78 3337 3860 3509 1 vdd
<< end >>
