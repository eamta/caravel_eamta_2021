magic
tech sky130A
magscale 1 2
timestamp 1616617991
<< error_p >>
rect -70 50 -10 5750
rect 10 50 70 5750
rect -70 -5750 -10 -50
rect 10 -5750 70 -50
<< metal3 >>
rect -6309 5722 -10 5750
rect -6309 78 -94 5722
rect -30 78 -10 5722
rect -6309 50 -10 78
rect 10 5722 6309 5750
rect 10 78 6225 5722
rect 6289 78 6309 5722
rect 10 50 6309 78
rect -6309 -78 -10 -50
rect -6309 -5722 -94 -78
rect -30 -5722 -10 -78
rect -6309 -5750 -10 -5722
rect 10 -78 6309 -50
rect 10 -5722 6225 -78
rect 6289 -5722 6309 -78
rect 10 -5750 6309 -5722
<< via3 >>
rect -94 78 -30 5722
rect 6225 78 6289 5722
rect -94 -5722 -30 -78
rect 6225 -5722 6289 -78
<< mimcap >>
rect -6209 5610 -209 5650
rect -6209 190 -6169 5610
rect -249 190 -209 5610
rect -6209 150 -209 190
rect 110 5610 6110 5650
rect 110 190 150 5610
rect 6070 190 6110 5610
rect 110 150 6110 190
rect -6209 -190 -209 -150
rect -6209 -5610 -6169 -190
rect -249 -5610 -209 -190
rect -6209 -5650 -209 -5610
rect 110 -190 6110 -150
rect 110 -5610 150 -190
rect 6070 -5610 6110 -190
rect 110 -5650 6110 -5610
<< mimcapcontact >>
rect -6169 190 -249 5610
rect 150 190 6070 5610
rect -6169 -5610 -249 -190
rect 150 -5610 6070 -190
<< metal4 >>
rect -3261 5611 -3157 5800
rect -141 5738 -37 5800
rect -141 5722 -14 5738
rect -6170 5610 -248 5611
rect -6170 190 -6169 5610
rect -249 190 -248 5610
rect -6170 189 -248 190
rect -3261 -189 -3157 189
rect -141 78 -94 5722
rect -30 78 -14 5722
rect 3058 5611 3162 5800
rect 6178 5738 6282 5800
rect 6178 5722 6305 5738
rect 149 5610 6071 5611
rect 149 190 150 5610
rect 6070 190 6071 5610
rect 149 189 6071 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -6170 -190 -248 -189
rect -6170 -5610 -6169 -190
rect -249 -5610 -248 -190
rect -6170 -5611 -248 -5610
rect -3261 -5800 -3157 -5611
rect -141 -5722 -94 -78
rect -30 -5722 -14 -78
rect 3058 -189 3162 189
rect 6178 78 6225 5722
rect 6289 78 6305 5722
rect 6178 62 6305 78
rect 6178 -62 6282 62
rect 6178 -78 6305 -62
rect 149 -190 6071 -189
rect 149 -5610 150 -190
rect 6070 -5610 6071 -190
rect 149 -5611 6071 -5610
rect -141 -5738 -14 -5722
rect -141 -5800 -37 -5738
rect 3058 -5800 3162 -5611
rect 6178 -5722 6225 -78
rect 6289 -5722 6305 -78
rect 6178 -5738 6305 -5722
rect 6178 -5800 6282 -5738
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 10 50 6210 5750
string parameters w 30 l 27.5 val 844.55 carea 1.00 cperi 0.17 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
