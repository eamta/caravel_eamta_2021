magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 383 2192 436 2193
rect 2099 2192 2152 2193
rect 3815 2192 3868 2193
rect 5531 2192 5584 2193
rect 365 2158 436 2192
rect 2081 2158 2152 2192
rect 3797 2158 3868 2192
rect 5513 2158 5584 2192
rect 366 2157 436 2158
rect 2082 2157 2152 2158
rect 3798 2157 3868 2158
rect 5514 2157 5584 2158
rect 383 2123 454 2157
rect 734 2123 769 2140
rect 191 1871 204 2018
rect 219 1899 232 2046
rect 196 1800 254 1806
rect 196 1766 208 1800
rect 196 1760 254 1766
rect 383 1717 453 2123
rect 735 2122 769 2123
rect 2099 2123 2170 2157
rect 2450 2123 2485 2140
rect 735 2086 805 2122
rect 2099 2096 2169 2123
rect 1912 2090 1970 2096
rect 1121 2086 1174 2087
rect 565 2055 623 2061
rect 565 2021 577 2055
rect 752 2052 823 2086
rect 1103 2052 1174 2086
rect 565 2015 623 2021
rect 50 1698 84 1716
rect 366 1698 453 1717
rect 565 1747 623 1753
rect 565 1713 577 1747
rect 752 1734 822 2052
rect 1104 2051 1174 2052
rect 1912 2056 1924 2090
rect 1121 2017 1192 2051
rect 1472 2017 1507 2051
rect 1912 2050 1970 2056
rect 1121 1990 1191 2017
rect 1473 1998 1507 2017
rect 934 1984 992 1990
rect 934 1950 946 1984
rect 934 1944 992 1950
rect 890 1734 930 1752
rect 996 1734 1036 1752
rect 1104 1735 1191 1990
rect 1303 1949 1361 1955
rect 1303 1915 1315 1949
rect 1303 1909 1361 1915
rect 1492 1735 1507 1998
rect 1526 1964 1561 1998
rect 1526 1735 1560 1964
rect 1730 1902 1912 2034
rect 1672 1896 1912 1902
rect 1672 1862 1684 1896
rect 1730 1891 1912 1896
rect 1730 1868 1926 1891
rect 1730 1862 1929 1868
rect 1672 1856 1929 1862
rect 1730 1838 1929 1856
rect 1956 1838 2014 1891
rect 2082 1873 2169 2096
rect 2451 2122 2485 2123
rect 3815 2123 3886 2157
rect 4166 2123 4201 2140
rect 2451 2086 2521 2122
rect 3815 2096 3885 2123
rect 3628 2090 3686 2096
rect 2837 2086 2890 2087
rect 2281 2055 2339 2061
rect 2281 2021 2293 2055
rect 2468 2052 2539 2086
rect 2819 2052 2890 2086
rect 2281 2015 2339 2021
rect 1730 1837 1912 1838
rect 1914 1837 1929 1838
rect 2082 1837 2281 1873
rect 1730 1803 2281 1837
rect 1728 1800 1970 1803
rect 1728 1769 1974 1800
rect 1728 1766 1929 1769
rect 1728 1760 1970 1766
rect 1728 1735 1929 1760
rect 2082 1753 2281 1803
rect 2082 1747 2339 1753
rect 2082 1741 2293 1747
rect 1104 1734 1929 1735
rect 565 1707 623 1713
rect 752 1698 1929 1734
rect 2041 1735 2293 1741
rect 2468 1735 2538 2052
rect 2820 2051 2890 2052
rect 3628 2056 3640 2090
rect 2837 2017 2908 2051
rect 3188 2017 3223 2051
rect 3628 2050 3686 2056
rect 2837 1990 2907 2017
rect 3189 1998 3223 2017
rect 2650 1984 2708 1990
rect 2650 1950 2662 1984
rect 2650 1944 2708 1950
rect 2041 1732 2053 1735
rect 2082 1734 2538 1735
rect 2606 1734 2646 1752
rect 2712 1734 2752 1752
rect 2820 1735 2907 1990
rect 3208 1735 3223 1998
rect 3242 1964 3277 1998
rect 3242 1735 3276 1964
rect 3446 1902 3628 2034
rect 3388 1896 3628 1902
rect 3388 1862 3400 1896
rect 3446 1891 3628 1896
rect 3446 1868 3642 1891
rect 3446 1862 3645 1868
rect 3388 1856 3645 1862
rect 3446 1838 3645 1856
rect 3672 1838 3730 1891
rect 3798 1873 3885 2096
rect 4167 2122 4201 2123
rect 5531 2123 5602 2157
rect 5882 2123 5917 2140
rect 4167 2086 4237 2122
rect 5531 2096 5601 2123
rect 5344 2090 5402 2096
rect 4553 2086 4606 2087
rect 3997 2055 4055 2061
rect 3997 2021 4009 2055
rect 4184 2052 4255 2086
rect 4535 2052 4606 2086
rect 3997 2015 4055 2021
rect 3446 1837 3628 1838
rect 3630 1837 3645 1838
rect 3798 1837 3997 1873
rect 3446 1803 3997 1837
rect 3446 1800 3686 1803
rect 3446 1769 3690 1800
rect 3446 1766 3645 1769
rect 3446 1760 3686 1766
rect 3446 1735 3645 1760
rect 3798 1753 3997 1803
rect 3798 1747 4055 1753
rect 3798 1741 4009 1747
rect 2820 1734 3645 1735
rect 2082 1732 3645 1734
rect 3757 1735 4009 1741
rect 4184 1735 4254 2052
rect 4536 2051 4606 2052
rect 5344 2056 5356 2090
rect 4553 2017 4624 2051
rect 4904 2017 4939 2051
rect 5344 2050 5402 2056
rect 4366 1984 4424 1990
rect 4366 1950 4378 1984
rect 4366 1944 4424 1950
rect 3757 1732 3769 1735
rect 3798 1734 4254 1735
rect 4322 1734 4362 1753
rect 4428 1734 4468 1753
rect 4553 1735 4623 2017
rect 4905 1998 4939 2017
rect 4735 1949 4793 1955
rect 4735 1915 4747 1949
rect 4735 1909 4793 1915
rect 4924 1735 4939 1998
rect 4958 1964 4993 1998
rect 4958 1735 4992 1964
rect 5162 1902 5344 2034
rect 5104 1896 5344 1902
rect 5104 1862 5116 1896
rect 5162 1891 5344 1896
rect 5162 1868 5358 1891
rect 5162 1862 5361 1868
rect 5104 1856 5361 1862
rect 5162 1838 5361 1856
rect 5388 1838 5446 1891
rect 5514 1873 5601 2096
rect 5883 2122 5917 2123
rect 5883 2086 5953 2122
rect 6269 2086 6322 2087
rect 5713 2055 5771 2061
rect 5713 2021 5725 2055
rect 5900 2052 5971 2086
rect 6251 2052 6322 2086
rect 5713 2015 5771 2021
rect 5162 1837 5344 1838
rect 5346 1837 5361 1838
rect 5514 1837 5713 1873
rect 5162 1803 5713 1837
rect 5162 1800 5402 1803
rect 5162 1769 5406 1800
rect 5162 1766 5361 1769
rect 5162 1760 5402 1766
rect 5162 1735 5361 1760
rect 5514 1753 5713 1803
rect 5514 1747 5771 1753
rect 5514 1741 5725 1747
rect 4553 1734 5361 1735
rect 3798 1732 5361 1734
rect 5473 1735 5725 1741
rect 5473 1732 5485 1735
rect 5514 1732 5725 1735
rect 2037 1701 3645 1732
rect 3753 1701 5361 1732
rect 5469 1713 5725 1732
rect 5900 1734 5970 2052
rect 6252 2051 6322 2052
rect 6269 2017 6340 2051
rect 6620 2017 6655 2051
rect 6082 1984 6140 1990
rect 6082 1950 6094 1984
rect 6082 1944 6140 1950
rect 6038 1734 6078 1752
rect 6144 1734 6184 1752
rect 6269 1734 6339 2017
rect 6621 1998 6655 2017
rect 6451 1949 6509 1955
rect 6451 1915 6463 1949
rect 6451 1909 6509 1915
rect 5469 1707 5771 1713
rect 5469 1701 5713 1707
rect 2041 1698 3645 1701
rect 3757 1698 5361 1701
rect 5473 1698 5713 1701
rect 50 1666 5713 1698
rect 50 1664 3344 1666
rect 3356 1664 3390 1666
rect 3444 1664 5713 1666
rect 383 1663 1929 1664
rect 2009 1663 2043 1664
rect 39 1628 264 1662
rect 319 1661 1929 1663
rect 1997 1661 2055 1663
rect 2063 1661 3277 1664
rect 319 1646 3277 1661
rect 3344 1646 5361 1664
rect 5531 1663 5713 1664
rect 319 1639 5361 1646
rect 5429 1639 5487 1663
rect 5517 1639 5713 1663
rect 319 1628 2000 1639
rect 383 1626 2000 1628
rect 383 1616 1942 1626
rect 382 1615 1942 1616
rect 49 1594 1942 1615
rect 2009 1597 2043 1639
rect 2055 1629 5361 1639
rect 2055 1627 3277 1629
rect 3446 1628 3645 1629
rect 2097 1624 3277 1627
rect 3487 1624 3658 1628
rect 2097 1597 3658 1624
rect 239 1592 1942 1594
rect 228 1587 1942 1592
rect 228 1581 280 1587
rect 364 1581 1942 1587
rect 365 1580 1942 1581
rect 382 1575 1942 1580
rect 1997 1589 2043 1597
rect 2082 1593 3658 1597
rect 3713 1627 3728 1629
rect 3815 1628 5361 1629
rect 3713 1618 3759 1627
rect 3713 1593 3721 1618
rect 3725 1593 3759 1618
rect 3815 1593 5374 1628
rect 1997 1588 2038 1589
rect 1997 1581 2037 1588
rect 1997 1575 2043 1581
rect 2082 1575 5374 1593
rect 5429 1575 5469 1593
rect 5531 1575 5713 1639
rect 5900 1630 6339 1734
rect 6407 1688 6447 1699
rect 6513 1688 6553 1699
rect 6640 1683 6655 1998
rect 6674 1964 6709 1998
rect 6674 1683 6708 1964
rect 6820 1896 6878 1902
rect 6820 1862 6832 1896
rect 6990 1873 7024 1891
rect 6820 1856 6878 1862
rect 6990 1837 7060 1873
rect 7007 1803 7078 1837
rect 7007 1736 7077 1803
rect 6941 1700 7077 1736
rect 7189 1735 7247 1741
rect 7189 1734 7201 1735
rect 7185 1701 7251 1734
rect 7189 1700 7247 1701
rect 6941 1683 7327 1700
rect 6429 1645 6531 1675
rect 6572 1666 7327 1683
rect 6572 1645 7077 1666
rect 7259 1663 7279 1666
rect 6369 1630 7077 1645
rect 7145 1641 7203 1663
rect 7233 1641 7291 1663
rect 5900 1628 7077 1630
rect 7157 1632 7195 1636
rect 7157 1629 7203 1632
rect 5900 1577 7090 1628
rect 7145 1623 7203 1629
rect 7145 1619 7207 1623
rect 7135 1598 7207 1619
rect 5834 1575 7090 1577
rect 7135 1575 7137 1577
rect 7145 1575 7207 1598
rect 7259 1593 7291 1641
rect 7251 1575 7291 1593
rect 7293 1575 7327 1666
rect 7359 1575 7381 1754
rect 382 1573 2311 1575
rect 49 1481 83 1573
rect 157 1519 169 1523
rect 365 1522 2311 1573
rect 2323 1522 2329 1563
rect 2498 1522 4027 1575
rect 4034 1522 4047 1544
rect 4050 1522 4097 1552
rect 4174 1522 4205 1548
rect 4208 1524 5713 1575
rect 5930 1541 7429 1575
rect 4208 1522 5743 1524
rect 5870 1522 7429 1541
rect 157 1513 181 1519
rect 195 1513 203 1519
rect 157 1501 175 1513
rect 157 1481 169 1501
rect 176 1481 181 1513
rect 191 1481 203 1513
rect 207 1481 253 1513
rect 365 1481 7429 1522
rect 1 1363 7429 1481
rect 7442 1452 7477 1486
rect 7757 1452 7792 1486
rect 1 1352 7363 1363
rect 1 1351 4653 1352
rect 1 1271 1221 1351
rect 1289 1350 1435 1351
rect 1298 1340 1435 1350
rect 1472 1340 1590 1351
rect 1298 1338 1590 1340
rect 1298 1323 1347 1338
rect 1291 1322 1347 1323
rect 1291 1312 1346 1322
rect 1355 1312 1367 1338
rect 1383 1337 1590 1338
rect 1383 1324 1457 1337
rect 1472 1336 1590 1337
rect 1462 1332 1590 1336
rect 1383 1312 1461 1324
rect 1270 1301 1461 1312
rect 1245 1297 1255 1301
rect 13 1205 486 1271
rect 520 1241 578 1271
rect 608 1241 617 1271
rect 520 1217 529 1241
rect 532 1229 567 1241
rect 625 1229 654 1271
rect 521 1205 529 1217
rect 533 1217 567 1229
rect 629 1223 654 1229
rect 626 1217 654 1223
rect 533 1205 579 1217
rect 629 1213 657 1217
rect 13 1156 491 1205
rect 499 1191 579 1205
rect 499 1186 567 1191
rect 578 1186 579 1191
rect 499 1170 579 1186
rect 595 1170 622 1176
rect 651 1170 657 1213
rect 663 1196 692 1271
rect 734 1222 1221 1271
rect 1233 1285 1266 1297
rect 1267 1295 1346 1301
rect 1355 1296 1461 1301
rect 1275 1285 1346 1295
rect 1347 1291 1461 1296
rect 1347 1285 1377 1291
rect 1233 1279 1377 1285
rect 1392 1290 1461 1291
rect 1392 1282 1457 1290
rect 1390 1279 1426 1282
rect 1233 1278 1426 1279
rect 1233 1275 1310 1278
rect 1327 1275 1404 1278
rect 1418 1275 1426 1278
rect 1428 1275 1457 1282
rect 1472 1275 1590 1332
rect 1605 1325 1619 1351
rect 1599 1275 1619 1325
rect 1633 1319 1647 1351
rect 1649 1328 1991 1351
rect 2036 1347 2328 1351
rect 2036 1344 2081 1347
rect 1649 1324 2028 1328
rect 2039 1324 2081 1344
rect 2121 1344 2166 1347
rect 2121 1340 2161 1344
rect 2215 1340 2275 1347
rect 2121 1337 2195 1340
rect 1649 1319 2081 1324
rect 1633 1301 2081 1319
rect 1633 1297 1647 1301
rect 1627 1285 1647 1297
rect 1667 1296 2081 1301
rect 2127 1336 2195 1337
rect 2215 1336 2283 1340
rect 2294 1336 2328 1347
rect 2127 1322 2207 1336
rect 2215 1324 2328 1336
rect 2351 1347 2369 1351
rect 2379 1347 4653 1351
rect 2351 1329 4653 1347
rect 4687 1341 7363 1352
rect 4685 1329 7363 1341
rect 2351 1325 4676 1329
rect 2237 1322 2328 1324
rect 2127 1296 2195 1322
rect 2239 1313 2328 1322
rect 2201 1298 2328 1313
rect 2239 1296 2328 1298
rect 1667 1294 2328 1296
rect 1667 1285 1792 1294
rect 1627 1283 1716 1285
rect 1724 1283 1729 1285
rect 1627 1279 1743 1283
rect 1627 1275 1749 1279
rect 1233 1269 1749 1275
rect 1233 1259 1667 1269
rect 1670 1259 1749 1269
rect 1752 1259 1792 1285
rect 1823 1283 2328 1294
rect 1233 1242 1792 1259
rect 1233 1241 1667 1242
rect 1670 1241 1792 1242
rect 1233 1222 1413 1241
rect 734 1201 1413 1222
rect 663 1179 709 1196
rect 499 1169 657 1170
rect 675 1169 709 1179
rect 734 1193 1398 1201
rect 734 1188 1404 1193
rect 734 1169 1221 1188
rect 499 1156 1221 1169
rect 13 1151 452 1156
rect 479 1155 487 1156
rect 453 1151 486 1152
rect 560 1151 1221 1156
rect 13 1128 499 1151
rect 545 1139 1221 1151
rect 1233 1139 1404 1188
rect 13 1116 452 1128
rect 453 1116 486 1128
rect 491 1116 499 1128
rect 541 1135 1221 1139
rect 541 1130 703 1135
rect 541 1116 605 1130
rect 617 1129 703 1130
rect 617 1120 663 1129
rect 13 1098 605 1116
rect 623 1102 663 1120
rect 683 1117 703 1129
rect 709 1133 1221 1135
rect 1229 1133 1404 1139
rect 1418 1133 1426 1241
rect 1472 1232 1590 1241
rect 1436 1207 1590 1232
rect 1452 1182 1590 1207
rect 1465 1177 1590 1182
rect 1467 1167 1590 1177
rect 1436 1165 1590 1167
rect 1427 1139 1590 1165
rect 1427 1133 1451 1139
rect 1455 1134 1590 1139
rect 1455 1133 1591 1134
rect 709 1131 1591 1133
rect 709 1130 1404 1131
rect 1417 1130 1591 1131
rect 709 1117 1591 1130
rect 1599 1117 1619 1241
rect 1625 1226 1667 1241
rect 1678 1238 1792 1241
rect 1678 1226 1746 1238
rect 1755 1229 1792 1238
rect 1797 1279 2328 1283
rect 1797 1260 1831 1279
rect 1835 1260 2328 1279
rect 1755 1226 1795 1229
rect 1625 1134 1673 1226
rect 1621 1129 1673 1134
rect 1678 1225 1795 1226
rect 1678 1216 1767 1225
rect 1678 1148 1782 1216
rect 1783 1149 1795 1225
rect 1797 1176 2328 1260
rect 1797 1149 1831 1176
rect 1835 1152 2328 1176
rect 1678 1129 1767 1148
rect 1783 1144 1831 1149
rect 1781 1133 1831 1144
rect 1621 1117 1767 1129
rect 683 1113 697 1117
rect 709 1114 1579 1117
rect 13 1082 552 1098
rect 13 1068 452 1082
rect 453 1068 487 1082
rect 491 1068 499 1082
rect 518 1068 552 1082
rect 571 1068 605 1098
rect 629 1068 663 1102
rect 704 1101 1579 1114
rect 695 1099 1579 1101
rect 672 1068 1224 1099
rect 13 1051 1224 1068
rect 135 1013 157 1016
rect 35 986 157 1013
rect 165 986 181 1051
rect 35 971 181 986
rect 202 1020 206 1051
rect 230 1039 237 1051
rect 291 1039 296 1051
rect 325 1048 411 1051
rect 418 1048 1224 1051
rect 225 1028 236 1039
rect 325 1035 1224 1048
rect 353 1034 1224 1035
rect 353 1030 428 1034
rect 353 1020 441 1030
rect 43 966 93 971
rect 101 966 123 971
rect 135 967 157 971
rect 168 967 169 971
rect 43 945 123 966
rect 43 932 93 945
rect 101 942 165 945
rect 101 933 195 942
rect 123 923 195 933
rect 202 928 236 1020
rect 348 1014 441 1020
rect 344 1001 441 1014
rect 353 995 441 1001
rect 344 992 441 995
rect 453 992 483 995
rect 344 986 483 992
rect 484 986 487 1034
rect 491 986 499 1034
rect 344 980 499 986
rect 353 971 499 980
rect 518 971 552 1034
rect 365 967 410 971
rect 392 964 410 967
rect 411 964 441 971
rect 453 967 483 971
rect 484 967 487 971
rect 411 961 434 964
rect 253 928 283 942
rect 202 923 295 928
rect 115 921 304 923
rect 331 921 350 937
rect 365 933 449 961
rect 365 928 450 933
rect 115 916 350 921
rect 123 903 350 916
rect 356 921 450 928
rect 453 921 477 967
rect 356 909 477 921
rect 518 914 529 971
rect 537 914 552 967
rect 356 903 467 909
rect 115 902 467 903
rect 115 900 362 902
rect 365 900 467 902
rect 115 893 467 900
rect 115 879 450 893
rect 115 874 365 879
rect 107 873 165 874
rect 173 873 253 874
rect 283 873 363 874
rect 392 873 452 879
rect 107 862 122 873
rect 173 862 236 873
rect 304 862 363 873
rect 69 828 246 862
rect 295 861 363 862
rect 404 868 452 873
rect 404 861 477 868
rect 295 852 477 861
rect 518 860 552 914
rect 571 860 605 1034
rect 629 1024 1224 1034
rect 1256 1025 1343 1099
rect 1418 1096 1426 1099
rect 1469 1096 1579 1099
rect 1580 1096 1619 1117
rect 1418 1092 1590 1096
rect 1411 1084 1590 1092
rect 1599 1089 1619 1096
rect 1411 1080 1593 1084
rect 1605 1080 1619 1089
rect 1625 1080 1767 1117
rect 1783 1081 1831 1133
rect 1786 1080 1831 1081
rect 1838 1089 2328 1152
rect 2345 1318 4676 1325
rect 2345 1297 4665 1318
rect 4685 1297 4711 1329
rect 4712 1297 7363 1329
rect 2345 1202 7363 1297
rect 7408 1202 7423 1363
rect 7442 1202 7476 1452
rect 7758 1433 7792 1452
rect 7588 1384 7646 1390
rect 7588 1350 7600 1384
rect 7588 1344 7646 1350
rect 2345 1167 7588 1202
rect 2345 1149 7602 1167
rect 7632 1149 7690 1167
rect 7777 1149 7792 1433
rect 7811 1399 7846 1433
rect 8126 1399 8161 1416
rect 7811 1149 7845 1399
rect 8127 1398 8161 1399
rect 8127 1362 8197 1398
rect 7957 1331 8015 1337
rect 7957 1297 7969 1331
rect 8144 1328 8215 1362
rect 8495 1328 8530 1362
rect 7957 1291 8015 1297
rect 8144 1186 8214 1328
rect 8496 1309 8530 1328
rect 8515 1266 8530 1309
rect 8326 1260 8384 1266
rect 8326 1226 8338 1260
rect 8326 1220 8384 1226
rect 7904 1149 8214 1186
rect 2345 1121 8214 1149
rect 1838 1080 2283 1089
rect 1411 1069 2283 1080
rect 1348 1030 1377 1064
rect 1411 1057 1621 1069
rect 1625 1057 2283 1069
rect 1423 1046 2283 1057
rect 1423 1034 1559 1046
rect 1393 1025 1559 1034
rect 1576 1025 1593 1046
rect 1605 1030 1619 1046
rect 1625 1045 1659 1046
rect 1678 1045 1746 1046
rect 1625 1025 1751 1045
rect 1786 1030 1831 1046
rect 629 1002 1221 1024
rect 629 983 669 1002
rect 709 1001 1221 1002
rect 685 986 1221 1001
rect 679 985 1221 986
rect 629 967 639 983
rect 651 971 669 983
rect 675 974 1221 985
rect 679 971 1221 974
rect 651 909 663 971
rect 675 968 1221 971
rect 675 945 731 968
rect 739 967 1221 968
rect 751 962 1221 967
rect 1256 1014 1364 1025
rect 1256 962 1343 1014
rect 1393 1013 1751 1025
rect 1792 1013 1831 1030
rect 1838 1014 2283 1046
rect 2294 1018 2328 1089
rect 2335 1117 8214 1121
rect 2335 1105 2362 1117
rect 2363 1105 8214 1117
rect 8260 1116 8290 1150
rect 2335 1091 8214 1105
rect 2335 1090 2362 1091
rect 2363 1090 8214 1091
rect 1838 1013 2280 1014
rect 1393 1011 2280 1013
rect 1411 997 1559 1011
rect 1576 997 1593 1011
rect 1625 997 1659 1011
rect 1667 997 2280 1011
rect 1362 983 1396 996
rect 1411 983 2280 997
rect 1346 971 1559 983
rect 1576 971 1593 983
rect 1346 967 1589 971
rect 1346 962 1381 967
rect 1385 962 1589 967
rect 751 945 1589 962
rect 679 918 731 945
rect 773 933 807 945
rect 673 861 731 918
rect 778 903 807 933
rect 812 944 845 945
rect 812 928 841 944
rect 847 928 878 945
rect 881 929 975 945
rect 1005 933 1088 945
rect 981 929 1088 933
rect 1123 937 1589 945
rect 1123 929 1188 937
rect 1203 929 1589 937
rect 812 903 819 928
rect 761 873 819 903
rect 856 877 862 928
rect 881 924 1027 929
rect 1035 928 1589 929
rect 881 917 1020 924
rect 1035 917 1188 928
rect 881 914 1015 917
rect 881 908 974 914
rect 975 908 1008 914
rect 884 905 921 908
rect 804 861 819 873
rect 887 873 921 905
rect 887 862 898 873
rect 629 860 731 861
rect 518 852 521 860
rect 107 759 108 828
rect 164 781 165 785
rect 202 781 241 828
rect 295 827 490 852
rect 119 759 241 781
rect 252 759 253 785
rect 295 765 363 827
rect 404 784 438 827
rect 450 788 490 827
rect 445 784 490 788
rect 491 806 521 852
rect 530 852 552 860
rect 564 852 731 860
rect 773 852 819 861
rect 530 839 731 852
rect 751 845 819 852
rect 906 851 921 873
rect 887 845 921 851
rect 751 839 921 845
rect 530 826 921 839
rect 530 806 605 826
rect 491 784 605 806
rect 404 781 472 784
rect 475 781 491 784
rect 499 781 567 784
rect 571 781 605 784
rect 404 765 605 781
rect 295 759 362 765
rect 107 753 362 759
rect 107 694 409 753
rect 410 749 605 765
rect 651 750 659 826
rect 663 821 921 826
rect 663 818 819 821
rect 673 817 819 818
rect 673 806 885 817
rect 717 802 719 806
rect 739 797 764 806
rect 785 802 885 806
rect 797 801 885 802
rect 791 797 885 801
rect 691 793 697 797
rect 679 750 703 793
rect 717 759 731 765
rect 739 759 885 797
rect 713 751 885 759
rect 713 750 865 751
rect 651 749 865 750
rect 410 700 420 749
rect 432 719 605 749
rect 679 745 703 749
rect 432 694 601 719
rect 194 668 195 694
rect 202 604 240 694
rect 260 681 267 694
rect 260 646 266 681
rect 282 668 283 694
rect 288 653 295 694
rect 288 646 294 653
rect 310 646 340 694
rect 344 687 387 694
rect 344 674 394 687
rect 432 674 478 694
rect 344 672 410 674
rect 432 672 493 674
rect 348 666 406 672
rect 345 646 432 666
rect 310 640 434 646
rect 444 640 493 672
rect 310 638 493 640
rect 264 625 294 638
rect 322 634 328 638
rect 264 604 328 625
rect 371 606 493 638
rect 518 666 601 694
rect 689 691 703 745
rect 713 725 763 749
rect 717 719 731 725
rect 887 717 921 821
rect 887 692 896 717
rect 444 604 490 606
rect 518 604 566 666
rect 571 656 601 666
rect 887 681 898 692
rect 906 681 921 717
rect 887 657 921 681
rect 940 873 1008 908
rect 940 764 975 873
rect 981 764 1008 873
rect 1042 871 1210 917
rect 1042 859 1188 871
rect 1211 868 1221 928
rect 1233 911 1290 928
rect 1239 905 1290 911
rect 1239 868 1249 905
rect 1100 846 1115 859
rect 1145 850 1148 859
rect 1132 846 1170 850
rect 1064 812 1069 846
rect 1100 828 1182 846
rect 1082 821 1182 828
rect 1082 818 1115 821
rect 1132 818 1182 821
rect 1082 778 1182 818
rect 1082 764 1115 778
rect 1123 772 1144 778
rect 940 750 1115 764
rect 1145 764 1148 778
rect 1151 764 1182 778
rect 1189 764 1203 766
rect 1256 765 1290 905
rect 1309 917 1343 928
rect 1346 917 1379 928
rect 1389 917 1412 928
rect 1423 924 1457 928
rect 1423 917 1446 924
rect 1309 861 1379 917
rect 1411 915 1446 917
rect 1477 916 1495 928
rect 1501 927 1589 928
rect 1499 916 1589 927
rect 1411 912 1451 915
rect 1477 912 1489 916
rect 1499 912 1577 916
rect 1423 908 1446 912
rect 1501 909 1559 912
rect 1625 909 1659 983
rect 1667 977 2280 983
rect 1678 966 2280 977
rect 1678 963 1749 966
rect 1678 919 1755 963
rect 1773 943 1777 966
rect 1785 943 2280 966
rect 2294 993 2329 1018
rect 2335 1010 8214 1090
rect 2335 997 6867 1010
rect 2294 974 2328 993
rect 2335 976 6498 997
rect 6540 996 6574 997
rect 6588 996 6627 997
rect 6540 980 6631 996
rect 2335 974 6494 976
rect 2294 959 2309 974
rect 1678 915 1743 919
rect 1773 918 2280 943
rect 2323 951 6494 974
rect 2323 943 6498 951
rect 2323 941 5354 943
rect 5433 941 5442 943
rect 2323 940 5386 941
rect 2363 931 5386 940
rect 1773 916 1820 918
rect 1797 915 1827 916
rect 1678 909 1712 915
rect 1820 909 1827 915
rect 1836 909 2280 918
rect 1501 907 2280 909
rect 1465 875 2280 907
rect 1465 865 1552 875
rect 1447 862 1552 865
rect 1625 862 1712 875
rect 1831 874 2280 875
rect 1823 869 2280 874
rect 2380 928 5386 931
rect 5390 930 5442 941
rect 5401 928 5431 930
rect 5452 928 5482 943
rect 2380 923 5482 928
rect 2380 921 2952 923
rect 2961 921 5482 923
rect 2380 907 5482 921
rect 2380 887 5354 907
rect 5355 902 5467 907
rect 2380 874 2831 887
rect 2861 881 5354 887
rect 2861 874 5415 881
rect 2380 870 2819 874
rect 1447 861 1712 862
rect 1309 765 1343 861
rect 1352 765 1379 861
rect 1393 839 1712 861
rect 1393 831 1517 839
rect 1393 827 1420 831
rect 1440 827 1517 831
rect 1460 825 1517 827
rect 1533 831 1539 839
rect 1533 827 1534 831
rect 1545 827 1551 839
rect 1552 828 1667 839
rect 1401 821 1529 825
rect 1460 815 1517 821
rect 1429 795 1501 797
rect 1533 795 1586 827
rect 1233 764 1291 765
rect 1145 750 1203 764
rect 1219 750 1291 764
rect 1309 763 1379 765
rect 1422 773 1586 795
rect 1422 763 1590 773
rect 1599 763 1615 773
rect 1625 763 1667 828
rect 1678 816 1712 839
rect 1722 829 1805 863
rect 1823 862 2301 869
rect 1823 852 2280 862
rect 2284 861 2301 862
rect 2318 852 2335 861
rect 2341 852 2376 861
rect 1823 839 2376 852
rect 2397 845 2581 870
rect 2397 839 2629 845
rect 1823 835 2397 839
rect 1823 829 2376 835
rect 1823 816 1824 829
rect 1835 827 2376 829
rect 2379 827 2410 835
rect 1835 816 2363 827
rect 1678 784 2363 816
rect 1678 782 2125 784
rect 1309 752 1393 763
rect 1309 750 1382 752
rect 940 749 1382 750
rect 940 710 974 749
rect 981 745 1008 749
rect 1153 716 1203 749
rect 1233 715 1291 749
rect 1309 735 1382 749
rect 1422 750 1667 763
rect 1672 757 1747 782
rect 1823 775 1868 782
rect 1672 753 1772 757
rect 1679 750 1772 753
rect 1422 749 1772 750
rect 1422 740 1621 749
rect 1627 740 1643 749
rect 1644 748 1667 749
rect 1738 748 1772 749
rect 1309 729 1344 735
rect 1422 729 1643 740
rect 940 681 975 710
rect 1104 699 1158 710
rect 1178 699 1230 710
rect 1115 687 1147 699
rect 1189 687 1219 699
rect 1275 695 1290 715
rect 1576 696 1590 729
rect 1115 681 1158 687
rect 940 676 1158 681
rect 1178 676 1230 687
rect 1280 676 1290 695
rect 1444 681 1459 696
rect 1575 681 1590 696
rect 571 623 600 656
rect 844 651 921 657
rect 844 646 855 651
rect 202 589 566 604
rect 610 600 615 646
rect 638 600 643 646
rect 906 642 921 651
rect 910 640 921 642
rect 1444 651 1502 681
rect 1532 651 1590 681
rect 655 623 880 640
rect 1444 636 1459 651
rect 1575 636 1590 651
rect 1599 646 1615 729
rect 1627 646 1643 729
rect 1823 706 1894 775
rect 1923 706 1957 782
rect 1967 757 1983 782
rect 2003 773 2125 782
rect 2149 777 2193 784
rect 1995 761 2057 773
rect 2127 772 2193 777
rect 2127 761 2195 772
rect 1995 757 2011 761
rect 2025 740 2079 761
rect 2011 706 2079 740
rect 2125 706 2195 761
rect 2246 771 2363 784
rect 2367 825 2368 827
rect 2379 825 2413 827
rect 2367 771 2413 825
rect 2507 821 2629 839
rect 2513 817 2581 821
rect 2513 801 2601 817
rect 2414 771 2425 797
rect 2467 773 2501 797
rect 2507 793 2601 801
rect 2444 771 2501 773
rect 2246 759 2295 771
rect 2268 740 2317 759
rect 2367 750 2502 771
rect 2513 750 2581 793
rect 2367 749 2581 750
rect 2685 750 2686 870
rect 2735 869 2737 870
rect 2763 869 2765 870
rect 2785 863 2819 870
rect 2873 863 2907 874
rect 2908 869 2913 874
rect 2918 863 2952 874
rect 2961 863 2995 874
rect 2785 829 2995 863
rect 2785 822 2819 829
rect 2785 761 2825 822
rect 2800 760 2825 761
rect 2828 764 2853 822
rect 2884 798 2907 829
rect 2873 788 2907 798
rect 2908 788 2913 822
rect 2873 782 2913 788
rect 2918 782 2952 829
rect 2873 764 2952 782
rect 2961 786 2995 829
rect 2996 815 5354 874
rect 5355 873 5389 874
rect 5355 862 5359 873
rect 5355 815 5389 862
rect 5409 815 5415 874
rect 5433 878 5467 902
rect 5433 815 5477 878
rect 2996 798 5477 815
rect 2828 760 2868 764
rect 2873 760 2956 764
rect 2961 760 2998 786
rect 3020 784 3100 798
rect 3010 766 3100 784
rect 3120 766 3154 798
rect 3200 793 3217 797
rect 3234 786 3268 798
rect 3287 786 3321 798
rect 3010 760 3095 766
rect 2800 754 3095 760
rect 3126 754 3154 766
rect 3166 764 3178 784
rect 3234 782 3236 786
rect 3249 782 3321 786
rect 3160 754 3188 764
rect 2800 750 3056 754
rect 3063 750 3095 754
rect 2685 749 3095 750
rect 3117 750 3188 754
rect 2249 706 2317 740
rect 2368 747 2425 749
rect 1823 695 1872 706
rect 1967 695 1983 701
rect 1995 695 2011 701
rect 2025 695 2057 706
rect 1823 694 2057 695
rect 2125 695 2193 706
rect 2268 695 2295 706
rect 2125 694 2295 695
rect 1732 646 1743 674
rect 1866 653 1872 694
rect 1967 681 1983 694
rect 1995 653 2011 694
rect 655 607 656 623
rect 880 607 906 623
rect 655 606 906 607
rect 1239 600 1361 606
rect 1689 600 1715 646
rect 1717 600 1743 646
rect 2049 605 2071 678
rect 2125 640 2159 694
rect 2161 690 2193 694
rect 2171 640 2225 666
rect 2087 607 2171 640
rect 2175 607 2193 640
rect 2199 607 2225 640
rect 2087 606 2225 607
rect 202 579 552 589
rect 202 570 293 579
rect 337 572 444 579
rect 478 572 531 579
rect 1267 572 1333 578
rect 1732 573 1743 600
rect 2053 589 2071 605
rect 2326 600 2331 646
rect 2354 600 2359 646
rect 2368 640 2402 747
rect 2444 723 2455 749
rect 2456 723 2490 749
rect 2800 745 2819 749
rect 2828 721 2868 749
rect 2873 748 2956 749
rect 2873 745 2907 748
rect 2916 721 2956 748
rect 2961 745 2995 749
rect 3007 745 3078 749
rect 2831 711 2868 721
rect 2831 696 2861 711
rect 2456 640 2490 674
rect 2502 640 2622 666
rect 2368 606 2622 640
rect 2822 651 2861 696
rect 2822 636 2837 651
rect 479 570 531 572
rect 260 551 266 570
rect 66 504 206 509
rect 240 504 266 528
rect 67 476 206 481
rect 240 476 294 500
rect 260 300 294 325
rect 328 300 362 325
rect 260 281 267 300
rect 294 297 295 300
rect 260 128 266 281
rect 192 104 266 128
rect 288 253 295 297
rect 328 272 334 297
rect 1967 281 1983 481
rect 1995 253 2011 509
rect 2368 423 2402 606
rect 2918 605 2956 721
rect 3007 707 3056 745
rect 3117 717 3136 750
rect 3145 748 3188 750
rect 3214 761 3321 782
rect 3214 760 3268 761
rect 3287 760 3321 761
rect 3214 750 3321 760
rect 3349 750 3355 798
rect 3363 781 5477 798
rect 3365 750 5354 781
rect 3214 749 5354 750
rect 3214 748 3268 749
rect 3287 748 3321 749
rect 3145 745 3192 748
rect 3007 701 3044 707
rect 2976 646 2982 701
rect 3004 696 3044 701
rect 3045 696 3056 707
rect 3004 651 3056 696
rect 3060 681 3103 707
rect 3126 701 3136 717
rect 3148 728 3192 745
rect 3148 716 3188 728
rect 3148 681 3164 716
rect 3060 673 3082 681
rect 3089 667 3122 674
rect 3004 646 3010 651
rect 3026 639 3056 651
rect 3148 651 3206 681
rect 3234 658 3321 748
rect 3349 745 3355 749
rect 3365 745 5354 749
rect 5355 745 5389 781
rect 5409 745 5415 781
rect 3433 726 3445 745
rect 3471 726 3491 745
rect 3433 720 3491 726
rect 3499 692 3519 745
rect 3539 712 3540 745
rect 3569 712 3585 745
rect 3603 712 3637 745
rect 3539 695 3637 712
rect 3639 711 3690 745
rect 3693 711 3699 745
rect 3718 740 3727 745
rect 3734 740 5281 745
rect 3718 711 5281 740
rect 3639 695 5281 711
rect 5354 695 5422 745
rect 3539 694 5422 695
rect 5437 694 5443 781
rect 5452 694 5477 781
rect 5486 868 5520 943
rect 5562 936 5634 943
rect 5639 936 5646 943
rect 5562 902 5646 936
rect 5688 930 6498 943
rect 5688 929 6494 930
rect 6506 929 6515 933
rect 5688 904 6498 929
rect 5562 893 5597 902
rect 5600 898 5634 902
rect 5688 898 5722 904
rect 5566 879 5597 893
rect 5628 879 5639 880
rect 5486 728 5511 868
rect 5821 861 5836 904
rect 5777 843 5836 861
rect 5777 827 5845 843
rect 5855 827 5889 904
rect 5994 893 6009 904
rect 5957 880 6009 893
rect 5957 874 6003 880
rect 5957 851 5999 874
rect 6059 868 6498 904
rect 6506 868 6527 929
rect 6059 851 6527 868
rect 5957 849 6003 851
rect 6095 849 6097 851
rect 6117 849 6163 851
rect 5969 845 6003 849
rect 5802 824 5889 827
rect 5593 762 5627 796
rect 5681 762 5715 796
rect 5802 762 5845 824
rect 5581 728 5727 762
rect 5740 728 5749 762
rect 5799 749 5845 762
rect 5821 745 5845 749
rect 5855 763 5889 824
rect 5899 763 5923 843
rect 5935 827 5939 839
rect 6123 821 6125 849
rect 5967 811 6033 817
rect 5983 797 6047 811
rect 5983 777 6059 797
rect 5983 767 6017 777
rect 6033 771 6059 777
rect 5855 749 5945 763
rect 5821 728 5836 745
rect 5855 711 5889 749
rect 5899 745 5923 749
rect 6033 743 6087 769
rect 6137 763 6163 849
rect 6171 763 6205 851
rect 6117 749 6205 763
rect 6137 745 6163 749
rect 6171 711 6205 749
rect 6217 761 6285 851
rect 6305 808 6378 851
rect 6305 761 6339 808
rect 6359 796 6378 808
rect 6384 834 6527 851
rect 6384 808 6466 834
rect 6384 796 6427 808
rect 6430 800 6466 808
rect 6447 796 6466 800
rect 6359 792 6372 796
rect 6384 792 6460 796
rect 6217 745 6258 761
rect 6332 745 6339 761
rect 6342 749 6345 792
rect 6384 774 6454 792
rect 6370 758 6373 764
rect 5855 694 5870 711
rect 5992 698 6044 709
rect 6003 694 6033 698
rect 3569 692 3585 694
rect 3551 690 3585 692
rect 3603 658 3637 694
rect 3639 690 3715 694
rect 3734 692 5263 694
rect 3656 688 3715 690
rect 3752 688 3953 692
rect 3656 677 3726 688
rect 3752 677 3964 688
rect 4103 666 5263 692
rect 5409 681 5415 694
rect 5855 681 6082 694
rect 6190 681 6205 711
rect 5855 675 6205 681
rect 3234 651 3348 658
rect 3517 656 3637 658
rect 3148 646 3163 651
rect 3089 639 3163 646
rect 2980 626 3010 639
rect 3038 636 3056 639
rect 3148 636 3206 639
rect 3038 635 3044 636
rect 2980 605 3044 626
rect 3160 605 3206 636
rect 3234 605 3282 651
rect 3287 624 3316 651
rect 3337 647 3348 651
rect 2918 580 3056 605
rect 3148 590 3282 605
rect 3405 600 3431 646
rect 3433 600 3459 646
rect 3622 643 3637 656
rect 3777 640 3833 666
rect 3863 640 3905 666
rect 3803 629 3874 640
rect 3894 629 3915 640
rect 3803 617 3827 629
rect 3833 617 3863 629
rect 3905 617 3915 629
rect 3803 607 3874 617
rect 3894 607 3915 617
rect 4042 607 4047 646
rect 4061 640 5263 666
rect 6224 656 6258 745
rect 6366 724 6373 758
rect 6381 749 6454 774
rect 6475 770 6498 834
rect 6475 768 6494 770
rect 6481 761 6494 768
rect 6506 749 6527 834
rect 6540 868 6574 980
rect 6588 970 6627 980
rect 6593 868 6627 970
rect 6656 936 6661 970
rect 6665 930 6668 976
rect 6693 911 6696 997
rect 6711 927 6727 997
rect 6739 995 6814 997
rect 6735 961 6755 995
rect 6780 961 6814 995
rect 6739 955 6814 961
rect 6780 930 6814 955
rect 6780 923 6783 930
rect 6799 927 6814 930
rect 6799 923 6829 927
rect 6724 908 6753 923
rect 6739 868 6753 908
rect 6780 868 6829 923
rect 6540 834 6829 868
rect 6381 724 6431 749
rect 6439 708 6469 749
rect 6506 745 6515 749
rect 6540 718 6574 834
rect 6540 681 6551 692
rect 6559 681 6574 718
rect 6540 656 6574 681
rect 6224 651 6304 656
rect 3803 606 3915 607
rect 3955 600 4047 607
rect 4070 600 4075 640
rect 4087 639 5263 640
rect 4087 607 4111 639
rect 4160 607 4338 639
rect 4442 636 4457 639
rect 4087 606 4338 607
rect 3148 580 3268 590
rect 4267 584 4294 591
rect 4472 586 5263 639
rect 5758 600 5763 646
rect 5786 600 5791 646
rect 6224 641 6239 651
rect 6293 645 6304 651
rect 6428 651 6574 656
rect 6428 645 6439 651
rect 6224 640 6235 641
rect 6559 622 6574 651
rect 6593 622 6627 834
rect 6707 827 6741 834
rect 6770 827 6783 834
rect 6795 827 6829 834
rect 6693 761 6741 827
rect 6781 761 6829 827
rect 6833 923 6867 997
rect 6833 781 6863 923
rect 6909 815 6943 1010
rect 6947 951 6977 1010
rect 7037 957 8214 1010
rect 6979 917 7037 923
rect 6975 883 6977 917
rect 6979 883 6991 917
rect 6979 877 7037 883
rect 6909 781 7087 815
rect 7168 781 7183 957
rect 7202 781 7236 957
rect 7406 930 8214 957
rect 7406 904 8210 930
rect 7348 864 7406 870
rect 7348 830 7360 864
rect 7348 824 7406 830
rect 6707 755 6741 761
rect 6795 755 6829 761
rect 6724 749 6739 755
rect 6724 743 6753 749
rect 6799 747 6829 755
rect 6739 665 6775 674
rect 6909 665 6943 781
rect 7202 747 7217 781
rect 7537 728 7552 904
rect 7571 728 7605 904
rect 7775 851 8210 904
rect 7717 811 7775 817
rect 7717 777 7729 811
rect 7717 771 7775 777
rect 7571 694 7586 728
rect 7906 675 7921 851
rect 7940 675 7974 851
rect 8146 800 8176 851
rect 8180 834 8210 851
rect 8256 868 8290 1116
rect 8294 1097 8324 1184
rect 8371 1097 8382 1131
rect 8496 1097 8530 1266
rect 8549 1275 8584 1309
rect 8549 1097 8583 1275
rect 8695 1207 8753 1213
rect 8695 1173 8707 1207
rect 8695 1167 8753 1173
rect 8865 1166 8899 1220
rect 8294 1063 8583 1097
rect 8629 1063 8659 1097
rect 8294 1004 8343 1063
rect 8304 976 8343 1004
rect 8496 1001 8530 1063
rect 8455 995 8530 1001
rect 8304 970 8384 976
rect 8309 936 8343 970
rect 8372 936 8377 970
rect 8451 961 8467 995
rect 8496 961 8530 995
rect 8455 955 8530 961
rect 8309 930 8384 936
rect 8496 930 8530 955
rect 8309 868 8343 930
rect 8496 923 8499 930
rect 8515 927 8530 930
rect 8515 923 8545 927
rect 8496 868 8545 923
rect 8256 834 8545 868
rect 8086 758 8144 764
rect 8086 724 8098 758
rect 8086 718 8144 724
rect 8256 718 8290 834
rect 6711 637 6775 646
rect 7940 641 7955 675
rect 8275 622 8290 718
rect 8309 622 8343 834
rect 8515 747 8545 834
rect 8549 877 8583 1063
rect 8549 781 8579 877
rect 8625 815 8659 1063
rect 8663 951 8693 1131
rect 8695 917 8753 923
rect 8691 883 8693 917
rect 8695 883 8707 917
rect 8695 877 8753 883
rect 8625 781 8803 815
rect 8884 781 8899 1166
rect 8918 1132 8953 1166
rect 9233 1132 9268 1166
rect 8918 781 8952 1132
rect 9234 1113 9268 1132
rect 9656 1116 9691 1150
rect 9064 1064 9122 1070
rect 9064 1030 9076 1064
rect 9064 1024 9122 1030
rect 9064 864 9122 870
rect 9064 830 9076 864
rect 9064 824 9122 830
rect 8455 705 8513 711
rect 8455 671 8467 705
rect 8455 665 8513 671
rect 8625 665 8659 781
rect 8918 747 8933 781
rect 9253 728 9268 1113
rect 9287 1079 9322 1113
rect 9287 728 9321 1079
rect 9433 1011 9491 1017
rect 9433 977 9445 1011
rect 9433 971 9491 977
rect 9433 811 9491 817
rect 9433 777 9445 811
rect 9433 771 9491 777
rect 9287 694 9302 728
rect 9622 675 9637 1113
rect 9656 675 9690 1116
rect 9802 1048 9860 1054
rect 9802 1014 9814 1048
rect 9802 1008 9860 1014
rect 9802 758 9860 764
rect 9802 724 9814 758
rect 9802 718 9860 724
rect 9656 641 9671 675
rect 6593 588 6608 622
rect 8309 588 8324 622
rect 2918 571 3009 580
rect 3195 571 3247 580
rect 3983 572 4049 579
rect 2976 552 2982 571
rect 4267 569 4296 584
rect 4239 556 4266 563
rect 4239 541 4268 556
rect 4841 533 5263 586
rect 2956 505 2982 529
rect 2956 477 3010 501
rect 5084 424 5118 533
rect 5187 412 5212 509
rect 5187 402 5206 412
rect 2742 323 2751 369
rect 2770 348 2779 397
rect 5215 384 5240 481
rect 5215 374 5234 384
rect 5187 365 5196 374
rect 2772 340 2779 348
rect 2922 326 2936 333
rect 2744 318 2751 323
rect 2894 298 2936 305
rect 2976 301 3010 326
rect 3044 301 3078 326
rect 4239 317 4266 325
rect 4267 317 4294 353
rect 5187 313 5198 365
rect 5187 308 5196 313
rect 288 128 294 253
rect 2551 169 2685 192
rect 2754 169 2757 221
rect 2525 141 2685 164
rect 2782 141 2785 249
rect 2976 129 2982 301
rect 288 117 334 128
rect 192 81 200 104
rect 220 89 362 100
rect 220 81 294 89
rect 200 76 294 81
rect 410 69 420 100
rect 438 69 448 128
rect 1755 69 1778 109
rect 1895 105 1967 109
rect 2908 105 2982 129
rect 3004 129 3010 298
rect 3044 273 3050 298
rect 5215 285 5226 374
rect 5215 281 5224 285
rect 5187 253 5224 277
rect 4218 147 4306 154
rect 3004 118 3050 129
rect 2936 90 3078 101
rect 1783 69 1806 81
rect 1867 77 1983 81
rect 2936 77 3010 90
rect 3126 70 3136 101
rect 3154 70 3164 129
rect 4442 128 4588 154
rect 4454 124 4488 128
rect 4542 124 4576 128
rect 4353 90 4610 100
rect 4353 66 4578 90
rect 5187 71 5206 109
rect 5215 71 5234 81
rect 6978 67 7013 101
rect 40 50 240 63
rect 2756 51 2956 64
rect 40 29 265 50
rect 370 35 434 50
rect 370 29 482 35
rect 557 29 676 35
rect 706 29 823 35
rect 2756 30 2981 51
rect 3086 36 3150 51
rect 4030 47 4065 65
rect 3086 30 3198 36
rect 3253 30 3392 36
rect 3422 30 3539 36
rect 3471 18 3474 24
rect 3499 18 3502 24
rect 3893 19 3928 47
rect 3989 19 4147 47
rect 3099 17 3521 18
rect 383 16 805 17
rect 50 -5 805 16
rect 2766 -3 3521 17
rect 240 -7 805 -5
rect 229 -12 805 -7
rect 229 -18 281 -12
rect 365 -18 805 -12
rect 366 -19 805 -18
rect 383 -26 805 -19
rect 50 -170 84 -26
rect 158 -80 170 -76
rect 158 -86 182 -80
rect 158 -132 170 -86
rect 136 -140 170 -132
rect 177 -140 182 -86
rect 192 -120 204 -86
rect 208 -120 254 -86
rect 366 -90 805 -26
rect 2758 -4 3521 -3
rect 2758 -25 2779 -4
rect 2956 -6 3521 -4
rect 3893 13 4147 19
rect 4228 29 4251 38
rect 4407 32 4490 62
rect 4568 32 4578 62
rect 2945 -11 3521 -6
rect 2945 -17 2997 -11
rect 3081 -17 3521 -11
rect 3082 -18 3521 -17
rect 3099 -25 3521 -18
rect 1121 -90 1543 -89
rect 136 -158 198 -140
rect 204 -148 270 -120
rect 366 -124 823 -90
rect 918 -124 1064 -90
rect 1103 -124 1543 -90
rect 1979 -99 1983 -28
rect 1972 -119 1983 -99
rect 252 -158 286 -154
rect 170 -163 210 -158
rect 240 -163 292 -158
rect 170 -170 198 -163
rect 83 -322 84 -170
rect 164 -196 198 -170
rect 252 -176 292 -163
rect 252 -182 286 -176
rect 248 -255 298 -217
rect 204 -296 246 -291
rect 266 -305 298 -255
rect 316 -289 320 -255
rect 50 -328 61 -322
rect 73 -328 84 -322
rect 204 -324 246 -319
rect 283 -320 298 -305
rect 366 -305 822 -124
rect 930 -154 964 -124
rect 1104 -142 1543 -124
rect 1550 -142 1590 -124
rect 2007 -127 2011 -56
rect 2382 -114 2470 -111
rect 2363 -126 2470 -114
rect 918 -158 1006 -154
rect 918 -170 1030 -158
rect 1104 -170 1912 -142
rect 2000 -146 2011 -127
rect 930 -174 964 -170
rect 1018 -174 1030 -170
rect 930 -208 996 -192
rect 1118 -213 1912 -170
rect 2417 -182 2423 -165
rect 1104 -226 1912 -213
rect 1093 -235 1912 -226
rect 2012 -210 2434 -182
rect 2730 -197 2751 -31
rect 2758 -112 2800 -25
rect 2874 -79 2886 -75
rect 2874 -85 2898 -79
rect 2912 -85 2920 -79
rect 2874 -95 2892 -85
rect 2874 -112 2886 -95
rect 2893 -112 2898 -85
rect 2908 -112 2920 -85
rect 2924 -91 2958 -85
rect 2924 -112 2970 -91
rect 3082 -112 3521 -25
rect 3524 -11 3733 -6
rect 3524 -35 3559 -11
rect 3692 -17 3733 -11
rect 3822 -17 3874 -6
rect 3692 -25 3722 -17
rect 3826 -25 3874 -17
rect 3580 -35 3874 -25
rect 3893 -31 3927 13
rect 4209 -8 4220 3
rect 4228 -8 4243 29
rect 3892 -35 3927 -31
rect 4001 -35 4014 -31
rect 3524 -40 3874 -35
rect 3524 -89 3558 -40
rect 3648 -85 3750 -74
rect 3644 -89 3754 -85
rect 3840 -88 3874 -40
rect 3880 -88 3928 -35
rect 4001 -55 4026 -35
rect 4001 -81 4014 -55
rect 4020 -81 4026 -55
rect 4001 -88 4026 -81
rect 4035 -88 4048 -55
rect 4051 -81 4098 -47
rect 4051 -88 4085 -81
rect 4175 -88 4206 -51
rect 4209 -88 4243 -8
rect 4262 -51 4296 29
rect 4380 28 4490 32
rect 4592 28 4627 38
rect 4380 22 4426 28
rect 4460 22 4494 28
rect 6609 14 6644 48
rect 4408 -2 4426 4
rect 4430 -2 4470 14
rect 4404 -6 4470 -2
rect 4578 -6 4589 5
rect 4420 -32 4454 -6
rect 4472 -32 4502 -6
rect 3837 -89 4259 -88
rect 2758 -146 3068 -112
rect 3070 -146 3521 -112
rect 2758 -165 2820 -146
rect 2752 -169 2820 -165
rect 2766 -208 2800 -169
rect 2810 -208 2820 -169
rect 2852 -157 2914 -146
rect 2920 -147 2986 -146
rect 2968 -157 3002 -153
rect 2852 -173 2854 -157
rect 2886 -162 2926 -157
rect 2956 -162 3014 -157
rect 2886 -169 2920 -162
rect 2880 -171 2920 -169
rect 2968 -171 3014 -162
rect 2012 -235 2451 -210
rect 2551 -231 2555 -212
rect 366 -316 377 -305
rect 383 -328 822 -305
rect 956 -328 964 -236
rect 1093 -248 2451 -235
rect 2523 -241 2527 -240
rect 2457 -248 2485 -244
rect 2517 -248 2527 -241
rect 978 -279 1021 -264
rect 978 -328 1006 -279
rect 1090 -294 1195 -248
rect 1090 -328 1191 -294
rect 1275 -295 1298 -248
rect 1303 -261 1326 -248
rect 1303 -267 1361 -261
rect 14 -403 453 -328
rect 521 -358 579 -328
rect 609 -358 618 -328
rect 521 -367 530 -358
rect 521 -382 545 -367
rect 627 -382 667 -376
rect 735 -377 1191 -328
rect 1259 -377 1267 -308
rect 1276 -377 1305 -304
rect 1391 -312 1399 -308
rect 1391 -320 1405 -312
rect 1372 -324 1405 -320
rect 1419 -324 1427 -280
rect 1473 -324 1507 -248
rect 1526 -324 1560 -248
rect 1735 -271 1776 -248
rect 1844 -271 1876 -248
rect 2048 -252 2083 -248
rect 1679 -285 1986 -271
rect 1679 -290 1995 -285
rect 1668 -303 1995 -290
rect 1998 -303 2011 -291
rect 2014 -303 2029 -271
rect 2048 -303 2082 -252
rect 2201 -301 2280 -286
rect 1668 -305 2281 -303
rect 1668 -314 1734 -305
rect 1679 -316 1713 -314
rect 1679 -320 1744 -316
rect 1756 -320 1776 -305
rect 1798 -320 1832 -316
rect 1842 -320 2281 -305
rect 14 -410 442 -403
rect 446 -410 453 -403
rect 14 -483 453 -410
rect 519 -413 530 -382
rect 735 -411 1195 -377
rect 1211 -388 1305 -377
rect 1222 -400 1252 -388
rect 1259 -400 1305 -388
rect 1211 -411 1305 -400
rect 561 -430 572 -413
rect 596 -429 623 -423
rect 577 -430 668 -429
rect 735 -430 1191 -411
rect 454 -483 487 -444
rect 561 -448 1191 -430
rect 546 -460 1191 -448
rect 1257 -421 1305 -411
rect 1310 -358 1405 -324
rect 1406 -358 1564 -324
rect 1310 -421 1344 -358
rect 1359 -421 1378 -358
rect 1391 -406 1399 -358
rect 1390 -421 1405 -406
rect 1257 -460 1344 -421
rect 1347 -455 1405 -421
rect 542 -464 1191 -460
rect 542 -469 651 -464
rect 542 -483 606 -469
rect 618 -479 651 -469
rect 14 -501 606 -483
rect 624 -497 651 -479
rect 735 -485 1191 -464
rect 705 -494 1191 -485
rect 1230 -476 1344 -460
rect 1359 -476 1405 -455
rect 1230 -492 1305 -476
rect 1230 -494 1298 -492
rect 1310 -494 1344 -476
rect 1358 -488 1405 -476
rect 1359 -492 1378 -488
rect 1390 -492 1393 -488
rect 14 -517 553 -501
rect 14 -531 453 -517
rect 454 -531 488 -517
rect 519 -531 553 -517
rect 572 -531 606 -501
rect 630 -501 649 -497
rect 705 -498 1225 -494
rect 630 -531 640 -501
rect 696 -531 1225 -498
rect 14 -548 1225 -531
rect 169 -632 170 -548
rect 178 -628 182 -548
rect 203 -571 237 -548
rect 366 -551 412 -548
rect 419 -551 1225 -548
rect 366 -554 1225 -551
rect 354 -565 1225 -554
rect 354 -569 429 -565
rect 203 -579 236 -571
rect 203 -691 237 -579
rect 354 -612 442 -569
rect 485 -612 488 -565
rect 354 -616 488 -612
rect 354 -628 500 -616
rect 519 -628 553 -565
rect 366 -632 400 -628
rect 412 -635 442 -628
rect 454 -632 473 -628
rect 485 -632 488 -628
rect 332 -666 351 -662
rect 338 -678 357 -666
rect 317 -681 357 -678
rect 200 -696 266 -691
rect 305 -696 357 -681
rect 203 -719 237 -696
rect 200 -724 267 -719
rect 203 -737 237 -724
rect 115 -771 237 -737
rect 305 -726 363 -696
rect 305 -731 357 -726
rect 366 -731 385 -638
rect 412 -654 435 -635
rect 405 -666 439 -662
rect 397 -669 451 -666
rect 426 -678 445 -669
rect 405 -681 445 -678
rect 405 -696 451 -681
rect 454 -690 473 -638
rect 393 -704 451 -696
rect 393 -726 453 -704
rect 305 -738 351 -731
rect 405 -738 453 -726
rect 519 -737 530 -628
rect 305 -741 462 -738
rect 203 -818 237 -771
rect 317 -772 462 -741
rect 173 -852 237 -818
rect 203 -995 241 -852
rect 261 -961 267 -778
rect 289 -816 295 -778
rect 317 -816 351 -772
rect 289 -834 351 -816
rect 405 -834 439 -772
rect 519 -814 530 -803
rect 289 -836 317 -834
rect 289 -852 295 -836
rect 314 -852 341 -846
rect 411 -850 439 -834
rect 451 -836 463 -816
rect 519 -818 521 -814
rect 538 -818 553 -632
rect 499 -836 553 -818
rect 445 -852 473 -836
rect 499 -852 567 -836
rect 572 -840 606 -565
rect 630 -632 640 -565
rect 714 -572 1225 -565
rect 714 -575 1191 -572
rect 1210 -575 1225 -572
rect 1257 -574 1344 -494
rect 1419 -507 1427 -358
rect 1473 -388 1507 -358
rect 1428 -426 1452 -392
rect 1466 -420 1507 -388
rect 1456 -426 1507 -420
rect 1428 -456 1507 -426
rect 1526 -388 1560 -358
rect 1526 -456 1568 -388
rect 1428 -460 1518 -456
rect 1428 -494 1452 -460
rect 1456 -466 1507 -460
rect 1473 -481 1507 -466
rect 1526 -481 1552 -456
rect 1473 -503 1560 -481
rect 1418 -515 1427 -507
rect 1455 -515 1560 -503
rect 1456 -519 1594 -515
rect 1349 -569 1378 -535
rect 652 -585 664 -575
rect 714 -582 1210 -575
rect 652 -587 670 -585
rect 732 -587 1210 -582
rect 648 -616 670 -587
rect 718 -598 1210 -587
rect 686 -609 1210 -598
rect 686 -613 698 -609
rect 680 -614 698 -613
rect 652 -628 670 -616
rect 676 -625 706 -614
rect 718 -616 1210 -609
rect 732 -625 1210 -616
rect 680 -628 720 -625
rect 652 -690 664 -628
rect 676 -654 720 -628
rect 740 -637 1210 -625
rect 1257 -585 1365 -574
rect 1424 -585 1560 -519
rect 1257 -637 1344 -585
rect 1363 -616 1397 -603
rect 1412 -616 1560 -585
rect 1347 -628 1560 -616
rect 1578 -628 1594 -519
rect 1606 -569 1620 -333
rect 1634 -348 1660 -324
rect 1645 -357 1660 -348
rect 1679 -330 1756 -320
rect 1786 -330 2281 -320
rect 1679 -332 1749 -330
rect 1679 -333 1744 -332
rect 1645 -361 1674 -357
rect 1628 -386 1674 -361
rect 1679 -373 1747 -333
rect 1755 -373 1768 -361
rect 1679 -386 1768 -373
rect 1628 -449 1768 -386
rect 1626 -529 1768 -449
rect 1783 -455 1796 -333
rect 1782 -466 1796 -455
rect 1798 -357 1832 -330
rect 1842 -357 2281 -330
rect 1798 -423 2281 -357
rect 1798 -466 1832 -423
rect 1783 -519 1832 -466
rect 1626 -545 1674 -529
rect 1626 -554 1660 -545
rect 1679 -554 1747 -529
rect 1755 -541 1768 -529
rect 1759 -545 1762 -541
rect 1626 -588 1752 -554
rect 1787 -569 1832 -519
rect 1347 -632 1578 -628
rect 1347 -637 1382 -632
rect 1386 -636 1578 -632
rect 1386 -637 1590 -636
rect 740 -654 1590 -637
rect 680 -666 698 -654
rect 680 -681 692 -666
rect 674 -696 692 -681
rect 674 -726 732 -696
rect 674 -741 689 -726
rect 740 -731 752 -654
rect 768 -696 808 -654
rect 813 -655 846 -654
rect 813 -671 842 -655
rect 854 -671 879 -654
rect 813 -696 820 -671
rect 762 -726 820 -696
rect 768 -731 780 -726
rect 805 -741 820 -726
rect 888 -726 922 -654
rect 888 -737 899 -726
rect 718 -840 776 -834
rect 572 -852 601 -840
rect 289 -872 341 -852
rect 289 -961 295 -872
rect 311 -958 341 -872
rect 349 -893 407 -887
rect 345 -927 388 -893
rect 433 -927 442 -852
rect 445 -872 477 -852
rect 445 -884 473 -872
rect 349 -933 407 -927
rect 519 -933 601 -852
rect 718 -874 730 -840
rect 718 -880 776 -874
rect 311 -961 335 -958
rect 261 -974 295 -961
rect 323 -965 329 -961
rect 261 -995 329 -974
rect 445 -995 491 -961
rect 519 -995 567 -933
rect 572 -976 601 -933
rect 907 -957 922 -726
rect 941 -889 975 -654
rect 1055 -666 1086 -654
rect 1131 -662 1590 -654
rect 1131 -671 1189 -662
rect 1211 -671 1590 -662
rect 1131 -728 1177 -671
rect 1131 -740 1163 -728
rect 1059 -778 1173 -753
rect 1087 -806 1145 -781
rect 1087 -821 1099 -806
rect 1087 -827 1145 -821
rect 1148 -833 1149 -821
rect 1257 -827 1291 -671
rect 1190 -837 1191 -833
rect 1257 -834 1268 -827
rect 1276 -834 1291 -827
rect 1257 -864 1291 -834
rect 1257 -875 1268 -864
rect 941 -923 976 -889
rect 1107 -900 1159 -889
rect 1179 -900 1231 -889
rect 1118 -912 1148 -900
rect 1190 -912 1220 -900
rect 1276 -904 1291 -864
rect 1310 -836 1344 -671
rect 1347 -682 1378 -671
rect 1390 -682 1413 -671
rect 1424 -675 1458 -671
rect 1424 -682 1447 -675
rect 1412 -684 1447 -682
rect 1478 -683 1496 -671
rect 1502 -672 1590 -671
rect 1500 -683 1590 -672
rect 1412 -687 1452 -684
rect 1478 -687 1490 -683
rect 1500 -687 1578 -683
rect 1424 -691 1447 -687
rect 1502 -690 1560 -687
rect 1626 -690 1660 -588
rect 1668 -622 1752 -588
rect 1793 -622 1832 -569
rect 1679 -636 1747 -622
rect 1798 -634 1832 -622
rect 1839 -428 2281 -423
rect 2381 -327 2550 -248
rect 2559 -261 2567 -251
rect 2766 -261 2820 -208
rect 2559 -267 2621 -261
rect 2559 -301 2575 -267
rect 2559 -307 2621 -301
rect 2559 -311 2567 -307
rect 2733 -327 2820 -261
rect 2880 -291 2914 -171
rect 2968 -175 3008 -171
rect 2968 -176 3002 -175
rect 2968 -180 3006 -176
rect 2968 -198 3012 -180
rect 2956 -214 3012 -198
rect 2928 -216 3012 -214
rect 3082 -185 3521 -146
rect 3524 -185 3558 -102
rect 3634 -123 3780 -89
rect 3822 -100 4259 -89
rect 3833 -123 4259 -100
rect 3646 -126 3766 -123
rect 3634 -142 3780 -126
rect 3634 -153 3714 -142
rect 3722 -153 3780 -142
rect 3634 -169 3780 -153
rect 3820 -141 4259 -123
rect 4260 -123 4296 -51
rect 4414 -36 4492 -32
rect 4414 -47 4472 -36
rect 4514 -46 4532 -36
rect 4414 -52 4470 -47
rect 4508 -48 4532 -46
rect 4414 -67 4460 -52
rect 4392 -86 4410 -70
rect 4422 -74 4460 -67
rect 4260 -141 4306 -123
rect 4388 -141 4410 -86
rect 4426 -126 4460 -74
rect 4464 -74 4498 -70
rect 4464 -141 4504 -74
rect 4508 -110 4536 -48
rect 4508 -122 4532 -110
rect 4514 -141 4532 -122
rect 4544 -126 4548 -28
rect 4578 -32 4590 -6
rect 4578 -122 4612 -32
rect 6240 -39 6275 -5
rect 5871 -92 5906 -58
rect 5098 -113 5186 -110
rect 4578 -141 4590 -122
rect 5079 -125 5186 -113
rect 3820 -169 4628 -141
rect 5502 -145 5537 -111
rect 3646 -173 3706 -169
rect 3734 -173 3768 -169
rect 3662 -176 3706 -173
rect 3638 -180 3706 -176
rect 3726 -180 3760 -176
rect 2928 -248 3014 -216
rect 2956 -260 3014 -248
rect 3032 -260 3036 -254
rect 2956 -264 3036 -260
rect 2956 -286 2976 -264
rect 2926 -291 2934 -287
rect 2880 -295 2934 -291
rect 2968 -288 2976 -286
rect 2982 -288 3036 -264
rect 2968 -295 3034 -288
rect 2880 -325 2940 -295
rect 2900 -327 2940 -325
rect 2962 -319 3034 -295
rect 2962 -325 3022 -319
rect 2962 -327 2968 -325
rect 2988 -327 3022 -325
rect 3082 -327 3558 -185
rect 3626 -191 3766 -180
rect 3631 -195 3766 -191
rect 3632 -197 3766 -195
rect 3820 -185 3826 -169
rect 3833 -185 4628 -169
rect 5133 -181 5139 -164
rect 3638 -207 3760 -197
rect 3646 -225 3746 -207
rect 3646 -237 3684 -225
rect 3692 -231 3708 -225
rect 3638 -240 3684 -237
rect 3714 -237 3746 -225
rect 3820 -234 4628 -185
rect 4728 -209 5150 -181
rect 4728 -234 5167 -209
rect 3714 -240 3760 -237
rect 3618 -258 3684 -240
rect 3618 -259 3638 -258
rect 3664 -263 3684 -258
rect 3706 -258 3760 -240
rect 3820 -247 5167 -234
rect 5173 -247 5201 -243
rect 5233 -247 5241 -240
rect 3706 -259 3726 -258
rect 3714 -263 3722 -259
rect 3606 -327 3612 -263
rect 3618 -296 3652 -275
rect 3632 -327 3652 -296
rect 3672 -302 3680 -263
rect 3694 -270 3722 -263
rect 3800 -270 4648 -247
rect 4764 -251 4799 -247
rect 3694 -274 3744 -270
rect 3694 -308 3750 -274
rect 3666 -327 3750 -308
rect 3800 -284 4702 -270
rect 3800 -302 4711 -284
rect 4730 -302 4745 -270
rect 4764 -302 4798 -251
rect 4917 -300 4996 -285
rect 3800 -327 4997 -302
rect 2381 -427 4997 -327
rect 5097 -319 5354 -247
rect 5097 -334 5365 -319
rect 1839 -482 2296 -428
rect 2381 -460 5012 -427
rect 5097 -459 5354 -334
rect 2364 -464 5012 -460
rect 1839 -634 2281 -482
rect 2324 -581 2350 -482
rect 2364 -499 4294 -464
rect 2364 -514 4279 -499
rect 2364 -517 4310 -514
rect 2364 -564 3941 -517
rect 2364 -611 3172 -564
rect 3201 -611 3204 -564
rect 2364 -615 3204 -611
rect 2364 -616 3216 -615
rect 1790 -636 2281 -634
rect 1679 -680 1756 -636
rect 1786 -680 2281 -636
rect 2336 -627 3216 -616
rect 3235 -627 3269 -564
rect 2336 -631 3189 -627
rect 3201 -631 3204 -627
rect 2336 -637 3172 -631
rect 2336 -650 3189 -637
rect 2364 -662 3189 -650
rect 1679 -684 1744 -680
rect 1798 -681 2281 -680
rect 1798 -684 1828 -681
rect 1679 -690 1713 -684
rect 1821 -690 1828 -684
rect 1837 -690 2281 -681
rect 1502 -709 2281 -690
rect 1526 -724 2281 -709
rect 1448 -738 1518 -734
rect 1626 -737 1660 -724
rect 1394 -768 1518 -738
rect 1553 -758 1660 -737
rect 1394 -772 1421 -768
rect 1441 -772 1518 -768
rect 1461 -784 1518 -772
rect 1423 -836 1564 -804
rect 1626 -836 1660 -758
rect 1679 -783 1713 -724
rect 1859 -730 2281 -724
rect 2381 -676 3189 -662
rect 2381 -729 2803 -676
rect 1723 -770 1806 -736
rect 1859 -737 2302 -730
rect 2919 -736 2953 -676
rect 3054 -677 3073 -676
rect 3033 -680 3073 -677
rect 1679 -792 1840 -783
rect 1859 -792 2281 -737
rect 2285 -738 2302 -737
rect 2319 -764 2336 -738
rect 2294 -772 2299 -764
rect 2831 -770 2953 -736
rect 3021 -695 3073 -680
rect 3021 -725 3079 -695
rect 3021 -730 3073 -725
rect 3082 -730 3101 -676
rect 3142 -677 3161 -676
rect 3121 -680 3161 -677
rect 3121 -695 3167 -680
rect 3170 -689 3189 -676
rect 3109 -703 3167 -695
rect 3109 -725 3169 -703
rect 3021 -737 3067 -730
rect 3121 -737 3169 -725
rect 3235 -736 3246 -627
rect 3021 -740 3178 -737
rect 1679 -813 2281 -792
rect 1679 -817 1927 -813
rect 1968 -817 2029 -813
rect 2919 -817 2953 -770
rect 3033 -771 3178 -740
rect 3033 -815 3067 -771
rect 1310 -847 1394 -836
rect 1423 -838 1591 -836
rect 1310 -864 1383 -847
rect 1310 -870 1406 -864
rect 1423 -870 1598 -838
rect 1645 -851 1660 -836
rect 1968 -842 1983 -817
rect 1996 -842 2011 -826
rect 2026 -842 2029 -826
rect 1739 -851 1773 -842
rect 1827 -851 1861 -842
rect 2038 -851 2063 -822
rect 2889 -851 2953 -817
rect 3011 -833 3067 -815
rect 3121 -833 3155 -771
rect 3235 -813 3246 -802
rect 3011 -835 3033 -833
rect 3030 -851 3057 -845
rect 3127 -849 3155 -833
rect 3167 -835 3179 -815
rect 3235 -817 3237 -813
rect 3254 -817 3269 -631
rect 3215 -835 3269 -817
rect 3161 -851 3189 -835
rect 3215 -851 3283 -835
rect 3288 -839 3322 -564
rect 3346 -631 3356 -564
rect 3430 -571 3941 -564
rect 3430 -574 3907 -571
rect 3926 -574 3941 -571
rect 3973 -573 4060 -517
rect 4172 -518 4310 -517
rect 4065 -568 4094 -534
rect 3368 -584 3380 -574
rect 3430 -581 3926 -574
rect 3368 -586 3386 -584
rect 3448 -586 3926 -581
rect 3364 -615 3386 -586
rect 3434 -597 3926 -586
rect 3402 -608 3926 -597
rect 3402 -612 3414 -608
rect 3396 -613 3414 -612
rect 3368 -627 3386 -615
rect 3392 -624 3422 -613
rect 3434 -615 3926 -608
rect 3448 -624 3926 -615
rect 3396 -627 3436 -624
rect 3368 -689 3380 -627
rect 3392 -653 3436 -627
rect 3456 -636 3926 -624
rect 3973 -584 4081 -573
rect 4140 -584 4276 -518
rect 3973 -636 4060 -584
rect 4079 -615 4113 -602
rect 4128 -615 4276 -584
rect 4063 -627 4276 -615
rect 4294 -627 4310 -518
rect 4342 -528 4484 -464
rect 4498 -465 4502 -464
rect 4503 -465 4512 -464
rect 4514 -465 4548 -464
rect 4342 -544 4390 -528
rect 4342 -553 4376 -544
rect 4395 -553 4463 -528
rect 4475 -540 4484 -528
rect 4475 -544 4478 -540
rect 4342 -587 4468 -553
rect 4503 -568 4548 -465
rect 4063 -631 4294 -627
rect 4063 -636 4098 -631
rect 4102 -635 4294 -631
rect 4102 -636 4306 -635
rect 3456 -653 4306 -636
rect 3396 -665 3414 -653
rect 3396 -680 3408 -665
rect 3390 -695 3408 -680
rect 3390 -725 3448 -695
rect 3390 -740 3405 -725
rect 3456 -730 3468 -653
rect 3484 -695 3524 -653
rect 3529 -654 3562 -653
rect 3529 -670 3558 -654
rect 3570 -670 3595 -653
rect 3529 -695 3536 -670
rect 3478 -725 3536 -695
rect 3484 -730 3496 -725
rect 3521 -740 3536 -725
rect 3604 -725 3638 -653
rect 3604 -736 3615 -725
rect 3434 -839 3492 -833
rect 3288 -851 3317 -839
rect 1107 -923 1159 -912
rect 1179 -923 1231 -912
rect 1968 -919 1983 -898
rect 1996 -947 2011 -898
rect 203 -1020 341 -995
rect 433 -1010 567 -995
rect 2919 -994 2957 -851
rect 3011 -866 3057 -851
rect 3005 -871 3057 -866
rect 2977 -960 2983 -894
rect 3005 -960 3011 -871
rect 3027 -957 3057 -871
rect 3065 -892 3123 -886
rect 3061 -926 3104 -892
rect 3149 -926 3158 -851
rect 3161 -871 3193 -851
rect 3161 -883 3189 -871
rect 3065 -932 3123 -926
rect 3235 -932 3317 -851
rect 3434 -873 3446 -839
rect 3471 -873 3492 -839
rect 3434 -879 3492 -873
rect 3499 -907 3520 -805
rect 3027 -960 3051 -957
rect 2977 -973 3011 -960
rect 3039 -964 3045 -960
rect 2977 -994 3045 -973
rect 3161 -994 3207 -960
rect 3235 -994 3283 -932
rect 3288 -975 3317 -932
rect 3623 -956 3638 -725
rect 3657 -776 3691 -653
rect 3771 -665 3802 -653
rect 3847 -661 4306 -653
rect 3847 -670 3905 -661
rect 3927 -670 4306 -661
rect 3847 -727 3893 -670
rect 3847 -739 3879 -727
rect 3657 -805 3699 -776
rect 3702 -777 3727 -776
rect 3775 -777 3889 -752
rect 3803 -805 3861 -780
rect 3657 -888 3691 -805
rect 3803 -820 3815 -805
rect 3803 -826 3861 -820
rect 3864 -832 3865 -820
rect 3973 -826 4007 -670
rect 3906 -836 3907 -832
rect 3973 -833 3984 -826
rect 3992 -833 4007 -826
rect 3973 -863 4007 -833
rect 3973 -874 3984 -863
rect 3657 -922 3692 -888
rect 3823 -899 3875 -888
rect 3895 -899 3947 -888
rect 3834 -911 3864 -899
rect 3906 -911 3936 -899
rect 3992 -903 4007 -863
rect 4026 -835 4060 -670
rect 4063 -681 4094 -670
rect 4106 -681 4129 -670
rect 4140 -674 4174 -670
rect 4140 -681 4163 -674
rect 4128 -683 4163 -681
rect 4194 -682 4212 -670
rect 4218 -671 4306 -670
rect 4216 -682 4306 -671
rect 4128 -686 4168 -683
rect 4194 -686 4206 -682
rect 4216 -686 4294 -682
rect 4140 -690 4163 -686
rect 4218 -689 4276 -686
rect 4342 -689 4376 -587
rect 4384 -621 4468 -587
rect 4509 -621 4548 -568
rect 4395 -635 4463 -621
rect 4514 -633 4548 -621
rect 4555 -481 5012 -464
rect 4555 -633 4997 -481
rect 5040 -580 5066 -481
rect 5080 -615 5354 -459
rect 4506 -635 4997 -633
rect 4395 -679 4472 -635
rect 4502 -679 4997 -635
rect 5052 -649 5354 -615
rect 5080 -661 5354 -649
rect 4395 -683 4460 -679
rect 4514 -680 4997 -679
rect 4514 -683 4544 -680
rect 4395 -689 4429 -683
rect 4537 -689 4544 -683
rect 4553 -689 4997 -680
rect 4218 -708 4997 -689
rect 4242 -723 4997 -708
rect 4164 -737 4234 -733
rect 4342 -736 4376 -723
rect 4110 -767 4234 -737
rect 4269 -757 4376 -736
rect 4110 -771 4137 -767
rect 4157 -771 4234 -767
rect 4177 -783 4234 -771
rect 4139 -835 4280 -803
rect 4342 -835 4376 -757
rect 4395 -782 4429 -723
rect 4575 -729 4997 -723
rect 5097 -728 5354 -661
rect 5468 -673 5483 -164
rect 5502 -605 5536 -145
rect 5648 -213 5706 -207
rect 5648 -247 5660 -213
rect 5648 -253 5706 -247
rect 5648 -503 5706 -497
rect 5648 -537 5660 -503
rect 5837 -530 5852 -111
rect 5871 -462 5905 -92
rect 5983 -231 6141 -204
rect 5979 -259 6025 -232
rect 6067 -259 6113 -232
rect 6017 -360 6075 -354
rect 6017 -394 6029 -360
rect 6017 -400 6075 -394
rect 5871 -496 5906 -462
rect 6206 -477 6221 -58
rect 6240 -409 6274 -39
rect 6386 -107 6444 -101
rect 6386 -141 6398 -107
rect 6386 -147 6444 -141
rect 6386 -307 6444 -301
rect 6386 -341 6398 -307
rect 6386 -347 6444 -341
rect 6240 -443 6275 -409
rect 6575 -443 6590 -5
rect 6609 -443 6643 14
rect 6755 -54 6813 -48
rect 6755 -88 6767 -54
rect 6755 -94 6813 -88
rect 6755 -344 6813 -338
rect 6755 -378 6767 -344
rect 6755 -384 6813 -378
rect 6609 -477 6624 -443
rect 6944 -461 6959 48
rect 6978 -393 7012 67
rect 7124 -1 7182 5
rect 7124 -35 7136 -1
rect 7124 -41 7182 -35
rect 7124 -291 7182 -285
rect 7124 -325 7136 -291
rect 7124 -331 7182 -325
rect 6978 -427 7013 -393
rect 5648 -543 5706 -537
rect 5502 -639 5537 -605
rect 4513 -735 5018 -729
rect 4439 -736 5018 -735
rect 4439 -748 4997 -736
rect 5001 -737 5018 -736
rect 4439 -769 4522 -748
rect 4395 -791 4556 -782
rect 4575 -791 4997 -748
rect 5035 -763 5052 -737
rect 5010 -771 5015 -763
rect 4395 -812 4997 -791
rect 4395 -816 4643 -812
rect 4688 -816 4745 -812
rect 4026 -846 4110 -835
rect 4139 -837 4307 -835
rect 4026 -863 4099 -846
rect 4026 -869 4122 -863
rect 4139 -869 4314 -837
rect 4361 -850 4376 -835
rect 4742 -841 4745 -825
rect 4455 -850 4489 -841
rect 4543 -850 4577 -841
rect 4754 -850 4779 -821
rect 5187 -827 5207 -777
rect 5215 -799 5235 -777
rect 3823 -922 3875 -911
rect 3895 -922 3947 -911
rect 5187 -947 5213 -827
rect 5215 -919 5241 -799
rect 433 -1020 553 -1010
rect 2919 -1019 3057 -994
rect 3149 -1009 3283 -994
rect 3149 -1019 3269 -1009
rect 4267 -1015 4295 -1008
rect 203 -1029 294 -1020
rect 480 -1029 532 -1020
rect 2919 -1028 3010 -1019
rect 3196 -1028 3248 -1019
rect 261 -1048 267 -1029
rect 2977 -1047 2983 -1028
rect 4267 -1031 4297 -1015
rect 4239 -1043 4267 -1036
rect 4239 -1059 4269 -1043
rect 2782 -1095 2819 -1072
rect 179 -1200 200 -1096
rect 207 -1228 228 -1096
rect 2754 -1123 2819 -1100
rect 207 -1274 295 -1267
rect 2743 -1276 2751 -1231
rect 2771 -1251 2779 -1203
rect 2773 -1259 2779 -1251
rect 2923 -1273 3011 -1266
rect 2745 -1287 2751 -1276
rect 179 -1302 267 -1295
rect 2895 -1301 2983 -1294
rect 261 -1495 267 -1302
rect 289 -1482 295 -1302
rect 2977 -1494 2983 -1301
rect 3005 -1481 3011 -1301
rect 2977 -1495 2982 -1494
rect 261 -1496 266 -1495
<< nwell >>
rect -107 1050 1084 1271
rect 1090 1272 2550 1351
rect 3799 1272 5354 1352
rect 1090 1050 5354 1272
rect -107 767 5354 1050
rect -107 366 1147 767
rect 1090 339 1147 366
rect 1148 367 5354 767
rect 1148 339 2550 367
rect 3805 340 5354 367
rect 1090 -327 2550 -248
rect 3800 -327 5354 -247
rect 1090 -328 5354 -327
rect -107 -803 5354 -328
rect -107 -804 3800 -803
rect 3806 -804 5354 -803
rect -107 -1232 5354 -804
rect -107 -1233 2550 -1232
rect 1090 -1260 2550 -1233
rect 3806 -1259 5354 -1232
<< pwell >>
rect 1084 1698 5353 1735
rect -107 1666 5353 1698
rect -107 1624 3277 1666
rect 3580 1624 5353 1666
rect -107 1352 5353 1624
rect -107 1351 3799 1352
rect -107 1271 1084 1351
rect 2550 1272 3799 1351
rect -107 339 1084 366
rect 2550 340 3800 367
rect 2550 339 5354 340
rect -107 259 5354 339
rect -107 256 2684 259
rect 3509 256 5354 259
rect -107 167 5354 256
rect -107 164 1905 167
rect 1957 164 5354 167
rect -107 -247 5354 164
rect -107 -248 3800 -247
rect -107 -328 1084 -248
rect 2550 -327 3800 -248
rect -107 -1260 1090 -1233
rect 2550 -1259 3806 -1232
rect 2550 -1260 5353 -1259
rect -107 -1605 5353 -1260
<< psubdiff >>
rect 319 1628 343 1663
rect 1201 1628 1225 1663
rect 1827 1626 1851 1661
rect 1976 1626 2000 1661
rect 2397 1629 2421 1664
rect 2558 1629 2582 1664
rect 3043 1629 3067 1664
rect 3923 1629 3947 1664
rect 4565 1629 4589 1663
rect 4672 1629 4696 1663
rect 5115 1630 5139 1664
rect 5321 1630 5345 1664
rect 557 29 581 63
rect 900 29 924 63
rect 3139 30 3163 64
rect 3253 30 3277 64
rect 3644 30 3668 64
rect 36 -1570 60 -1536
rect 292 -1570 316 -1536
rect 552 -1571 576 -1536
rect 1397 -1571 1421 -1536
rect 2405 -1571 2429 -1535
rect 2981 -1571 3005 -1535
rect 3268 -1570 3292 -1536
rect 3605 -1570 3629 -1536
rect 3741 -1570 3765 -1536
rect 3877 -1570 3901 -1536
<< nsubdiff >>
rect 564 826 603 860
rect 690 826 724 860
<< psubdiffcont >>
rect 343 1628 1201 1663
rect 1851 1626 1976 1661
rect 2421 1629 2558 1664
rect 3067 1629 3923 1664
rect 4589 1629 4672 1663
rect 5139 1630 5321 1664
rect 581 29 900 63
rect 3277 30 3644 64
rect 60 -1570 292 -1536
rect 576 -1571 1397 -1536
rect 2429 -1571 2981 -1535
rect 3292 -1570 3605 -1536
rect 3765 -1570 3877 -1536
<< nsubdiffcont >>
rect 603 826 690 860
<< poly >>
rect 1118 808 1148 1311
rect 640 381 706 397
rect 640 347 656 381
rect 690 366 706 381
rect 690 347 1006 366
rect 640 336 1006 347
rect 640 331 676 336
rect 976 -80 1006 336
rect 1118 339 1147 808
rect 3356 382 3422 398
rect 3356 348 3372 382
rect 3406 367 3422 382
rect 3406 348 3722 367
rect 1118 -294 1148 339
rect 3356 337 3722 348
rect 3356 332 3392 337
rect 3692 -21 3722 337
rect 3833 323 3863 325
rect 3833 307 3899 323
rect 3833 273 3849 307
rect 3883 273 3899 307
rect 3833 257 3899 273
rect 3833 -240 3863 257
<< polycont >>
rect 656 347 690 381
rect 3372 348 3406 382
rect 3849 273 3883 307
<< locali >>
rect 640 381 706 397
rect 640 347 656 381
rect 690 347 706 381
rect 640 331 706 347
rect 3356 382 3422 398
rect 3356 348 3372 382
rect 3406 348 3422 382
rect 3356 332 3422 348
rect 3833 307 3899 323
rect 3833 273 3849 307
rect 3883 273 3899 307
rect 3833 257 3899 273
<< viali >>
rect 319 1628 343 1663
rect 343 1628 1201 1663
rect 1201 1628 1225 1663
rect 1827 1626 1851 1661
rect 1851 1626 1976 1661
rect 1976 1626 2000 1661
rect 2397 1629 2421 1664
rect 2421 1629 2558 1664
rect 2558 1629 2582 1664
rect 3043 1629 3067 1664
rect 3067 1629 3923 1664
rect 3923 1629 3947 1664
rect 4565 1629 4589 1663
rect 4589 1629 4672 1663
rect 4672 1629 4696 1663
rect 5115 1630 5139 1664
rect 5139 1630 5321 1664
rect 5321 1630 5345 1664
rect 564 826 603 860
rect 603 826 690 860
rect 690 826 724 860
rect 656 347 690 381
rect 3372 348 3406 382
rect 3849 273 3883 307
rect 557 29 581 63
rect 581 29 900 63
rect 900 29 924 63
rect 3253 30 3277 64
rect 3277 30 3644 64
rect 3644 30 3668 64
rect 36 -1570 60 -1536
rect 60 -1570 292 -1536
rect 292 -1570 316 -1536
rect 552 -1571 576 -1536
rect 576 -1571 1397 -1536
rect 1397 -1571 1421 -1536
rect 2405 -1571 2429 -1535
rect 2429 -1571 2981 -1535
rect 2981 -1571 3005 -1535
rect 3268 -1570 3292 -1536
rect 3292 -1570 3605 -1536
rect 3605 -1570 3629 -1536
rect 3741 -1570 3765 -1536
rect 3765 -1570 3877 -1536
rect 3877 -1570 3901 -1536
<< metal1 >>
rect 307 1668 1237 1669
rect 53 1667 2011 1668
rect 53 1663 2012 1667
rect 53 1662 319 1663
rect 53 1628 65 1662
rect 307 1628 319 1662
rect 1225 1662 2012 1663
rect 1225 1628 1237 1662
rect 1815 1661 2012 1662
rect 1815 1628 1827 1661
rect 53 1626 1827 1628
rect 2000 1626 2012 1661
rect 53 1622 2012 1626
rect 2385 1664 2594 1670
rect 3031 1669 3959 1670
rect 2385 1629 2397 1664
rect 2582 1629 2594 1664
rect 2385 1623 2594 1629
rect 1815 1620 2012 1622
rect 2599 1617 2609 1669
rect 2661 1664 3959 1669
rect 2661 1663 3043 1664
rect 2661 1629 2742 1663
rect 2768 1629 2780 1663
rect 3031 1629 3043 1663
rect 3947 1629 3959 1664
rect 2661 1623 3959 1629
rect 3969 1664 5357 1670
rect 3969 1630 3981 1664
rect 4553 1663 4708 1664
rect 4553 1630 4565 1663
rect 3969 1629 4565 1630
rect 4696 1630 4708 1663
rect 5103 1630 5115 1664
rect 5345 1630 5357 1664
rect 4696 1629 5357 1630
rect 3969 1624 5357 1629
rect 4553 1623 4708 1624
rect 2661 1622 2768 1623
rect 2661 1617 2671 1622
rect 2551 1403 2556 1437
rect 5270 1404 5271 1438
rect -62 816 -52 868
rect 0 816 10 868
rect 480 866 665 868
rect 480 862 736 866
rect 480 826 492 862
rect 552 860 736 862
rect 552 826 564 860
rect 724 826 736 860
rect 480 820 736 826
rect 2546 821 2723 869
rect 3190 863 3377 869
rect 3190 827 3202 863
rect 3365 827 3377 863
rect 3190 821 3377 827
rect 4456 863 4582 869
rect 4456 829 4468 863
rect 4570 829 4582 863
rect 4456 823 4582 829
rect 4949 824 4959 869
rect 604 381 706 397
rect 565 367 571 373
rect 604 367 656 381
rect 565 365 656 367
rect 640 347 656 365
rect 690 347 706 381
rect 3320 382 3422 398
rect 3320 367 3372 382
rect 640 331 706 347
rect 2431 323 2718 358
rect 3356 348 3372 367
rect 3406 348 3422 382
rect 3356 332 3422 348
rect 2674 318 2718 323
rect 0 69 200 200
rect 1918 157 1952 306
rect 2674 266 2684 318
rect 2736 266 2746 318
rect 3833 307 3899 323
rect 3833 304 3849 307
rect 3353 273 3849 304
rect 3883 273 3899 307
rect 3353 270 3899 273
rect 3353 221 3387 270
rect 3833 257 3899 270
rect 2685 169 2695 221
rect 2747 169 2757 221
rect 3332 169 3342 221
rect 3394 169 3404 221
rect 3447 186 3457 238
rect 3509 220 3519 238
rect 3699 220 3709 233
rect 3509 186 3709 220
rect 3699 181 3709 186
rect 3761 181 3771 233
rect 2685 164 2747 169
rect 2525 163 2747 164
rect 1895 105 1905 157
rect 1957 105 1967 157
rect 2525 111 2535 163
rect 2587 130 2747 163
rect 2587 111 2597 130
rect 0 63 1088 69
rect 0 29 200 63
rect 489 29 501 63
rect 545 29 557 63
rect 924 29 936 63
rect 1076 29 1088 63
rect 0 23 1088 29
rect 1190 63 2486 69
rect 1190 29 1202 63
rect 2474 29 2486 63
rect 1190 23 2486 29
rect 0 0 200 23
rect 2599 18 2609 74
rect 2661 70 2671 74
rect 2661 64 3813 70
rect 2661 30 2747 64
rect 3127 30 3139 64
rect 3241 30 3253 64
rect 3668 30 3680 64
rect 3801 30 3813 64
rect 2661 24 3813 30
rect 4089 64 5253 70
rect 4089 30 4101 64
rect 5241 30 5253 64
rect 4089 24 5253 30
rect 2661 18 2671 24
rect 2555 -196 2556 -162
rect 5271 -195 5272 -161
rect 0 -400 200 -200
rect -62 -780 -52 -728
rect 0 -800 200 -600
rect 494 -737 633 -731
rect 494 -773 506 -737
rect 621 -773 633 -737
rect 494 -779 633 -773
rect 2549 -778 2731 -730
rect 3219 -736 3342 -730
rect 3219 -772 3231 -736
rect 3330 -772 3342 -736
rect 3219 -778 3342 -772
rect 0 -1200 200 -1000
rect 2819 -1100 2829 -1091
rect 2684 -1134 2829 -1100
rect 2684 -1242 2718 -1134
rect 2819 -1143 2829 -1134
rect 2881 -1143 2891 -1091
rect 3323 -1232 3324 -1201
rect 2411 -1276 2718 -1242
rect 0 -1530 200 -1400
rect 557 -1486 567 -1434
rect 619 -1486 629 -1434
rect 2590 -1466 2600 -1414
rect 2652 -1466 2662 -1414
rect 2599 -1529 2652 -1466
rect 2661 -1529 2671 -1525
rect 2393 -1530 3017 -1529
rect 0 -1535 5302 -1530
rect 0 -1536 2405 -1535
rect 0 -1570 36 -1536
rect 316 -1570 328 -1536
rect 540 -1570 552 -1536
rect 0 -1571 552 -1570
rect 1421 -1570 1433 -1536
rect 2393 -1570 2405 -1536
rect 1421 -1571 2405 -1570
rect 3005 -1536 5302 -1535
rect 3005 -1570 3017 -1536
rect 3256 -1570 3268 -1536
rect 3629 -1570 3641 -1536
rect 3729 -1570 3741 -1536
rect 3901 -1570 3913 -1536
rect 4144 -1570 4156 -1536
rect 5162 -1570 5174 -1536
rect 5290 -1570 5302 -1536
rect 3005 -1571 5302 -1570
rect 0 -1576 5302 -1571
rect 0 -1600 200 -1576
rect 540 -1577 1433 -1576
rect 2393 -1577 3017 -1576
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
<< via1 >>
rect 2609 1617 2661 1669
rect -52 816 0 868
rect 2684 266 2736 318
rect 2695 169 2747 221
rect 3342 169 3394 221
rect 3457 186 3509 238
rect 3709 181 3761 233
rect 1905 105 1957 157
rect 2535 111 2587 163
rect 2609 18 2661 74
rect -52 -780 0 -728
rect 2829 -1143 2881 -1091
rect 567 -1486 619 -1434
rect 2600 -1466 2652 -1414
<< metal2 >>
rect 2609 1669 2661 1679
rect 2609 1611 2661 1617
rect 2615 1607 2661 1611
rect 33 1207 35 1259
rect -52 868 0 878
rect -52 806 0 816
rect -52 -718 -18 806
rect 382 464 387 516
rect 1905 157 1957 164
rect 2535 163 2587 173
rect 1957 111 2535 129
rect 1957 105 2587 111
rect 1905 101 2587 105
rect 1905 95 2572 101
rect 1905 90 1957 95
rect 2615 84 2649 1607
rect 5179 1298 5180 1350
rect 2684 318 2736 328
rect 2736 266 3509 293
rect 2684 259 3509 266
rect 3457 238 3509 259
rect 2695 221 2747 231
rect 3342 221 3394 231
rect 2747 176 3342 210
rect 2695 159 2747 169
rect 3457 176 3509 186
rect 3342 159 3394 169
rect 3544 131 3579 532
rect 3709 233 3761 243
rect 3761 193 3839 227
rect 5315 204 5349 208
rect 3709 171 3761 181
rect 5146 168 5349 204
rect 2689 97 3579 131
rect 2615 74 2661 84
rect 2600 18 2609 74
rect 2600 8 2661 18
rect 34 -392 35 -340
rect -52 -728 0 -718
rect -52 -790 0 -780
rect 2600 -1404 2634 8
rect 2600 -1414 2652 -1404
rect 567 -1434 619 -1424
rect 2600 -1476 2652 -1466
rect 567 -1496 619 -1486
rect 588 -1514 619 -1496
rect 2689 -1514 2723 97
rect 5180 -301 5181 -249
rect 2829 -1091 2881 -1081
rect 2881 -1143 2949 -1109
rect 2829 -1153 2881 -1143
rect 2915 -1372 2949 -1143
rect 5315 -1325 5349 168
rect 2915 -1406 3895 -1372
rect 5315 -1402 5350 -1325
rect 5138 -1436 5350 -1402
rect 588 -1548 2723 -1514
use xor_lede  x3
timestamp 1624053917
transform 1 0 835 0 1 569
box -220 -2000 4428 1165
use xor_lede  x6
timestamp 1624053917
transform 1 0 2551 0 1 569
box -220 -2000 4428 1165
use bitc  bitc_1
timestamp 1624053917
transform 1 0 3799 0 1 11
box -1084 -1506 3564 3689
use bitc  bitc_3
timestamp 1624053917
transform 1 0 3800 0 1 -1588
box -1084 -1506 3564 3689
use bitc  bitc_2
timestamp 1624053917
transform 1 0 1084 0 1 -1589
box -1084 -1506 3564 3689
use bitc  bitc_0
timestamp 1624053917
transform 1 0 1083 0 1 10
box -1084 -1506 3564 3689
use xor_lede  x9
timestamp 1624053917
transform 1 0 4267 0 1 569
box -220 -2000 4428 1165
use xor_lede  x12
timestamp 1624053917
transform 1 0 5983 0 1 569
box -220 -2000 4428 1165
use and_lede  x2
timestamp 1624053917
transform 1 0 67 0 1 1081
box -67 -2000 2214 1147
use and_lede  x5
timestamp 1624053917
transform 1 0 1783 0 1 1081
box -67 -2000 2214 1147
use and_lede  x8
timestamp 1624053917
transform 1 0 3499 0 1 1081
box -67 -2000 2214 1147
use and_lede  x11
timestamp 1624053917
transform 1 0 5215 0 1 1081
box -67 -2000 2214 1147
<< labels >>
rlabel metal2 384 464 387 516 1 CE
rlabel metal2 33 1207 35 1259 1 Q0
rlabel metal2 34 -392 35 -340 1 Q1
rlabel metal2 5179 1298 5180 1350 1 Q2
rlabel metal2 5180 -301 5181 -249 1 Q3
rlabel metal1 2555 1403 2556 1437 1 Q0n
rlabel metal1 2555 -196 2556 -162 1 Q1n
rlabel metal1 5270 1404 5271 1438 1 Q2n
rlabel metal1 5271 -195 5272 -161 1 Q3n
rlabel metal1 3323 -1232 3324 -1201 1 Sout3
rlabel metal2 2600 -1414 2634 18 1 vss!
rlabel pwell 3741 -1570 3901 -1536 1 vss!
rlabel nwell 603 826 690 860 1 vdd!
rlabel metal1 1106 1288 1183 1359 1 CLK
rlabel metal1 2411 -1276 2718 -1242 1 CLR
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Q0
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 CE
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Q0n
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Q1
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Q1n
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Q2
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Q2n
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 Q3
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 Q3n
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 Sout3
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 vss
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 vdd
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 CLR
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 CLK
port 14 nsew
<< end >>
