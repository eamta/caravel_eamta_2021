magic
tech sky130A
magscale 1 2
timestamp 1620951170
<< metal1 >>
rect -1668 877 2296 910
rect -29 574 2003 607
rect -429 573 12 574
rect -1529 541 12 573
rect -1529 381 -1494 541
rect -434 517 -368 541
rect 1967 540 2003 574
rect -434 513 -383 517
rect -1282 493 -1212 499
rect -1282 481 -1276 493
rect -1409 447 -1276 481
rect -1282 435 -1276 447
rect -1218 481 -1212 493
rect -418 488 -383 513
rect 120 512 190 518
rect -1218 447 -518 481
rect 120 454 126 512
rect 184 454 190 512
rect 120 448 190 454
rect -1218 435 -1212 447
rect -1282 429 -1212 435
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect -552 373 -518 447
rect -552 339 -296 373
rect -49 342 223 373
rect 810 367 880 373
rect -49 266 -18 342
rect 810 309 816 367
rect 874 309 880 367
rect 810 303 880 309
rect 1967 305 2002 540
rect 2226 318 2296 324
rect 2226 305 2232 318
rect -542 235 -18 266
rect 1967 271 2232 305
rect -542 184 -511 235
rect 1967 185 2002 271
rect 2226 260 2232 271
rect 2290 260 2296 318
rect 2226 254 2296 260
rect -1668 0 2296 33
<< via1 >>
rect -1276 435 -1218 493
rect 126 454 184 512
rect -1110 352 -1052 410
rect 816 309 874 367
rect 2232 260 2290 318
<< metal2 >>
rect 120 512 190 910
rect -1282 493 -1212 498
rect -1282 435 -1276 493
rect -1218 435 -1212 493
rect -1282 429 -1212 435
rect 120 454 126 512
rect 184 454 190 512
rect -1116 410 -1046 416
rect -1116 352 -1110 410
rect -1052 352 -1046 410
rect -1116 346 -1046 352
rect 120 0 190 454
rect 810 367 880 910
rect 810 309 816 367
rect 874 309 880 367
rect 810 0 880 309
rect 2226 318 2296 324
rect 2226 260 2232 318
rect 2290 260 2296 318
rect 2226 254 2296 260
use and  and_0
timestamp 1620950905
transform 1 0 -1632 0 1 344
box -36 -344 582 566
use xor  xor_0
timestamp 1620674245
transform 1 0 -1756 0 1 102
box 706 -102 1756 808
use dffc  dffc_0
timestamp 1620659937
transform 1 0 66 0 1 106
box -66 -106 2230 804
<< labels >>
rlabel metal2 845 910 845 910 1 CLR
rlabel metal2 2296 288 2296 288 3 Dn
rlabel metal2 157 910 157 910 1 CLK
rlabel metal2 -1246 498 -1246 498 1 CE
rlabel metal2 -1081 346 -1081 346 5 Sout
rlabel metal1 260 910 260 910 1 VDD
rlabel metal1 226 0 226 0 5 VSS
rlabel metal1 15 16 15 16 5 VSS
rlabel space 15 852 15 852 5 VDD
<< end >>
