magic
tech sky130A
timestamp 1616191617
<< nwell >>
rect 1539 1212 1676 1213
rect 608 891 961 1211
rect 1533 893 2935 1212
<< pwell >>
rect 606 415 1786 836
rect 2776 -54 2804 -16
<< poly >>
rect 892 1268 935 1281
rect 892 1250 905 1268
rect 922 1250 935 1268
rect 892 1238 935 1250
rect 1571 1180 1590 1181
rect 2556 1180 2576 1181
rect 1571 1155 2576 1180
rect 1571 1093 1590 1155
rect 1277 1070 1590 1093
rect 765 848 807 876
rect 765 831 779 848
rect 796 831 807 848
rect 856 846 982 876
rect 1114 867 1145 876
rect 1114 849 1122 867
rect 1139 849 1145 867
rect 1114 837 1145 849
rect 1567 869 1593 870
rect 1567 839 1598 869
rect 765 808 807 831
rect 1567 384 1593 839
rect 2556 773 2576 1155
rect 2556 743 2612 773
rect 2597 708 2612 743
rect 2597 704 2637 708
rect 2597 679 2667 704
rect 1538 352 1618 384
rect 1538 314 1558 352
rect 1598 314 1618 352
rect 1538 289 1618 314
rect 2748 151 2774 157
rect 2719 119 2799 151
rect 2719 81 2739 119
rect 2779 81 2799 119
rect 2719 56 2799 81
rect 2484 -25 2507 56
rect 2752 -25 2775 56
rect 2484 -48 2776 -25
<< polycont >>
rect 905 1250 922 1268
rect 779 831 796 848
rect 1122 849 1139 867
rect 1558 314 1598 352
rect 2739 81 2779 119
<< locali >>
rect 897 1271 928 1278
rect 897 1244 900 1271
rect 925 1244 928 1271
rect 897 1238 928 1244
rect 1114 870 1145 877
rect 767 856 805 858
rect 767 823 770 856
rect 802 823 805 856
rect 1114 843 1117 870
rect 1142 843 1145 870
rect 1114 837 1145 843
rect 767 819 805 823
rect 1537 370 1618 371
rect 1537 302 1545 370
rect 1611 302 1618 370
rect 2718 137 2799 138
rect 2718 69 2726 137
rect 2792 69 2799 137
<< viali >>
rect 900 1268 925 1271
rect 900 1250 905 1268
rect 905 1250 922 1268
rect 922 1250 925 1268
rect 900 1244 925 1250
rect 770 848 802 856
rect 770 831 779 848
rect 779 831 796 848
rect 796 831 802 848
rect 770 823 802 831
rect 1117 867 1142 870
rect 1117 849 1122 867
rect 1122 849 1139 867
rect 1139 849 1142 867
rect 1117 843 1142 849
rect 1545 352 1611 370
rect 1545 314 1558 352
rect 1558 314 1598 352
rect 1598 314 1611 352
rect 1545 298 1611 314
rect 2726 119 2792 137
rect 2726 81 2739 119
rect 2739 81 2779 119
rect 2779 81 2792 119
rect 2726 65 2792 81
<< metal1 >>
rect 847 1276 936 1281
rect 847 1239 897 1276
rect 892 1238 897 1239
rect 929 1239 936 1276
rect 929 1238 935 1239
rect 608 1104 931 1210
rect 1114 875 1145 876
rect 545 848 627 871
rect 767 856 805 863
rect 767 854 770 856
rect 802 854 805 856
rect 766 825 770 854
rect 802 825 806 854
rect 1109 837 1114 875
rect 1146 837 1151 875
rect 767 823 770 825
rect 802 823 805 825
rect 767 817 805 823
rect 1548 800 1566 820
rect 1536 742 1566 800
rect 1548 651 1566 742
rect 2529 655 2534 696
rect 2563 655 2568 696
rect 1548 610 1717 651
rect 1538 370 1618 384
rect 1538 298 1545 370
rect 1611 298 1618 370
rect 1538 289 1618 298
rect 2719 137 2799 151
rect 2719 65 2726 137
rect 2792 65 2799 137
rect 2719 56 2799 65
<< via1 >>
rect 897 1271 929 1276
rect 897 1244 900 1271
rect 900 1244 925 1271
rect 925 1244 929 1271
rect 897 1238 929 1244
rect 771 825 801 854
rect 1114 870 1146 875
rect 1114 843 1117 870
rect 1117 843 1142 870
rect 1142 843 1146 870
rect 1114 837 1146 843
rect 2534 655 2563 696
rect 1545 298 1611 370
rect 2726 65 2792 137
<< metal2 >>
rect 847 1276 936 1281
rect 847 1239 897 1276
rect 892 1238 897 1239
rect 929 1239 936 1276
rect 929 1238 935 1239
rect 904 869 924 1238
rect 1109 875 1146 880
rect 1109 869 1114 875
rect 779 866 1114 869
rect 769 854 1114 866
rect 769 840 771 854
rect 801 837 1114 854
rect 1146 837 1150 851
rect 801 835 1142 837
rect 771 820 801 825
rect 2534 696 2563 701
rect 2534 650 2563 655
rect 1545 370 1611 375
rect 1545 293 1611 298
rect 2726 137 2792 142
rect 2726 60 2792 65
use and  and_0
timestamp 1616191617
transform -1 0 918 0 1 893
box 0 -319 312 304
use xor2  xor2_0
timestamp 1616170071
transform -1 0 1538 0 1 893
box -26 -454 618 319
use dffc  dffc_0
timestamp 1616191617
transform 1 0 2027 0 1 396
box -433 -545 907 731
<< end >>
