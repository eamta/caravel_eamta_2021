magic
tech sky130A
magscale 1 2
timestamp 1619111721
<< pwell >>
rect -759 -630 759 630
<< nmos >>
rect -563 -420 -473 420
rect -415 -420 -325 420
rect -267 -420 -177 420
rect -119 -420 -29 420
rect 29 -420 119 420
rect 177 -420 267 420
rect 325 -420 415 420
rect 473 -420 563 420
<< ndiff >>
rect -621 408 -563 420
rect -621 -408 -609 408
rect -575 -408 -563 408
rect -621 -420 -563 -408
rect -473 408 -415 420
rect -473 -408 -461 408
rect -427 -408 -415 408
rect -473 -420 -415 -408
rect -325 408 -267 420
rect -325 -408 -313 408
rect -279 -408 -267 408
rect -325 -420 -267 -408
rect -177 408 -119 420
rect -177 -408 -165 408
rect -131 -408 -119 408
rect -177 -420 -119 -408
rect -29 408 29 420
rect -29 -408 -17 408
rect 17 -408 29 408
rect -29 -420 29 -408
rect 119 408 177 420
rect 119 -408 131 408
rect 165 -408 177 408
rect 119 -420 177 -408
rect 267 408 325 420
rect 267 -408 279 408
rect 313 -408 325 408
rect 267 -420 325 -408
rect 415 408 473 420
rect 415 -408 427 408
rect 461 -408 473 408
rect 415 -420 473 -408
rect 563 408 621 420
rect 563 -408 575 408
rect 609 -408 621 408
rect 563 -420 621 -408
<< ndiffc >>
rect -609 -408 -575 408
rect -461 -408 -427 408
rect -313 -408 -279 408
rect -165 -408 -131 408
rect -17 -408 17 408
rect 131 -408 165 408
rect 279 -408 313 408
rect 427 -408 461 408
rect 575 -408 609 408
<< psubdiff >>
rect -723 560 -627 594
rect 627 560 723 594
rect -723 498 -689 560
rect 689 498 723 560
rect -723 -560 -689 -498
rect 689 -560 723 -498
rect -723 -594 -627 -560
rect 627 -594 723 -560
<< psubdiffcont >>
rect -627 560 627 594
rect -723 -498 -689 498
rect 689 -498 723 498
rect -627 -594 627 -560
<< poly >>
rect -563 492 -473 508
rect -563 458 -547 492
rect -489 458 -473 492
rect -563 420 -473 458
rect -415 492 -325 508
rect -415 458 -399 492
rect -341 458 -325 492
rect -415 420 -325 458
rect -267 492 -177 508
rect -267 458 -251 492
rect -193 458 -177 492
rect -267 420 -177 458
rect -119 492 -29 508
rect -119 458 -103 492
rect -45 458 -29 492
rect -119 420 -29 458
rect 29 492 119 508
rect 29 458 45 492
rect 103 458 119 492
rect 29 420 119 458
rect 177 492 267 508
rect 177 458 193 492
rect 251 458 267 492
rect 177 420 267 458
rect 325 492 415 508
rect 325 458 341 492
rect 399 458 415 492
rect 325 420 415 458
rect 473 492 563 508
rect 473 458 489 492
rect 547 458 563 492
rect 473 420 563 458
rect -563 -458 -473 -420
rect -563 -492 -547 -458
rect -489 -492 -473 -458
rect -563 -508 -473 -492
rect -415 -458 -325 -420
rect -415 -492 -399 -458
rect -341 -492 -325 -458
rect -415 -508 -325 -492
rect -267 -458 -177 -420
rect -267 -492 -251 -458
rect -193 -492 -177 -458
rect -267 -508 -177 -492
rect -119 -458 -29 -420
rect -119 -492 -103 -458
rect -45 -492 -29 -458
rect -119 -508 -29 -492
rect 29 -458 119 -420
rect 29 -492 45 -458
rect 103 -492 119 -458
rect 29 -508 119 -492
rect 177 -458 267 -420
rect 177 -492 193 -458
rect 251 -492 267 -458
rect 177 -508 267 -492
rect 325 -458 415 -420
rect 325 -492 341 -458
rect 399 -492 415 -458
rect 325 -508 415 -492
rect 473 -458 563 -420
rect 473 -492 489 -458
rect 547 -492 563 -458
rect 473 -508 563 -492
<< polycont >>
rect -547 458 -489 492
rect -399 458 -341 492
rect -251 458 -193 492
rect -103 458 -45 492
rect 45 458 103 492
rect 193 458 251 492
rect 341 458 399 492
rect 489 458 547 492
rect -547 -492 -489 -458
rect -399 -492 -341 -458
rect -251 -492 -193 -458
rect -103 -492 -45 -458
rect 45 -492 103 -458
rect 193 -492 251 -458
rect 341 -492 399 -458
rect 489 -492 547 -458
<< locali >>
rect -723 560 -627 594
rect 627 560 723 594
rect -723 498 -689 560
rect 689 498 723 560
rect -563 458 -547 492
rect -489 458 -473 492
rect -415 458 -399 492
rect -341 458 -325 492
rect -267 458 -251 492
rect -193 458 -177 492
rect -119 458 -103 492
rect -45 458 -29 492
rect 29 458 45 492
rect 103 458 119 492
rect 177 458 193 492
rect 251 458 267 492
rect 325 458 341 492
rect 399 458 415 492
rect 473 458 489 492
rect 547 458 563 492
rect -609 408 -575 424
rect -609 -424 -575 -408
rect -461 408 -427 424
rect -461 -424 -427 -408
rect -313 408 -279 424
rect -313 -424 -279 -408
rect -165 408 -131 424
rect -165 -424 -131 -408
rect -17 408 17 424
rect -17 -424 17 -408
rect 131 408 165 424
rect 131 -424 165 -408
rect 279 408 313 424
rect 279 -424 313 -408
rect 427 408 461 424
rect 427 -424 461 -408
rect 575 408 609 424
rect 575 -424 609 -408
rect -563 -492 -547 -458
rect -489 -492 -473 -458
rect -415 -492 -399 -458
rect -341 -492 -325 -458
rect -267 -492 -251 -458
rect -193 -492 -177 -458
rect -119 -492 -103 -458
rect -45 -492 -29 -458
rect 29 -492 45 -458
rect 103 -492 119 -458
rect 177 -492 193 -458
rect 251 -492 267 -458
rect 325 -492 341 -458
rect 399 -492 415 -458
rect 473 -492 489 -458
rect 547 -492 563 -458
rect -723 -560 -689 -498
rect 689 -560 723 -498
rect -723 -594 -627 -560
rect 627 -594 723 -560
<< viali >>
rect -547 458 -489 492
rect -399 458 -341 492
rect -251 458 -193 492
rect -103 458 -45 492
rect 45 458 103 492
rect 193 458 251 492
rect 341 458 399 492
rect 489 458 547 492
rect -609 -408 -575 408
rect -461 -408 -427 408
rect -313 -408 -279 408
rect -165 -408 -131 408
rect -17 -408 17 408
rect 131 -408 165 408
rect 279 -408 313 408
rect 427 -408 461 408
rect 575 -408 609 408
rect -547 -492 -489 -458
rect -399 -492 -341 -458
rect -251 -492 -193 -458
rect -103 -492 -45 -458
rect 45 -492 103 -458
rect 193 -492 251 -458
rect 341 -492 399 -458
rect 489 -492 547 -458
<< metal1 >>
rect -559 492 -477 498
rect -559 458 -547 492
rect -489 458 -477 492
rect -559 452 -477 458
rect -411 492 -329 498
rect -411 458 -399 492
rect -341 458 -329 492
rect -411 452 -329 458
rect -263 492 -181 498
rect -263 458 -251 492
rect -193 458 -181 492
rect -263 452 -181 458
rect -115 492 -33 498
rect -115 458 -103 492
rect -45 458 -33 492
rect -115 452 -33 458
rect 33 492 115 498
rect 33 458 45 492
rect 103 458 115 492
rect 33 452 115 458
rect 181 492 263 498
rect 181 458 193 492
rect 251 458 263 492
rect 181 452 263 458
rect 329 492 411 498
rect 329 458 341 492
rect 399 458 411 492
rect 329 452 411 458
rect 477 492 559 498
rect 477 458 489 492
rect 547 458 559 492
rect 477 452 559 458
rect -615 408 -569 420
rect -615 -408 -609 408
rect -575 -408 -569 408
rect -615 -420 -569 -408
rect -467 408 -421 420
rect -467 -408 -461 408
rect -427 -408 -421 408
rect -467 -420 -421 -408
rect -319 408 -273 420
rect -319 -408 -313 408
rect -279 -408 -273 408
rect -319 -420 -273 -408
rect -171 408 -125 420
rect -171 -408 -165 408
rect -131 -408 -125 408
rect -171 -420 -125 -408
rect -23 408 23 420
rect -23 -408 -17 408
rect 17 -408 23 408
rect -23 -420 23 -408
rect 125 408 171 420
rect 125 -408 131 408
rect 165 -408 171 408
rect 125 -420 171 -408
rect 273 408 319 420
rect 273 -408 279 408
rect 313 -408 319 408
rect 273 -420 319 -408
rect 421 408 467 420
rect 421 -408 427 408
rect 461 -408 467 408
rect 421 -420 467 -408
rect 569 408 615 420
rect 569 -408 575 408
rect 609 -408 615 408
rect 569 -420 615 -408
rect -559 -458 -477 -452
rect -559 -492 -547 -458
rect -489 -492 -477 -458
rect -559 -498 -477 -492
rect -411 -458 -329 -452
rect -411 -492 -399 -458
rect -341 -492 -329 -458
rect -411 -498 -329 -492
rect -263 -458 -181 -452
rect -263 -492 -251 -458
rect -193 -492 -181 -458
rect -263 -498 -181 -492
rect -115 -458 -33 -452
rect -115 -492 -103 -458
rect -45 -492 -33 -458
rect -115 -498 -33 -492
rect 33 -458 115 -452
rect 33 -492 45 -458
rect 103 -492 115 -458
rect 33 -498 115 -492
rect 181 -458 263 -452
rect 181 -492 193 -458
rect 251 -492 263 -458
rect 181 -498 263 -492
rect 329 -458 411 -452
rect 329 -492 341 -458
rect 399 -492 411 -458
rect 329 -498 411 -492
rect 477 -458 559 -452
rect 477 -492 489 -458
rect 547 -492 559 -458
rect 477 -498 559 -492
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -706 -577 706 577
string parameters w 4.2 l 0.45 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
