magic
tech sky130A
magscale 1 2
timestamp 1616195620
<< nwell >>
rect -36 663 470 764
<< psubdiff >>
rect 18 -30 42 4
rect 430 -30 454 4
<< nsubdiff >>
rect 131 694 186 728
rect 322 694 380 728
<< psubdiffcont >>
rect 42 -30 430 4
<< nsubdiffcont >>
rect 186 694 322 728
<< poly >>
rect 58 322 88 396
rect 146 336 176 402
rect 238 354 304 370
rect 346 354 376 398
rect -36 310 88 322
rect -36 276 -19 310
rect 15 276 88 310
rect -36 266 88 276
rect 130 326 196 336
rect 130 292 146 326
rect 180 292 196 326
rect 238 320 254 354
rect 288 320 376 354
rect 238 303 304 320
rect 130 275 196 292
rect 58 244 88 266
rect 146 245 176 275
rect 58 215 88 223
rect 146 211 176 223
rect 346 174 376 320
<< polycont >>
rect -19 276 15 310
rect 146 292 180 326
rect 254 320 288 354
<< locali >>
rect -35 276 -19 310
rect 15 276 31 310
rect 130 292 146 326
rect 180 292 196 326
rect 238 320 254 354
rect 288 320 304 354
<< viali >>
rect 130 694 186 728
rect 186 694 322 728
rect 322 694 380 728
rect 130 693 380 694
rect -19 276 15 310
rect 146 292 180 326
rect 254 320 288 354
rect 17 4 454 5
rect 17 -30 42 4
rect 42 -30 430 4
rect 430 -30 454 4
<< metal1 >>
rect -36 728 470 764
rect -36 693 130 728
rect 380 693 470 728
rect -36 644 470 693
rect 6 544 52 644
rect 100 446 134 590
rect 182 571 228 644
rect 294 600 340 644
rect 100 434 140 446
rect 94 422 140 434
rect 400 428 428 459
rect 94 408 145 422
rect 95 401 145 408
rect 117 394 145 401
rect 117 393 296 394
rect -36 370 88 373
rect 117 370 302 393
rect 382 370 428 424
rect -36 345 89 370
rect 117 365 304 370
rect -36 310 33 317
rect -36 276 -19 310
rect 15 276 33 310
rect 61 316 89 345
rect 238 354 304 365
rect 130 326 196 334
rect 130 316 146 326
rect 61 292 146 316
rect 180 292 196 326
rect 238 320 254 354
rect 288 320 304 354
rect 238 306 304 320
rect 242 303 304 306
rect 61 288 196 292
rect 130 278 196 288
rect -36 268 33 276
rect 206 233 228 236
rect 261 233 304 303
rect 100 157 134 206
rect 182 205 184 213
rect 206 205 304 233
rect 189 192 304 205
rect 382 236 470 370
rect 189 189 228 192
rect 6 23 52 95
rect 100 59 140 157
rect 182 59 228 157
rect 382 147 428 236
rect 294 23 340 63
rect -36 5 470 23
rect -36 -30 17 5
rect 454 -30 470 5
rect -36 -36 470 -30
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_2
timestamp 1614978561
transform 1 0 361 0 1 512
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_0
timestamp 1614978561
transform 1 0 73 0 1 512
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5AYHFE  sky130_fd_pr__pfet_01v8_5AYHFE_1
timestamp 1614978561
transform 1 0 161 0 1 512
box -109 -152 109 152
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615298455
transform 1 0 361 0 1 104
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_0
timestamp 1614978561
transform 1 0 73 0 1 148
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_P8KVP3  sky130_fd_pr__nfet_01v8_P8KVP3_1
timestamp 1614978561
transform 1 0 161 0 1 148
box -73 -116 73 116
<< labels >>
rlabel metal1 -36 345 88 373 1 vb
rlabel metal1 -36 268 -19 317 1 va
rlabel nwell 130 693 380 728 1 vdd
rlabel metal1 17 -30 454 5 1 vss
rlabel metal1 382 236 470 370 1 out
<< end >>
