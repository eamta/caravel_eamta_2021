magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 298 1095 333 1112
rect 299 1094 333 1095
rect 299 1058 369 1094
rect 129 1027 187 1033
rect 129 993 141 1027
rect 316 1024 387 1058
rect 667 1024 702 1058
rect 129 987 187 993
rect 316 852 386 1024
rect 668 1005 702 1024
rect 498 956 556 962
rect 498 922 510 956
rect 498 916 556 922
rect 687 852 702 1005
rect 721 971 756 1005
rect 1036 971 1071 1005
rect 721 852 755 971
rect 1037 952 1071 971
rect 867 903 925 909
rect 867 869 879 903
rect 867 863 925 869
rect 85 782 231 816
rect -17 727 17 781
rect 63 738 83 776
rect 85 768 125 781
rect 85 766 140 768
rect 103 762 131 765
rect 143 749 167 782
rect 219 778 231 781
rect 183 766 231 778
rect 141 731 205 749
rect 243 738 253 776
rect 316 765 990 852
rect 49 727 51 731
rect 137 728 205 731
rect 141 727 205 728
rect 12 617 17 727
rect 37 617 71 727
rect 94 719 205 727
rect 125 685 205 719
rect 125 669 183 685
rect 168 654 183 669
rect 265 651 283 731
rect 249 617 283 651
rect 299 617 990 765
rect 37 583 183 617
rect 237 583 990 617
rect 137 543 171 583
rect 316 494 990 583
rect 685 485 990 494
rect 721 477 818 485
rect 1056 477 1071 952
rect 1090 918 1125 952
rect 1405 918 1440 952
rect 1090 477 1124 918
rect 1406 899 1440 918
rect 1792 899 1845 900
rect 1236 850 1294 856
rect 1236 816 1248 850
rect 1236 810 1294 816
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1090 443 1105 477
rect 1425 424 1440 899
rect 1459 865 1494 899
rect 1774 865 1845 899
rect 1459 424 1493 865
rect 1775 864 1845 865
rect 1792 830 1863 864
rect 2143 830 2178 864
rect 1605 797 1663 803
rect 1605 763 1617 797
rect 1605 757 1663 763
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 830
rect 2144 811 2178 830
rect 1974 762 2032 768
rect 1974 728 1986 762
rect 1974 722 2032 728
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2163 318 2178 811
rect 2197 777 2232 811
rect 2197 318 2231 777
rect 2343 709 2401 715
rect 2343 675 2355 709
rect 2513 686 2547 704
rect 2343 669 2401 675
rect 2513 650 2583 686
rect 2530 616 2601 650
rect 2881 616 2916 650
rect 3304 633 3339 651
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2530 265 2600 616
rect 2882 597 2916 616
rect 3268 618 3339 633
rect 3619 618 3654 652
rect 2712 548 2770 554
rect 2712 514 2724 548
rect 2712 508 2770 514
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
rect 2901 212 2916 597
rect 2935 563 2970 597
rect 2935 212 2969 563
rect 3081 495 3139 501
rect 3081 461 3093 495
rect 3081 455 3139 461
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2935 178 2950 212
rect 3268 159 3338 618
rect 3620 599 3654 618
rect 3450 550 3508 556
rect 3450 516 3462 550
rect 3450 510 3508 516
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3268 123 3321 159
rect 3639 106 3654 599
rect 3673 565 3708 599
rect 3988 565 4023 599
rect 3673 106 3707 565
rect 3989 546 4023 565
rect 3819 497 3877 503
rect 3819 463 3831 497
rect 3819 457 3877 463
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4008 53 4023 546
rect 4042 512 4077 546
rect 4042 53 4076 512
rect 4188 444 4246 450
rect 4188 410 4200 444
rect 4188 404 4246 410
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
<< nwell >>
rect -96 745 990 852
rect -96 741 4 745
rect 208 744 990 745
rect -96 485 3 741
rect 207 670 990 744
rect 883 485 990 670
<< psubdiff >>
rect -60 -17 58 17
rect 824 -17 954 17
<< nsubdiff >>
rect -60 782 389 816
rect 595 782 954 816
<< psubdiffcont >>
rect 58 -17 824 17
<< nsubdiffcont >>
rect 389 782 595 816
<< poly >>
rect 95 502 125 521
rect 295 516 325 526
rect 589 521 777 523
rect 275 502 341 516
rect 95 500 341 502
rect 95 468 291 500
rect 95 300 125 468
rect 275 466 291 468
rect 325 466 341 500
rect 275 450 341 466
rect 275 393 341 408
rect 383 393 413 521
rect 275 392 413 393
rect 275 358 292 392
rect 326 358 413 392
rect 275 342 341 358
rect 95 270 325 300
rect 383 277 413 358
rect 471 431 501 521
rect 559 489 807 521
rect 631 432 697 447
rect 631 431 698 432
rect 471 397 648 431
rect 682 397 719 431
rect 471 277 501 397
rect 631 381 697 397
rect 777 362 807 489
rect 777 346 862 362
rect 777 339 812 346
rect 559 312 812 339
rect 846 312 862 346
rect 559 305 862 312
rect 559 277 589 305
rect 777 296 862 305
rect 95 187 125 270
rect 777 187 807 296
<< polycont >>
rect 291 466 325 500
rect 292 358 326 392
rect 648 397 682 431
rect 812 312 846 346
<< locali >>
rect -60 782 389 816
rect 595 782 954 816
rect 275 466 291 500
rect 325 466 341 500
rect 631 397 648 431
rect 682 397 698 431
rect 275 358 292 392
rect 326 358 342 392
rect 796 312 812 346
rect 846 312 862 346
rect -60 -17 58 17
rect 824 -17 954 17
<< viali >>
rect 389 782 595 816
rect 291 466 325 500
rect 648 397 682 431
rect 292 358 326 392
rect 812 312 846 346
rect 58 -17 824 17
<< metal1 >>
rect -2 816 905 822
rect -2 782 389 816
rect 595 782 905 816
rect -2 776 905 782
rect 49 727 83 776
rect 243 727 289 776
rect 331 719 553 747
rect 595 727 641 776
rect 819 726 853 776
rect 417 676 469 686
rect 406 633 417 667
rect 469 633 479 667
rect 417 614 469 624
rect 137 392 171 547
rect 265 450 275 516
rect 341 450 351 516
rect 275 392 341 408
rect 137 358 292 392
rect 326 358 341 392
rect 137 200 171 358
rect 275 342 341 358
rect 425 307 459 547
rect 513 543 547 547
rect 631 431 697 447
rect 731 431 765 547
rect 631 397 648 431
rect 682 397 765 431
rect 631 381 697 397
rect 337 279 459 307
rect 507 279 697 307
rect 337 251 371 279
rect 507 251 553 279
rect 0 23 200 200
rect 669 23 697 279
rect 731 161 765 397
rect 796 361 862 362
rect 796 305 812 361
rect 868 305 878 361
rect 796 296 862 305
rect 819 23 853 71
rect -2 17 905 23
rect -2 -17 58 17
rect 824 -17 905 17
rect -2 -23 905 -17
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
<< via1 >>
rect 417 624 469 676
rect 275 500 341 516
rect 275 466 291 500
rect 291 466 325 500
rect 325 466 341 500
rect 275 450 341 466
rect 812 346 868 361
rect 812 312 846 346
rect 846 312 868 346
rect 812 305 868 312
<< metal2 >>
rect 406 624 417 676
rect 469 624 479 676
rect 275 516 341 526
rect 275 440 341 450
rect 812 361 868 371
rect 812 295 868 305
<< comment >>
rect 10 799 602 800
rect 816 799 893 800
rect 10 1 11 799
rect 892 1 893 799
rect 10 0 893 1
use sky130_fd_pr__nfet_01v8_NNQ2PV  sky130_fd_pr__nfet_01v8_NNQ2PV_0
timestamp 1615600491
transform 1 0 110 0 1 116
box -73 -71 73 71
use nmos_900_derecha  nmos_900_derecha_0
timestamp 1615566114
transform 1 0 310 0 1 167
box -73 -122 73 110
use nmos_900_dos  nmos_900_dos_1
timestamp 1615566114
transform 1 0 486 0 1 167
box -73 -122 73 110
use nmos_900_dos  nmos_900_dos_0
timestamp 1615566114
transform 1 0 398 0 1 167
box -73 -122 73 110
use nmos_900_izquierda  nmos_900_izquierda_0
timestamp 1615566114
transform 1 0 574 0 1 167
box -73 -122 73 110
use sky130_fd_pr__nfet_01v8_NNQ2PV  sky130_fd_pr__nfet_01v8_NNQ2PV_1
timestamp 1615600491
transform 1 0 792 0 1 116
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_L9ESED  XM7
timestamp 1624053917
transform 1 0 1634 0 1 635
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_XSLFBL  XM10
timestamp 1624053917
transform 1 0 2372 0 1 538
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM8
timestamp 1624053917
transform 1 0 2003 0 1 591
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 3479 0 1 379
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM11
timestamp 1624053917
transform 1 0 3110 0 1 378
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 2741 0 1 431
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM3
timestamp 1624053917
transform 1 0 4217 0 1 273
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 3848 0 1 326
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_1
timestamp 1615568138
transform 1 0 310 0 1 637
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_0
timestamp 1615568138
transform 1 0 110 0 1 637
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_2
timestamp 1615568138
transform 1 0 574 0 1 637
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_3
timestamp 1615568138
transform 1 0 792 0 1 637
box -109 -152 109 152
use pmos_900_derecho  pmos_900_derecho_0
timestamp 1615566114
transform 1 0 289 0 1 485
box 0 0 218 286
use pmos_900_izquierdo  pmos_900_izquierdo_0
timestamp 1615566114
transform 1 0 377 0 1 485
box 0 0 218 286
use sky130_fd_pr__nfet_01v8_L9ESED  XM6
timestamp 1624053917
transform 1 0 896 0 1 741
box -211 -300 211 300
use sky130_fd_pr__nfet_01v8_L9ESED  XM4
timestamp 1624053917
transform 1 0 527 0 1 794
box -211 -300 211 300
use sky130_fd_pr__pfet_01v8_XSLFBL  XM0
timestamp 1624053917
transform 1 0 158 0 1 856
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_L9ESED  XM5
timestamp 1624053917
transform 1 0 1265 0 1 688
box -211 -300 211 300
<< labels >>
rlabel metal2 275 450 341 516 1 A
rlabel metal1 347 -18 408 16 1 vss
rlabel metal2 812 305 868 361 1 B
rlabel nwell 86 782 816 816 1 vdd
rlabel via1 417 624 469 676 3 Z
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Z
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 A
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 B
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vss
port 5 nsew
<< end >>
