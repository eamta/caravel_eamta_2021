magic
tech sky130A
magscale 1 2
timestamp 1615920820
<< nwell >>
rect -4223 -3003 4223 3003
<< pmos >>
rect -4129 1541 -3989 2941
rect -3931 1541 -3791 2941
rect -3733 1541 -3593 2941
rect -3535 1541 -3395 2941
rect -3337 1541 -3197 2941
rect -3139 1541 -2999 2941
rect -2941 1541 -2801 2941
rect -2743 1541 -2603 2941
rect -2545 1541 -2405 2941
rect -2347 1541 -2207 2941
rect -2149 1541 -2009 2941
rect -1951 1541 -1811 2941
rect -1753 1541 -1613 2941
rect -1555 1541 -1415 2941
rect -1357 1541 -1217 2941
rect -1159 1541 -1019 2941
rect -961 1541 -821 2941
rect -763 1541 -623 2941
rect -565 1541 -425 2941
rect -367 1541 -227 2941
rect -169 1541 -29 2941
rect 29 1541 169 2941
rect 227 1541 367 2941
rect 425 1541 565 2941
rect 623 1541 763 2941
rect 821 1541 961 2941
rect 1019 1541 1159 2941
rect 1217 1541 1357 2941
rect 1415 1541 1555 2941
rect 1613 1541 1753 2941
rect 1811 1541 1951 2941
rect 2009 1541 2149 2941
rect 2207 1541 2347 2941
rect 2405 1541 2545 2941
rect 2603 1541 2743 2941
rect 2801 1541 2941 2941
rect 2999 1541 3139 2941
rect 3197 1541 3337 2941
rect 3395 1541 3535 2941
rect 3593 1541 3733 2941
rect 3791 1541 3931 2941
rect 3989 1541 4129 2941
rect -4129 47 -3989 1447
rect -3931 47 -3791 1447
rect -3733 47 -3593 1447
rect -3535 47 -3395 1447
rect -3337 47 -3197 1447
rect -3139 47 -2999 1447
rect -2941 47 -2801 1447
rect -2743 47 -2603 1447
rect -2545 47 -2405 1447
rect -2347 47 -2207 1447
rect -2149 47 -2009 1447
rect -1951 47 -1811 1447
rect -1753 47 -1613 1447
rect -1555 47 -1415 1447
rect -1357 47 -1217 1447
rect -1159 47 -1019 1447
rect -961 47 -821 1447
rect -763 47 -623 1447
rect -565 47 -425 1447
rect -367 47 -227 1447
rect -169 47 -29 1447
rect 29 47 169 1447
rect 227 47 367 1447
rect 425 47 565 1447
rect 623 47 763 1447
rect 821 47 961 1447
rect 1019 47 1159 1447
rect 1217 47 1357 1447
rect 1415 47 1555 1447
rect 1613 47 1753 1447
rect 1811 47 1951 1447
rect 2009 47 2149 1447
rect 2207 47 2347 1447
rect 2405 47 2545 1447
rect 2603 47 2743 1447
rect 2801 47 2941 1447
rect 2999 47 3139 1447
rect 3197 47 3337 1447
rect 3395 47 3535 1447
rect 3593 47 3733 1447
rect 3791 47 3931 1447
rect 3989 47 4129 1447
rect -4129 -1447 -3989 -47
rect -3931 -1447 -3791 -47
rect -3733 -1447 -3593 -47
rect -3535 -1447 -3395 -47
rect -3337 -1447 -3197 -47
rect -3139 -1447 -2999 -47
rect -2941 -1447 -2801 -47
rect -2743 -1447 -2603 -47
rect -2545 -1447 -2405 -47
rect -2347 -1447 -2207 -47
rect -2149 -1447 -2009 -47
rect -1951 -1447 -1811 -47
rect -1753 -1447 -1613 -47
rect -1555 -1447 -1415 -47
rect -1357 -1447 -1217 -47
rect -1159 -1447 -1019 -47
rect -961 -1447 -821 -47
rect -763 -1447 -623 -47
rect -565 -1447 -425 -47
rect -367 -1447 -227 -47
rect -169 -1447 -29 -47
rect 29 -1447 169 -47
rect 227 -1447 367 -47
rect 425 -1447 565 -47
rect 623 -1447 763 -47
rect 821 -1447 961 -47
rect 1019 -1447 1159 -47
rect 1217 -1447 1357 -47
rect 1415 -1447 1555 -47
rect 1613 -1447 1753 -47
rect 1811 -1447 1951 -47
rect 2009 -1447 2149 -47
rect 2207 -1447 2347 -47
rect 2405 -1447 2545 -47
rect 2603 -1447 2743 -47
rect 2801 -1447 2941 -47
rect 2999 -1447 3139 -47
rect 3197 -1447 3337 -47
rect 3395 -1447 3535 -47
rect 3593 -1447 3733 -47
rect 3791 -1447 3931 -47
rect 3989 -1447 4129 -47
rect -4129 -2941 -3989 -1541
rect -3931 -2941 -3791 -1541
rect -3733 -2941 -3593 -1541
rect -3535 -2941 -3395 -1541
rect -3337 -2941 -3197 -1541
rect -3139 -2941 -2999 -1541
rect -2941 -2941 -2801 -1541
rect -2743 -2941 -2603 -1541
rect -2545 -2941 -2405 -1541
rect -2347 -2941 -2207 -1541
rect -2149 -2941 -2009 -1541
rect -1951 -2941 -1811 -1541
rect -1753 -2941 -1613 -1541
rect -1555 -2941 -1415 -1541
rect -1357 -2941 -1217 -1541
rect -1159 -2941 -1019 -1541
rect -961 -2941 -821 -1541
rect -763 -2941 -623 -1541
rect -565 -2941 -425 -1541
rect -367 -2941 -227 -1541
rect -169 -2941 -29 -1541
rect 29 -2941 169 -1541
rect 227 -2941 367 -1541
rect 425 -2941 565 -1541
rect 623 -2941 763 -1541
rect 821 -2941 961 -1541
rect 1019 -2941 1159 -1541
rect 1217 -2941 1357 -1541
rect 1415 -2941 1555 -1541
rect 1613 -2941 1753 -1541
rect 1811 -2941 1951 -1541
rect 2009 -2941 2149 -1541
rect 2207 -2941 2347 -1541
rect 2405 -2941 2545 -1541
rect 2603 -2941 2743 -1541
rect 2801 -2941 2941 -1541
rect 2999 -2941 3139 -1541
rect 3197 -2941 3337 -1541
rect 3395 -2941 3535 -1541
rect 3593 -2941 3733 -1541
rect 3791 -2941 3931 -1541
rect 3989 -2941 4129 -1541
<< pdiff >>
rect -4187 2929 -4129 2941
rect -4187 1553 -4175 2929
rect -4141 1553 -4129 2929
rect -4187 1541 -4129 1553
rect -3989 2929 -3931 2941
rect -3989 1553 -3977 2929
rect -3943 1553 -3931 2929
rect -3989 1541 -3931 1553
rect -3791 2929 -3733 2941
rect -3791 1553 -3779 2929
rect -3745 1553 -3733 2929
rect -3791 1541 -3733 1553
rect -3593 2929 -3535 2941
rect -3593 1553 -3581 2929
rect -3547 1553 -3535 2929
rect -3593 1541 -3535 1553
rect -3395 2929 -3337 2941
rect -3395 1553 -3383 2929
rect -3349 1553 -3337 2929
rect -3395 1541 -3337 1553
rect -3197 2929 -3139 2941
rect -3197 1553 -3185 2929
rect -3151 1553 -3139 2929
rect -3197 1541 -3139 1553
rect -2999 2929 -2941 2941
rect -2999 1553 -2987 2929
rect -2953 1553 -2941 2929
rect -2999 1541 -2941 1553
rect -2801 2929 -2743 2941
rect -2801 1553 -2789 2929
rect -2755 1553 -2743 2929
rect -2801 1541 -2743 1553
rect -2603 2929 -2545 2941
rect -2603 1553 -2591 2929
rect -2557 1553 -2545 2929
rect -2603 1541 -2545 1553
rect -2405 2929 -2347 2941
rect -2405 1553 -2393 2929
rect -2359 1553 -2347 2929
rect -2405 1541 -2347 1553
rect -2207 2929 -2149 2941
rect -2207 1553 -2195 2929
rect -2161 1553 -2149 2929
rect -2207 1541 -2149 1553
rect -2009 2929 -1951 2941
rect -2009 1553 -1997 2929
rect -1963 1553 -1951 2929
rect -2009 1541 -1951 1553
rect -1811 2929 -1753 2941
rect -1811 1553 -1799 2929
rect -1765 1553 -1753 2929
rect -1811 1541 -1753 1553
rect -1613 2929 -1555 2941
rect -1613 1553 -1601 2929
rect -1567 1553 -1555 2929
rect -1613 1541 -1555 1553
rect -1415 2929 -1357 2941
rect -1415 1553 -1403 2929
rect -1369 1553 -1357 2929
rect -1415 1541 -1357 1553
rect -1217 2929 -1159 2941
rect -1217 1553 -1205 2929
rect -1171 1553 -1159 2929
rect -1217 1541 -1159 1553
rect -1019 2929 -961 2941
rect -1019 1553 -1007 2929
rect -973 1553 -961 2929
rect -1019 1541 -961 1553
rect -821 2929 -763 2941
rect -821 1553 -809 2929
rect -775 1553 -763 2929
rect -821 1541 -763 1553
rect -623 2929 -565 2941
rect -623 1553 -611 2929
rect -577 1553 -565 2929
rect -623 1541 -565 1553
rect -425 2929 -367 2941
rect -425 1553 -413 2929
rect -379 1553 -367 2929
rect -425 1541 -367 1553
rect -227 2929 -169 2941
rect -227 1553 -215 2929
rect -181 1553 -169 2929
rect -227 1541 -169 1553
rect -29 2929 29 2941
rect -29 1553 -17 2929
rect 17 1553 29 2929
rect -29 1541 29 1553
rect 169 2929 227 2941
rect 169 1553 181 2929
rect 215 1553 227 2929
rect 169 1541 227 1553
rect 367 2929 425 2941
rect 367 1553 379 2929
rect 413 1553 425 2929
rect 367 1541 425 1553
rect 565 2929 623 2941
rect 565 1553 577 2929
rect 611 1553 623 2929
rect 565 1541 623 1553
rect 763 2929 821 2941
rect 763 1553 775 2929
rect 809 1553 821 2929
rect 763 1541 821 1553
rect 961 2929 1019 2941
rect 961 1553 973 2929
rect 1007 1553 1019 2929
rect 961 1541 1019 1553
rect 1159 2929 1217 2941
rect 1159 1553 1171 2929
rect 1205 1553 1217 2929
rect 1159 1541 1217 1553
rect 1357 2929 1415 2941
rect 1357 1553 1369 2929
rect 1403 1553 1415 2929
rect 1357 1541 1415 1553
rect 1555 2929 1613 2941
rect 1555 1553 1567 2929
rect 1601 1553 1613 2929
rect 1555 1541 1613 1553
rect 1753 2929 1811 2941
rect 1753 1553 1765 2929
rect 1799 1553 1811 2929
rect 1753 1541 1811 1553
rect 1951 2929 2009 2941
rect 1951 1553 1963 2929
rect 1997 1553 2009 2929
rect 1951 1541 2009 1553
rect 2149 2929 2207 2941
rect 2149 1553 2161 2929
rect 2195 1553 2207 2929
rect 2149 1541 2207 1553
rect 2347 2929 2405 2941
rect 2347 1553 2359 2929
rect 2393 1553 2405 2929
rect 2347 1541 2405 1553
rect 2545 2929 2603 2941
rect 2545 1553 2557 2929
rect 2591 1553 2603 2929
rect 2545 1541 2603 1553
rect 2743 2929 2801 2941
rect 2743 1553 2755 2929
rect 2789 1553 2801 2929
rect 2743 1541 2801 1553
rect 2941 2929 2999 2941
rect 2941 1553 2953 2929
rect 2987 1553 2999 2929
rect 2941 1541 2999 1553
rect 3139 2929 3197 2941
rect 3139 1553 3151 2929
rect 3185 1553 3197 2929
rect 3139 1541 3197 1553
rect 3337 2929 3395 2941
rect 3337 1553 3349 2929
rect 3383 1553 3395 2929
rect 3337 1541 3395 1553
rect 3535 2929 3593 2941
rect 3535 1553 3547 2929
rect 3581 1553 3593 2929
rect 3535 1541 3593 1553
rect 3733 2929 3791 2941
rect 3733 1553 3745 2929
rect 3779 1553 3791 2929
rect 3733 1541 3791 1553
rect 3931 2929 3989 2941
rect 3931 1553 3943 2929
rect 3977 1553 3989 2929
rect 3931 1541 3989 1553
rect 4129 2929 4187 2941
rect 4129 1553 4141 2929
rect 4175 1553 4187 2929
rect 4129 1541 4187 1553
rect -4187 1435 -4129 1447
rect -4187 59 -4175 1435
rect -4141 59 -4129 1435
rect -4187 47 -4129 59
rect -3989 1435 -3931 1447
rect -3989 59 -3977 1435
rect -3943 59 -3931 1435
rect -3989 47 -3931 59
rect -3791 1435 -3733 1447
rect -3791 59 -3779 1435
rect -3745 59 -3733 1435
rect -3791 47 -3733 59
rect -3593 1435 -3535 1447
rect -3593 59 -3581 1435
rect -3547 59 -3535 1435
rect -3593 47 -3535 59
rect -3395 1435 -3337 1447
rect -3395 59 -3383 1435
rect -3349 59 -3337 1435
rect -3395 47 -3337 59
rect -3197 1435 -3139 1447
rect -3197 59 -3185 1435
rect -3151 59 -3139 1435
rect -3197 47 -3139 59
rect -2999 1435 -2941 1447
rect -2999 59 -2987 1435
rect -2953 59 -2941 1435
rect -2999 47 -2941 59
rect -2801 1435 -2743 1447
rect -2801 59 -2789 1435
rect -2755 59 -2743 1435
rect -2801 47 -2743 59
rect -2603 1435 -2545 1447
rect -2603 59 -2591 1435
rect -2557 59 -2545 1435
rect -2603 47 -2545 59
rect -2405 1435 -2347 1447
rect -2405 59 -2393 1435
rect -2359 59 -2347 1435
rect -2405 47 -2347 59
rect -2207 1435 -2149 1447
rect -2207 59 -2195 1435
rect -2161 59 -2149 1435
rect -2207 47 -2149 59
rect -2009 1435 -1951 1447
rect -2009 59 -1997 1435
rect -1963 59 -1951 1435
rect -2009 47 -1951 59
rect -1811 1435 -1753 1447
rect -1811 59 -1799 1435
rect -1765 59 -1753 1435
rect -1811 47 -1753 59
rect -1613 1435 -1555 1447
rect -1613 59 -1601 1435
rect -1567 59 -1555 1435
rect -1613 47 -1555 59
rect -1415 1435 -1357 1447
rect -1415 59 -1403 1435
rect -1369 59 -1357 1435
rect -1415 47 -1357 59
rect -1217 1435 -1159 1447
rect -1217 59 -1205 1435
rect -1171 59 -1159 1435
rect -1217 47 -1159 59
rect -1019 1435 -961 1447
rect -1019 59 -1007 1435
rect -973 59 -961 1435
rect -1019 47 -961 59
rect -821 1435 -763 1447
rect -821 59 -809 1435
rect -775 59 -763 1435
rect -821 47 -763 59
rect -623 1435 -565 1447
rect -623 59 -611 1435
rect -577 59 -565 1435
rect -623 47 -565 59
rect -425 1435 -367 1447
rect -425 59 -413 1435
rect -379 59 -367 1435
rect -425 47 -367 59
rect -227 1435 -169 1447
rect -227 59 -215 1435
rect -181 59 -169 1435
rect -227 47 -169 59
rect -29 1435 29 1447
rect -29 59 -17 1435
rect 17 59 29 1435
rect -29 47 29 59
rect 169 1435 227 1447
rect 169 59 181 1435
rect 215 59 227 1435
rect 169 47 227 59
rect 367 1435 425 1447
rect 367 59 379 1435
rect 413 59 425 1435
rect 367 47 425 59
rect 565 1435 623 1447
rect 565 59 577 1435
rect 611 59 623 1435
rect 565 47 623 59
rect 763 1435 821 1447
rect 763 59 775 1435
rect 809 59 821 1435
rect 763 47 821 59
rect 961 1435 1019 1447
rect 961 59 973 1435
rect 1007 59 1019 1435
rect 961 47 1019 59
rect 1159 1435 1217 1447
rect 1159 59 1171 1435
rect 1205 59 1217 1435
rect 1159 47 1217 59
rect 1357 1435 1415 1447
rect 1357 59 1369 1435
rect 1403 59 1415 1435
rect 1357 47 1415 59
rect 1555 1435 1613 1447
rect 1555 59 1567 1435
rect 1601 59 1613 1435
rect 1555 47 1613 59
rect 1753 1435 1811 1447
rect 1753 59 1765 1435
rect 1799 59 1811 1435
rect 1753 47 1811 59
rect 1951 1435 2009 1447
rect 1951 59 1963 1435
rect 1997 59 2009 1435
rect 1951 47 2009 59
rect 2149 1435 2207 1447
rect 2149 59 2161 1435
rect 2195 59 2207 1435
rect 2149 47 2207 59
rect 2347 1435 2405 1447
rect 2347 59 2359 1435
rect 2393 59 2405 1435
rect 2347 47 2405 59
rect 2545 1435 2603 1447
rect 2545 59 2557 1435
rect 2591 59 2603 1435
rect 2545 47 2603 59
rect 2743 1435 2801 1447
rect 2743 59 2755 1435
rect 2789 59 2801 1435
rect 2743 47 2801 59
rect 2941 1435 2999 1447
rect 2941 59 2953 1435
rect 2987 59 2999 1435
rect 2941 47 2999 59
rect 3139 1435 3197 1447
rect 3139 59 3151 1435
rect 3185 59 3197 1435
rect 3139 47 3197 59
rect 3337 1435 3395 1447
rect 3337 59 3349 1435
rect 3383 59 3395 1435
rect 3337 47 3395 59
rect 3535 1435 3593 1447
rect 3535 59 3547 1435
rect 3581 59 3593 1435
rect 3535 47 3593 59
rect 3733 1435 3791 1447
rect 3733 59 3745 1435
rect 3779 59 3791 1435
rect 3733 47 3791 59
rect 3931 1435 3989 1447
rect 3931 59 3943 1435
rect 3977 59 3989 1435
rect 3931 47 3989 59
rect 4129 1435 4187 1447
rect 4129 59 4141 1435
rect 4175 59 4187 1435
rect 4129 47 4187 59
rect -4187 -59 -4129 -47
rect -4187 -1435 -4175 -59
rect -4141 -1435 -4129 -59
rect -4187 -1447 -4129 -1435
rect -3989 -59 -3931 -47
rect -3989 -1435 -3977 -59
rect -3943 -1435 -3931 -59
rect -3989 -1447 -3931 -1435
rect -3791 -59 -3733 -47
rect -3791 -1435 -3779 -59
rect -3745 -1435 -3733 -59
rect -3791 -1447 -3733 -1435
rect -3593 -59 -3535 -47
rect -3593 -1435 -3581 -59
rect -3547 -1435 -3535 -59
rect -3593 -1447 -3535 -1435
rect -3395 -59 -3337 -47
rect -3395 -1435 -3383 -59
rect -3349 -1435 -3337 -59
rect -3395 -1447 -3337 -1435
rect -3197 -59 -3139 -47
rect -3197 -1435 -3185 -59
rect -3151 -1435 -3139 -59
rect -3197 -1447 -3139 -1435
rect -2999 -59 -2941 -47
rect -2999 -1435 -2987 -59
rect -2953 -1435 -2941 -59
rect -2999 -1447 -2941 -1435
rect -2801 -59 -2743 -47
rect -2801 -1435 -2789 -59
rect -2755 -1435 -2743 -59
rect -2801 -1447 -2743 -1435
rect -2603 -59 -2545 -47
rect -2603 -1435 -2591 -59
rect -2557 -1435 -2545 -59
rect -2603 -1447 -2545 -1435
rect -2405 -59 -2347 -47
rect -2405 -1435 -2393 -59
rect -2359 -1435 -2347 -59
rect -2405 -1447 -2347 -1435
rect -2207 -59 -2149 -47
rect -2207 -1435 -2195 -59
rect -2161 -1435 -2149 -59
rect -2207 -1447 -2149 -1435
rect -2009 -59 -1951 -47
rect -2009 -1435 -1997 -59
rect -1963 -1435 -1951 -59
rect -2009 -1447 -1951 -1435
rect -1811 -59 -1753 -47
rect -1811 -1435 -1799 -59
rect -1765 -1435 -1753 -59
rect -1811 -1447 -1753 -1435
rect -1613 -59 -1555 -47
rect -1613 -1435 -1601 -59
rect -1567 -1435 -1555 -59
rect -1613 -1447 -1555 -1435
rect -1415 -59 -1357 -47
rect -1415 -1435 -1403 -59
rect -1369 -1435 -1357 -59
rect -1415 -1447 -1357 -1435
rect -1217 -59 -1159 -47
rect -1217 -1435 -1205 -59
rect -1171 -1435 -1159 -59
rect -1217 -1447 -1159 -1435
rect -1019 -59 -961 -47
rect -1019 -1435 -1007 -59
rect -973 -1435 -961 -59
rect -1019 -1447 -961 -1435
rect -821 -59 -763 -47
rect -821 -1435 -809 -59
rect -775 -1435 -763 -59
rect -821 -1447 -763 -1435
rect -623 -59 -565 -47
rect -623 -1435 -611 -59
rect -577 -1435 -565 -59
rect -623 -1447 -565 -1435
rect -425 -59 -367 -47
rect -425 -1435 -413 -59
rect -379 -1435 -367 -59
rect -425 -1447 -367 -1435
rect -227 -59 -169 -47
rect -227 -1435 -215 -59
rect -181 -1435 -169 -59
rect -227 -1447 -169 -1435
rect -29 -59 29 -47
rect -29 -1435 -17 -59
rect 17 -1435 29 -59
rect -29 -1447 29 -1435
rect 169 -59 227 -47
rect 169 -1435 181 -59
rect 215 -1435 227 -59
rect 169 -1447 227 -1435
rect 367 -59 425 -47
rect 367 -1435 379 -59
rect 413 -1435 425 -59
rect 367 -1447 425 -1435
rect 565 -59 623 -47
rect 565 -1435 577 -59
rect 611 -1435 623 -59
rect 565 -1447 623 -1435
rect 763 -59 821 -47
rect 763 -1435 775 -59
rect 809 -1435 821 -59
rect 763 -1447 821 -1435
rect 961 -59 1019 -47
rect 961 -1435 973 -59
rect 1007 -1435 1019 -59
rect 961 -1447 1019 -1435
rect 1159 -59 1217 -47
rect 1159 -1435 1171 -59
rect 1205 -1435 1217 -59
rect 1159 -1447 1217 -1435
rect 1357 -59 1415 -47
rect 1357 -1435 1369 -59
rect 1403 -1435 1415 -59
rect 1357 -1447 1415 -1435
rect 1555 -59 1613 -47
rect 1555 -1435 1567 -59
rect 1601 -1435 1613 -59
rect 1555 -1447 1613 -1435
rect 1753 -59 1811 -47
rect 1753 -1435 1765 -59
rect 1799 -1435 1811 -59
rect 1753 -1447 1811 -1435
rect 1951 -59 2009 -47
rect 1951 -1435 1963 -59
rect 1997 -1435 2009 -59
rect 1951 -1447 2009 -1435
rect 2149 -59 2207 -47
rect 2149 -1435 2161 -59
rect 2195 -1435 2207 -59
rect 2149 -1447 2207 -1435
rect 2347 -59 2405 -47
rect 2347 -1435 2359 -59
rect 2393 -1435 2405 -59
rect 2347 -1447 2405 -1435
rect 2545 -59 2603 -47
rect 2545 -1435 2557 -59
rect 2591 -1435 2603 -59
rect 2545 -1447 2603 -1435
rect 2743 -59 2801 -47
rect 2743 -1435 2755 -59
rect 2789 -1435 2801 -59
rect 2743 -1447 2801 -1435
rect 2941 -59 2999 -47
rect 2941 -1435 2953 -59
rect 2987 -1435 2999 -59
rect 2941 -1447 2999 -1435
rect 3139 -59 3197 -47
rect 3139 -1435 3151 -59
rect 3185 -1435 3197 -59
rect 3139 -1447 3197 -1435
rect 3337 -59 3395 -47
rect 3337 -1435 3349 -59
rect 3383 -1435 3395 -59
rect 3337 -1447 3395 -1435
rect 3535 -59 3593 -47
rect 3535 -1435 3547 -59
rect 3581 -1435 3593 -59
rect 3535 -1447 3593 -1435
rect 3733 -59 3791 -47
rect 3733 -1435 3745 -59
rect 3779 -1435 3791 -59
rect 3733 -1447 3791 -1435
rect 3931 -59 3989 -47
rect 3931 -1435 3943 -59
rect 3977 -1435 3989 -59
rect 3931 -1447 3989 -1435
rect 4129 -59 4187 -47
rect 4129 -1435 4141 -59
rect 4175 -1435 4187 -59
rect 4129 -1447 4187 -1435
rect -4187 -1553 -4129 -1541
rect -4187 -2929 -4175 -1553
rect -4141 -2929 -4129 -1553
rect -4187 -2941 -4129 -2929
rect -3989 -1553 -3931 -1541
rect -3989 -2929 -3977 -1553
rect -3943 -2929 -3931 -1553
rect -3989 -2941 -3931 -2929
rect -3791 -1553 -3733 -1541
rect -3791 -2929 -3779 -1553
rect -3745 -2929 -3733 -1553
rect -3791 -2941 -3733 -2929
rect -3593 -1553 -3535 -1541
rect -3593 -2929 -3581 -1553
rect -3547 -2929 -3535 -1553
rect -3593 -2941 -3535 -2929
rect -3395 -1553 -3337 -1541
rect -3395 -2929 -3383 -1553
rect -3349 -2929 -3337 -1553
rect -3395 -2941 -3337 -2929
rect -3197 -1553 -3139 -1541
rect -3197 -2929 -3185 -1553
rect -3151 -2929 -3139 -1553
rect -3197 -2941 -3139 -2929
rect -2999 -1553 -2941 -1541
rect -2999 -2929 -2987 -1553
rect -2953 -2929 -2941 -1553
rect -2999 -2941 -2941 -2929
rect -2801 -1553 -2743 -1541
rect -2801 -2929 -2789 -1553
rect -2755 -2929 -2743 -1553
rect -2801 -2941 -2743 -2929
rect -2603 -1553 -2545 -1541
rect -2603 -2929 -2591 -1553
rect -2557 -2929 -2545 -1553
rect -2603 -2941 -2545 -2929
rect -2405 -1553 -2347 -1541
rect -2405 -2929 -2393 -1553
rect -2359 -2929 -2347 -1553
rect -2405 -2941 -2347 -2929
rect -2207 -1553 -2149 -1541
rect -2207 -2929 -2195 -1553
rect -2161 -2929 -2149 -1553
rect -2207 -2941 -2149 -2929
rect -2009 -1553 -1951 -1541
rect -2009 -2929 -1997 -1553
rect -1963 -2929 -1951 -1553
rect -2009 -2941 -1951 -2929
rect -1811 -1553 -1753 -1541
rect -1811 -2929 -1799 -1553
rect -1765 -2929 -1753 -1553
rect -1811 -2941 -1753 -2929
rect -1613 -1553 -1555 -1541
rect -1613 -2929 -1601 -1553
rect -1567 -2929 -1555 -1553
rect -1613 -2941 -1555 -2929
rect -1415 -1553 -1357 -1541
rect -1415 -2929 -1403 -1553
rect -1369 -2929 -1357 -1553
rect -1415 -2941 -1357 -2929
rect -1217 -1553 -1159 -1541
rect -1217 -2929 -1205 -1553
rect -1171 -2929 -1159 -1553
rect -1217 -2941 -1159 -2929
rect -1019 -1553 -961 -1541
rect -1019 -2929 -1007 -1553
rect -973 -2929 -961 -1553
rect -1019 -2941 -961 -2929
rect -821 -1553 -763 -1541
rect -821 -2929 -809 -1553
rect -775 -2929 -763 -1553
rect -821 -2941 -763 -2929
rect -623 -1553 -565 -1541
rect -623 -2929 -611 -1553
rect -577 -2929 -565 -1553
rect -623 -2941 -565 -2929
rect -425 -1553 -367 -1541
rect -425 -2929 -413 -1553
rect -379 -2929 -367 -1553
rect -425 -2941 -367 -2929
rect -227 -1553 -169 -1541
rect -227 -2929 -215 -1553
rect -181 -2929 -169 -1553
rect -227 -2941 -169 -2929
rect -29 -1553 29 -1541
rect -29 -2929 -17 -1553
rect 17 -2929 29 -1553
rect -29 -2941 29 -2929
rect 169 -1553 227 -1541
rect 169 -2929 181 -1553
rect 215 -2929 227 -1553
rect 169 -2941 227 -2929
rect 367 -1553 425 -1541
rect 367 -2929 379 -1553
rect 413 -2929 425 -1553
rect 367 -2941 425 -2929
rect 565 -1553 623 -1541
rect 565 -2929 577 -1553
rect 611 -2929 623 -1553
rect 565 -2941 623 -2929
rect 763 -1553 821 -1541
rect 763 -2929 775 -1553
rect 809 -2929 821 -1553
rect 763 -2941 821 -2929
rect 961 -1553 1019 -1541
rect 961 -2929 973 -1553
rect 1007 -2929 1019 -1553
rect 961 -2941 1019 -2929
rect 1159 -1553 1217 -1541
rect 1159 -2929 1171 -1553
rect 1205 -2929 1217 -1553
rect 1159 -2941 1217 -2929
rect 1357 -1553 1415 -1541
rect 1357 -2929 1369 -1553
rect 1403 -2929 1415 -1553
rect 1357 -2941 1415 -2929
rect 1555 -1553 1613 -1541
rect 1555 -2929 1567 -1553
rect 1601 -2929 1613 -1553
rect 1555 -2941 1613 -2929
rect 1753 -1553 1811 -1541
rect 1753 -2929 1765 -1553
rect 1799 -2929 1811 -1553
rect 1753 -2941 1811 -2929
rect 1951 -1553 2009 -1541
rect 1951 -2929 1963 -1553
rect 1997 -2929 2009 -1553
rect 1951 -2941 2009 -2929
rect 2149 -1553 2207 -1541
rect 2149 -2929 2161 -1553
rect 2195 -2929 2207 -1553
rect 2149 -2941 2207 -2929
rect 2347 -1553 2405 -1541
rect 2347 -2929 2359 -1553
rect 2393 -2929 2405 -1553
rect 2347 -2941 2405 -2929
rect 2545 -1553 2603 -1541
rect 2545 -2929 2557 -1553
rect 2591 -2929 2603 -1553
rect 2545 -2941 2603 -2929
rect 2743 -1553 2801 -1541
rect 2743 -2929 2755 -1553
rect 2789 -2929 2801 -1553
rect 2743 -2941 2801 -2929
rect 2941 -1553 2999 -1541
rect 2941 -2929 2953 -1553
rect 2987 -2929 2999 -1553
rect 2941 -2941 2999 -2929
rect 3139 -1553 3197 -1541
rect 3139 -2929 3151 -1553
rect 3185 -2929 3197 -1553
rect 3139 -2941 3197 -2929
rect 3337 -1553 3395 -1541
rect 3337 -2929 3349 -1553
rect 3383 -2929 3395 -1553
rect 3337 -2941 3395 -2929
rect 3535 -1553 3593 -1541
rect 3535 -2929 3547 -1553
rect 3581 -2929 3593 -1553
rect 3535 -2941 3593 -2929
rect 3733 -1553 3791 -1541
rect 3733 -2929 3745 -1553
rect 3779 -2929 3791 -1553
rect 3733 -2941 3791 -2929
rect 3931 -1553 3989 -1541
rect 3931 -2929 3943 -1553
rect 3977 -2929 3989 -1553
rect 3931 -2941 3989 -2929
rect 4129 -1553 4187 -1541
rect 4129 -2929 4141 -1553
rect 4175 -2929 4187 -1553
rect 4129 -2941 4187 -2929
<< pdiffc >>
rect -4175 1553 -4141 2929
rect -3977 1553 -3943 2929
rect -3779 1553 -3745 2929
rect -3581 1553 -3547 2929
rect -3383 1553 -3349 2929
rect -3185 1553 -3151 2929
rect -2987 1553 -2953 2929
rect -2789 1553 -2755 2929
rect -2591 1553 -2557 2929
rect -2393 1553 -2359 2929
rect -2195 1553 -2161 2929
rect -1997 1553 -1963 2929
rect -1799 1553 -1765 2929
rect -1601 1553 -1567 2929
rect -1403 1553 -1369 2929
rect -1205 1553 -1171 2929
rect -1007 1553 -973 2929
rect -809 1553 -775 2929
rect -611 1553 -577 2929
rect -413 1553 -379 2929
rect -215 1553 -181 2929
rect -17 1553 17 2929
rect 181 1553 215 2929
rect 379 1553 413 2929
rect 577 1553 611 2929
rect 775 1553 809 2929
rect 973 1553 1007 2929
rect 1171 1553 1205 2929
rect 1369 1553 1403 2929
rect 1567 1553 1601 2929
rect 1765 1553 1799 2929
rect 1963 1553 1997 2929
rect 2161 1553 2195 2929
rect 2359 1553 2393 2929
rect 2557 1553 2591 2929
rect 2755 1553 2789 2929
rect 2953 1553 2987 2929
rect 3151 1553 3185 2929
rect 3349 1553 3383 2929
rect 3547 1553 3581 2929
rect 3745 1553 3779 2929
rect 3943 1553 3977 2929
rect 4141 1553 4175 2929
rect -4175 59 -4141 1435
rect -3977 59 -3943 1435
rect -3779 59 -3745 1435
rect -3581 59 -3547 1435
rect -3383 59 -3349 1435
rect -3185 59 -3151 1435
rect -2987 59 -2953 1435
rect -2789 59 -2755 1435
rect -2591 59 -2557 1435
rect -2393 59 -2359 1435
rect -2195 59 -2161 1435
rect -1997 59 -1963 1435
rect -1799 59 -1765 1435
rect -1601 59 -1567 1435
rect -1403 59 -1369 1435
rect -1205 59 -1171 1435
rect -1007 59 -973 1435
rect -809 59 -775 1435
rect -611 59 -577 1435
rect -413 59 -379 1435
rect -215 59 -181 1435
rect -17 59 17 1435
rect 181 59 215 1435
rect 379 59 413 1435
rect 577 59 611 1435
rect 775 59 809 1435
rect 973 59 1007 1435
rect 1171 59 1205 1435
rect 1369 59 1403 1435
rect 1567 59 1601 1435
rect 1765 59 1799 1435
rect 1963 59 1997 1435
rect 2161 59 2195 1435
rect 2359 59 2393 1435
rect 2557 59 2591 1435
rect 2755 59 2789 1435
rect 2953 59 2987 1435
rect 3151 59 3185 1435
rect 3349 59 3383 1435
rect 3547 59 3581 1435
rect 3745 59 3779 1435
rect 3943 59 3977 1435
rect 4141 59 4175 1435
rect -4175 -1435 -4141 -59
rect -3977 -1435 -3943 -59
rect -3779 -1435 -3745 -59
rect -3581 -1435 -3547 -59
rect -3383 -1435 -3349 -59
rect -3185 -1435 -3151 -59
rect -2987 -1435 -2953 -59
rect -2789 -1435 -2755 -59
rect -2591 -1435 -2557 -59
rect -2393 -1435 -2359 -59
rect -2195 -1435 -2161 -59
rect -1997 -1435 -1963 -59
rect -1799 -1435 -1765 -59
rect -1601 -1435 -1567 -59
rect -1403 -1435 -1369 -59
rect -1205 -1435 -1171 -59
rect -1007 -1435 -973 -59
rect -809 -1435 -775 -59
rect -611 -1435 -577 -59
rect -413 -1435 -379 -59
rect -215 -1435 -181 -59
rect -17 -1435 17 -59
rect 181 -1435 215 -59
rect 379 -1435 413 -59
rect 577 -1435 611 -59
rect 775 -1435 809 -59
rect 973 -1435 1007 -59
rect 1171 -1435 1205 -59
rect 1369 -1435 1403 -59
rect 1567 -1435 1601 -59
rect 1765 -1435 1799 -59
rect 1963 -1435 1997 -59
rect 2161 -1435 2195 -59
rect 2359 -1435 2393 -59
rect 2557 -1435 2591 -59
rect 2755 -1435 2789 -59
rect 2953 -1435 2987 -59
rect 3151 -1435 3185 -59
rect 3349 -1435 3383 -59
rect 3547 -1435 3581 -59
rect 3745 -1435 3779 -59
rect 3943 -1435 3977 -59
rect 4141 -1435 4175 -59
rect -4175 -2929 -4141 -1553
rect -3977 -2929 -3943 -1553
rect -3779 -2929 -3745 -1553
rect -3581 -2929 -3547 -1553
rect -3383 -2929 -3349 -1553
rect -3185 -2929 -3151 -1553
rect -2987 -2929 -2953 -1553
rect -2789 -2929 -2755 -1553
rect -2591 -2929 -2557 -1553
rect -2393 -2929 -2359 -1553
rect -2195 -2929 -2161 -1553
rect -1997 -2929 -1963 -1553
rect -1799 -2929 -1765 -1553
rect -1601 -2929 -1567 -1553
rect -1403 -2929 -1369 -1553
rect -1205 -2929 -1171 -1553
rect -1007 -2929 -973 -1553
rect -809 -2929 -775 -1553
rect -611 -2929 -577 -1553
rect -413 -2929 -379 -1553
rect -215 -2929 -181 -1553
rect -17 -2929 17 -1553
rect 181 -2929 215 -1553
rect 379 -2929 413 -1553
rect 577 -2929 611 -1553
rect 775 -2929 809 -1553
rect 973 -2929 1007 -1553
rect 1171 -2929 1205 -1553
rect 1369 -2929 1403 -1553
rect 1567 -2929 1601 -1553
rect 1765 -2929 1799 -1553
rect 1963 -2929 1997 -1553
rect 2161 -2929 2195 -1553
rect 2359 -2929 2393 -1553
rect 2557 -2929 2591 -1553
rect 2755 -2929 2789 -1553
rect 2953 -2929 2987 -1553
rect 3151 -2929 3185 -1553
rect 3349 -2929 3383 -1553
rect 3547 -2929 3581 -1553
rect 3745 -2929 3779 -1553
rect 3943 -2929 3977 -1553
rect 4141 -2929 4175 -1553
<< poly >>
rect -4129 2941 -3989 2967
rect -3931 2941 -3791 2967
rect -3733 2941 -3593 2967
rect -3535 2941 -3395 2967
rect -3337 2941 -3197 2967
rect -3139 2941 -2999 2967
rect -2941 2941 -2801 2967
rect -2743 2941 -2603 2967
rect -2545 2941 -2405 2967
rect -2347 2941 -2207 2967
rect -2149 2941 -2009 2967
rect -1951 2941 -1811 2967
rect -1753 2941 -1613 2967
rect -1555 2941 -1415 2967
rect -1357 2941 -1217 2967
rect -1159 2941 -1019 2967
rect -961 2941 -821 2967
rect -763 2941 -623 2967
rect -565 2941 -425 2967
rect -367 2941 -227 2967
rect -169 2941 -29 2967
rect 29 2941 169 2967
rect 227 2941 367 2967
rect 425 2941 565 2967
rect 623 2941 763 2967
rect 821 2941 961 2967
rect 1019 2941 1159 2967
rect 1217 2941 1357 2967
rect 1415 2941 1555 2967
rect 1613 2941 1753 2967
rect 1811 2941 1951 2967
rect 2009 2941 2149 2967
rect 2207 2941 2347 2967
rect 2405 2941 2545 2967
rect 2603 2941 2743 2967
rect 2801 2941 2941 2967
rect 2999 2941 3139 2967
rect 3197 2941 3337 2967
rect 3395 2941 3535 2967
rect 3593 2941 3733 2967
rect 3791 2941 3931 2967
rect 3989 2941 4129 2967
rect -4129 1515 -3989 1541
rect -3931 1515 -3791 1541
rect -3733 1515 -3593 1541
rect -3535 1515 -3395 1541
rect -3337 1515 -3197 1541
rect -3139 1515 -2999 1541
rect -2941 1515 -2801 1541
rect -2743 1515 -2603 1541
rect -2545 1515 -2405 1541
rect -2347 1515 -2207 1541
rect -2149 1515 -2009 1541
rect -1951 1515 -1811 1541
rect -1753 1515 -1613 1541
rect -1555 1515 -1415 1541
rect -1357 1515 -1217 1541
rect -1159 1515 -1019 1541
rect -961 1515 -821 1541
rect -763 1515 -623 1541
rect -565 1515 -425 1541
rect -367 1515 -227 1541
rect -169 1515 -29 1541
rect 29 1515 169 1541
rect 227 1515 367 1541
rect 425 1515 565 1541
rect 623 1515 763 1541
rect 821 1515 961 1541
rect 1019 1515 1159 1541
rect 1217 1515 1357 1541
rect 1415 1515 1555 1541
rect 1613 1515 1753 1541
rect 1811 1515 1951 1541
rect 2009 1515 2149 1541
rect 2207 1515 2347 1541
rect 2405 1515 2545 1541
rect 2603 1515 2743 1541
rect 2801 1515 2941 1541
rect 2999 1515 3139 1541
rect 3197 1515 3337 1541
rect 3395 1515 3535 1541
rect 3593 1515 3733 1541
rect 3791 1515 3931 1541
rect 3989 1515 4129 1541
rect -4129 1447 -3989 1473
rect -3931 1447 -3791 1473
rect -3733 1447 -3593 1473
rect -3535 1447 -3395 1473
rect -3337 1447 -3197 1473
rect -3139 1447 -2999 1473
rect -2941 1447 -2801 1473
rect -2743 1447 -2603 1473
rect -2545 1447 -2405 1473
rect -2347 1447 -2207 1473
rect -2149 1447 -2009 1473
rect -1951 1447 -1811 1473
rect -1753 1447 -1613 1473
rect -1555 1447 -1415 1473
rect -1357 1447 -1217 1473
rect -1159 1447 -1019 1473
rect -961 1447 -821 1473
rect -763 1447 -623 1473
rect -565 1447 -425 1473
rect -367 1447 -227 1473
rect -169 1447 -29 1473
rect 29 1447 169 1473
rect 227 1447 367 1473
rect 425 1447 565 1473
rect 623 1447 763 1473
rect 821 1447 961 1473
rect 1019 1447 1159 1473
rect 1217 1447 1357 1473
rect 1415 1447 1555 1473
rect 1613 1447 1753 1473
rect 1811 1447 1951 1473
rect 2009 1447 2149 1473
rect 2207 1447 2347 1473
rect 2405 1447 2545 1473
rect 2603 1447 2743 1473
rect 2801 1447 2941 1473
rect 2999 1447 3139 1473
rect 3197 1447 3337 1473
rect 3395 1447 3535 1473
rect 3593 1447 3733 1473
rect 3791 1447 3931 1473
rect 3989 1447 4129 1473
rect -4129 21 -3989 47
rect -3931 21 -3791 47
rect -3733 21 -3593 47
rect -3535 21 -3395 47
rect -3337 21 -3197 47
rect -3139 21 -2999 47
rect -2941 21 -2801 47
rect -2743 21 -2603 47
rect -2545 21 -2405 47
rect -2347 21 -2207 47
rect -2149 21 -2009 47
rect -1951 21 -1811 47
rect -1753 21 -1613 47
rect -1555 21 -1415 47
rect -1357 21 -1217 47
rect -1159 21 -1019 47
rect -961 21 -821 47
rect -763 21 -623 47
rect -565 21 -425 47
rect -367 21 -227 47
rect -169 21 -29 47
rect 29 21 169 47
rect 227 21 367 47
rect 425 21 565 47
rect 623 21 763 47
rect 821 21 961 47
rect 1019 21 1159 47
rect 1217 21 1357 47
rect 1415 21 1555 47
rect 1613 21 1753 47
rect 1811 21 1951 47
rect 2009 21 2149 47
rect 2207 21 2347 47
rect 2405 21 2545 47
rect 2603 21 2743 47
rect 2801 21 2941 47
rect 2999 21 3139 47
rect 3197 21 3337 47
rect 3395 21 3535 47
rect 3593 21 3733 47
rect 3791 21 3931 47
rect 3989 21 4129 47
rect -4129 -47 -3989 -21
rect -3931 -47 -3791 -21
rect -3733 -47 -3593 -21
rect -3535 -47 -3395 -21
rect -3337 -47 -3197 -21
rect -3139 -47 -2999 -21
rect -2941 -47 -2801 -21
rect -2743 -47 -2603 -21
rect -2545 -47 -2405 -21
rect -2347 -47 -2207 -21
rect -2149 -47 -2009 -21
rect -1951 -47 -1811 -21
rect -1753 -47 -1613 -21
rect -1555 -47 -1415 -21
rect -1357 -47 -1217 -21
rect -1159 -47 -1019 -21
rect -961 -47 -821 -21
rect -763 -47 -623 -21
rect -565 -47 -425 -21
rect -367 -47 -227 -21
rect -169 -47 -29 -21
rect 29 -47 169 -21
rect 227 -47 367 -21
rect 425 -47 565 -21
rect 623 -47 763 -21
rect 821 -47 961 -21
rect 1019 -47 1159 -21
rect 1217 -47 1357 -21
rect 1415 -47 1555 -21
rect 1613 -47 1753 -21
rect 1811 -47 1951 -21
rect 2009 -47 2149 -21
rect 2207 -47 2347 -21
rect 2405 -47 2545 -21
rect 2603 -47 2743 -21
rect 2801 -47 2941 -21
rect 2999 -47 3139 -21
rect 3197 -47 3337 -21
rect 3395 -47 3535 -21
rect 3593 -47 3733 -21
rect 3791 -47 3931 -21
rect 3989 -47 4129 -21
rect -4129 -1473 -3989 -1447
rect -3931 -1473 -3791 -1447
rect -3733 -1473 -3593 -1447
rect -3535 -1473 -3395 -1447
rect -3337 -1473 -3197 -1447
rect -3139 -1473 -2999 -1447
rect -2941 -1473 -2801 -1447
rect -2743 -1473 -2603 -1447
rect -2545 -1473 -2405 -1447
rect -2347 -1473 -2207 -1447
rect -2149 -1473 -2009 -1447
rect -1951 -1473 -1811 -1447
rect -1753 -1473 -1613 -1447
rect -1555 -1473 -1415 -1447
rect -1357 -1473 -1217 -1447
rect -1159 -1473 -1019 -1447
rect -961 -1473 -821 -1447
rect -763 -1473 -623 -1447
rect -565 -1473 -425 -1447
rect -367 -1473 -227 -1447
rect -169 -1473 -29 -1447
rect 29 -1473 169 -1447
rect 227 -1473 367 -1447
rect 425 -1473 565 -1447
rect 623 -1473 763 -1447
rect 821 -1473 961 -1447
rect 1019 -1473 1159 -1447
rect 1217 -1473 1357 -1447
rect 1415 -1473 1555 -1447
rect 1613 -1473 1753 -1447
rect 1811 -1473 1951 -1447
rect 2009 -1473 2149 -1447
rect 2207 -1473 2347 -1447
rect 2405 -1473 2545 -1447
rect 2603 -1473 2743 -1447
rect 2801 -1473 2941 -1447
rect 2999 -1473 3139 -1447
rect 3197 -1473 3337 -1447
rect 3395 -1473 3535 -1447
rect 3593 -1473 3733 -1447
rect 3791 -1473 3931 -1447
rect 3989 -1473 4129 -1447
rect -4129 -1541 -3989 -1515
rect -3931 -1541 -3791 -1515
rect -3733 -1541 -3593 -1515
rect -3535 -1541 -3395 -1515
rect -3337 -1541 -3197 -1515
rect -3139 -1541 -2999 -1515
rect -2941 -1541 -2801 -1515
rect -2743 -1541 -2603 -1515
rect -2545 -1541 -2405 -1515
rect -2347 -1541 -2207 -1515
rect -2149 -1541 -2009 -1515
rect -1951 -1541 -1811 -1515
rect -1753 -1541 -1613 -1515
rect -1555 -1541 -1415 -1515
rect -1357 -1541 -1217 -1515
rect -1159 -1541 -1019 -1515
rect -961 -1541 -821 -1515
rect -763 -1541 -623 -1515
rect -565 -1541 -425 -1515
rect -367 -1541 -227 -1515
rect -169 -1541 -29 -1515
rect 29 -1541 169 -1515
rect 227 -1541 367 -1515
rect 425 -1541 565 -1515
rect 623 -1541 763 -1515
rect 821 -1541 961 -1515
rect 1019 -1541 1159 -1515
rect 1217 -1541 1357 -1515
rect 1415 -1541 1555 -1515
rect 1613 -1541 1753 -1515
rect 1811 -1541 1951 -1515
rect 2009 -1541 2149 -1515
rect 2207 -1541 2347 -1515
rect 2405 -1541 2545 -1515
rect 2603 -1541 2743 -1515
rect 2801 -1541 2941 -1515
rect 2999 -1541 3139 -1515
rect 3197 -1541 3337 -1515
rect 3395 -1541 3535 -1515
rect 3593 -1541 3733 -1515
rect 3791 -1541 3931 -1515
rect 3989 -1541 4129 -1515
rect -4129 -2967 -3989 -2941
rect -3931 -2967 -3791 -2941
rect -3733 -2967 -3593 -2941
rect -3535 -2967 -3395 -2941
rect -3337 -2967 -3197 -2941
rect -3139 -2967 -2999 -2941
rect -2941 -2967 -2801 -2941
rect -2743 -2967 -2603 -2941
rect -2545 -2967 -2405 -2941
rect -2347 -2967 -2207 -2941
rect -2149 -2967 -2009 -2941
rect -1951 -2967 -1811 -2941
rect -1753 -2967 -1613 -2941
rect -1555 -2967 -1415 -2941
rect -1357 -2967 -1217 -2941
rect -1159 -2967 -1019 -2941
rect -961 -2967 -821 -2941
rect -763 -2967 -623 -2941
rect -565 -2967 -425 -2941
rect -367 -2967 -227 -2941
rect -169 -2967 -29 -2941
rect 29 -2967 169 -2941
rect 227 -2967 367 -2941
rect 425 -2967 565 -2941
rect 623 -2967 763 -2941
rect 821 -2967 961 -2941
rect 1019 -2967 1159 -2941
rect 1217 -2967 1357 -2941
rect 1415 -2967 1555 -2941
rect 1613 -2967 1753 -2941
rect 1811 -2967 1951 -2941
rect 2009 -2967 2149 -2941
rect 2207 -2967 2347 -2941
rect 2405 -2967 2545 -2941
rect 2603 -2967 2743 -2941
rect 2801 -2967 2941 -2941
rect 2999 -2967 3139 -2941
rect 3197 -2967 3337 -2941
rect 3395 -2967 3535 -2941
rect 3593 -2967 3733 -2941
rect 3791 -2967 3931 -2941
rect 3989 -2967 4129 -2941
<< locali >>
rect -4175 2929 -4141 2945
rect -4175 1537 -4141 1553
rect -3977 2929 -3943 2945
rect -3977 1537 -3943 1553
rect -3779 2929 -3745 2945
rect -3779 1537 -3745 1553
rect -3581 2929 -3547 2945
rect -3581 1537 -3547 1553
rect -3383 2929 -3349 2945
rect -3383 1537 -3349 1553
rect -3185 2929 -3151 2945
rect -3185 1537 -3151 1553
rect -2987 2929 -2953 2945
rect -2987 1537 -2953 1553
rect -2789 2929 -2755 2945
rect -2789 1537 -2755 1553
rect -2591 2929 -2557 2945
rect -2591 1537 -2557 1553
rect -2393 2929 -2359 2945
rect -2393 1537 -2359 1553
rect -2195 2929 -2161 2945
rect -2195 1537 -2161 1553
rect -1997 2929 -1963 2945
rect -1997 1537 -1963 1553
rect -1799 2929 -1765 2945
rect -1799 1537 -1765 1553
rect -1601 2929 -1567 2945
rect -1601 1537 -1567 1553
rect -1403 2929 -1369 2945
rect -1403 1537 -1369 1553
rect -1205 2929 -1171 2945
rect -1205 1537 -1171 1553
rect -1007 2929 -973 2945
rect -1007 1537 -973 1553
rect -809 2929 -775 2945
rect -809 1537 -775 1553
rect -611 2929 -577 2945
rect -611 1537 -577 1553
rect -413 2929 -379 2945
rect -413 1537 -379 1553
rect -215 2929 -181 2945
rect -215 1537 -181 1553
rect -17 2929 17 2945
rect -17 1537 17 1553
rect 181 2929 215 2945
rect 181 1537 215 1553
rect 379 2929 413 2945
rect 379 1537 413 1553
rect 577 2929 611 2945
rect 577 1537 611 1553
rect 775 2929 809 2945
rect 775 1537 809 1553
rect 973 2929 1007 2945
rect 973 1537 1007 1553
rect 1171 2929 1205 2945
rect 1171 1537 1205 1553
rect 1369 2929 1403 2945
rect 1369 1537 1403 1553
rect 1567 2929 1601 2945
rect 1567 1537 1601 1553
rect 1765 2929 1799 2945
rect 1765 1537 1799 1553
rect 1963 2929 1997 2945
rect 1963 1537 1997 1553
rect 2161 2929 2195 2945
rect 2161 1537 2195 1553
rect 2359 2929 2393 2945
rect 2359 1537 2393 1553
rect 2557 2929 2591 2945
rect 2557 1537 2591 1553
rect 2755 2929 2789 2945
rect 2755 1537 2789 1553
rect 2953 2929 2987 2945
rect 2953 1537 2987 1553
rect 3151 2929 3185 2945
rect 3151 1537 3185 1553
rect 3349 2929 3383 2945
rect 3349 1537 3383 1553
rect 3547 2929 3581 2945
rect 3547 1537 3581 1553
rect 3745 2929 3779 2945
rect 3745 1537 3779 1553
rect 3943 2929 3977 2945
rect 3943 1537 3977 1553
rect 4141 2929 4175 2945
rect 4141 1537 4175 1553
rect -4175 1435 -4141 1451
rect -4175 43 -4141 59
rect -3977 1435 -3943 1451
rect -3977 43 -3943 59
rect -3779 1435 -3745 1451
rect -3779 43 -3745 59
rect -3581 1435 -3547 1451
rect -3581 43 -3547 59
rect -3383 1435 -3349 1451
rect -3383 43 -3349 59
rect -3185 1435 -3151 1451
rect -3185 43 -3151 59
rect -2987 1435 -2953 1451
rect -2987 43 -2953 59
rect -2789 1435 -2755 1451
rect -2789 43 -2755 59
rect -2591 1435 -2557 1451
rect -2591 43 -2557 59
rect -2393 1435 -2359 1451
rect -2393 43 -2359 59
rect -2195 1435 -2161 1451
rect -2195 43 -2161 59
rect -1997 1435 -1963 1451
rect -1997 43 -1963 59
rect -1799 1435 -1765 1451
rect -1799 43 -1765 59
rect -1601 1435 -1567 1451
rect -1601 43 -1567 59
rect -1403 1435 -1369 1451
rect -1403 43 -1369 59
rect -1205 1435 -1171 1451
rect -1205 43 -1171 59
rect -1007 1435 -973 1451
rect -1007 43 -973 59
rect -809 1435 -775 1451
rect -809 43 -775 59
rect -611 1435 -577 1451
rect -611 43 -577 59
rect -413 1435 -379 1451
rect -413 43 -379 59
rect -215 1435 -181 1451
rect -215 43 -181 59
rect -17 1435 17 1451
rect -17 43 17 59
rect 181 1435 215 1451
rect 181 43 215 59
rect 379 1435 413 1451
rect 379 43 413 59
rect 577 1435 611 1451
rect 577 43 611 59
rect 775 1435 809 1451
rect 775 43 809 59
rect 973 1435 1007 1451
rect 973 43 1007 59
rect 1171 1435 1205 1451
rect 1171 43 1205 59
rect 1369 1435 1403 1451
rect 1369 43 1403 59
rect 1567 1435 1601 1451
rect 1567 43 1601 59
rect 1765 1435 1799 1451
rect 1765 43 1799 59
rect 1963 1435 1997 1451
rect 1963 43 1997 59
rect 2161 1435 2195 1451
rect 2161 43 2195 59
rect 2359 1435 2393 1451
rect 2359 43 2393 59
rect 2557 1435 2591 1451
rect 2557 43 2591 59
rect 2755 1435 2789 1451
rect 2755 43 2789 59
rect 2953 1435 2987 1451
rect 2953 43 2987 59
rect 3151 1435 3185 1451
rect 3151 43 3185 59
rect 3349 1435 3383 1451
rect 3349 43 3383 59
rect 3547 1435 3581 1451
rect 3547 43 3581 59
rect 3745 1435 3779 1451
rect 3745 43 3779 59
rect 3943 1435 3977 1451
rect 3943 43 3977 59
rect 4141 1435 4175 1451
rect 4141 43 4175 59
rect -4175 -59 -4141 -43
rect -4175 -1451 -4141 -1435
rect -3977 -59 -3943 -43
rect -3977 -1451 -3943 -1435
rect -3779 -59 -3745 -43
rect -3779 -1451 -3745 -1435
rect -3581 -59 -3547 -43
rect -3581 -1451 -3547 -1435
rect -3383 -59 -3349 -43
rect -3383 -1451 -3349 -1435
rect -3185 -59 -3151 -43
rect -3185 -1451 -3151 -1435
rect -2987 -59 -2953 -43
rect -2987 -1451 -2953 -1435
rect -2789 -59 -2755 -43
rect -2789 -1451 -2755 -1435
rect -2591 -59 -2557 -43
rect -2591 -1451 -2557 -1435
rect -2393 -59 -2359 -43
rect -2393 -1451 -2359 -1435
rect -2195 -59 -2161 -43
rect -2195 -1451 -2161 -1435
rect -1997 -59 -1963 -43
rect -1997 -1451 -1963 -1435
rect -1799 -59 -1765 -43
rect -1799 -1451 -1765 -1435
rect -1601 -59 -1567 -43
rect -1601 -1451 -1567 -1435
rect -1403 -59 -1369 -43
rect -1403 -1451 -1369 -1435
rect -1205 -59 -1171 -43
rect -1205 -1451 -1171 -1435
rect -1007 -59 -973 -43
rect -1007 -1451 -973 -1435
rect -809 -59 -775 -43
rect -809 -1451 -775 -1435
rect -611 -59 -577 -43
rect -611 -1451 -577 -1435
rect -413 -59 -379 -43
rect -413 -1451 -379 -1435
rect -215 -59 -181 -43
rect -215 -1451 -181 -1435
rect -17 -59 17 -43
rect -17 -1451 17 -1435
rect 181 -59 215 -43
rect 181 -1451 215 -1435
rect 379 -59 413 -43
rect 379 -1451 413 -1435
rect 577 -59 611 -43
rect 577 -1451 611 -1435
rect 775 -59 809 -43
rect 775 -1451 809 -1435
rect 973 -59 1007 -43
rect 973 -1451 1007 -1435
rect 1171 -59 1205 -43
rect 1171 -1451 1205 -1435
rect 1369 -59 1403 -43
rect 1369 -1451 1403 -1435
rect 1567 -59 1601 -43
rect 1567 -1451 1601 -1435
rect 1765 -59 1799 -43
rect 1765 -1451 1799 -1435
rect 1963 -59 1997 -43
rect 1963 -1451 1997 -1435
rect 2161 -59 2195 -43
rect 2161 -1451 2195 -1435
rect 2359 -59 2393 -43
rect 2359 -1451 2393 -1435
rect 2557 -59 2591 -43
rect 2557 -1451 2591 -1435
rect 2755 -59 2789 -43
rect 2755 -1451 2789 -1435
rect 2953 -59 2987 -43
rect 2953 -1451 2987 -1435
rect 3151 -59 3185 -43
rect 3151 -1451 3185 -1435
rect 3349 -59 3383 -43
rect 3349 -1451 3383 -1435
rect 3547 -59 3581 -43
rect 3547 -1451 3581 -1435
rect 3745 -59 3779 -43
rect 3745 -1451 3779 -1435
rect 3943 -59 3977 -43
rect 3943 -1451 3977 -1435
rect 4141 -59 4175 -43
rect 4141 -1451 4175 -1435
rect -4175 -1553 -4141 -1537
rect -4175 -2945 -4141 -2929
rect -3977 -1553 -3943 -1537
rect -3977 -2945 -3943 -2929
rect -3779 -1553 -3745 -1537
rect -3779 -2945 -3745 -2929
rect -3581 -1553 -3547 -1537
rect -3581 -2945 -3547 -2929
rect -3383 -1553 -3349 -1537
rect -3383 -2945 -3349 -2929
rect -3185 -1553 -3151 -1537
rect -3185 -2945 -3151 -2929
rect -2987 -1553 -2953 -1537
rect -2987 -2945 -2953 -2929
rect -2789 -1553 -2755 -1537
rect -2789 -2945 -2755 -2929
rect -2591 -1553 -2557 -1537
rect -2591 -2945 -2557 -2929
rect -2393 -1553 -2359 -1537
rect -2393 -2945 -2359 -2929
rect -2195 -1553 -2161 -1537
rect -2195 -2945 -2161 -2929
rect -1997 -1553 -1963 -1537
rect -1997 -2945 -1963 -2929
rect -1799 -1553 -1765 -1537
rect -1799 -2945 -1765 -2929
rect -1601 -1553 -1567 -1537
rect -1601 -2945 -1567 -2929
rect -1403 -1553 -1369 -1537
rect -1403 -2945 -1369 -2929
rect -1205 -1553 -1171 -1537
rect -1205 -2945 -1171 -2929
rect -1007 -1553 -973 -1537
rect -1007 -2945 -973 -2929
rect -809 -1553 -775 -1537
rect -809 -2945 -775 -2929
rect -611 -1553 -577 -1537
rect -611 -2945 -577 -2929
rect -413 -1553 -379 -1537
rect -413 -2945 -379 -2929
rect -215 -1553 -181 -1537
rect -215 -2945 -181 -2929
rect -17 -1553 17 -1537
rect -17 -2945 17 -2929
rect 181 -1553 215 -1537
rect 181 -2945 215 -2929
rect 379 -1553 413 -1537
rect 379 -2945 413 -2929
rect 577 -1553 611 -1537
rect 577 -2945 611 -2929
rect 775 -1553 809 -1537
rect 775 -2945 809 -2929
rect 973 -1553 1007 -1537
rect 973 -2945 1007 -2929
rect 1171 -1553 1205 -1537
rect 1171 -2945 1205 -2929
rect 1369 -1553 1403 -1537
rect 1369 -2945 1403 -2929
rect 1567 -1553 1601 -1537
rect 1567 -2945 1601 -2929
rect 1765 -1553 1799 -1537
rect 1765 -2945 1799 -2929
rect 1963 -1553 1997 -1537
rect 1963 -2945 1997 -2929
rect 2161 -1553 2195 -1537
rect 2161 -2945 2195 -2929
rect 2359 -1553 2393 -1537
rect 2359 -2945 2393 -2929
rect 2557 -1553 2591 -1537
rect 2557 -2945 2591 -2929
rect 2755 -1553 2789 -1537
rect 2755 -2945 2789 -2929
rect 2953 -1553 2987 -1537
rect 2953 -2945 2987 -2929
rect 3151 -1553 3185 -1537
rect 3151 -2945 3185 -2929
rect 3349 -1553 3383 -1537
rect 3349 -2945 3383 -2929
rect 3547 -1553 3581 -1537
rect 3547 -2945 3581 -2929
rect 3745 -1553 3779 -1537
rect 3745 -2945 3779 -2929
rect 3943 -1553 3977 -1537
rect 3943 -2945 3977 -2929
rect 4141 -1553 4175 -1537
rect 4141 -2945 4175 -2929
<< viali >>
rect -4175 1553 -4141 2929
rect -3977 1553 -3943 2929
rect -3779 1553 -3745 2929
rect -3581 1553 -3547 2929
rect -3383 1553 -3349 2929
rect -3185 1553 -3151 2929
rect -2987 1553 -2953 2929
rect -2789 1553 -2755 2929
rect -2591 1553 -2557 2929
rect -2393 1553 -2359 2929
rect -2195 1553 -2161 2929
rect -1997 1553 -1963 2929
rect -1799 1553 -1765 2929
rect -1601 1553 -1567 2929
rect -1403 1553 -1369 2929
rect -1205 1553 -1171 2929
rect -1007 1553 -973 2929
rect -809 1553 -775 2929
rect -611 1553 -577 2929
rect -413 1553 -379 2929
rect -215 1553 -181 2929
rect -17 1553 17 2929
rect 181 1553 215 2929
rect 379 1553 413 2929
rect 577 1553 611 2929
rect 775 1553 809 2929
rect 973 1553 1007 2929
rect 1171 1553 1205 2929
rect 1369 1553 1403 2929
rect 1567 1553 1601 2929
rect 1765 1553 1799 2929
rect 1963 1553 1997 2929
rect 2161 1553 2195 2929
rect 2359 1553 2393 2929
rect 2557 1553 2591 2929
rect 2755 1553 2789 2929
rect 2953 1553 2987 2929
rect 3151 1553 3185 2929
rect 3349 1553 3383 2929
rect 3547 1553 3581 2929
rect 3745 1553 3779 2929
rect 3943 1553 3977 2929
rect 4141 1553 4175 2929
rect -4175 59 -4141 1435
rect -3977 59 -3943 1435
rect -3779 59 -3745 1435
rect -3581 59 -3547 1435
rect -3383 59 -3349 1435
rect -3185 59 -3151 1435
rect -2987 59 -2953 1435
rect -2789 59 -2755 1435
rect -2591 59 -2557 1435
rect -2393 59 -2359 1435
rect -2195 59 -2161 1435
rect -1997 59 -1963 1435
rect -1799 59 -1765 1435
rect -1601 59 -1567 1435
rect -1403 59 -1369 1435
rect -1205 59 -1171 1435
rect -1007 59 -973 1435
rect -809 59 -775 1435
rect -611 59 -577 1435
rect -413 59 -379 1435
rect -215 59 -181 1435
rect -17 59 17 1435
rect 181 59 215 1435
rect 379 59 413 1435
rect 577 59 611 1435
rect 775 59 809 1435
rect 973 59 1007 1435
rect 1171 59 1205 1435
rect 1369 59 1403 1435
rect 1567 59 1601 1435
rect 1765 59 1799 1435
rect 1963 59 1997 1435
rect 2161 59 2195 1435
rect 2359 59 2393 1435
rect 2557 59 2591 1435
rect 2755 59 2789 1435
rect 2953 59 2987 1435
rect 3151 59 3185 1435
rect 3349 59 3383 1435
rect 3547 59 3581 1435
rect 3745 59 3779 1435
rect 3943 59 3977 1435
rect 4141 59 4175 1435
rect -4175 -1435 -4141 -59
rect -3977 -1435 -3943 -59
rect -3779 -1435 -3745 -59
rect -3581 -1435 -3547 -59
rect -3383 -1435 -3349 -59
rect -3185 -1435 -3151 -59
rect -2987 -1435 -2953 -59
rect -2789 -1435 -2755 -59
rect -2591 -1435 -2557 -59
rect -2393 -1435 -2359 -59
rect -2195 -1435 -2161 -59
rect -1997 -1435 -1963 -59
rect -1799 -1435 -1765 -59
rect -1601 -1435 -1567 -59
rect -1403 -1435 -1369 -59
rect -1205 -1435 -1171 -59
rect -1007 -1435 -973 -59
rect -809 -1435 -775 -59
rect -611 -1435 -577 -59
rect -413 -1435 -379 -59
rect -215 -1435 -181 -59
rect -17 -1435 17 -59
rect 181 -1435 215 -59
rect 379 -1435 413 -59
rect 577 -1435 611 -59
rect 775 -1435 809 -59
rect 973 -1435 1007 -59
rect 1171 -1435 1205 -59
rect 1369 -1435 1403 -59
rect 1567 -1435 1601 -59
rect 1765 -1435 1799 -59
rect 1963 -1435 1997 -59
rect 2161 -1435 2195 -59
rect 2359 -1435 2393 -59
rect 2557 -1435 2591 -59
rect 2755 -1435 2789 -59
rect 2953 -1435 2987 -59
rect 3151 -1435 3185 -59
rect 3349 -1435 3383 -59
rect 3547 -1435 3581 -59
rect 3745 -1435 3779 -59
rect 3943 -1435 3977 -59
rect 4141 -1435 4175 -59
rect -4175 -2929 -4141 -1553
rect -3977 -2929 -3943 -1553
rect -3779 -2929 -3745 -1553
rect -3581 -2929 -3547 -1553
rect -3383 -2929 -3349 -1553
rect -3185 -2929 -3151 -1553
rect -2987 -2929 -2953 -1553
rect -2789 -2929 -2755 -1553
rect -2591 -2929 -2557 -1553
rect -2393 -2929 -2359 -1553
rect -2195 -2929 -2161 -1553
rect -1997 -2929 -1963 -1553
rect -1799 -2929 -1765 -1553
rect -1601 -2929 -1567 -1553
rect -1403 -2929 -1369 -1553
rect -1205 -2929 -1171 -1553
rect -1007 -2929 -973 -1553
rect -809 -2929 -775 -1553
rect -611 -2929 -577 -1553
rect -413 -2929 -379 -1553
rect -215 -2929 -181 -1553
rect -17 -2929 17 -1553
rect 181 -2929 215 -1553
rect 379 -2929 413 -1553
rect 577 -2929 611 -1553
rect 775 -2929 809 -1553
rect 973 -2929 1007 -1553
rect 1171 -2929 1205 -1553
rect 1369 -2929 1403 -1553
rect 1567 -2929 1601 -1553
rect 1765 -2929 1799 -1553
rect 1963 -2929 1997 -1553
rect 2161 -2929 2195 -1553
rect 2359 -2929 2393 -1553
rect 2557 -2929 2591 -1553
rect 2755 -2929 2789 -1553
rect 2953 -2929 2987 -1553
rect 3151 -2929 3185 -1553
rect 3349 -2929 3383 -1553
rect 3547 -2929 3581 -1553
rect 3745 -2929 3779 -1553
rect 3943 -2929 3977 -1553
rect 4141 -2929 4175 -1553
<< metal1 >>
rect -4181 2929 -4135 2941
rect -4181 1553 -4175 2929
rect -4141 1553 -4135 2929
rect -4181 1541 -4135 1553
rect -3983 2929 -3937 2941
rect -3983 1553 -3977 2929
rect -3943 1553 -3937 2929
rect -3983 1541 -3937 1553
rect -3785 2929 -3739 2941
rect -3785 1553 -3779 2929
rect -3745 1553 -3739 2929
rect -3785 1541 -3739 1553
rect -3587 2929 -3541 2941
rect -3587 1553 -3581 2929
rect -3547 1553 -3541 2929
rect -3587 1541 -3541 1553
rect -3389 2929 -3343 2941
rect -3389 1553 -3383 2929
rect -3349 1553 -3343 2929
rect -3389 1541 -3343 1553
rect -3191 2929 -3145 2941
rect -3191 1553 -3185 2929
rect -3151 1553 -3145 2929
rect -3191 1541 -3145 1553
rect -2993 2929 -2947 2941
rect -2993 1553 -2987 2929
rect -2953 1553 -2947 2929
rect -2993 1541 -2947 1553
rect -2795 2929 -2749 2941
rect -2795 1553 -2789 2929
rect -2755 1553 -2749 2929
rect -2795 1541 -2749 1553
rect -2597 2929 -2551 2941
rect -2597 1553 -2591 2929
rect -2557 1553 -2551 2929
rect -2597 1541 -2551 1553
rect -2399 2929 -2353 2941
rect -2399 1553 -2393 2929
rect -2359 1553 -2353 2929
rect -2399 1541 -2353 1553
rect -2201 2929 -2155 2941
rect -2201 1553 -2195 2929
rect -2161 1553 -2155 2929
rect -2201 1541 -2155 1553
rect -2003 2929 -1957 2941
rect -2003 1553 -1997 2929
rect -1963 1553 -1957 2929
rect -2003 1541 -1957 1553
rect -1805 2929 -1759 2941
rect -1805 1553 -1799 2929
rect -1765 1553 -1759 2929
rect -1805 1541 -1759 1553
rect -1607 2929 -1561 2941
rect -1607 1553 -1601 2929
rect -1567 1553 -1561 2929
rect -1607 1541 -1561 1553
rect -1409 2929 -1363 2941
rect -1409 1553 -1403 2929
rect -1369 1553 -1363 2929
rect -1409 1541 -1363 1553
rect -1211 2929 -1165 2941
rect -1211 1553 -1205 2929
rect -1171 1553 -1165 2929
rect -1211 1541 -1165 1553
rect -1013 2929 -967 2941
rect -1013 1553 -1007 2929
rect -973 1553 -967 2929
rect -1013 1541 -967 1553
rect -815 2929 -769 2941
rect -815 1553 -809 2929
rect -775 1553 -769 2929
rect -815 1541 -769 1553
rect -617 2929 -571 2941
rect -617 1553 -611 2929
rect -577 1553 -571 2929
rect -617 1541 -571 1553
rect -419 2929 -373 2941
rect -419 1553 -413 2929
rect -379 1553 -373 2929
rect -419 1541 -373 1553
rect -221 2929 -175 2941
rect -221 1553 -215 2929
rect -181 1553 -175 2929
rect -221 1541 -175 1553
rect -23 2929 23 2941
rect -23 1553 -17 2929
rect 17 1553 23 2929
rect -23 1541 23 1553
rect 175 2929 221 2941
rect 175 1553 181 2929
rect 215 1553 221 2929
rect 175 1541 221 1553
rect 373 2929 419 2941
rect 373 1553 379 2929
rect 413 1553 419 2929
rect 373 1541 419 1553
rect 571 2929 617 2941
rect 571 1553 577 2929
rect 611 1553 617 2929
rect 571 1541 617 1553
rect 769 2929 815 2941
rect 769 1553 775 2929
rect 809 1553 815 2929
rect 769 1541 815 1553
rect 967 2929 1013 2941
rect 967 1553 973 2929
rect 1007 1553 1013 2929
rect 967 1541 1013 1553
rect 1165 2929 1211 2941
rect 1165 1553 1171 2929
rect 1205 1553 1211 2929
rect 1165 1541 1211 1553
rect 1363 2929 1409 2941
rect 1363 1553 1369 2929
rect 1403 1553 1409 2929
rect 1363 1541 1409 1553
rect 1561 2929 1607 2941
rect 1561 1553 1567 2929
rect 1601 1553 1607 2929
rect 1561 1541 1607 1553
rect 1759 2929 1805 2941
rect 1759 1553 1765 2929
rect 1799 1553 1805 2929
rect 1759 1541 1805 1553
rect 1957 2929 2003 2941
rect 1957 1553 1963 2929
rect 1997 1553 2003 2929
rect 1957 1541 2003 1553
rect 2155 2929 2201 2941
rect 2155 1553 2161 2929
rect 2195 1553 2201 2929
rect 2155 1541 2201 1553
rect 2353 2929 2399 2941
rect 2353 1553 2359 2929
rect 2393 1553 2399 2929
rect 2353 1541 2399 1553
rect 2551 2929 2597 2941
rect 2551 1553 2557 2929
rect 2591 1553 2597 2929
rect 2551 1541 2597 1553
rect 2749 2929 2795 2941
rect 2749 1553 2755 2929
rect 2789 1553 2795 2929
rect 2749 1541 2795 1553
rect 2947 2929 2993 2941
rect 2947 1553 2953 2929
rect 2987 1553 2993 2929
rect 2947 1541 2993 1553
rect 3145 2929 3191 2941
rect 3145 1553 3151 2929
rect 3185 1553 3191 2929
rect 3145 1541 3191 1553
rect 3343 2929 3389 2941
rect 3343 1553 3349 2929
rect 3383 1553 3389 2929
rect 3343 1541 3389 1553
rect 3541 2929 3587 2941
rect 3541 1553 3547 2929
rect 3581 1553 3587 2929
rect 3541 1541 3587 1553
rect 3739 2929 3785 2941
rect 3739 1553 3745 2929
rect 3779 1553 3785 2929
rect 3739 1541 3785 1553
rect 3937 2929 3983 2941
rect 3937 1553 3943 2929
rect 3977 1553 3983 2929
rect 3937 1541 3983 1553
rect 4135 2929 4181 2941
rect 4135 1553 4141 2929
rect 4175 1553 4181 2929
rect 4135 1541 4181 1553
rect -4181 1435 -4135 1447
rect -4181 59 -4175 1435
rect -4141 59 -4135 1435
rect -4181 47 -4135 59
rect -3983 1435 -3937 1447
rect -3983 59 -3977 1435
rect -3943 59 -3937 1435
rect -3983 47 -3937 59
rect -3785 1435 -3739 1447
rect -3785 59 -3779 1435
rect -3745 59 -3739 1435
rect -3785 47 -3739 59
rect -3587 1435 -3541 1447
rect -3587 59 -3581 1435
rect -3547 59 -3541 1435
rect -3587 47 -3541 59
rect -3389 1435 -3343 1447
rect -3389 59 -3383 1435
rect -3349 59 -3343 1435
rect -3389 47 -3343 59
rect -3191 1435 -3145 1447
rect -3191 59 -3185 1435
rect -3151 59 -3145 1435
rect -3191 47 -3145 59
rect -2993 1435 -2947 1447
rect -2993 59 -2987 1435
rect -2953 59 -2947 1435
rect -2993 47 -2947 59
rect -2795 1435 -2749 1447
rect -2795 59 -2789 1435
rect -2755 59 -2749 1435
rect -2795 47 -2749 59
rect -2597 1435 -2551 1447
rect -2597 59 -2591 1435
rect -2557 59 -2551 1435
rect -2597 47 -2551 59
rect -2399 1435 -2353 1447
rect -2399 59 -2393 1435
rect -2359 59 -2353 1435
rect -2399 47 -2353 59
rect -2201 1435 -2155 1447
rect -2201 59 -2195 1435
rect -2161 59 -2155 1435
rect -2201 47 -2155 59
rect -2003 1435 -1957 1447
rect -2003 59 -1997 1435
rect -1963 59 -1957 1435
rect -2003 47 -1957 59
rect -1805 1435 -1759 1447
rect -1805 59 -1799 1435
rect -1765 59 -1759 1435
rect -1805 47 -1759 59
rect -1607 1435 -1561 1447
rect -1607 59 -1601 1435
rect -1567 59 -1561 1435
rect -1607 47 -1561 59
rect -1409 1435 -1363 1447
rect -1409 59 -1403 1435
rect -1369 59 -1363 1435
rect -1409 47 -1363 59
rect -1211 1435 -1165 1447
rect -1211 59 -1205 1435
rect -1171 59 -1165 1435
rect -1211 47 -1165 59
rect -1013 1435 -967 1447
rect -1013 59 -1007 1435
rect -973 59 -967 1435
rect -1013 47 -967 59
rect -815 1435 -769 1447
rect -815 59 -809 1435
rect -775 59 -769 1435
rect -815 47 -769 59
rect -617 1435 -571 1447
rect -617 59 -611 1435
rect -577 59 -571 1435
rect -617 47 -571 59
rect -419 1435 -373 1447
rect -419 59 -413 1435
rect -379 59 -373 1435
rect -419 47 -373 59
rect -221 1435 -175 1447
rect -221 59 -215 1435
rect -181 59 -175 1435
rect -221 47 -175 59
rect -23 1435 23 1447
rect -23 59 -17 1435
rect 17 59 23 1435
rect -23 47 23 59
rect 175 1435 221 1447
rect 175 59 181 1435
rect 215 59 221 1435
rect 175 47 221 59
rect 373 1435 419 1447
rect 373 59 379 1435
rect 413 59 419 1435
rect 373 47 419 59
rect 571 1435 617 1447
rect 571 59 577 1435
rect 611 59 617 1435
rect 571 47 617 59
rect 769 1435 815 1447
rect 769 59 775 1435
rect 809 59 815 1435
rect 769 47 815 59
rect 967 1435 1013 1447
rect 967 59 973 1435
rect 1007 59 1013 1435
rect 967 47 1013 59
rect 1165 1435 1211 1447
rect 1165 59 1171 1435
rect 1205 59 1211 1435
rect 1165 47 1211 59
rect 1363 1435 1409 1447
rect 1363 59 1369 1435
rect 1403 59 1409 1435
rect 1363 47 1409 59
rect 1561 1435 1607 1447
rect 1561 59 1567 1435
rect 1601 59 1607 1435
rect 1561 47 1607 59
rect 1759 1435 1805 1447
rect 1759 59 1765 1435
rect 1799 59 1805 1435
rect 1759 47 1805 59
rect 1957 1435 2003 1447
rect 1957 59 1963 1435
rect 1997 59 2003 1435
rect 1957 47 2003 59
rect 2155 1435 2201 1447
rect 2155 59 2161 1435
rect 2195 59 2201 1435
rect 2155 47 2201 59
rect 2353 1435 2399 1447
rect 2353 59 2359 1435
rect 2393 59 2399 1435
rect 2353 47 2399 59
rect 2551 1435 2597 1447
rect 2551 59 2557 1435
rect 2591 59 2597 1435
rect 2551 47 2597 59
rect 2749 1435 2795 1447
rect 2749 59 2755 1435
rect 2789 59 2795 1435
rect 2749 47 2795 59
rect 2947 1435 2993 1447
rect 2947 59 2953 1435
rect 2987 59 2993 1435
rect 2947 47 2993 59
rect 3145 1435 3191 1447
rect 3145 59 3151 1435
rect 3185 59 3191 1435
rect 3145 47 3191 59
rect 3343 1435 3389 1447
rect 3343 59 3349 1435
rect 3383 59 3389 1435
rect 3343 47 3389 59
rect 3541 1435 3587 1447
rect 3541 59 3547 1435
rect 3581 59 3587 1435
rect 3541 47 3587 59
rect 3739 1435 3785 1447
rect 3739 59 3745 1435
rect 3779 59 3785 1435
rect 3739 47 3785 59
rect 3937 1435 3983 1447
rect 3937 59 3943 1435
rect 3977 59 3983 1435
rect 3937 47 3983 59
rect 4135 1435 4181 1447
rect 4135 59 4141 1435
rect 4175 59 4181 1435
rect 4135 47 4181 59
rect -4181 -59 -4135 -47
rect -4181 -1435 -4175 -59
rect -4141 -1435 -4135 -59
rect -4181 -1447 -4135 -1435
rect -3983 -59 -3937 -47
rect -3983 -1435 -3977 -59
rect -3943 -1435 -3937 -59
rect -3983 -1447 -3937 -1435
rect -3785 -59 -3739 -47
rect -3785 -1435 -3779 -59
rect -3745 -1435 -3739 -59
rect -3785 -1447 -3739 -1435
rect -3587 -59 -3541 -47
rect -3587 -1435 -3581 -59
rect -3547 -1435 -3541 -59
rect -3587 -1447 -3541 -1435
rect -3389 -59 -3343 -47
rect -3389 -1435 -3383 -59
rect -3349 -1435 -3343 -59
rect -3389 -1447 -3343 -1435
rect -3191 -59 -3145 -47
rect -3191 -1435 -3185 -59
rect -3151 -1435 -3145 -59
rect -3191 -1447 -3145 -1435
rect -2993 -59 -2947 -47
rect -2993 -1435 -2987 -59
rect -2953 -1435 -2947 -59
rect -2993 -1447 -2947 -1435
rect -2795 -59 -2749 -47
rect -2795 -1435 -2789 -59
rect -2755 -1435 -2749 -59
rect -2795 -1447 -2749 -1435
rect -2597 -59 -2551 -47
rect -2597 -1435 -2591 -59
rect -2557 -1435 -2551 -59
rect -2597 -1447 -2551 -1435
rect -2399 -59 -2353 -47
rect -2399 -1435 -2393 -59
rect -2359 -1435 -2353 -59
rect -2399 -1447 -2353 -1435
rect -2201 -59 -2155 -47
rect -2201 -1435 -2195 -59
rect -2161 -1435 -2155 -59
rect -2201 -1447 -2155 -1435
rect -2003 -59 -1957 -47
rect -2003 -1435 -1997 -59
rect -1963 -1435 -1957 -59
rect -2003 -1447 -1957 -1435
rect -1805 -59 -1759 -47
rect -1805 -1435 -1799 -59
rect -1765 -1435 -1759 -59
rect -1805 -1447 -1759 -1435
rect -1607 -59 -1561 -47
rect -1607 -1435 -1601 -59
rect -1567 -1435 -1561 -59
rect -1607 -1447 -1561 -1435
rect -1409 -59 -1363 -47
rect -1409 -1435 -1403 -59
rect -1369 -1435 -1363 -59
rect -1409 -1447 -1363 -1435
rect -1211 -59 -1165 -47
rect -1211 -1435 -1205 -59
rect -1171 -1435 -1165 -59
rect -1211 -1447 -1165 -1435
rect -1013 -59 -967 -47
rect -1013 -1435 -1007 -59
rect -973 -1435 -967 -59
rect -1013 -1447 -967 -1435
rect -815 -59 -769 -47
rect -815 -1435 -809 -59
rect -775 -1435 -769 -59
rect -815 -1447 -769 -1435
rect -617 -59 -571 -47
rect -617 -1435 -611 -59
rect -577 -1435 -571 -59
rect -617 -1447 -571 -1435
rect -419 -59 -373 -47
rect -419 -1435 -413 -59
rect -379 -1435 -373 -59
rect -419 -1447 -373 -1435
rect -221 -59 -175 -47
rect -221 -1435 -215 -59
rect -181 -1435 -175 -59
rect -221 -1447 -175 -1435
rect -23 -59 23 -47
rect -23 -1435 -17 -59
rect 17 -1435 23 -59
rect -23 -1447 23 -1435
rect 175 -59 221 -47
rect 175 -1435 181 -59
rect 215 -1435 221 -59
rect 175 -1447 221 -1435
rect 373 -59 419 -47
rect 373 -1435 379 -59
rect 413 -1435 419 -59
rect 373 -1447 419 -1435
rect 571 -59 617 -47
rect 571 -1435 577 -59
rect 611 -1435 617 -59
rect 571 -1447 617 -1435
rect 769 -59 815 -47
rect 769 -1435 775 -59
rect 809 -1435 815 -59
rect 769 -1447 815 -1435
rect 967 -59 1013 -47
rect 967 -1435 973 -59
rect 1007 -1435 1013 -59
rect 967 -1447 1013 -1435
rect 1165 -59 1211 -47
rect 1165 -1435 1171 -59
rect 1205 -1435 1211 -59
rect 1165 -1447 1211 -1435
rect 1363 -59 1409 -47
rect 1363 -1435 1369 -59
rect 1403 -1435 1409 -59
rect 1363 -1447 1409 -1435
rect 1561 -59 1607 -47
rect 1561 -1435 1567 -59
rect 1601 -1435 1607 -59
rect 1561 -1447 1607 -1435
rect 1759 -59 1805 -47
rect 1759 -1435 1765 -59
rect 1799 -1435 1805 -59
rect 1759 -1447 1805 -1435
rect 1957 -59 2003 -47
rect 1957 -1435 1963 -59
rect 1997 -1435 2003 -59
rect 1957 -1447 2003 -1435
rect 2155 -59 2201 -47
rect 2155 -1435 2161 -59
rect 2195 -1435 2201 -59
rect 2155 -1447 2201 -1435
rect 2353 -59 2399 -47
rect 2353 -1435 2359 -59
rect 2393 -1435 2399 -59
rect 2353 -1447 2399 -1435
rect 2551 -59 2597 -47
rect 2551 -1435 2557 -59
rect 2591 -1435 2597 -59
rect 2551 -1447 2597 -1435
rect 2749 -59 2795 -47
rect 2749 -1435 2755 -59
rect 2789 -1435 2795 -59
rect 2749 -1447 2795 -1435
rect 2947 -59 2993 -47
rect 2947 -1435 2953 -59
rect 2987 -1435 2993 -59
rect 2947 -1447 2993 -1435
rect 3145 -59 3191 -47
rect 3145 -1435 3151 -59
rect 3185 -1435 3191 -59
rect 3145 -1447 3191 -1435
rect 3343 -59 3389 -47
rect 3343 -1435 3349 -59
rect 3383 -1435 3389 -59
rect 3343 -1447 3389 -1435
rect 3541 -59 3587 -47
rect 3541 -1435 3547 -59
rect 3581 -1435 3587 -59
rect 3541 -1447 3587 -1435
rect 3739 -59 3785 -47
rect 3739 -1435 3745 -59
rect 3779 -1435 3785 -59
rect 3739 -1447 3785 -1435
rect 3937 -59 3983 -47
rect 3937 -1435 3943 -59
rect 3977 -1435 3983 -59
rect 3937 -1447 3983 -1435
rect 4135 -59 4181 -47
rect 4135 -1435 4141 -59
rect 4175 -1435 4181 -59
rect 4135 -1447 4181 -1435
rect -4181 -1553 -4135 -1541
rect -4181 -2929 -4175 -1553
rect -4141 -2929 -4135 -1553
rect -4181 -2941 -4135 -2929
rect -3983 -1553 -3937 -1541
rect -3983 -2929 -3977 -1553
rect -3943 -2929 -3937 -1553
rect -3983 -2941 -3937 -2929
rect -3785 -1553 -3739 -1541
rect -3785 -2929 -3779 -1553
rect -3745 -2929 -3739 -1553
rect -3785 -2941 -3739 -2929
rect -3587 -1553 -3541 -1541
rect -3587 -2929 -3581 -1553
rect -3547 -2929 -3541 -1553
rect -3587 -2941 -3541 -2929
rect -3389 -1553 -3343 -1541
rect -3389 -2929 -3383 -1553
rect -3349 -2929 -3343 -1553
rect -3389 -2941 -3343 -2929
rect -3191 -1553 -3145 -1541
rect -3191 -2929 -3185 -1553
rect -3151 -2929 -3145 -1553
rect -3191 -2941 -3145 -2929
rect -2993 -1553 -2947 -1541
rect -2993 -2929 -2987 -1553
rect -2953 -2929 -2947 -1553
rect -2993 -2941 -2947 -2929
rect -2795 -1553 -2749 -1541
rect -2795 -2929 -2789 -1553
rect -2755 -2929 -2749 -1553
rect -2795 -2941 -2749 -2929
rect -2597 -1553 -2551 -1541
rect -2597 -2929 -2591 -1553
rect -2557 -2929 -2551 -1553
rect -2597 -2941 -2551 -2929
rect -2399 -1553 -2353 -1541
rect -2399 -2929 -2393 -1553
rect -2359 -2929 -2353 -1553
rect -2399 -2941 -2353 -2929
rect -2201 -1553 -2155 -1541
rect -2201 -2929 -2195 -1553
rect -2161 -2929 -2155 -1553
rect -2201 -2941 -2155 -2929
rect -2003 -1553 -1957 -1541
rect -2003 -2929 -1997 -1553
rect -1963 -2929 -1957 -1553
rect -2003 -2941 -1957 -2929
rect -1805 -1553 -1759 -1541
rect -1805 -2929 -1799 -1553
rect -1765 -2929 -1759 -1553
rect -1805 -2941 -1759 -2929
rect -1607 -1553 -1561 -1541
rect -1607 -2929 -1601 -1553
rect -1567 -2929 -1561 -1553
rect -1607 -2941 -1561 -2929
rect -1409 -1553 -1363 -1541
rect -1409 -2929 -1403 -1553
rect -1369 -2929 -1363 -1553
rect -1409 -2941 -1363 -2929
rect -1211 -1553 -1165 -1541
rect -1211 -2929 -1205 -1553
rect -1171 -2929 -1165 -1553
rect -1211 -2941 -1165 -2929
rect -1013 -1553 -967 -1541
rect -1013 -2929 -1007 -1553
rect -973 -2929 -967 -1553
rect -1013 -2941 -967 -2929
rect -815 -1553 -769 -1541
rect -815 -2929 -809 -1553
rect -775 -2929 -769 -1553
rect -815 -2941 -769 -2929
rect -617 -1553 -571 -1541
rect -617 -2929 -611 -1553
rect -577 -2929 -571 -1553
rect -617 -2941 -571 -2929
rect -419 -1553 -373 -1541
rect -419 -2929 -413 -1553
rect -379 -2929 -373 -1553
rect -419 -2941 -373 -2929
rect -221 -1553 -175 -1541
rect -221 -2929 -215 -1553
rect -181 -2929 -175 -1553
rect -221 -2941 -175 -2929
rect -23 -1553 23 -1541
rect -23 -2929 -17 -1553
rect 17 -2929 23 -1553
rect -23 -2941 23 -2929
rect 175 -1553 221 -1541
rect 175 -2929 181 -1553
rect 215 -2929 221 -1553
rect 175 -2941 221 -2929
rect 373 -1553 419 -1541
rect 373 -2929 379 -1553
rect 413 -2929 419 -1553
rect 373 -2941 419 -2929
rect 571 -1553 617 -1541
rect 571 -2929 577 -1553
rect 611 -2929 617 -1553
rect 571 -2941 617 -2929
rect 769 -1553 815 -1541
rect 769 -2929 775 -1553
rect 809 -2929 815 -1553
rect 769 -2941 815 -2929
rect 967 -1553 1013 -1541
rect 967 -2929 973 -1553
rect 1007 -2929 1013 -1553
rect 967 -2941 1013 -2929
rect 1165 -1553 1211 -1541
rect 1165 -2929 1171 -1553
rect 1205 -2929 1211 -1553
rect 1165 -2941 1211 -2929
rect 1363 -1553 1409 -1541
rect 1363 -2929 1369 -1553
rect 1403 -2929 1409 -1553
rect 1363 -2941 1409 -2929
rect 1561 -1553 1607 -1541
rect 1561 -2929 1567 -1553
rect 1601 -2929 1607 -1553
rect 1561 -2941 1607 -2929
rect 1759 -1553 1805 -1541
rect 1759 -2929 1765 -1553
rect 1799 -2929 1805 -1553
rect 1759 -2941 1805 -2929
rect 1957 -1553 2003 -1541
rect 1957 -2929 1963 -1553
rect 1997 -2929 2003 -1553
rect 1957 -2941 2003 -2929
rect 2155 -1553 2201 -1541
rect 2155 -2929 2161 -1553
rect 2195 -2929 2201 -1553
rect 2155 -2941 2201 -2929
rect 2353 -1553 2399 -1541
rect 2353 -2929 2359 -1553
rect 2393 -2929 2399 -1553
rect 2353 -2941 2399 -2929
rect 2551 -1553 2597 -1541
rect 2551 -2929 2557 -1553
rect 2591 -2929 2597 -1553
rect 2551 -2941 2597 -2929
rect 2749 -1553 2795 -1541
rect 2749 -2929 2755 -1553
rect 2789 -2929 2795 -1553
rect 2749 -2941 2795 -2929
rect 2947 -1553 2993 -1541
rect 2947 -2929 2953 -1553
rect 2987 -2929 2993 -1553
rect 2947 -2941 2993 -2929
rect 3145 -1553 3191 -1541
rect 3145 -2929 3151 -1553
rect 3185 -2929 3191 -1553
rect 3145 -2941 3191 -2929
rect 3343 -1553 3389 -1541
rect 3343 -2929 3349 -1553
rect 3383 -2929 3389 -1553
rect 3343 -2941 3389 -2929
rect 3541 -1553 3587 -1541
rect 3541 -2929 3547 -1553
rect 3581 -2929 3587 -1553
rect 3541 -2941 3587 -2929
rect 3739 -1553 3785 -1541
rect 3739 -2929 3745 -1553
rect 3779 -2929 3785 -1553
rect 3739 -2941 3785 -2929
rect 3937 -1553 3983 -1541
rect 3937 -2929 3943 -1553
rect 3977 -2929 3983 -1553
rect 3937 -2941 3983 -2929
rect 4135 -1553 4181 -1541
rect 4135 -2929 4141 -1553
rect 4175 -2929 4181 -1553
rect 4135 -2941 4181 -2929
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 4 nf 42 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
