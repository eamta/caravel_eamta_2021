magic
tech sky130A
magscale 1 2
timestamp 1624338677
<< nwell >>
rect 56 972 3586 1174
rect 3506 544 3586 972
rect 3508 -922 3586 -494
rect 56 -1196 3586 -922
<< poly >>
rect -158 40 -128 1174
rect -86 148 -56 1174
rect 3024 1144 3560 1174
rect 3492 760 3550 788
rect 3426 734 3550 760
rect -86 132 16 148
rect -86 98 -34 132
rect 0 112 16 132
rect 0 98 76 112
rect -86 82 76 98
rect -158 10 70 40
rect -158 -1196 -128 10
rect -86 -48 82 -32
rect -86 -82 -34 -48
rect 0 -62 82 -48
rect 0 -82 16 -62
rect -86 -98 16 -82
rect -86 -1196 -56 -98
rect 3520 -540 3550 734
rect 3520 -556 3586 -540
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 3520 -606 3586 -590
rect 3490 -736 3560 -702
rect 3426 -756 3560 -736
rect 3422 -842 3488 -826
rect 3422 -876 3438 -842
rect 3472 -876 3488 -842
rect 3422 -892 3488 -876
rect 3422 -896 3452 -892
rect 3024 -926 3452 -896
rect 3530 -1196 3560 -756
<< polycont >>
rect -34 98 0 132
rect -34 -82 0 -48
rect 3536 -590 3570 -556
rect 3438 -876 3472 -842
<< locali >>
rect -50 98 -34 132
rect 0 98 16 132
rect -50 -82 -34 -48
rect 0 -82 16 -48
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 3422 -876 3438 -842
rect 3472 -876 3488 -842
<< viali >>
rect -34 98 0 132
rect -34 -82 0 -48
rect 3536 -590 3570 -556
rect 3438 -876 3472 -842
<< metal1 >>
rect 56 972 3586 1174
rect -50 132 16 148
rect -50 98 -34 132
rect 0 98 16 132
rect -50 82 16 98
rect -34 -32 0 82
rect -50 -48 16 -32
rect -50 -82 -34 -48
rect 0 -82 16 -48
rect -50 -98 16 -82
rect 58 -156 3586 206
rect 3520 -556 3586 -540
rect 3520 -590 3536 -556
rect 3570 -590 3586 -556
rect 3520 -606 3586 -590
rect 3520 -826 3554 -606
rect 3422 -842 3554 -826
rect 3422 -876 3438 -842
rect 3472 -860 3554 -842
rect 3472 -876 3488 -860
rect 3422 -892 3488 -876
rect 56 -1196 3586 -922
<< metal2 >>
rect 2946 364 2998 416
rect 2946 -366 2998 -314
use c1b  c1b_1
timestamp 1624338677
transform 1 0 58 0 -1 -68
box -72 -108 3457 1056
use c1b  c1b_0
timestamp 1624338677
transform 1 0 58 0 1 118
box -72 -108 3457 1056
<< labels >>
rlabel metal2 2946 364 2998 416 1 b0
rlabel metal2 2946 -366 2998 -314 1 b1
rlabel poly -150 1154 -134 1170 1 clr
rlabel poly -78 1154 -62 1170 1 clk
rlabel metal1 3476 0 3506 58 1 vss
rlabel metal1 924 -996 966 -968 1 vdd
rlabel metal1 3466 992 3496 1050 1 vdd
rlabel poly -78 -54 -62 -38 1 clk
rlabel poly 3540 1152 3552 1168 1 ce
rlabel poly 3538 -916 3554 -874 1 out
<< end >>
