magic
tech sky130A
magscale 1 2
timestamp 1616600406
<< error_p >>
rect -5713 381 -5655 387
rect -5481 381 -5423 387
rect -5249 381 -5191 387
rect -5017 381 -4959 387
rect -4785 381 -4727 387
rect -4553 381 -4495 387
rect -4321 381 -4263 387
rect -4089 381 -4031 387
rect -3857 381 -3799 387
rect -3625 381 -3567 387
rect -3393 381 -3335 387
rect -3161 381 -3103 387
rect -2929 381 -2871 387
rect -2697 381 -2639 387
rect -2465 381 -2407 387
rect -2233 381 -2175 387
rect -2001 381 -1943 387
rect -1769 381 -1711 387
rect -1537 381 -1479 387
rect -1305 381 -1247 387
rect -1073 381 -1015 387
rect -841 381 -783 387
rect -609 381 -551 387
rect -377 381 -319 387
rect -145 381 -87 387
rect 87 381 145 387
rect 319 381 377 387
rect 551 381 609 387
rect 783 381 841 387
rect 1015 381 1073 387
rect 1247 381 1305 387
rect 1479 381 1537 387
rect 1711 381 1769 387
rect 1943 381 2001 387
rect 2175 381 2233 387
rect 2407 381 2465 387
rect 2639 381 2697 387
rect 2871 381 2929 387
rect 3103 381 3161 387
rect 3335 381 3393 387
rect 3567 381 3625 387
rect 3799 381 3857 387
rect 4031 381 4089 387
rect 4263 381 4321 387
rect 4495 381 4553 387
rect 4727 381 4785 387
rect 4959 381 5017 387
rect 5191 381 5249 387
rect 5423 381 5481 387
rect 5655 381 5713 387
rect -5713 347 -5701 381
rect -5481 347 -5469 381
rect -5249 347 -5237 381
rect -5017 347 -5005 381
rect -4785 347 -4773 381
rect -4553 347 -4541 381
rect -4321 347 -4309 381
rect -4089 347 -4077 381
rect -3857 347 -3845 381
rect -3625 347 -3613 381
rect -3393 347 -3381 381
rect -3161 347 -3149 381
rect -2929 347 -2917 381
rect -2697 347 -2685 381
rect -2465 347 -2453 381
rect -2233 347 -2221 381
rect -2001 347 -1989 381
rect -1769 347 -1757 381
rect -1537 347 -1525 381
rect -1305 347 -1293 381
rect -1073 347 -1061 381
rect -841 347 -829 381
rect -609 347 -597 381
rect -377 347 -365 381
rect -145 347 -133 381
rect 87 347 99 381
rect 319 347 331 381
rect 551 347 563 381
rect 783 347 795 381
rect 1015 347 1027 381
rect 1247 347 1259 381
rect 1479 347 1491 381
rect 1711 347 1723 381
rect 1943 347 1955 381
rect 2175 347 2187 381
rect 2407 347 2419 381
rect 2639 347 2651 381
rect 2871 347 2883 381
rect 3103 347 3115 381
rect 3335 347 3347 381
rect 3567 347 3579 381
rect 3799 347 3811 381
rect 4031 347 4043 381
rect 4263 347 4275 381
rect 4495 347 4507 381
rect 4727 347 4739 381
rect 4959 347 4971 381
rect 5191 347 5203 381
rect 5423 347 5435 381
rect 5655 347 5667 381
rect -5713 341 -5655 347
rect -5481 341 -5423 347
rect -5249 341 -5191 347
rect -5017 341 -4959 347
rect -4785 341 -4727 347
rect -4553 341 -4495 347
rect -4321 341 -4263 347
rect -4089 341 -4031 347
rect -3857 341 -3799 347
rect -3625 341 -3567 347
rect -3393 341 -3335 347
rect -3161 341 -3103 347
rect -2929 341 -2871 347
rect -2697 341 -2639 347
rect -2465 341 -2407 347
rect -2233 341 -2175 347
rect -2001 341 -1943 347
rect -1769 341 -1711 347
rect -1537 341 -1479 347
rect -1305 341 -1247 347
rect -1073 341 -1015 347
rect -841 341 -783 347
rect -609 341 -551 347
rect -377 341 -319 347
rect -145 341 -87 347
rect 87 341 145 347
rect 319 341 377 347
rect 551 341 609 347
rect 783 341 841 347
rect 1015 341 1073 347
rect 1247 341 1305 347
rect 1479 341 1537 347
rect 1711 341 1769 347
rect 1943 341 2001 347
rect 2175 341 2233 347
rect 2407 341 2465 347
rect 2639 341 2697 347
rect 2871 341 2929 347
rect 3103 341 3161 347
rect 3335 341 3393 347
rect 3567 341 3625 347
rect 3799 341 3857 347
rect 4031 341 4089 347
rect 4263 341 4321 347
rect 4495 341 4553 347
rect 4727 341 4785 347
rect 4959 341 5017 347
rect 5191 341 5249 347
rect 5423 341 5481 347
rect 5655 341 5713 347
rect -5713 -347 -5655 -341
rect -5481 -347 -5423 -341
rect -5249 -347 -5191 -341
rect -5017 -347 -4959 -341
rect -4785 -347 -4727 -341
rect -4553 -347 -4495 -341
rect -4321 -347 -4263 -341
rect -4089 -347 -4031 -341
rect -3857 -347 -3799 -341
rect -3625 -347 -3567 -341
rect -3393 -347 -3335 -341
rect -3161 -347 -3103 -341
rect -2929 -347 -2871 -341
rect -2697 -347 -2639 -341
rect -2465 -347 -2407 -341
rect -2233 -347 -2175 -341
rect -2001 -347 -1943 -341
rect -1769 -347 -1711 -341
rect -1537 -347 -1479 -341
rect -1305 -347 -1247 -341
rect -1073 -347 -1015 -341
rect -841 -347 -783 -341
rect -609 -347 -551 -341
rect -377 -347 -319 -341
rect -145 -347 -87 -341
rect 87 -347 145 -341
rect 319 -347 377 -341
rect 551 -347 609 -341
rect 783 -347 841 -341
rect 1015 -347 1073 -341
rect 1247 -347 1305 -341
rect 1479 -347 1537 -341
rect 1711 -347 1769 -341
rect 1943 -347 2001 -341
rect 2175 -347 2233 -341
rect 2407 -347 2465 -341
rect 2639 -347 2697 -341
rect 2871 -347 2929 -341
rect 3103 -347 3161 -341
rect 3335 -347 3393 -341
rect 3567 -347 3625 -341
rect 3799 -347 3857 -341
rect 4031 -347 4089 -341
rect 4263 -347 4321 -341
rect 4495 -347 4553 -341
rect 4727 -347 4785 -341
rect 4959 -347 5017 -341
rect 5191 -347 5249 -341
rect 5423 -347 5481 -341
rect 5655 -347 5713 -341
rect -5713 -381 -5701 -347
rect -5481 -381 -5469 -347
rect -5249 -381 -5237 -347
rect -5017 -381 -5005 -347
rect -4785 -381 -4773 -347
rect -4553 -381 -4541 -347
rect -4321 -381 -4309 -347
rect -4089 -381 -4077 -347
rect -3857 -381 -3845 -347
rect -3625 -381 -3613 -347
rect -3393 -381 -3381 -347
rect -3161 -381 -3149 -347
rect -2929 -381 -2917 -347
rect -2697 -381 -2685 -347
rect -2465 -381 -2453 -347
rect -2233 -381 -2221 -347
rect -2001 -381 -1989 -347
rect -1769 -381 -1757 -347
rect -1537 -381 -1525 -347
rect -1305 -381 -1293 -347
rect -1073 -381 -1061 -347
rect -841 -381 -829 -347
rect -609 -381 -597 -347
rect -377 -381 -365 -347
rect -145 -381 -133 -347
rect 87 -381 99 -347
rect 319 -381 331 -347
rect 551 -381 563 -347
rect 783 -381 795 -347
rect 1015 -381 1027 -347
rect 1247 -381 1259 -347
rect 1479 -381 1491 -347
rect 1711 -381 1723 -347
rect 1943 -381 1955 -347
rect 2175 -381 2187 -347
rect 2407 -381 2419 -347
rect 2639 -381 2651 -347
rect 2871 -381 2883 -347
rect 3103 -381 3115 -347
rect 3335 -381 3347 -347
rect 3567 -381 3579 -347
rect 3799 -381 3811 -347
rect 4031 -381 4043 -347
rect 4263 -381 4275 -347
rect 4495 -381 4507 -347
rect 4727 -381 4739 -347
rect 4959 -381 4971 -347
rect 5191 -381 5203 -347
rect 5423 -381 5435 -347
rect 5655 -381 5667 -347
rect -5713 -387 -5655 -381
rect -5481 -387 -5423 -381
rect -5249 -387 -5191 -381
rect -5017 -387 -4959 -381
rect -4785 -387 -4727 -381
rect -4553 -387 -4495 -381
rect -4321 -387 -4263 -381
rect -4089 -387 -4031 -381
rect -3857 -387 -3799 -381
rect -3625 -387 -3567 -381
rect -3393 -387 -3335 -381
rect -3161 -387 -3103 -381
rect -2929 -387 -2871 -381
rect -2697 -387 -2639 -381
rect -2465 -387 -2407 -381
rect -2233 -387 -2175 -381
rect -2001 -387 -1943 -381
rect -1769 -387 -1711 -381
rect -1537 -387 -1479 -381
rect -1305 -387 -1247 -381
rect -1073 -387 -1015 -381
rect -841 -387 -783 -381
rect -609 -387 -551 -381
rect -377 -387 -319 -381
rect -145 -387 -87 -381
rect 87 -387 145 -381
rect 319 -387 377 -381
rect 551 -387 609 -381
rect 783 -387 841 -381
rect 1015 -387 1073 -381
rect 1247 -387 1305 -381
rect 1479 -387 1537 -381
rect 1711 -387 1769 -381
rect 1943 -387 2001 -381
rect 2175 -387 2233 -381
rect 2407 -387 2465 -381
rect 2639 -387 2697 -381
rect 2871 -387 2929 -381
rect 3103 -387 3161 -381
rect 3335 -387 3393 -381
rect 3567 -387 3625 -381
rect 3799 -387 3857 -381
rect 4031 -387 4089 -381
rect 4263 -387 4321 -381
rect 4495 -387 4553 -381
rect 4727 -387 4785 -381
rect 4959 -387 5017 -381
rect 5191 -387 5249 -381
rect 5423 -387 5481 -381
rect 5655 -387 5713 -381
<< nwell >>
rect -5910 -519 5910 519
<< pmos >>
rect -5714 -300 -5654 300
rect -5482 -300 -5422 300
rect -5250 -300 -5190 300
rect -5018 -300 -4958 300
rect -4786 -300 -4726 300
rect -4554 -300 -4494 300
rect -4322 -300 -4262 300
rect -4090 -300 -4030 300
rect -3858 -300 -3798 300
rect -3626 -300 -3566 300
rect -3394 -300 -3334 300
rect -3162 -300 -3102 300
rect -2930 -300 -2870 300
rect -2698 -300 -2638 300
rect -2466 -300 -2406 300
rect -2234 -300 -2174 300
rect -2002 -300 -1942 300
rect -1770 -300 -1710 300
rect -1538 -300 -1478 300
rect -1306 -300 -1246 300
rect -1074 -300 -1014 300
rect -842 -300 -782 300
rect -610 -300 -550 300
rect -378 -300 -318 300
rect -146 -300 -86 300
rect 86 -300 146 300
rect 318 -300 378 300
rect 550 -300 610 300
rect 782 -300 842 300
rect 1014 -300 1074 300
rect 1246 -300 1306 300
rect 1478 -300 1538 300
rect 1710 -300 1770 300
rect 1942 -300 2002 300
rect 2174 -300 2234 300
rect 2406 -300 2466 300
rect 2638 -300 2698 300
rect 2870 -300 2930 300
rect 3102 -300 3162 300
rect 3334 -300 3394 300
rect 3566 -300 3626 300
rect 3798 -300 3858 300
rect 4030 -300 4090 300
rect 4262 -300 4322 300
rect 4494 -300 4554 300
rect 4726 -300 4786 300
rect 4958 -300 5018 300
rect 5190 -300 5250 300
rect 5422 -300 5482 300
rect 5654 -300 5714 300
<< pdiff >>
rect -5772 288 -5714 300
rect -5772 -288 -5760 288
rect -5726 -288 -5714 288
rect -5772 -300 -5714 -288
rect -5654 288 -5596 300
rect -5654 -288 -5642 288
rect -5608 -288 -5596 288
rect -5654 -300 -5596 -288
rect -5540 288 -5482 300
rect -5540 -288 -5528 288
rect -5494 -288 -5482 288
rect -5540 -300 -5482 -288
rect -5422 288 -5364 300
rect -5422 -288 -5410 288
rect -5376 -288 -5364 288
rect -5422 -300 -5364 -288
rect -5308 288 -5250 300
rect -5308 -288 -5296 288
rect -5262 -288 -5250 288
rect -5308 -300 -5250 -288
rect -5190 288 -5132 300
rect -5190 -288 -5178 288
rect -5144 -288 -5132 288
rect -5190 -300 -5132 -288
rect -5076 288 -5018 300
rect -5076 -288 -5064 288
rect -5030 -288 -5018 288
rect -5076 -300 -5018 -288
rect -4958 288 -4900 300
rect -4958 -288 -4946 288
rect -4912 -288 -4900 288
rect -4958 -300 -4900 -288
rect -4844 288 -4786 300
rect -4844 -288 -4832 288
rect -4798 -288 -4786 288
rect -4844 -300 -4786 -288
rect -4726 288 -4668 300
rect -4726 -288 -4714 288
rect -4680 -288 -4668 288
rect -4726 -300 -4668 -288
rect -4612 288 -4554 300
rect -4612 -288 -4600 288
rect -4566 -288 -4554 288
rect -4612 -300 -4554 -288
rect -4494 288 -4436 300
rect -4494 -288 -4482 288
rect -4448 -288 -4436 288
rect -4494 -300 -4436 -288
rect -4380 288 -4322 300
rect -4380 -288 -4368 288
rect -4334 -288 -4322 288
rect -4380 -300 -4322 -288
rect -4262 288 -4204 300
rect -4262 -288 -4250 288
rect -4216 -288 -4204 288
rect -4262 -300 -4204 -288
rect -4148 288 -4090 300
rect -4148 -288 -4136 288
rect -4102 -288 -4090 288
rect -4148 -300 -4090 -288
rect -4030 288 -3972 300
rect -4030 -288 -4018 288
rect -3984 -288 -3972 288
rect -4030 -300 -3972 -288
rect -3916 288 -3858 300
rect -3916 -288 -3904 288
rect -3870 -288 -3858 288
rect -3916 -300 -3858 -288
rect -3798 288 -3740 300
rect -3798 -288 -3786 288
rect -3752 -288 -3740 288
rect -3798 -300 -3740 -288
rect -3684 288 -3626 300
rect -3684 -288 -3672 288
rect -3638 -288 -3626 288
rect -3684 -300 -3626 -288
rect -3566 288 -3508 300
rect -3566 -288 -3554 288
rect -3520 -288 -3508 288
rect -3566 -300 -3508 -288
rect -3452 288 -3394 300
rect -3452 -288 -3440 288
rect -3406 -288 -3394 288
rect -3452 -300 -3394 -288
rect -3334 288 -3276 300
rect -3334 -288 -3322 288
rect -3288 -288 -3276 288
rect -3334 -300 -3276 -288
rect -3220 288 -3162 300
rect -3220 -288 -3208 288
rect -3174 -288 -3162 288
rect -3220 -300 -3162 -288
rect -3102 288 -3044 300
rect -3102 -288 -3090 288
rect -3056 -288 -3044 288
rect -3102 -300 -3044 -288
rect -2988 288 -2930 300
rect -2988 -288 -2976 288
rect -2942 -288 -2930 288
rect -2988 -300 -2930 -288
rect -2870 288 -2812 300
rect -2870 -288 -2858 288
rect -2824 -288 -2812 288
rect -2870 -300 -2812 -288
rect -2756 288 -2698 300
rect -2756 -288 -2744 288
rect -2710 -288 -2698 288
rect -2756 -300 -2698 -288
rect -2638 288 -2580 300
rect -2638 -288 -2626 288
rect -2592 -288 -2580 288
rect -2638 -300 -2580 -288
rect -2524 288 -2466 300
rect -2524 -288 -2512 288
rect -2478 -288 -2466 288
rect -2524 -300 -2466 -288
rect -2406 288 -2348 300
rect -2406 -288 -2394 288
rect -2360 -288 -2348 288
rect -2406 -300 -2348 -288
rect -2292 288 -2234 300
rect -2292 -288 -2280 288
rect -2246 -288 -2234 288
rect -2292 -300 -2234 -288
rect -2174 288 -2116 300
rect -2174 -288 -2162 288
rect -2128 -288 -2116 288
rect -2174 -300 -2116 -288
rect -2060 288 -2002 300
rect -2060 -288 -2048 288
rect -2014 -288 -2002 288
rect -2060 -300 -2002 -288
rect -1942 288 -1884 300
rect -1942 -288 -1930 288
rect -1896 -288 -1884 288
rect -1942 -300 -1884 -288
rect -1828 288 -1770 300
rect -1828 -288 -1816 288
rect -1782 -288 -1770 288
rect -1828 -300 -1770 -288
rect -1710 288 -1652 300
rect -1710 -288 -1698 288
rect -1664 -288 -1652 288
rect -1710 -300 -1652 -288
rect -1596 288 -1538 300
rect -1596 -288 -1584 288
rect -1550 -288 -1538 288
rect -1596 -300 -1538 -288
rect -1478 288 -1420 300
rect -1478 -288 -1466 288
rect -1432 -288 -1420 288
rect -1478 -300 -1420 -288
rect -1364 288 -1306 300
rect -1364 -288 -1352 288
rect -1318 -288 -1306 288
rect -1364 -300 -1306 -288
rect -1246 288 -1188 300
rect -1246 -288 -1234 288
rect -1200 -288 -1188 288
rect -1246 -300 -1188 -288
rect -1132 288 -1074 300
rect -1132 -288 -1120 288
rect -1086 -288 -1074 288
rect -1132 -300 -1074 -288
rect -1014 288 -956 300
rect -1014 -288 -1002 288
rect -968 -288 -956 288
rect -1014 -300 -956 -288
rect -900 288 -842 300
rect -900 -288 -888 288
rect -854 -288 -842 288
rect -900 -300 -842 -288
rect -782 288 -724 300
rect -782 -288 -770 288
rect -736 -288 -724 288
rect -782 -300 -724 -288
rect -668 288 -610 300
rect -668 -288 -656 288
rect -622 -288 -610 288
rect -668 -300 -610 -288
rect -550 288 -492 300
rect -550 -288 -538 288
rect -504 -288 -492 288
rect -550 -300 -492 -288
rect -436 288 -378 300
rect -436 -288 -424 288
rect -390 -288 -378 288
rect -436 -300 -378 -288
rect -318 288 -260 300
rect -318 -288 -306 288
rect -272 -288 -260 288
rect -318 -300 -260 -288
rect -204 288 -146 300
rect -204 -288 -192 288
rect -158 -288 -146 288
rect -204 -300 -146 -288
rect -86 288 -28 300
rect -86 -288 -74 288
rect -40 -288 -28 288
rect -86 -300 -28 -288
rect 28 288 86 300
rect 28 -288 40 288
rect 74 -288 86 288
rect 28 -300 86 -288
rect 146 288 204 300
rect 146 -288 158 288
rect 192 -288 204 288
rect 146 -300 204 -288
rect 260 288 318 300
rect 260 -288 272 288
rect 306 -288 318 288
rect 260 -300 318 -288
rect 378 288 436 300
rect 378 -288 390 288
rect 424 -288 436 288
rect 378 -300 436 -288
rect 492 288 550 300
rect 492 -288 504 288
rect 538 -288 550 288
rect 492 -300 550 -288
rect 610 288 668 300
rect 610 -288 622 288
rect 656 -288 668 288
rect 610 -300 668 -288
rect 724 288 782 300
rect 724 -288 736 288
rect 770 -288 782 288
rect 724 -300 782 -288
rect 842 288 900 300
rect 842 -288 854 288
rect 888 -288 900 288
rect 842 -300 900 -288
rect 956 288 1014 300
rect 956 -288 968 288
rect 1002 -288 1014 288
rect 956 -300 1014 -288
rect 1074 288 1132 300
rect 1074 -288 1086 288
rect 1120 -288 1132 288
rect 1074 -300 1132 -288
rect 1188 288 1246 300
rect 1188 -288 1200 288
rect 1234 -288 1246 288
rect 1188 -300 1246 -288
rect 1306 288 1364 300
rect 1306 -288 1318 288
rect 1352 -288 1364 288
rect 1306 -300 1364 -288
rect 1420 288 1478 300
rect 1420 -288 1432 288
rect 1466 -288 1478 288
rect 1420 -300 1478 -288
rect 1538 288 1596 300
rect 1538 -288 1550 288
rect 1584 -288 1596 288
rect 1538 -300 1596 -288
rect 1652 288 1710 300
rect 1652 -288 1664 288
rect 1698 -288 1710 288
rect 1652 -300 1710 -288
rect 1770 288 1828 300
rect 1770 -288 1782 288
rect 1816 -288 1828 288
rect 1770 -300 1828 -288
rect 1884 288 1942 300
rect 1884 -288 1896 288
rect 1930 -288 1942 288
rect 1884 -300 1942 -288
rect 2002 288 2060 300
rect 2002 -288 2014 288
rect 2048 -288 2060 288
rect 2002 -300 2060 -288
rect 2116 288 2174 300
rect 2116 -288 2128 288
rect 2162 -288 2174 288
rect 2116 -300 2174 -288
rect 2234 288 2292 300
rect 2234 -288 2246 288
rect 2280 -288 2292 288
rect 2234 -300 2292 -288
rect 2348 288 2406 300
rect 2348 -288 2360 288
rect 2394 -288 2406 288
rect 2348 -300 2406 -288
rect 2466 288 2524 300
rect 2466 -288 2478 288
rect 2512 -288 2524 288
rect 2466 -300 2524 -288
rect 2580 288 2638 300
rect 2580 -288 2592 288
rect 2626 -288 2638 288
rect 2580 -300 2638 -288
rect 2698 288 2756 300
rect 2698 -288 2710 288
rect 2744 -288 2756 288
rect 2698 -300 2756 -288
rect 2812 288 2870 300
rect 2812 -288 2824 288
rect 2858 -288 2870 288
rect 2812 -300 2870 -288
rect 2930 288 2988 300
rect 2930 -288 2942 288
rect 2976 -288 2988 288
rect 2930 -300 2988 -288
rect 3044 288 3102 300
rect 3044 -288 3056 288
rect 3090 -288 3102 288
rect 3044 -300 3102 -288
rect 3162 288 3220 300
rect 3162 -288 3174 288
rect 3208 -288 3220 288
rect 3162 -300 3220 -288
rect 3276 288 3334 300
rect 3276 -288 3288 288
rect 3322 -288 3334 288
rect 3276 -300 3334 -288
rect 3394 288 3452 300
rect 3394 -288 3406 288
rect 3440 -288 3452 288
rect 3394 -300 3452 -288
rect 3508 288 3566 300
rect 3508 -288 3520 288
rect 3554 -288 3566 288
rect 3508 -300 3566 -288
rect 3626 288 3684 300
rect 3626 -288 3638 288
rect 3672 -288 3684 288
rect 3626 -300 3684 -288
rect 3740 288 3798 300
rect 3740 -288 3752 288
rect 3786 -288 3798 288
rect 3740 -300 3798 -288
rect 3858 288 3916 300
rect 3858 -288 3870 288
rect 3904 -288 3916 288
rect 3858 -300 3916 -288
rect 3972 288 4030 300
rect 3972 -288 3984 288
rect 4018 -288 4030 288
rect 3972 -300 4030 -288
rect 4090 288 4148 300
rect 4090 -288 4102 288
rect 4136 -288 4148 288
rect 4090 -300 4148 -288
rect 4204 288 4262 300
rect 4204 -288 4216 288
rect 4250 -288 4262 288
rect 4204 -300 4262 -288
rect 4322 288 4380 300
rect 4322 -288 4334 288
rect 4368 -288 4380 288
rect 4322 -300 4380 -288
rect 4436 288 4494 300
rect 4436 -288 4448 288
rect 4482 -288 4494 288
rect 4436 -300 4494 -288
rect 4554 288 4612 300
rect 4554 -288 4566 288
rect 4600 -288 4612 288
rect 4554 -300 4612 -288
rect 4668 288 4726 300
rect 4668 -288 4680 288
rect 4714 -288 4726 288
rect 4668 -300 4726 -288
rect 4786 288 4844 300
rect 4786 -288 4798 288
rect 4832 -288 4844 288
rect 4786 -300 4844 -288
rect 4900 288 4958 300
rect 4900 -288 4912 288
rect 4946 -288 4958 288
rect 4900 -300 4958 -288
rect 5018 288 5076 300
rect 5018 -288 5030 288
rect 5064 -288 5076 288
rect 5018 -300 5076 -288
rect 5132 288 5190 300
rect 5132 -288 5144 288
rect 5178 -288 5190 288
rect 5132 -300 5190 -288
rect 5250 288 5308 300
rect 5250 -288 5262 288
rect 5296 -288 5308 288
rect 5250 -300 5308 -288
rect 5364 288 5422 300
rect 5364 -288 5376 288
rect 5410 -288 5422 288
rect 5364 -300 5422 -288
rect 5482 288 5540 300
rect 5482 -288 5494 288
rect 5528 -288 5540 288
rect 5482 -300 5540 -288
rect 5596 288 5654 300
rect 5596 -288 5608 288
rect 5642 -288 5654 288
rect 5596 -300 5654 -288
rect 5714 288 5772 300
rect 5714 -288 5726 288
rect 5760 -288 5772 288
rect 5714 -300 5772 -288
<< pdiffc >>
rect -5760 -288 -5726 288
rect -5642 -288 -5608 288
rect -5528 -288 -5494 288
rect -5410 -288 -5376 288
rect -5296 -288 -5262 288
rect -5178 -288 -5144 288
rect -5064 -288 -5030 288
rect -4946 -288 -4912 288
rect -4832 -288 -4798 288
rect -4714 -288 -4680 288
rect -4600 -288 -4566 288
rect -4482 -288 -4448 288
rect -4368 -288 -4334 288
rect -4250 -288 -4216 288
rect -4136 -288 -4102 288
rect -4018 -288 -3984 288
rect -3904 -288 -3870 288
rect -3786 -288 -3752 288
rect -3672 -288 -3638 288
rect -3554 -288 -3520 288
rect -3440 -288 -3406 288
rect -3322 -288 -3288 288
rect -3208 -288 -3174 288
rect -3090 -288 -3056 288
rect -2976 -288 -2942 288
rect -2858 -288 -2824 288
rect -2744 -288 -2710 288
rect -2626 -288 -2592 288
rect -2512 -288 -2478 288
rect -2394 -288 -2360 288
rect -2280 -288 -2246 288
rect -2162 -288 -2128 288
rect -2048 -288 -2014 288
rect -1930 -288 -1896 288
rect -1816 -288 -1782 288
rect -1698 -288 -1664 288
rect -1584 -288 -1550 288
rect -1466 -288 -1432 288
rect -1352 -288 -1318 288
rect -1234 -288 -1200 288
rect -1120 -288 -1086 288
rect -1002 -288 -968 288
rect -888 -288 -854 288
rect -770 -288 -736 288
rect -656 -288 -622 288
rect -538 -288 -504 288
rect -424 -288 -390 288
rect -306 -288 -272 288
rect -192 -288 -158 288
rect -74 -288 -40 288
rect 40 -288 74 288
rect 158 -288 192 288
rect 272 -288 306 288
rect 390 -288 424 288
rect 504 -288 538 288
rect 622 -288 656 288
rect 736 -288 770 288
rect 854 -288 888 288
rect 968 -288 1002 288
rect 1086 -288 1120 288
rect 1200 -288 1234 288
rect 1318 -288 1352 288
rect 1432 -288 1466 288
rect 1550 -288 1584 288
rect 1664 -288 1698 288
rect 1782 -288 1816 288
rect 1896 -288 1930 288
rect 2014 -288 2048 288
rect 2128 -288 2162 288
rect 2246 -288 2280 288
rect 2360 -288 2394 288
rect 2478 -288 2512 288
rect 2592 -288 2626 288
rect 2710 -288 2744 288
rect 2824 -288 2858 288
rect 2942 -288 2976 288
rect 3056 -288 3090 288
rect 3174 -288 3208 288
rect 3288 -288 3322 288
rect 3406 -288 3440 288
rect 3520 -288 3554 288
rect 3638 -288 3672 288
rect 3752 -288 3786 288
rect 3870 -288 3904 288
rect 3984 -288 4018 288
rect 4102 -288 4136 288
rect 4216 -288 4250 288
rect 4334 -288 4368 288
rect 4448 -288 4482 288
rect 4566 -288 4600 288
rect 4680 -288 4714 288
rect 4798 -288 4832 288
rect 4912 -288 4946 288
rect 5030 -288 5064 288
rect 5144 -288 5178 288
rect 5262 -288 5296 288
rect 5376 -288 5410 288
rect 5494 -288 5528 288
rect 5608 -288 5642 288
rect 5726 -288 5760 288
<< nsubdiff >>
rect -5874 449 -5778 483
rect 5778 449 5874 483
rect -5874 387 -5840 449
rect 5840 387 5874 449
rect -5874 -449 -5840 -387
rect 5840 -449 5874 -387
rect -5874 -483 -5778 -449
rect 5778 -483 5874 -449
<< nsubdiffcont >>
rect -5778 449 5778 483
rect -5874 -387 -5840 387
rect 5840 -387 5874 387
rect -5778 -483 5778 -449
<< poly >>
rect -5717 381 -5651 397
rect -5717 347 -5701 381
rect -5667 347 -5651 381
rect -5717 331 -5651 347
rect -5485 381 -5419 397
rect -5485 347 -5469 381
rect -5435 347 -5419 381
rect -5485 331 -5419 347
rect -5253 381 -5187 397
rect -5253 347 -5237 381
rect -5203 347 -5187 381
rect -5253 331 -5187 347
rect -5021 381 -4955 397
rect -5021 347 -5005 381
rect -4971 347 -4955 381
rect -5021 331 -4955 347
rect -4789 381 -4723 397
rect -4789 347 -4773 381
rect -4739 347 -4723 381
rect -4789 331 -4723 347
rect -4557 381 -4491 397
rect -4557 347 -4541 381
rect -4507 347 -4491 381
rect -4557 331 -4491 347
rect -4325 381 -4259 397
rect -4325 347 -4309 381
rect -4275 347 -4259 381
rect -4325 331 -4259 347
rect -4093 381 -4027 397
rect -4093 347 -4077 381
rect -4043 347 -4027 381
rect -4093 331 -4027 347
rect -3861 381 -3795 397
rect -3861 347 -3845 381
rect -3811 347 -3795 381
rect -3861 331 -3795 347
rect -3629 381 -3563 397
rect -3629 347 -3613 381
rect -3579 347 -3563 381
rect -3629 331 -3563 347
rect -3397 381 -3331 397
rect -3397 347 -3381 381
rect -3347 347 -3331 381
rect -3397 331 -3331 347
rect -3165 381 -3099 397
rect -3165 347 -3149 381
rect -3115 347 -3099 381
rect -3165 331 -3099 347
rect -2933 381 -2867 397
rect -2933 347 -2917 381
rect -2883 347 -2867 381
rect -2933 331 -2867 347
rect -2701 381 -2635 397
rect -2701 347 -2685 381
rect -2651 347 -2635 381
rect -2701 331 -2635 347
rect -2469 381 -2403 397
rect -2469 347 -2453 381
rect -2419 347 -2403 381
rect -2469 331 -2403 347
rect -2237 381 -2171 397
rect -2237 347 -2221 381
rect -2187 347 -2171 381
rect -2237 331 -2171 347
rect -2005 381 -1939 397
rect -2005 347 -1989 381
rect -1955 347 -1939 381
rect -2005 331 -1939 347
rect -1773 381 -1707 397
rect -1773 347 -1757 381
rect -1723 347 -1707 381
rect -1773 331 -1707 347
rect -1541 381 -1475 397
rect -1541 347 -1525 381
rect -1491 347 -1475 381
rect -1541 331 -1475 347
rect -1309 381 -1243 397
rect -1309 347 -1293 381
rect -1259 347 -1243 381
rect -1309 331 -1243 347
rect -1077 381 -1011 397
rect -1077 347 -1061 381
rect -1027 347 -1011 381
rect -1077 331 -1011 347
rect -845 381 -779 397
rect -845 347 -829 381
rect -795 347 -779 381
rect -845 331 -779 347
rect -613 381 -547 397
rect -613 347 -597 381
rect -563 347 -547 381
rect -613 331 -547 347
rect -381 381 -315 397
rect -381 347 -365 381
rect -331 347 -315 381
rect -381 331 -315 347
rect -149 381 -83 397
rect -149 347 -133 381
rect -99 347 -83 381
rect -149 331 -83 347
rect 83 381 149 397
rect 83 347 99 381
rect 133 347 149 381
rect 83 331 149 347
rect 315 381 381 397
rect 315 347 331 381
rect 365 347 381 381
rect 315 331 381 347
rect 547 381 613 397
rect 547 347 563 381
rect 597 347 613 381
rect 547 331 613 347
rect 779 381 845 397
rect 779 347 795 381
rect 829 347 845 381
rect 779 331 845 347
rect 1011 381 1077 397
rect 1011 347 1027 381
rect 1061 347 1077 381
rect 1011 331 1077 347
rect 1243 381 1309 397
rect 1243 347 1259 381
rect 1293 347 1309 381
rect 1243 331 1309 347
rect 1475 381 1541 397
rect 1475 347 1491 381
rect 1525 347 1541 381
rect 1475 331 1541 347
rect 1707 381 1773 397
rect 1707 347 1723 381
rect 1757 347 1773 381
rect 1707 331 1773 347
rect 1939 381 2005 397
rect 1939 347 1955 381
rect 1989 347 2005 381
rect 1939 331 2005 347
rect 2171 381 2237 397
rect 2171 347 2187 381
rect 2221 347 2237 381
rect 2171 331 2237 347
rect 2403 381 2469 397
rect 2403 347 2419 381
rect 2453 347 2469 381
rect 2403 331 2469 347
rect 2635 381 2701 397
rect 2635 347 2651 381
rect 2685 347 2701 381
rect 2635 331 2701 347
rect 2867 381 2933 397
rect 2867 347 2883 381
rect 2917 347 2933 381
rect 2867 331 2933 347
rect 3099 381 3165 397
rect 3099 347 3115 381
rect 3149 347 3165 381
rect 3099 331 3165 347
rect 3331 381 3397 397
rect 3331 347 3347 381
rect 3381 347 3397 381
rect 3331 331 3397 347
rect 3563 381 3629 397
rect 3563 347 3579 381
rect 3613 347 3629 381
rect 3563 331 3629 347
rect 3795 381 3861 397
rect 3795 347 3811 381
rect 3845 347 3861 381
rect 3795 331 3861 347
rect 4027 381 4093 397
rect 4027 347 4043 381
rect 4077 347 4093 381
rect 4027 331 4093 347
rect 4259 381 4325 397
rect 4259 347 4275 381
rect 4309 347 4325 381
rect 4259 331 4325 347
rect 4491 381 4557 397
rect 4491 347 4507 381
rect 4541 347 4557 381
rect 4491 331 4557 347
rect 4723 381 4789 397
rect 4723 347 4739 381
rect 4773 347 4789 381
rect 4723 331 4789 347
rect 4955 381 5021 397
rect 4955 347 4971 381
rect 5005 347 5021 381
rect 4955 331 5021 347
rect 5187 381 5253 397
rect 5187 347 5203 381
rect 5237 347 5253 381
rect 5187 331 5253 347
rect 5419 381 5485 397
rect 5419 347 5435 381
rect 5469 347 5485 381
rect 5419 331 5485 347
rect 5651 381 5717 397
rect 5651 347 5667 381
rect 5701 347 5717 381
rect 5651 331 5717 347
rect -5714 300 -5654 331
rect -5482 300 -5422 331
rect -5250 300 -5190 331
rect -5018 300 -4958 331
rect -4786 300 -4726 331
rect -4554 300 -4494 331
rect -4322 300 -4262 331
rect -4090 300 -4030 331
rect -3858 300 -3798 331
rect -3626 300 -3566 331
rect -3394 300 -3334 331
rect -3162 300 -3102 331
rect -2930 300 -2870 331
rect -2698 300 -2638 331
rect -2466 300 -2406 331
rect -2234 300 -2174 331
rect -2002 300 -1942 331
rect -1770 300 -1710 331
rect -1538 300 -1478 331
rect -1306 300 -1246 331
rect -1074 300 -1014 331
rect -842 300 -782 331
rect -610 300 -550 331
rect -378 300 -318 331
rect -146 300 -86 331
rect 86 300 146 331
rect 318 300 378 331
rect 550 300 610 331
rect 782 300 842 331
rect 1014 300 1074 331
rect 1246 300 1306 331
rect 1478 300 1538 331
rect 1710 300 1770 331
rect 1942 300 2002 331
rect 2174 300 2234 331
rect 2406 300 2466 331
rect 2638 300 2698 331
rect 2870 300 2930 331
rect 3102 300 3162 331
rect 3334 300 3394 331
rect 3566 300 3626 331
rect 3798 300 3858 331
rect 4030 300 4090 331
rect 4262 300 4322 331
rect 4494 300 4554 331
rect 4726 300 4786 331
rect 4958 300 5018 331
rect 5190 300 5250 331
rect 5422 300 5482 331
rect 5654 300 5714 331
rect -5714 -331 -5654 -300
rect -5482 -331 -5422 -300
rect -5250 -331 -5190 -300
rect -5018 -331 -4958 -300
rect -4786 -331 -4726 -300
rect -4554 -331 -4494 -300
rect -4322 -331 -4262 -300
rect -4090 -331 -4030 -300
rect -3858 -331 -3798 -300
rect -3626 -331 -3566 -300
rect -3394 -331 -3334 -300
rect -3162 -331 -3102 -300
rect -2930 -331 -2870 -300
rect -2698 -331 -2638 -300
rect -2466 -331 -2406 -300
rect -2234 -331 -2174 -300
rect -2002 -331 -1942 -300
rect -1770 -331 -1710 -300
rect -1538 -331 -1478 -300
rect -1306 -331 -1246 -300
rect -1074 -331 -1014 -300
rect -842 -331 -782 -300
rect -610 -331 -550 -300
rect -378 -331 -318 -300
rect -146 -331 -86 -300
rect 86 -331 146 -300
rect 318 -331 378 -300
rect 550 -331 610 -300
rect 782 -331 842 -300
rect 1014 -331 1074 -300
rect 1246 -331 1306 -300
rect 1478 -331 1538 -300
rect 1710 -331 1770 -300
rect 1942 -331 2002 -300
rect 2174 -331 2234 -300
rect 2406 -331 2466 -300
rect 2638 -331 2698 -300
rect 2870 -331 2930 -300
rect 3102 -331 3162 -300
rect 3334 -331 3394 -300
rect 3566 -331 3626 -300
rect 3798 -331 3858 -300
rect 4030 -331 4090 -300
rect 4262 -331 4322 -300
rect 4494 -331 4554 -300
rect 4726 -331 4786 -300
rect 4958 -331 5018 -300
rect 5190 -331 5250 -300
rect 5422 -331 5482 -300
rect 5654 -331 5714 -300
rect -5717 -347 -5651 -331
rect -5717 -381 -5701 -347
rect -5667 -381 -5651 -347
rect -5717 -397 -5651 -381
rect -5485 -347 -5419 -331
rect -5485 -381 -5469 -347
rect -5435 -381 -5419 -347
rect -5485 -397 -5419 -381
rect -5253 -347 -5187 -331
rect -5253 -381 -5237 -347
rect -5203 -381 -5187 -347
rect -5253 -397 -5187 -381
rect -5021 -347 -4955 -331
rect -5021 -381 -5005 -347
rect -4971 -381 -4955 -347
rect -5021 -397 -4955 -381
rect -4789 -347 -4723 -331
rect -4789 -381 -4773 -347
rect -4739 -381 -4723 -347
rect -4789 -397 -4723 -381
rect -4557 -347 -4491 -331
rect -4557 -381 -4541 -347
rect -4507 -381 -4491 -347
rect -4557 -397 -4491 -381
rect -4325 -347 -4259 -331
rect -4325 -381 -4309 -347
rect -4275 -381 -4259 -347
rect -4325 -397 -4259 -381
rect -4093 -347 -4027 -331
rect -4093 -381 -4077 -347
rect -4043 -381 -4027 -347
rect -4093 -397 -4027 -381
rect -3861 -347 -3795 -331
rect -3861 -381 -3845 -347
rect -3811 -381 -3795 -347
rect -3861 -397 -3795 -381
rect -3629 -347 -3563 -331
rect -3629 -381 -3613 -347
rect -3579 -381 -3563 -347
rect -3629 -397 -3563 -381
rect -3397 -347 -3331 -331
rect -3397 -381 -3381 -347
rect -3347 -381 -3331 -347
rect -3397 -397 -3331 -381
rect -3165 -347 -3099 -331
rect -3165 -381 -3149 -347
rect -3115 -381 -3099 -347
rect -3165 -397 -3099 -381
rect -2933 -347 -2867 -331
rect -2933 -381 -2917 -347
rect -2883 -381 -2867 -347
rect -2933 -397 -2867 -381
rect -2701 -347 -2635 -331
rect -2701 -381 -2685 -347
rect -2651 -381 -2635 -347
rect -2701 -397 -2635 -381
rect -2469 -347 -2403 -331
rect -2469 -381 -2453 -347
rect -2419 -381 -2403 -347
rect -2469 -397 -2403 -381
rect -2237 -347 -2171 -331
rect -2237 -381 -2221 -347
rect -2187 -381 -2171 -347
rect -2237 -397 -2171 -381
rect -2005 -347 -1939 -331
rect -2005 -381 -1989 -347
rect -1955 -381 -1939 -347
rect -2005 -397 -1939 -381
rect -1773 -347 -1707 -331
rect -1773 -381 -1757 -347
rect -1723 -381 -1707 -347
rect -1773 -397 -1707 -381
rect -1541 -347 -1475 -331
rect -1541 -381 -1525 -347
rect -1491 -381 -1475 -347
rect -1541 -397 -1475 -381
rect -1309 -347 -1243 -331
rect -1309 -381 -1293 -347
rect -1259 -381 -1243 -347
rect -1309 -397 -1243 -381
rect -1077 -347 -1011 -331
rect -1077 -381 -1061 -347
rect -1027 -381 -1011 -347
rect -1077 -397 -1011 -381
rect -845 -347 -779 -331
rect -845 -381 -829 -347
rect -795 -381 -779 -347
rect -845 -397 -779 -381
rect -613 -347 -547 -331
rect -613 -381 -597 -347
rect -563 -381 -547 -347
rect -613 -397 -547 -381
rect -381 -347 -315 -331
rect -381 -381 -365 -347
rect -331 -381 -315 -347
rect -381 -397 -315 -381
rect -149 -347 -83 -331
rect -149 -381 -133 -347
rect -99 -381 -83 -347
rect -149 -397 -83 -381
rect 83 -347 149 -331
rect 83 -381 99 -347
rect 133 -381 149 -347
rect 83 -397 149 -381
rect 315 -347 381 -331
rect 315 -381 331 -347
rect 365 -381 381 -347
rect 315 -397 381 -381
rect 547 -347 613 -331
rect 547 -381 563 -347
rect 597 -381 613 -347
rect 547 -397 613 -381
rect 779 -347 845 -331
rect 779 -381 795 -347
rect 829 -381 845 -347
rect 779 -397 845 -381
rect 1011 -347 1077 -331
rect 1011 -381 1027 -347
rect 1061 -381 1077 -347
rect 1011 -397 1077 -381
rect 1243 -347 1309 -331
rect 1243 -381 1259 -347
rect 1293 -381 1309 -347
rect 1243 -397 1309 -381
rect 1475 -347 1541 -331
rect 1475 -381 1491 -347
rect 1525 -381 1541 -347
rect 1475 -397 1541 -381
rect 1707 -347 1773 -331
rect 1707 -381 1723 -347
rect 1757 -381 1773 -347
rect 1707 -397 1773 -381
rect 1939 -347 2005 -331
rect 1939 -381 1955 -347
rect 1989 -381 2005 -347
rect 1939 -397 2005 -381
rect 2171 -347 2237 -331
rect 2171 -381 2187 -347
rect 2221 -381 2237 -347
rect 2171 -397 2237 -381
rect 2403 -347 2469 -331
rect 2403 -381 2419 -347
rect 2453 -381 2469 -347
rect 2403 -397 2469 -381
rect 2635 -347 2701 -331
rect 2635 -381 2651 -347
rect 2685 -381 2701 -347
rect 2635 -397 2701 -381
rect 2867 -347 2933 -331
rect 2867 -381 2883 -347
rect 2917 -381 2933 -347
rect 2867 -397 2933 -381
rect 3099 -347 3165 -331
rect 3099 -381 3115 -347
rect 3149 -381 3165 -347
rect 3099 -397 3165 -381
rect 3331 -347 3397 -331
rect 3331 -381 3347 -347
rect 3381 -381 3397 -347
rect 3331 -397 3397 -381
rect 3563 -347 3629 -331
rect 3563 -381 3579 -347
rect 3613 -381 3629 -347
rect 3563 -397 3629 -381
rect 3795 -347 3861 -331
rect 3795 -381 3811 -347
rect 3845 -381 3861 -347
rect 3795 -397 3861 -381
rect 4027 -347 4093 -331
rect 4027 -381 4043 -347
rect 4077 -381 4093 -347
rect 4027 -397 4093 -381
rect 4259 -347 4325 -331
rect 4259 -381 4275 -347
rect 4309 -381 4325 -347
rect 4259 -397 4325 -381
rect 4491 -347 4557 -331
rect 4491 -381 4507 -347
rect 4541 -381 4557 -347
rect 4491 -397 4557 -381
rect 4723 -347 4789 -331
rect 4723 -381 4739 -347
rect 4773 -381 4789 -347
rect 4723 -397 4789 -381
rect 4955 -347 5021 -331
rect 4955 -381 4971 -347
rect 5005 -381 5021 -347
rect 4955 -397 5021 -381
rect 5187 -347 5253 -331
rect 5187 -381 5203 -347
rect 5237 -381 5253 -347
rect 5187 -397 5253 -381
rect 5419 -347 5485 -331
rect 5419 -381 5435 -347
rect 5469 -381 5485 -347
rect 5419 -397 5485 -381
rect 5651 -347 5717 -331
rect 5651 -381 5667 -347
rect 5701 -381 5717 -347
rect 5651 -397 5717 -381
<< polycont >>
rect -5701 347 -5667 381
rect -5469 347 -5435 381
rect -5237 347 -5203 381
rect -5005 347 -4971 381
rect -4773 347 -4739 381
rect -4541 347 -4507 381
rect -4309 347 -4275 381
rect -4077 347 -4043 381
rect -3845 347 -3811 381
rect -3613 347 -3579 381
rect -3381 347 -3347 381
rect -3149 347 -3115 381
rect -2917 347 -2883 381
rect -2685 347 -2651 381
rect -2453 347 -2419 381
rect -2221 347 -2187 381
rect -1989 347 -1955 381
rect -1757 347 -1723 381
rect -1525 347 -1491 381
rect -1293 347 -1259 381
rect -1061 347 -1027 381
rect -829 347 -795 381
rect -597 347 -563 381
rect -365 347 -331 381
rect -133 347 -99 381
rect 99 347 133 381
rect 331 347 365 381
rect 563 347 597 381
rect 795 347 829 381
rect 1027 347 1061 381
rect 1259 347 1293 381
rect 1491 347 1525 381
rect 1723 347 1757 381
rect 1955 347 1989 381
rect 2187 347 2221 381
rect 2419 347 2453 381
rect 2651 347 2685 381
rect 2883 347 2917 381
rect 3115 347 3149 381
rect 3347 347 3381 381
rect 3579 347 3613 381
rect 3811 347 3845 381
rect 4043 347 4077 381
rect 4275 347 4309 381
rect 4507 347 4541 381
rect 4739 347 4773 381
rect 4971 347 5005 381
rect 5203 347 5237 381
rect 5435 347 5469 381
rect 5667 347 5701 381
rect -5701 -381 -5667 -347
rect -5469 -381 -5435 -347
rect -5237 -381 -5203 -347
rect -5005 -381 -4971 -347
rect -4773 -381 -4739 -347
rect -4541 -381 -4507 -347
rect -4309 -381 -4275 -347
rect -4077 -381 -4043 -347
rect -3845 -381 -3811 -347
rect -3613 -381 -3579 -347
rect -3381 -381 -3347 -347
rect -3149 -381 -3115 -347
rect -2917 -381 -2883 -347
rect -2685 -381 -2651 -347
rect -2453 -381 -2419 -347
rect -2221 -381 -2187 -347
rect -1989 -381 -1955 -347
rect -1757 -381 -1723 -347
rect -1525 -381 -1491 -347
rect -1293 -381 -1259 -347
rect -1061 -381 -1027 -347
rect -829 -381 -795 -347
rect -597 -381 -563 -347
rect -365 -381 -331 -347
rect -133 -381 -99 -347
rect 99 -381 133 -347
rect 331 -381 365 -347
rect 563 -381 597 -347
rect 795 -381 829 -347
rect 1027 -381 1061 -347
rect 1259 -381 1293 -347
rect 1491 -381 1525 -347
rect 1723 -381 1757 -347
rect 1955 -381 1989 -347
rect 2187 -381 2221 -347
rect 2419 -381 2453 -347
rect 2651 -381 2685 -347
rect 2883 -381 2917 -347
rect 3115 -381 3149 -347
rect 3347 -381 3381 -347
rect 3579 -381 3613 -347
rect 3811 -381 3845 -347
rect 4043 -381 4077 -347
rect 4275 -381 4309 -347
rect 4507 -381 4541 -347
rect 4739 -381 4773 -347
rect 4971 -381 5005 -347
rect 5203 -381 5237 -347
rect 5435 -381 5469 -347
rect 5667 -381 5701 -347
<< locali >>
rect -5874 449 -5778 483
rect 5778 449 5874 483
rect -5874 387 -5840 449
rect 5840 387 5874 449
rect -5717 347 -5701 381
rect -5667 347 -5651 381
rect -5485 347 -5469 381
rect -5435 347 -5419 381
rect -5253 347 -5237 381
rect -5203 347 -5187 381
rect -5021 347 -5005 381
rect -4971 347 -4955 381
rect -4789 347 -4773 381
rect -4739 347 -4723 381
rect -4557 347 -4541 381
rect -4507 347 -4491 381
rect -4325 347 -4309 381
rect -4275 347 -4259 381
rect -4093 347 -4077 381
rect -4043 347 -4027 381
rect -3861 347 -3845 381
rect -3811 347 -3795 381
rect -3629 347 -3613 381
rect -3579 347 -3563 381
rect -3397 347 -3381 381
rect -3347 347 -3331 381
rect -3165 347 -3149 381
rect -3115 347 -3099 381
rect -2933 347 -2917 381
rect -2883 347 -2867 381
rect -2701 347 -2685 381
rect -2651 347 -2635 381
rect -2469 347 -2453 381
rect -2419 347 -2403 381
rect -2237 347 -2221 381
rect -2187 347 -2171 381
rect -2005 347 -1989 381
rect -1955 347 -1939 381
rect -1773 347 -1757 381
rect -1723 347 -1707 381
rect -1541 347 -1525 381
rect -1491 347 -1475 381
rect -1309 347 -1293 381
rect -1259 347 -1243 381
rect -1077 347 -1061 381
rect -1027 347 -1011 381
rect -845 347 -829 381
rect -795 347 -779 381
rect -613 347 -597 381
rect -563 347 -547 381
rect -381 347 -365 381
rect -331 347 -315 381
rect -149 347 -133 381
rect -99 347 -83 381
rect 83 347 99 381
rect 133 347 149 381
rect 315 347 331 381
rect 365 347 381 381
rect 547 347 563 381
rect 597 347 613 381
rect 779 347 795 381
rect 829 347 845 381
rect 1011 347 1027 381
rect 1061 347 1077 381
rect 1243 347 1259 381
rect 1293 347 1309 381
rect 1475 347 1491 381
rect 1525 347 1541 381
rect 1707 347 1723 381
rect 1757 347 1773 381
rect 1939 347 1955 381
rect 1989 347 2005 381
rect 2171 347 2187 381
rect 2221 347 2237 381
rect 2403 347 2419 381
rect 2453 347 2469 381
rect 2635 347 2651 381
rect 2685 347 2701 381
rect 2867 347 2883 381
rect 2917 347 2933 381
rect 3099 347 3115 381
rect 3149 347 3165 381
rect 3331 347 3347 381
rect 3381 347 3397 381
rect 3563 347 3579 381
rect 3613 347 3629 381
rect 3795 347 3811 381
rect 3845 347 3861 381
rect 4027 347 4043 381
rect 4077 347 4093 381
rect 4259 347 4275 381
rect 4309 347 4325 381
rect 4491 347 4507 381
rect 4541 347 4557 381
rect 4723 347 4739 381
rect 4773 347 4789 381
rect 4955 347 4971 381
rect 5005 347 5021 381
rect 5187 347 5203 381
rect 5237 347 5253 381
rect 5419 347 5435 381
rect 5469 347 5485 381
rect 5651 347 5667 381
rect 5701 347 5717 381
rect -5760 288 -5726 304
rect -5760 -304 -5726 -288
rect -5642 288 -5608 304
rect -5642 -304 -5608 -288
rect -5528 288 -5494 304
rect -5528 -304 -5494 -288
rect -5410 288 -5376 304
rect -5410 -304 -5376 -288
rect -5296 288 -5262 304
rect -5296 -304 -5262 -288
rect -5178 288 -5144 304
rect -5178 -304 -5144 -288
rect -5064 288 -5030 304
rect -5064 -304 -5030 -288
rect -4946 288 -4912 304
rect -4946 -304 -4912 -288
rect -4832 288 -4798 304
rect -4832 -304 -4798 -288
rect -4714 288 -4680 304
rect -4714 -304 -4680 -288
rect -4600 288 -4566 304
rect -4600 -304 -4566 -288
rect -4482 288 -4448 304
rect -4482 -304 -4448 -288
rect -4368 288 -4334 304
rect -4368 -304 -4334 -288
rect -4250 288 -4216 304
rect -4250 -304 -4216 -288
rect -4136 288 -4102 304
rect -4136 -304 -4102 -288
rect -4018 288 -3984 304
rect -4018 -304 -3984 -288
rect -3904 288 -3870 304
rect -3904 -304 -3870 -288
rect -3786 288 -3752 304
rect -3786 -304 -3752 -288
rect -3672 288 -3638 304
rect -3672 -304 -3638 -288
rect -3554 288 -3520 304
rect -3554 -304 -3520 -288
rect -3440 288 -3406 304
rect -3440 -304 -3406 -288
rect -3322 288 -3288 304
rect -3322 -304 -3288 -288
rect -3208 288 -3174 304
rect -3208 -304 -3174 -288
rect -3090 288 -3056 304
rect -3090 -304 -3056 -288
rect -2976 288 -2942 304
rect -2976 -304 -2942 -288
rect -2858 288 -2824 304
rect -2858 -304 -2824 -288
rect -2744 288 -2710 304
rect -2744 -304 -2710 -288
rect -2626 288 -2592 304
rect -2626 -304 -2592 -288
rect -2512 288 -2478 304
rect -2512 -304 -2478 -288
rect -2394 288 -2360 304
rect -2394 -304 -2360 -288
rect -2280 288 -2246 304
rect -2280 -304 -2246 -288
rect -2162 288 -2128 304
rect -2162 -304 -2128 -288
rect -2048 288 -2014 304
rect -2048 -304 -2014 -288
rect -1930 288 -1896 304
rect -1930 -304 -1896 -288
rect -1816 288 -1782 304
rect -1816 -304 -1782 -288
rect -1698 288 -1664 304
rect -1698 -304 -1664 -288
rect -1584 288 -1550 304
rect -1584 -304 -1550 -288
rect -1466 288 -1432 304
rect -1466 -304 -1432 -288
rect -1352 288 -1318 304
rect -1352 -304 -1318 -288
rect -1234 288 -1200 304
rect -1234 -304 -1200 -288
rect -1120 288 -1086 304
rect -1120 -304 -1086 -288
rect -1002 288 -968 304
rect -1002 -304 -968 -288
rect -888 288 -854 304
rect -888 -304 -854 -288
rect -770 288 -736 304
rect -770 -304 -736 -288
rect -656 288 -622 304
rect -656 -304 -622 -288
rect -538 288 -504 304
rect -538 -304 -504 -288
rect -424 288 -390 304
rect -424 -304 -390 -288
rect -306 288 -272 304
rect -306 -304 -272 -288
rect -192 288 -158 304
rect -192 -304 -158 -288
rect -74 288 -40 304
rect -74 -304 -40 -288
rect 40 288 74 304
rect 40 -304 74 -288
rect 158 288 192 304
rect 158 -304 192 -288
rect 272 288 306 304
rect 272 -304 306 -288
rect 390 288 424 304
rect 390 -304 424 -288
rect 504 288 538 304
rect 504 -304 538 -288
rect 622 288 656 304
rect 622 -304 656 -288
rect 736 288 770 304
rect 736 -304 770 -288
rect 854 288 888 304
rect 854 -304 888 -288
rect 968 288 1002 304
rect 968 -304 1002 -288
rect 1086 288 1120 304
rect 1086 -304 1120 -288
rect 1200 288 1234 304
rect 1200 -304 1234 -288
rect 1318 288 1352 304
rect 1318 -304 1352 -288
rect 1432 288 1466 304
rect 1432 -304 1466 -288
rect 1550 288 1584 304
rect 1550 -304 1584 -288
rect 1664 288 1698 304
rect 1664 -304 1698 -288
rect 1782 288 1816 304
rect 1782 -304 1816 -288
rect 1896 288 1930 304
rect 1896 -304 1930 -288
rect 2014 288 2048 304
rect 2014 -304 2048 -288
rect 2128 288 2162 304
rect 2128 -304 2162 -288
rect 2246 288 2280 304
rect 2246 -304 2280 -288
rect 2360 288 2394 304
rect 2360 -304 2394 -288
rect 2478 288 2512 304
rect 2478 -304 2512 -288
rect 2592 288 2626 304
rect 2592 -304 2626 -288
rect 2710 288 2744 304
rect 2710 -304 2744 -288
rect 2824 288 2858 304
rect 2824 -304 2858 -288
rect 2942 288 2976 304
rect 2942 -304 2976 -288
rect 3056 288 3090 304
rect 3056 -304 3090 -288
rect 3174 288 3208 304
rect 3174 -304 3208 -288
rect 3288 288 3322 304
rect 3288 -304 3322 -288
rect 3406 288 3440 304
rect 3406 -304 3440 -288
rect 3520 288 3554 304
rect 3520 -304 3554 -288
rect 3638 288 3672 304
rect 3638 -304 3672 -288
rect 3752 288 3786 304
rect 3752 -304 3786 -288
rect 3870 288 3904 304
rect 3870 -304 3904 -288
rect 3984 288 4018 304
rect 3984 -304 4018 -288
rect 4102 288 4136 304
rect 4102 -304 4136 -288
rect 4216 288 4250 304
rect 4216 -304 4250 -288
rect 4334 288 4368 304
rect 4334 -304 4368 -288
rect 4448 288 4482 304
rect 4448 -304 4482 -288
rect 4566 288 4600 304
rect 4566 -304 4600 -288
rect 4680 288 4714 304
rect 4680 -304 4714 -288
rect 4798 288 4832 304
rect 4798 -304 4832 -288
rect 4912 288 4946 304
rect 4912 -304 4946 -288
rect 5030 288 5064 304
rect 5030 -304 5064 -288
rect 5144 288 5178 304
rect 5144 -304 5178 -288
rect 5262 288 5296 304
rect 5262 -304 5296 -288
rect 5376 288 5410 304
rect 5376 -304 5410 -288
rect 5494 288 5528 304
rect 5494 -304 5528 -288
rect 5608 288 5642 304
rect 5608 -304 5642 -288
rect 5726 288 5760 304
rect 5726 -304 5760 -288
rect -5717 -381 -5701 -347
rect -5667 -381 -5651 -347
rect -5485 -381 -5469 -347
rect -5435 -381 -5419 -347
rect -5253 -381 -5237 -347
rect -5203 -381 -5187 -347
rect -5021 -381 -5005 -347
rect -4971 -381 -4955 -347
rect -4789 -381 -4773 -347
rect -4739 -381 -4723 -347
rect -4557 -381 -4541 -347
rect -4507 -381 -4491 -347
rect -4325 -381 -4309 -347
rect -4275 -381 -4259 -347
rect -4093 -381 -4077 -347
rect -4043 -381 -4027 -347
rect -3861 -381 -3845 -347
rect -3811 -381 -3795 -347
rect -3629 -381 -3613 -347
rect -3579 -381 -3563 -347
rect -3397 -381 -3381 -347
rect -3347 -381 -3331 -347
rect -3165 -381 -3149 -347
rect -3115 -381 -3099 -347
rect -2933 -381 -2917 -347
rect -2883 -381 -2867 -347
rect -2701 -381 -2685 -347
rect -2651 -381 -2635 -347
rect -2469 -381 -2453 -347
rect -2419 -381 -2403 -347
rect -2237 -381 -2221 -347
rect -2187 -381 -2171 -347
rect -2005 -381 -1989 -347
rect -1955 -381 -1939 -347
rect -1773 -381 -1757 -347
rect -1723 -381 -1707 -347
rect -1541 -381 -1525 -347
rect -1491 -381 -1475 -347
rect -1309 -381 -1293 -347
rect -1259 -381 -1243 -347
rect -1077 -381 -1061 -347
rect -1027 -381 -1011 -347
rect -845 -381 -829 -347
rect -795 -381 -779 -347
rect -613 -381 -597 -347
rect -563 -381 -547 -347
rect -381 -381 -365 -347
rect -331 -381 -315 -347
rect -149 -381 -133 -347
rect -99 -381 -83 -347
rect 83 -381 99 -347
rect 133 -381 149 -347
rect 315 -381 331 -347
rect 365 -381 381 -347
rect 547 -381 563 -347
rect 597 -381 613 -347
rect 779 -381 795 -347
rect 829 -381 845 -347
rect 1011 -381 1027 -347
rect 1061 -381 1077 -347
rect 1243 -381 1259 -347
rect 1293 -381 1309 -347
rect 1475 -381 1491 -347
rect 1525 -381 1541 -347
rect 1707 -381 1723 -347
rect 1757 -381 1773 -347
rect 1939 -381 1955 -347
rect 1989 -381 2005 -347
rect 2171 -381 2187 -347
rect 2221 -381 2237 -347
rect 2403 -381 2419 -347
rect 2453 -381 2469 -347
rect 2635 -381 2651 -347
rect 2685 -381 2701 -347
rect 2867 -381 2883 -347
rect 2917 -381 2933 -347
rect 3099 -381 3115 -347
rect 3149 -381 3165 -347
rect 3331 -381 3347 -347
rect 3381 -381 3397 -347
rect 3563 -381 3579 -347
rect 3613 -381 3629 -347
rect 3795 -381 3811 -347
rect 3845 -381 3861 -347
rect 4027 -381 4043 -347
rect 4077 -381 4093 -347
rect 4259 -381 4275 -347
rect 4309 -381 4325 -347
rect 4491 -381 4507 -347
rect 4541 -381 4557 -347
rect 4723 -381 4739 -347
rect 4773 -381 4789 -347
rect 4955 -381 4971 -347
rect 5005 -381 5021 -347
rect 5187 -381 5203 -347
rect 5237 -381 5253 -347
rect 5419 -381 5435 -347
rect 5469 -381 5485 -347
rect 5651 -381 5667 -347
rect 5701 -381 5717 -347
rect -5874 -449 -5840 -387
rect 5840 -449 5874 -387
rect -5874 -483 -5778 -449
rect 5778 -483 5874 -449
<< viali >>
rect -5701 347 -5667 381
rect -5469 347 -5435 381
rect -5237 347 -5203 381
rect -5005 347 -4971 381
rect -4773 347 -4739 381
rect -4541 347 -4507 381
rect -4309 347 -4275 381
rect -4077 347 -4043 381
rect -3845 347 -3811 381
rect -3613 347 -3579 381
rect -3381 347 -3347 381
rect -3149 347 -3115 381
rect -2917 347 -2883 381
rect -2685 347 -2651 381
rect -2453 347 -2419 381
rect -2221 347 -2187 381
rect -1989 347 -1955 381
rect -1757 347 -1723 381
rect -1525 347 -1491 381
rect -1293 347 -1259 381
rect -1061 347 -1027 381
rect -829 347 -795 381
rect -597 347 -563 381
rect -365 347 -331 381
rect -133 347 -99 381
rect 99 347 133 381
rect 331 347 365 381
rect 563 347 597 381
rect 795 347 829 381
rect 1027 347 1061 381
rect 1259 347 1293 381
rect 1491 347 1525 381
rect 1723 347 1757 381
rect 1955 347 1989 381
rect 2187 347 2221 381
rect 2419 347 2453 381
rect 2651 347 2685 381
rect 2883 347 2917 381
rect 3115 347 3149 381
rect 3347 347 3381 381
rect 3579 347 3613 381
rect 3811 347 3845 381
rect 4043 347 4077 381
rect 4275 347 4309 381
rect 4507 347 4541 381
rect 4739 347 4773 381
rect 4971 347 5005 381
rect 5203 347 5237 381
rect 5435 347 5469 381
rect 5667 347 5701 381
rect -5760 -288 -5726 288
rect -5642 -288 -5608 288
rect -5528 -288 -5494 288
rect -5410 -288 -5376 288
rect -5296 -288 -5262 288
rect -5178 -288 -5144 288
rect -5064 -288 -5030 288
rect -4946 -288 -4912 288
rect -4832 -288 -4798 288
rect -4714 -288 -4680 288
rect -4600 -288 -4566 288
rect -4482 -288 -4448 288
rect -4368 -288 -4334 288
rect -4250 -288 -4216 288
rect -4136 -288 -4102 288
rect -4018 -288 -3984 288
rect -3904 -288 -3870 288
rect -3786 -288 -3752 288
rect -3672 -288 -3638 288
rect -3554 -288 -3520 288
rect -3440 -288 -3406 288
rect -3322 -288 -3288 288
rect -3208 -288 -3174 288
rect -3090 -288 -3056 288
rect -2976 -288 -2942 288
rect -2858 -288 -2824 288
rect -2744 -288 -2710 288
rect -2626 -288 -2592 288
rect -2512 -288 -2478 288
rect -2394 -288 -2360 288
rect -2280 -288 -2246 288
rect -2162 -288 -2128 288
rect -2048 -288 -2014 288
rect -1930 -288 -1896 288
rect -1816 -288 -1782 288
rect -1698 -288 -1664 288
rect -1584 -288 -1550 288
rect -1466 -288 -1432 288
rect -1352 -288 -1318 288
rect -1234 -288 -1200 288
rect -1120 -288 -1086 288
rect -1002 -288 -968 288
rect -888 -288 -854 288
rect -770 -288 -736 288
rect -656 -288 -622 288
rect -538 -288 -504 288
rect -424 -288 -390 288
rect -306 -288 -272 288
rect -192 -288 -158 288
rect -74 -288 -40 288
rect 40 -288 74 288
rect 158 -288 192 288
rect 272 -288 306 288
rect 390 -288 424 288
rect 504 -288 538 288
rect 622 -288 656 288
rect 736 -288 770 288
rect 854 -288 888 288
rect 968 -288 1002 288
rect 1086 -288 1120 288
rect 1200 -288 1234 288
rect 1318 -288 1352 288
rect 1432 -288 1466 288
rect 1550 -288 1584 288
rect 1664 -288 1698 288
rect 1782 -288 1816 288
rect 1896 -288 1930 288
rect 2014 -288 2048 288
rect 2128 -288 2162 288
rect 2246 -288 2280 288
rect 2360 -288 2394 288
rect 2478 -288 2512 288
rect 2592 -288 2626 288
rect 2710 -288 2744 288
rect 2824 -288 2858 288
rect 2942 -288 2976 288
rect 3056 -288 3090 288
rect 3174 -288 3208 288
rect 3288 -288 3322 288
rect 3406 -288 3440 288
rect 3520 -288 3554 288
rect 3638 -288 3672 288
rect 3752 -288 3786 288
rect 3870 -288 3904 288
rect 3984 -288 4018 288
rect 4102 -288 4136 288
rect 4216 -288 4250 288
rect 4334 -288 4368 288
rect 4448 -288 4482 288
rect 4566 -288 4600 288
rect 4680 -288 4714 288
rect 4798 -288 4832 288
rect 4912 -288 4946 288
rect 5030 -288 5064 288
rect 5144 -288 5178 288
rect 5262 -288 5296 288
rect 5376 -288 5410 288
rect 5494 -288 5528 288
rect 5608 -288 5642 288
rect 5726 -288 5760 288
rect -5701 -381 -5667 -347
rect -5469 -381 -5435 -347
rect -5237 -381 -5203 -347
rect -5005 -381 -4971 -347
rect -4773 -381 -4739 -347
rect -4541 -381 -4507 -347
rect -4309 -381 -4275 -347
rect -4077 -381 -4043 -347
rect -3845 -381 -3811 -347
rect -3613 -381 -3579 -347
rect -3381 -381 -3347 -347
rect -3149 -381 -3115 -347
rect -2917 -381 -2883 -347
rect -2685 -381 -2651 -347
rect -2453 -381 -2419 -347
rect -2221 -381 -2187 -347
rect -1989 -381 -1955 -347
rect -1757 -381 -1723 -347
rect -1525 -381 -1491 -347
rect -1293 -381 -1259 -347
rect -1061 -381 -1027 -347
rect -829 -381 -795 -347
rect -597 -381 -563 -347
rect -365 -381 -331 -347
rect -133 -381 -99 -347
rect 99 -381 133 -347
rect 331 -381 365 -347
rect 563 -381 597 -347
rect 795 -381 829 -347
rect 1027 -381 1061 -347
rect 1259 -381 1293 -347
rect 1491 -381 1525 -347
rect 1723 -381 1757 -347
rect 1955 -381 1989 -347
rect 2187 -381 2221 -347
rect 2419 -381 2453 -347
rect 2651 -381 2685 -347
rect 2883 -381 2917 -347
rect 3115 -381 3149 -347
rect 3347 -381 3381 -347
rect 3579 -381 3613 -347
rect 3811 -381 3845 -347
rect 4043 -381 4077 -347
rect 4275 -381 4309 -347
rect 4507 -381 4541 -347
rect 4739 -381 4773 -347
rect 4971 -381 5005 -347
rect 5203 -381 5237 -347
rect 5435 -381 5469 -347
rect 5667 -381 5701 -347
<< metal1 >>
rect -5713 381 -5655 387
rect -5713 347 -5701 381
rect -5667 347 -5655 381
rect -5713 341 -5655 347
rect -5481 381 -5423 387
rect -5481 347 -5469 381
rect -5435 347 -5423 381
rect -5481 341 -5423 347
rect -5249 381 -5191 387
rect -5249 347 -5237 381
rect -5203 347 -5191 381
rect -5249 341 -5191 347
rect -5017 381 -4959 387
rect -5017 347 -5005 381
rect -4971 347 -4959 381
rect -5017 341 -4959 347
rect -4785 381 -4727 387
rect -4785 347 -4773 381
rect -4739 347 -4727 381
rect -4785 341 -4727 347
rect -4553 381 -4495 387
rect -4553 347 -4541 381
rect -4507 347 -4495 381
rect -4553 341 -4495 347
rect -4321 381 -4263 387
rect -4321 347 -4309 381
rect -4275 347 -4263 381
rect -4321 341 -4263 347
rect -4089 381 -4031 387
rect -4089 347 -4077 381
rect -4043 347 -4031 381
rect -4089 341 -4031 347
rect -3857 381 -3799 387
rect -3857 347 -3845 381
rect -3811 347 -3799 381
rect -3857 341 -3799 347
rect -3625 381 -3567 387
rect -3625 347 -3613 381
rect -3579 347 -3567 381
rect -3625 341 -3567 347
rect -3393 381 -3335 387
rect -3393 347 -3381 381
rect -3347 347 -3335 381
rect -3393 341 -3335 347
rect -3161 381 -3103 387
rect -3161 347 -3149 381
rect -3115 347 -3103 381
rect -3161 341 -3103 347
rect -2929 381 -2871 387
rect -2929 347 -2917 381
rect -2883 347 -2871 381
rect -2929 341 -2871 347
rect -2697 381 -2639 387
rect -2697 347 -2685 381
rect -2651 347 -2639 381
rect -2697 341 -2639 347
rect -2465 381 -2407 387
rect -2465 347 -2453 381
rect -2419 347 -2407 381
rect -2465 341 -2407 347
rect -2233 381 -2175 387
rect -2233 347 -2221 381
rect -2187 347 -2175 381
rect -2233 341 -2175 347
rect -2001 381 -1943 387
rect -2001 347 -1989 381
rect -1955 347 -1943 381
rect -2001 341 -1943 347
rect -1769 381 -1711 387
rect -1769 347 -1757 381
rect -1723 347 -1711 381
rect -1769 341 -1711 347
rect -1537 381 -1479 387
rect -1537 347 -1525 381
rect -1491 347 -1479 381
rect -1537 341 -1479 347
rect -1305 381 -1247 387
rect -1305 347 -1293 381
rect -1259 347 -1247 381
rect -1305 341 -1247 347
rect -1073 381 -1015 387
rect -1073 347 -1061 381
rect -1027 347 -1015 381
rect -1073 341 -1015 347
rect -841 381 -783 387
rect -841 347 -829 381
rect -795 347 -783 381
rect -841 341 -783 347
rect -609 381 -551 387
rect -609 347 -597 381
rect -563 347 -551 381
rect -609 341 -551 347
rect -377 381 -319 387
rect -377 347 -365 381
rect -331 347 -319 381
rect -377 341 -319 347
rect -145 381 -87 387
rect -145 347 -133 381
rect -99 347 -87 381
rect -145 341 -87 347
rect 87 381 145 387
rect 87 347 99 381
rect 133 347 145 381
rect 87 341 145 347
rect 319 381 377 387
rect 319 347 331 381
rect 365 347 377 381
rect 319 341 377 347
rect 551 381 609 387
rect 551 347 563 381
rect 597 347 609 381
rect 551 341 609 347
rect 783 381 841 387
rect 783 347 795 381
rect 829 347 841 381
rect 783 341 841 347
rect 1015 381 1073 387
rect 1015 347 1027 381
rect 1061 347 1073 381
rect 1015 341 1073 347
rect 1247 381 1305 387
rect 1247 347 1259 381
rect 1293 347 1305 381
rect 1247 341 1305 347
rect 1479 381 1537 387
rect 1479 347 1491 381
rect 1525 347 1537 381
rect 1479 341 1537 347
rect 1711 381 1769 387
rect 1711 347 1723 381
rect 1757 347 1769 381
rect 1711 341 1769 347
rect 1943 381 2001 387
rect 1943 347 1955 381
rect 1989 347 2001 381
rect 1943 341 2001 347
rect 2175 381 2233 387
rect 2175 347 2187 381
rect 2221 347 2233 381
rect 2175 341 2233 347
rect 2407 381 2465 387
rect 2407 347 2419 381
rect 2453 347 2465 381
rect 2407 341 2465 347
rect 2639 381 2697 387
rect 2639 347 2651 381
rect 2685 347 2697 381
rect 2639 341 2697 347
rect 2871 381 2929 387
rect 2871 347 2883 381
rect 2917 347 2929 381
rect 2871 341 2929 347
rect 3103 381 3161 387
rect 3103 347 3115 381
rect 3149 347 3161 381
rect 3103 341 3161 347
rect 3335 381 3393 387
rect 3335 347 3347 381
rect 3381 347 3393 381
rect 3335 341 3393 347
rect 3567 381 3625 387
rect 3567 347 3579 381
rect 3613 347 3625 381
rect 3567 341 3625 347
rect 3799 381 3857 387
rect 3799 347 3811 381
rect 3845 347 3857 381
rect 3799 341 3857 347
rect 4031 381 4089 387
rect 4031 347 4043 381
rect 4077 347 4089 381
rect 4031 341 4089 347
rect 4263 381 4321 387
rect 4263 347 4275 381
rect 4309 347 4321 381
rect 4263 341 4321 347
rect 4495 381 4553 387
rect 4495 347 4507 381
rect 4541 347 4553 381
rect 4495 341 4553 347
rect 4727 381 4785 387
rect 4727 347 4739 381
rect 4773 347 4785 381
rect 4727 341 4785 347
rect 4959 381 5017 387
rect 4959 347 4971 381
rect 5005 347 5017 381
rect 4959 341 5017 347
rect 5191 381 5249 387
rect 5191 347 5203 381
rect 5237 347 5249 381
rect 5191 341 5249 347
rect 5423 381 5481 387
rect 5423 347 5435 381
rect 5469 347 5481 381
rect 5423 341 5481 347
rect 5655 381 5713 387
rect 5655 347 5667 381
rect 5701 347 5713 381
rect 5655 341 5713 347
rect -5766 288 -5720 300
rect -5766 -288 -5760 288
rect -5726 -288 -5720 288
rect -5766 -300 -5720 -288
rect -5648 288 -5602 300
rect -5648 -288 -5642 288
rect -5608 -288 -5602 288
rect -5648 -300 -5602 -288
rect -5534 288 -5488 300
rect -5534 -288 -5528 288
rect -5494 -288 -5488 288
rect -5534 -300 -5488 -288
rect -5416 288 -5370 300
rect -5416 -288 -5410 288
rect -5376 -288 -5370 288
rect -5416 -300 -5370 -288
rect -5302 288 -5256 300
rect -5302 -288 -5296 288
rect -5262 -288 -5256 288
rect -5302 -300 -5256 -288
rect -5184 288 -5138 300
rect -5184 -288 -5178 288
rect -5144 -288 -5138 288
rect -5184 -300 -5138 -288
rect -5070 288 -5024 300
rect -5070 -288 -5064 288
rect -5030 -288 -5024 288
rect -5070 -300 -5024 -288
rect -4952 288 -4906 300
rect -4952 -288 -4946 288
rect -4912 -288 -4906 288
rect -4952 -300 -4906 -288
rect -4838 288 -4792 300
rect -4838 -288 -4832 288
rect -4798 -288 -4792 288
rect -4838 -300 -4792 -288
rect -4720 288 -4674 300
rect -4720 -288 -4714 288
rect -4680 -288 -4674 288
rect -4720 -300 -4674 -288
rect -4606 288 -4560 300
rect -4606 -288 -4600 288
rect -4566 -288 -4560 288
rect -4606 -300 -4560 -288
rect -4488 288 -4442 300
rect -4488 -288 -4482 288
rect -4448 -288 -4442 288
rect -4488 -300 -4442 -288
rect -4374 288 -4328 300
rect -4374 -288 -4368 288
rect -4334 -288 -4328 288
rect -4374 -300 -4328 -288
rect -4256 288 -4210 300
rect -4256 -288 -4250 288
rect -4216 -288 -4210 288
rect -4256 -300 -4210 -288
rect -4142 288 -4096 300
rect -4142 -288 -4136 288
rect -4102 -288 -4096 288
rect -4142 -300 -4096 -288
rect -4024 288 -3978 300
rect -4024 -288 -4018 288
rect -3984 -288 -3978 288
rect -4024 -300 -3978 -288
rect -3910 288 -3864 300
rect -3910 -288 -3904 288
rect -3870 -288 -3864 288
rect -3910 -300 -3864 -288
rect -3792 288 -3746 300
rect -3792 -288 -3786 288
rect -3752 -288 -3746 288
rect -3792 -300 -3746 -288
rect -3678 288 -3632 300
rect -3678 -288 -3672 288
rect -3638 -288 -3632 288
rect -3678 -300 -3632 -288
rect -3560 288 -3514 300
rect -3560 -288 -3554 288
rect -3520 -288 -3514 288
rect -3560 -300 -3514 -288
rect -3446 288 -3400 300
rect -3446 -288 -3440 288
rect -3406 -288 -3400 288
rect -3446 -300 -3400 -288
rect -3328 288 -3282 300
rect -3328 -288 -3322 288
rect -3288 -288 -3282 288
rect -3328 -300 -3282 -288
rect -3214 288 -3168 300
rect -3214 -288 -3208 288
rect -3174 -288 -3168 288
rect -3214 -300 -3168 -288
rect -3096 288 -3050 300
rect -3096 -288 -3090 288
rect -3056 -288 -3050 288
rect -3096 -300 -3050 -288
rect -2982 288 -2936 300
rect -2982 -288 -2976 288
rect -2942 -288 -2936 288
rect -2982 -300 -2936 -288
rect -2864 288 -2818 300
rect -2864 -288 -2858 288
rect -2824 -288 -2818 288
rect -2864 -300 -2818 -288
rect -2750 288 -2704 300
rect -2750 -288 -2744 288
rect -2710 -288 -2704 288
rect -2750 -300 -2704 -288
rect -2632 288 -2586 300
rect -2632 -288 -2626 288
rect -2592 -288 -2586 288
rect -2632 -300 -2586 -288
rect -2518 288 -2472 300
rect -2518 -288 -2512 288
rect -2478 -288 -2472 288
rect -2518 -300 -2472 -288
rect -2400 288 -2354 300
rect -2400 -288 -2394 288
rect -2360 -288 -2354 288
rect -2400 -300 -2354 -288
rect -2286 288 -2240 300
rect -2286 -288 -2280 288
rect -2246 -288 -2240 288
rect -2286 -300 -2240 -288
rect -2168 288 -2122 300
rect -2168 -288 -2162 288
rect -2128 -288 -2122 288
rect -2168 -300 -2122 -288
rect -2054 288 -2008 300
rect -2054 -288 -2048 288
rect -2014 -288 -2008 288
rect -2054 -300 -2008 -288
rect -1936 288 -1890 300
rect -1936 -288 -1930 288
rect -1896 -288 -1890 288
rect -1936 -300 -1890 -288
rect -1822 288 -1776 300
rect -1822 -288 -1816 288
rect -1782 -288 -1776 288
rect -1822 -300 -1776 -288
rect -1704 288 -1658 300
rect -1704 -288 -1698 288
rect -1664 -288 -1658 288
rect -1704 -300 -1658 -288
rect -1590 288 -1544 300
rect -1590 -288 -1584 288
rect -1550 -288 -1544 288
rect -1590 -300 -1544 -288
rect -1472 288 -1426 300
rect -1472 -288 -1466 288
rect -1432 -288 -1426 288
rect -1472 -300 -1426 -288
rect -1358 288 -1312 300
rect -1358 -288 -1352 288
rect -1318 -288 -1312 288
rect -1358 -300 -1312 -288
rect -1240 288 -1194 300
rect -1240 -288 -1234 288
rect -1200 -288 -1194 288
rect -1240 -300 -1194 -288
rect -1126 288 -1080 300
rect -1126 -288 -1120 288
rect -1086 -288 -1080 288
rect -1126 -300 -1080 -288
rect -1008 288 -962 300
rect -1008 -288 -1002 288
rect -968 -288 -962 288
rect -1008 -300 -962 -288
rect -894 288 -848 300
rect -894 -288 -888 288
rect -854 -288 -848 288
rect -894 -300 -848 -288
rect -776 288 -730 300
rect -776 -288 -770 288
rect -736 -288 -730 288
rect -776 -300 -730 -288
rect -662 288 -616 300
rect -662 -288 -656 288
rect -622 -288 -616 288
rect -662 -300 -616 -288
rect -544 288 -498 300
rect -544 -288 -538 288
rect -504 -288 -498 288
rect -544 -300 -498 -288
rect -430 288 -384 300
rect -430 -288 -424 288
rect -390 -288 -384 288
rect -430 -300 -384 -288
rect -312 288 -266 300
rect -312 -288 -306 288
rect -272 -288 -266 288
rect -312 -300 -266 -288
rect -198 288 -152 300
rect -198 -288 -192 288
rect -158 -288 -152 288
rect -198 -300 -152 -288
rect -80 288 -34 300
rect -80 -288 -74 288
rect -40 -288 -34 288
rect -80 -300 -34 -288
rect 34 288 80 300
rect 34 -288 40 288
rect 74 -288 80 288
rect 34 -300 80 -288
rect 152 288 198 300
rect 152 -288 158 288
rect 192 -288 198 288
rect 152 -300 198 -288
rect 266 288 312 300
rect 266 -288 272 288
rect 306 -288 312 288
rect 266 -300 312 -288
rect 384 288 430 300
rect 384 -288 390 288
rect 424 -288 430 288
rect 384 -300 430 -288
rect 498 288 544 300
rect 498 -288 504 288
rect 538 -288 544 288
rect 498 -300 544 -288
rect 616 288 662 300
rect 616 -288 622 288
rect 656 -288 662 288
rect 616 -300 662 -288
rect 730 288 776 300
rect 730 -288 736 288
rect 770 -288 776 288
rect 730 -300 776 -288
rect 848 288 894 300
rect 848 -288 854 288
rect 888 -288 894 288
rect 848 -300 894 -288
rect 962 288 1008 300
rect 962 -288 968 288
rect 1002 -288 1008 288
rect 962 -300 1008 -288
rect 1080 288 1126 300
rect 1080 -288 1086 288
rect 1120 -288 1126 288
rect 1080 -300 1126 -288
rect 1194 288 1240 300
rect 1194 -288 1200 288
rect 1234 -288 1240 288
rect 1194 -300 1240 -288
rect 1312 288 1358 300
rect 1312 -288 1318 288
rect 1352 -288 1358 288
rect 1312 -300 1358 -288
rect 1426 288 1472 300
rect 1426 -288 1432 288
rect 1466 -288 1472 288
rect 1426 -300 1472 -288
rect 1544 288 1590 300
rect 1544 -288 1550 288
rect 1584 -288 1590 288
rect 1544 -300 1590 -288
rect 1658 288 1704 300
rect 1658 -288 1664 288
rect 1698 -288 1704 288
rect 1658 -300 1704 -288
rect 1776 288 1822 300
rect 1776 -288 1782 288
rect 1816 -288 1822 288
rect 1776 -300 1822 -288
rect 1890 288 1936 300
rect 1890 -288 1896 288
rect 1930 -288 1936 288
rect 1890 -300 1936 -288
rect 2008 288 2054 300
rect 2008 -288 2014 288
rect 2048 -288 2054 288
rect 2008 -300 2054 -288
rect 2122 288 2168 300
rect 2122 -288 2128 288
rect 2162 -288 2168 288
rect 2122 -300 2168 -288
rect 2240 288 2286 300
rect 2240 -288 2246 288
rect 2280 -288 2286 288
rect 2240 -300 2286 -288
rect 2354 288 2400 300
rect 2354 -288 2360 288
rect 2394 -288 2400 288
rect 2354 -300 2400 -288
rect 2472 288 2518 300
rect 2472 -288 2478 288
rect 2512 -288 2518 288
rect 2472 -300 2518 -288
rect 2586 288 2632 300
rect 2586 -288 2592 288
rect 2626 -288 2632 288
rect 2586 -300 2632 -288
rect 2704 288 2750 300
rect 2704 -288 2710 288
rect 2744 -288 2750 288
rect 2704 -300 2750 -288
rect 2818 288 2864 300
rect 2818 -288 2824 288
rect 2858 -288 2864 288
rect 2818 -300 2864 -288
rect 2936 288 2982 300
rect 2936 -288 2942 288
rect 2976 -288 2982 288
rect 2936 -300 2982 -288
rect 3050 288 3096 300
rect 3050 -288 3056 288
rect 3090 -288 3096 288
rect 3050 -300 3096 -288
rect 3168 288 3214 300
rect 3168 -288 3174 288
rect 3208 -288 3214 288
rect 3168 -300 3214 -288
rect 3282 288 3328 300
rect 3282 -288 3288 288
rect 3322 -288 3328 288
rect 3282 -300 3328 -288
rect 3400 288 3446 300
rect 3400 -288 3406 288
rect 3440 -288 3446 288
rect 3400 -300 3446 -288
rect 3514 288 3560 300
rect 3514 -288 3520 288
rect 3554 -288 3560 288
rect 3514 -300 3560 -288
rect 3632 288 3678 300
rect 3632 -288 3638 288
rect 3672 -288 3678 288
rect 3632 -300 3678 -288
rect 3746 288 3792 300
rect 3746 -288 3752 288
rect 3786 -288 3792 288
rect 3746 -300 3792 -288
rect 3864 288 3910 300
rect 3864 -288 3870 288
rect 3904 -288 3910 288
rect 3864 -300 3910 -288
rect 3978 288 4024 300
rect 3978 -288 3984 288
rect 4018 -288 4024 288
rect 3978 -300 4024 -288
rect 4096 288 4142 300
rect 4096 -288 4102 288
rect 4136 -288 4142 288
rect 4096 -300 4142 -288
rect 4210 288 4256 300
rect 4210 -288 4216 288
rect 4250 -288 4256 288
rect 4210 -300 4256 -288
rect 4328 288 4374 300
rect 4328 -288 4334 288
rect 4368 -288 4374 288
rect 4328 -300 4374 -288
rect 4442 288 4488 300
rect 4442 -288 4448 288
rect 4482 -288 4488 288
rect 4442 -300 4488 -288
rect 4560 288 4606 300
rect 4560 -288 4566 288
rect 4600 -288 4606 288
rect 4560 -300 4606 -288
rect 4674 288 4720 300
rect 4674 -288 4680 288
rect 4714 -288 4720 288
rect 4674 -300 4720 -288
rect 4792 288 4838 300
rect 4792 -288 4798 288
rect 4832 -288 4838 288
rect 4792 -300 4838 -288
rect 4906 288 4952 300
rect 4906 -288 4912 288
rect 4946 -288 4952 288
rect 4906 -300 4952 -288
rect 5024 288 5070 300
rect 5024 -288 5030 288
rect 5064 -288 5070 288
rect 5024 -300 5070 -288
rect 5138 288 5184 300
rect 5138 -288 5144 288
rect 5178 -288 5184 288
rect 5138 -300 5184 -288
rect 5256 288 5302 300
rect 5256 -288 5262 288
rect 5296 -288 5302 288
rect 5256 -300 5302 -288
rect 5370 288 5416 300
rect 5370 -288 5376 288
rect 5410 -288 5416 288
rect 5370 -300 5416 -288
rect 5488 288 5534 300
rect 5488 -288 5494 288
rect 5528 -288 5534 288
rect 5488 -300 5534 -288
rect 5602 288 5648 300
rect 5602 -288 5608 288
rect 5642 -288 5648 288
rect 5602 -300 5648 -288
rect 5720 288 5766 300
rect 5720 -288 5726 288
rect 5760 -288 5766 288
rect 5720 -300 5766 -288
rect -5713 -347 -5655 -341
rect -5713 -381 -5701 -347
rect -5667 -381 -5655 -347
rect -5713 -387 -5655 -381
rect -5481 -347 -5423 -341
rect -5481 -381 -5469 -347
rect -5435 -381 -5423 -347
rect -5481 -387 -5423 -381
rect -5249 -347 -5191 -341
rect -5249 -381 -5237 -347
rect -5203 -381 -5191 -347
rect -5249 -387 -5191 -381
rect -5017 -347 -4959 -341
rect -5017 -381 -5005 -347
rect -4971 -381 -4959 -347
rect -5017 -387 -4959 -381
rect -4785 -347 -4727 -341
rect -4785 -381 -4773 -347
rect -4739 -381 -4727 -347
rect -4785 -387 -4727 -381
rect -4553 -347 -4495 -341
rect -4553 -381 -4541 -347
rect -4507 -381 -4495 -347
rect -4553 -387 -4495 -381
rect -4321 -347 -4263 -341
rect -4321 -381 -4309 -347
rect -4275 -381 -4263 -347
rect -4321 -387 -4263 -381
rect -4089 -347 -4031 -341
rect -4089 -381 -4077 -347
rect -4043 -381 -4031 -347
rect -4089 -387 -4031 -381
rect -3857 -347 -3799 -341
rect -3857 -381 -3845 -347
rect -3811 -381 -3799 -347
rect -3857 -387 -3799 -381
rect -3625 -347 -3567 -341
rect -3625 -381 -3613 -347
rect -3579 -381 -3567 -347
rect -3625 -387 -3567 -381
rect -3393 -347 -3335 -341
rect -3393 -381 -3381 -347
rect -3347 -381 -3335 -347
rect -3393 -387 -3335 -381
rect -3161 -347 -3103 -341
rect -3161 -381 -3149 -347
rect -3115 -381 -3103 -347
rect -3161 -387 -3103 -381
rect -2929 -347 -2871 -341
rect -2929 -381 -2917 -347
rect -2883 -381 -2871 -347
rect -2929 -387 -2871 -381
rect -2697 -347 -2639 -341
rect -2697 -381 -2685 -347
rect -2651 -381 -2639 -347
rect -2697 -387 -2639 -381
rect -2465 -347 -2407 -341
rect -2465 -381 -2453 -347
rect -2419 -381 -2407 -347
rect -2465 -387 -2407 -381
rect -2233 -347 -2175 -341
rect -2233 -381 -2221 -347
rect -2187 -381 -2175 -347
rect -2233 -387 -2175 -381
rect -2001 -347 -1943 -341
rect -2001 -381 -1989 -347
rect -1955 -381 -1943 -347
rect -2001 -387 -1943 -381
rect -1769 -347 -1711 -341
rect -1769 -381 -1757 -347
rect -1723 -381 -1711 -347
rect -1769 -387 -1711 -381
rect -1537 -347 -1479 -341
rect -1537 -381 -1525 -347
rect -1491 -381 -1479 -347
rect -1537 -387 -1479 -381
rect -1305 -347 -1247 -341
rect -1305 -381 -1293 -347
rect -1259 -381 -1247 -347
rect -1305 -387 -1247 -381
rect -1073 -347 -1015 -341
rect -1073 -381 -1061 -347
rect -1027 -381 -1015 -347
rect -1073 -387 -1015 -381
rect -841 -347 -783 -341
rect -841 -381 -829 -347
rect -795 -381 -783 -347
rect -841 -387 -783 -381
rect -609 -347 -551 -341
rect -609 -381 -597 -347
rect -563 -381 -551 -347
rect -609 -387 -551 -381
rect -377 -347 -319 -341
rect -377 -381 -365 -347
rect -331 -381 -319 -347
rect -377 -387 -319 -381
rect -145 -347 -87 -341
rect -145 -381 -133 -347
rect -99 -381 -87 -347
rect -145 -387 -87 -381
rect 87 -347 145 -341
rect 87 -381 99 -347
rect 133 -381 145 -347
rect 87 -387 145 -381
rect 319 -347 377 -341
rect 319 -381 331 -347
rect 365 -381 377 -347
rect 319 -387 377 -381
rect 551 -347 609 -341
rect 551 -381 563 -347
rect 597 -381 609 -347
rect 551 -387 609 -381
rect 783 -347 841 -341
rect 783 -381 795 -347
rect 829 -381 841 -347
rect 783 -387 841 -381
rect 1015 -347 1073 -341
rect 1015 -381 1027 -347
rect 1061 -381 1073 -347
rect 1015 -387 1073 -381
rect 1247 -347 1305 -341
rect 1247 -381 1259 -347
rect 1293 -381 1305 -347
rect 1247 -387 1305 -381
rect 1479 -347 1537 -341
rect 1479 -381 1491 -347
rect 1525 -381 1537 -347
rect 1479 -387 1537 -381
rect 1711 -347 1769 -341
rect 1711 -381 1723 -347
rect 1757 -381 1769 -347
rect 1711 -387 1769 -381
rect 1943 -347 2001 -341
rect 1943 -381 1955 -347
rect 1989 -381 2001 -347
rect 1943 -387 2001 -381
rect 2175 -347 2233 -341
rect 2175 -381 2187 -347
rect 2221 -381 2233 -347
rect 2175 -387 2233 -381
rect 2407 -347 2465 -341
rect 2407 -381 2419 -347
rect 2453 -381 2465 -347
rect 2407 -387 2465 -381
rect 2639 -347 2697 -341
rect 2639 -381 2651 -347
rect 2685 -381 2697 -347
rect 2639 -387 2697 -381
rect 2871 -347 2929 -341
rect 2871 -381 2883 -347
rect 2917 -381 2929 -347
rect 2871 -387 2929 -381
rect 3103 -347 3161 -341
rect 3103 -381 3115 -347
rect 3149 -381 3161 -347
rect 3103 -387 3161 -381
rect 3335 -347 3393 -341
rect 3335 -381 3347 -347
rect 3381 -381 3393 -347
rect 3335 -387 3393 -381
rect 3567 -347 3625 -341
rect 3567 -381 3579 -347
rect 3613 -381 3625 -347
rect 3567 -387 3625 -381
rect 3799 -347 3857 -341
rect 3799 -381 3811 -347
rect 3845 -381 3857 -347
rect 3799 -387 3857 -381
rect 4031 -347 4089 -341
rect 4031 -381 4043 -347
rect 4077 -381 4089 -347
rect 4031 -387 4089 -381
rect 4263 -347 4321 -341
rect 4263 -381 4275 -347
rect 4309 -381 4321 -347
rect 4263 -387 4321 -381
rect 4495 -347 4553 -341
rect 4495 -381 4507 -347
rect 4541 -381 4553 -347
rect 4495 -387 4553 -381
rect 4727 -347 4785 -341
rect 4727 -381 4739 -347
rect 4773 -381 4785 -347
rect 4727 -387 4785 -381
rect 4959 -347 5017 -341
rect 4959 -381 4971 -347
rect 5005 -381 5017 -347
rect 4959 -387 5017 -381
rect 5191 -347 5249 -341
rect 5191 -381 5203 -347
rect 5237 -381 5249 -347
rect 5191 -387 5249 -381
rect 5423 -347 5481 -341
rect 5423 -381 5435 -347
rect 5469 -381 5481 -347
rect 5423 -387 5481 -381
rect 5655 -347 5713 -341
rect 5655 -381 5667 -347
rect 5701 -381 5713 -347
rect 5655 -387 5713 -381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -5857 -466 5857 466
string parameters w 3 l 0.3 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
