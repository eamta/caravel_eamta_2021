magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 2116 2223 2232 2226
rect 3590 2223 3706 2226
rect 5064 2223 5180 2226
rect 6538 2223 6654 2226
rect 8012 2223 8128 2226
rect 9486 2223 9602 2226
rect 2126 2221 2192 2223
rect 3600 2221 3666 2223
rect 5074 2221 5140 2223
rect 6548 2221 6614 2223
rect 8022 2221 8088 2223
rect 9496 2221 9562 2223
rect 2088 2195 2204 2198
rect 3562 2195 3678 2198
rect 5036 2195 5152 2198
rect 6510 2195 6626 2198
rect 7984 2195 8100 2198
rect 9458 2195 9574 2198
rect 2098 2193 2204 2195
rect 3572 2193 3678 2195
rect 5046 2193 5152 2195
rect 6520 2193 6626 2195
rect 7994 2193 8100 2195
rect 9468 2193 9574 2195
rect 190 2133 210 2141
rect 1664 2133 1684 2141
rect 3138 2133 3158 2141
rect 4612 2133 4632 2141
rect 6086 2133 6106 2141
rect 7560 2133 7580 2141
rect 9034 2133 9054 2141
rect 668 1970 675 2075
rect 696 1983 703 2047
rect 10848 1998 10987 2004
rect 2142 1970 2149 1998
rect 2170 1983 2177 1998
rect 3616 1970 3623 1998
rect 3644 1983 3651 1998
rect 5090 1970 5097 1998
rect 5118 1983 5125 1998
rect 6564 1970 6571 1998
rect 6592 1983 6599 1998
rect 8038 1970 8045 1998
rect 8066 1983 8073 1998
rect 9512 1970 9519 1998
rect 9540 1983 9547 1998
rect 10851 1970 10959 1976
rect 36 1831 70 1841
rect 352 1831 386 1841
rect 36 1823 386 1831
rect 1510 1831 1544 1841
rect 1826 1831 1860 1841
rect 1510 1823 1860 1831
rect 2984 1831 3018 1841
rect 3300 1831 3334 1841
rect 2984 1823 3334 1831
rect 4458 1831 4492 1841
rect 4774 1831 4808 1841
rect 4458 1823 4808 1831
rect 5932 1831 5966 1841
rect 6248 1831 6282 1841
rect 5932 1823 6282 1831
rect 7406 1831 7440 1841
rect 7722 1831 7756 1841
rect 7406 1823 7756 1831
rect 8880 1831 8914 1841
rect 9196 1831 9230 1841
rect 8880 1823 9230 1831
rect 0 1761 422 1823
rect 1474 1761 1896 1823
rect 2948 1761 3370 1823
rect 4422 1761 4844 1823
rect 5896 1761 6318 1823
rect 7370 1761 7792 1823
rect 8844 1761 9266 1823
rect 11024 1766 11048 1798
rect 11052 1794 11076 1826
rect 2182 1598 2204 1620
rect 3656 1598 3678 1620
rect 5130 1598 5152 1620
rect 6604 1598 6626 1620
rect 8078 1598 8100 1620
rect 9552 1598 9574 1620
rect 2182 1570 2198 1592
rect 3656 1570 3672 1592
rect 5130 1570 5146 1592
rect 6604 1570 6620 1592
rect 8078 1570 8094 1592
rect 9552 1570 9568 1592
rect 194 1355 228 1389
rect 1511 1382 1544 1400
rect 1668 1382 1702 1389
rect 1932 1382 1966 1400
rect 2034 1382 2072 1399
rect 2246 1382 2284 1399
rect 2985 1382 3018 1400
rect 3142 1382 3176 1389
rect 3406 1382 3440 1400
rect 3508 1382 3546 1399
rect 3720 1382 3758 1399
rect 4459 1382 4492 1400
rect 4616 1382 4650 1389
rect 4880 1382 4914 1400
rect 4982 1382 5020 1399
rect 5194 1382 5232 1399
rect 5933 1382 5966 1400
rect 6090 1382 6124 1389
rect 6354 1382 6388 1400
rect 6456 1382 6494 1399
rect 6668 1382 6706 1399
rect 7407 1382 7440 1400
rect 7564 1382 7598 1389
rect 7828 1382 7862 1400
rect 7930 1382 7968 1399
rect 8142 1382 8180 1399
rect 8881 1382 8914 1400
rect 9038 1382 9072 1389
rect 9302 1382 9336 1400
rect 9404 1382 9442 1399
rect 9616 1382 9654 1399
rect 1511 1346 2374 1382
rect 2985 1346 3848 1382
rect 4459 1346 5322 1382
rect 5933 1346 6796 1382
rect 7407 1346 8270 1382
rect 8881 1346 9744 1382
rect 70 1320 352 1321
rect 1162 1301 1190 1327
rect 1232 1301 1298 1327
rect 1404 1295 1438 1327
rect 1507 1320 1510 1327
rect 1529 1311 2374 1346
rect 1196 1287 1332 1293
rect 70 1286 352 1287
rect 132 1227 290 1286
rect 1196 1276 1404 1287
rect 1473 1286 1510 1293
rect 791 1259 1404 1276
rect 1529 1276 2386 1311
rect 2636 1301 2664 1327
rect 2706 1301 2772 1327
rect 2878 1295 2912 1327
rect 2981 1320 2984 1327
rect 3003 1311 3848 1346
rect 2670 1287 2806 1293
rect 2670 1276 2878 1287
rect 2947 1286 2984 1293
rect 1529 1259 2878 1276
rect 3003 1276 3860 1311
rect 4110 1301 4138 1327
rect 4180 1301 4246 1327
rect 4352 1295 4386 1327
rect 4455 1320 4458 1327
rect 4477 1311 5322 1346
rect 4144 1287 4280 1293
rect 4144 1276 4352 1287
rect 4421 1286 4458 1293
rect 3003 1259 4352 1276
rect 4477 1276 5334 1311
rect 5584 1301 5612 1327
rect 5654 1301 5720 1327
rect 5826 1295 5860 1327
rect 5929 1320 5932 1327
rect 5951 1311 6796 1346
rect 5618 1287 5754 1293
rect 5618 1276 5826 1287
rect 5895 1286 5932 1293
rect 4477 1259 5826 1276
rect 5951 1276 6808 1311
rect 7058 1301 7086 1327
rect 7128 1301 7194 1327
rect 7300 1295 7334 1327
rect 7403 1320 7406 1327
rect 7425 1311 8270 1346
rect 7092 1287 7228 1293
rect 7092 1276 7300 1287
rect 7369 1286 7406 1293
rect 5951 1259 7300 1276
rect 7425 1276 8282 1311
rect 8532 1301 8560 1327
rect 8602 1301 8668 1327
rect 8774 1295 8808 1327
rect 8877 1320 8880 1327
rect 8899 1311 9744 1346
rect 8566 1287 8702 1293
rect 8566 1276 8774 1287
rect 8843 1286 8880 1293
rect 7425 1259 8774 1276
rect 8899 1276 9756 1311
rect 10006 1301 10034 1327
rect 10076 1301 10142 1327
rect 10248 1295 10282 1327
rect 10040 1287 10176 1293
rect 10040 1276 10248 1287
rect 8899 1259 10248 1276
rect 458 1233 492 1241
rect 791 1233 1230 1259
rect 1529 1233 2704 1259
rect 3003 1233 4178 1259
rect 4477 1233 5652 1259
rect 5951 1233 7126 1259
rect 7425 1233 8600 1259
rect 8899 1233 10074 1259
rect 458 1199 1213 1233
rect 1230 1229 1404 1233
rect 1230 1225 1426 1229
rect 1304 1199 1438 1225
rect 1529 1199 2687 1233
rect 2704 1229 2878 1233
rect 2704 1225 2900 1229
rect 2778 1199 2912 1225
rect 3003 1199 4161 1233
rect 4178 1229 4352 1233
rect 4178 1225 4374 1229
rect 4252 1199 4386 1225
rect 4477 1199 5635 1233
rect 5652 1229 5826 1233
rect 5652 1225 5848 1229
rect 5726 1199 5860 1225
rect 5951 1199 7109 1233
rect 7126 1229 7300 1233
rect 7126 1225 7322 1229
rect 7200 1199 7334 1225
rect 7425 1199 8583 1233
rect 8600 1229 8774 1233
rect 8600 1225 8796 1229
rect 8674 1199 8808 1225
rect 8899 1199 10057 1233
rect 10074 1229 10248 1233
rect 10074 1225 10270 1229
rect 10148 1199 10282 1225
rect 791 1187 1230 1199
rect 458 1165 1230 1187
rect 1338 1165 1404 1191
rect 791 1163 1230 1165
rect 604 1085 662 1091
rect 604 1051 616 1085
rect 604 1045 662 1051
rect 791 704 861 1163
rect 973 806 1031 812
rect 973 772 985 806
rect 973 766 1031 772
rect 791 670 862 704
rect 1160 670 1230 1163
rect 1529 1163 2704 1199
rect 2812 1165 2878 1191
rect 1276 1130 1466 1138
rect 1304 1102 1350 1110
rect 1392 1102 1438 1110
rect 1529 810 1599 1163
rect 1896 1161 2336 1163
rect 1896 921 2337 1161
rect 1711 912 1769 918
rect 1711 878 1723 912
rect 1711 872 1769 878
rect 1896 869 2336 921
rect 1896 851 2337 869
rect 1529 776 1600 810
rect 1896 789 2373 851
rect 1896 776 1966 789
rect 1529 740 1582 776
rect 1896 740 1951 776
rect 791 634 844 670
rect 1160 634 1213 670
rect 1342 619 1400 625
rect 1342 585 1354 619
rect 1342 579 1400 585
rect 1732 544 1751 546
rect 604 513 662 519
rect 604 479 616 513
rect 604 473 662 479
rect 1953 411 1966 776
rect 1987 781 2020 789
rect 2034 781 2180 789
rect 2248 781 2373 789
rect 1987 522 2021 781
rect 2034 670 2075 781
rect 2111 729 2134 747
rect 2179 744 2180 760
rect 2165 729 2180 744
rect 2111 713 2180 729
rect 2129 679 2202 713
rect 2265 686 2373 781
rect 2447 806 2505 812
rect 2447 772 2459 806
rect 2447 766 2505 772
rect 2034 660 2080 670
rect 2129 663 2180 679
rect 2034 560 2086 660
rect 2134 648 2180 663
rect 2101 632 2114 636
rect 2095 631 2114 632
rect 2134 632 2177 648
rect 2189 632 2202 636
rect 2092 620 2122 631
rect 2134 620 2174 632
rect 2095 572 2174 620
rect 2095 560 2135 572
rect 2155 560 2174 572
rect 2183 620 2202 632
rect 2214 632 2223 636
rect 2248 634 2373 686
rect 2634 670 2704 1163
rect 3003 1163 4178 1199
rect 4286 1165 4352 1191
rect 2750 1130 2940 1138
rect 2778 1102 2824 1110
rect 2866 1102 2912 1110
rect 3003 810 3073 1163
rect 3370 1161 3810 1163
rect 3370 921 3811 1161
rect 3185 912 3243 918
rect 3185 878 3197 912
rect 3185 872 3243 878
rect 3370 869 3810 921
rect 3370 851 3811 869
rect 3003 776 3074 810
rect 3370 789 3847 851
rect 3370 776 3440 789
rect 3003 740 3056 776
rect 3370 740 3425 776
rect 2634 634 2687 670
rect 2046 556 2055 560
rect 2067 556 2080 560
rect 2092 547 2148 560
rect 2155 556 2168 560
rect 2092 544 2158 547
rect 1987 445 2020 522
rect 2089 479 2158 544
rect 2183 534 2206 620
rect 2183 532 2202 534
rect 2189 522 2202 532
rect 2089 464 2147 479
rect 2214 465 2235 632
rect 2195 464 2235 465
rect 2248 464 2282 634
rect 2087 463 2140 464
rect 2147 463 2177 464
rect 2214 460 2223 464
rect 1987 411 2021 445
rect 2248 426 2257 464
rect 2145 411 2179 417
rect 2028 377 2055 411
rect 2118 400 2206 411
rect 2129 388 2195 400
rect 2269 388 2282 464
rect 2118 377 2206 388
rect 2303 377 2336 634
rect 2816 619 2874 625
rect 2816 585 2828 619
rect 2816 579 2874 585
rect 3393 493 3409 569
rect 3427 548 3440 776
rect 3461 781 3494 789
rect 3508 781 3654 789
rect 3722 781 3847 789
rect 3421 546 3446 548
rect 3421 520 3449 546
rect 3461 522 3495 781
rect 3508 670 3549 781
rect 3585 729 3608 747
rect 3653 744 3654 760
rect 3639 729 3654 744
rect 3585 713 3654 729
rect 3603 679 3676 713
rect 3739 686 3847 781
rect 3921 806 3979 812
rect 3921 772 3933 806
rect 3921 766 3979 772
rect 3508 660 3554 670
rect 3603 663 3654 679
rect 3508 560 3560 660
rect 3608 648 3654 663
rect 3575 632 3588 636
rect 3569 631 3588 632
rect 3608 632 3651 648
rect 3663 632 3676 636
rect 3566 620 3596 631
rect 3608 620 3648 632
rect 3569 572 3648 620
rect 3569 560 3609 572
rect 3629 560 3648 572
rect 3657 620 3676 632
rect 3688 632 3697 636
rect 3722 634 3847 686
rect 4108 670 4178 1163
rect 4477 1163 5652 1199
rect 5760 1165 5826 1191
rect 4224 1130 4414 1138
rect 4252 1102 4298 1110
rect 4340 1102 4386 1110
rect 4477 810 4547 1163
rect 4844 1161 5284 1163
rect 4844 921 5285 1161
rect 4659 912 4717 918
rect 4659 878 4671 912
rect 4659 872 4717 878
rect 4844 869 5284 921
rect 4844 851 5285 869
rect 4477 776 4548 810
rect 4844 789 5321 851
rect 4844 776 4914 789
rect 4477 740 4530 776
rect 4844 740 4899 776
rect 4108 634 4161 670
rect 3520 556 3529 560
rect 3541 556 3554 560
rect 3566 547 3622 560
rect 3629 556 3642 560
rect 3566 544 3632 547
rect 3427 411 3440 520
rect 3461 445 3494 522
rect 3563 479 3632 544
rect 3657 534 3680 620
rect 3657 532 3676 534
rect 3663 522 3676 532
rect 3563 464 3621 479
rect 3688 465 3709 632
rect 3669 464 3709 465
rect 3722 464 3756 634
rect 3561 463 3614 464
rect 3621 463 3651 464
rect 3688 460 3697 464
rect 3461 411 3495 445
rect 3722 426 3731 464
rect 3619 411 3653 417
rect 3502 377 3529 411
rect 3592 400 3680 411
rect 3603 388 3669 400
rect 3743 388 3756 464
rect 3592 377 3680 388
rect 3777 377 3810 634
rect 4290 619 4348 625
rect 4290 585 4302 619
rect 4290 579 4348 585
rect 4901 411 4914 776
rect 4935 781 4968 789
rect 4982 781 5128 789
rect 5196 781 5321 789
rect 4935 522 4969 781
rect 4982 670 5023 781
rect 5059 729 5082 747
rect 5127 744 5128 760
rect 5113 729 5128 744
rect 5059 713 5128 729
rect 5077 679 5150 713
rect 5213 686 5321 781
rect 5395 806 5453 812
rect 5395 772 5407 806
rect 5395 766 5453 772
rect 4982 660 5028 670
rect 5077 663 5128 679
rect 4982 560 5034 660
rect 5082 648 5128 663
rect 5049 632 5062 636
rect 5043 631 5062 632
rect 5082 632 5125 648
rect 5137 632 5150 636
rect 5040 620 5070 631
rect 5082 620 5122 632
rect 5043 572 5122 620
rect 5043 569 5083 572
rect 5043 560 5096 569
rect 4994 556 5003 560
rect 5015 556 5028 560
rect 5040 547 5096 560
rect 5103 560 5122 572
rect 5131 620 5150 632
rect 5162 632 5171 636
rect 5196 634 5321 686
rect 5582 670 5652 1163
rect 5951 1163 7126 1199
rect 7234 1165 7300 1191
rect 5698 1130 5888 1138
rect 5726 1102 5772 1110
rect 5814 1102 5860 1110
rect 5951 810 6021 1163
rect 6318 1161 6758 1163
rect 6318 921 6759 1161
rect 6133 912 6191 918
rect 6133 878 6145 912
rect 6133 872 6191 878
rect 6318 869 6758 921
rect 6318 851 6759 869
rect 5951 776 6022 810
rect 6318 789 6795 851
rect 6318 776 6388 789
rect 5951 740 6004 776
rect 6318 740 6373 776
rect 5582 634 5635 670
rect 5103 556 5116 560
rect 5131 547 5154 620
rect 5040 544 5154 547
rect 5037 534 5154 544
rect 5037 532 5150 534
rect 4935 445 4968 522
rect 5037 519 5134 532
rect 5137 522 5150 532
rect 5037 479 5106 519
rect 5037 464 5095 479
rect 5162 465 5183 632
rect 5143 464 5183 465
rect 5196 464 5230 634
rect 5035 463 5088 464
rect 5095 463 5125 464
rect 5162 460 5171 464
rect 4935 411 4969 445
rect 5093 411 5127 445
rect 5196 426 5205 464
rect 4976 377 5003 411
rect 5066 400 5161 411
rect 5077 388 5161 400
rect 5217 388 5230 464
rect 5066 383 5161 388
rect 5066 377 5154 383
rect 5251 377 5284 634
rect 5764 619 5822 625
rect 5764 585 5776 619
rect 5764 579 5822 585
rect 6375 411 6388 776
rect 6409 781 6442 789
rect 6456 781 6602 789
rect 6670 781 6795 789
rect 6409 522 6443 781
rect 6456 670 6497 781
rect 6533 729 6556 747
rect 6601 744 6602 760
rect 6587 729 6602 744
rect 6533 713 6602 729
rect 6551 679 6624 713
rect 6687 686 6795 781
rect 6869 806 6927 812
rect 6869 772 6881 806
rect 6869 766 6927 772
rect 6456 660 6502 670
rect 6551 663 6602 679
rect 6456 560 6508 660
rect 6556 648 6602 663
rect 6523 632 6536 636
rect 6517 631 6536 632
rect 6556 632 6599 648
rect 6611 632 6624 636
rect 6514 620 6544 631
rect 6556 620 6596 632
rect 6517 572 6596 620
rect 6517 560 6557 572
rect 6577 560 6596 572
rect 6605 620 6624 632
rect 6636 632 6645 636
rect 6670 634 6795 686
rect 7056 670 7126 1163
rect 7425 1163 8600 1199
rect 8708 1165 8774 1191
rect 7172 1130 7362 1138
rect 7200 1102 7246 1110
rect 7288 1102 7334 1110
rect 7425 810 7495 1163
rect 7792 1161 8232 1163
rect 7792 921 8233 1161
rect 7607 912 7665 918
rect 7607 878 7619 912
rect 7607 872 7665 878
rect 7792 869 8232 921
rect 7792 851 8233 869
rect 7425 776 7496 810
rect 7792 789 8269 851
rect 7792 776 7862 789
rect 7425 740 7478 776
rect 7792 740 7847 776
rect 7056 634 7109 670
rect 6468 556 6477 560
rect 6489 556 6502 560
rect 6514 547 6570 560
rect 6577 556 6590 560
rect 6514 544 6580 547
rect 6409 445 6442 522
rect 6511 479 6580 544
rect 6605 534 6628 620
rect 6605 532 6624 534
rect 6611 522 6624 532
rect 6511 464 6569 479
rect 6636 465 6657 632
rect 6617 464 6657 465
rect 6670 464 6704 634
rect 6509 463 6562 464
rect 6569 463 6599 464
rect 6636 460 6645 464
rect 6409 411 6443 445
rect 6670 426 6679 464
rect 6567 411 6601 417
rect 6450 377 6477 411
rect 6540 400 6628 411
rect 6551 388 6617 400
rect 6691 388 6704 464
rect 6540 377 6628 388
rect 6725 377 6758 634
rect 7238 619 7296 625
rect 7238 585 7250 619
rect 7238 579 7296 585
rect 6762 493 6786 569
rect 6790 546 6815 548
rect 6790 520 6818 546
rect 7849 411 7862 776
rect 7883 781 7916 789
rect 7930 781 8076 789
rect 8144 781 8269 789
rect 7883 522 7917 781
rect 7930 670 7971 781
rect 8007 729 8030 747
rect 8075 744 8076 760
rect 8061 729 8076 744
rect 8007 713 8076 729
rect 8025 679 8098 713
rect 8161 686 8269 781
rect 8343 806 8401 812
rect 8343 772 8355 806
rect 8343 766 8401 772
rect 7930 660 7976 670
rect 8025 663 8076 679
rect 7930 560 7982 660
rect 8030 648 8076 663
rect 7997 632 8010 636
rect 7991 631 8010 632
rect 8030 632 8073 648
rect 8085 632 8098 636
rect 7988 620 8018 631
rect 8030 620 8070 632
rect 7991 572 8070 620
rect 7991 560 8031 572
rect 8051 560 8070 572
rect 8079 620 8098 632
rect 8110 632 8119 636
rect 8144 634 8269 686
rect 8530 670 8600 1163
rect 8899 1163 10074 1199
rect 10186 1191 10244 1197
rect 10182 1165 10248 1191
rect 8646 1130 8836 1138
rect 8674 1102 8720 1110
rect 8762 1102 8808 1110
rect 8899 810 8969 1163
rect 9266 1161 9706 1163
rect 9266 921 9707 1161
rect 9817 1138 9875 1144
rect 9817 1104 9829 1138
rect 9817 1098 9875 1104
rect 9081 912 9139 918
rect 9081 878 9093 912
rect 9081 872 9139 878
rect 9266 869 9706 921
rect 9266 851 9707 869
rect 8899 776 8970 810
rect 9266 789 9743 851
rect 9266 776 9336 789
rect 8899 740 8952 776
rect 9266 740 9321 776
rect 8530 634 8583 670
rect 7942 556 7951 560
rect 7963 556 7976 560
rect 7988 547 8044 560
rect 8051 556 8064 560
rect 7988 544 8054 547
rect 7883 445 7916 522
rect 7985 479 8054 544
rect 8079 534 8102 620
rect 8079 532 8098 534
rect 8085 522 8098 532
rect 7985 464 8043 479
rect 8110 465 8131 632
rect 8091 464 8131 465
rect 8144 464 8178 634
rect 7983 463 8036 464
rect 8043 463 8073 464
rect 8110 460 8119 464
rect 7883 411 7917 445
rect 8144 426 8153 464
rect 8041 411 8075 417
rect 7924 377 7951 411
rect 8014 400 8102 411
rect 8025 388 8091 400
rect 8165 388 8178 464
rect 8014 377 8102 388
rect 8199 377 8232 634
rect 8712 619 8770 625
rect 8712 585 8724 619
rect 8712 579 8770 585
rect 8453 493 8474 568
rect 8481 540 8506 542
rect 8481 514 8509 540
rect 9323 411 9336 776
rect 9357 781 9390 789
rect 9404 781 9550 789
rect 9618 781 9743 789
rect 9357 522 9391 781
rect 9404 670 9445 781
rect 9481 729 9504 747
rect 9549 744 9550 760
rect 9535 729 9550 744
rect 9481 713 9550 729
rect 9499 679 9572 713
rect 9635 686 9743 781
rect 9817 806 9875 812
rect 9817 772 9829 806
rect 9817 766 9875 772
rect 9404 660 9450 670
rect 9499 663 9550 679
rect 9404 560 9456 660
rect 9504 648 9550 663
rect 9471 632 9484 636
rect 9465 631 9484 632
rect 9504 632 9547 648
rect 9559 632 9572 636
rect 9462 620 9492 631
rect 9504 620 9544 632
rect 9465 572 9544 620
rect 9465 560 9505 572
rect 9525 560 9544 572
rect 9553 620 9572 632
rect 9584 632 9593 636
rect 9618 634 9743 686
rect 10004 670 10074 1163
rect 10186 1157 10198 1165
rect 10186 1151 10244 1157
rect 10373 1147 10722 1382
rect 10795 1214 10939 1218
rect 10848 1198 10939 1214
rect 10985 1214 11217 1218
rect 10985 1198 11048 1214
rect 10767 1186 10939 1190
rect 10820 1170 10939 1186
rect 10985 1186 11245 1190
rect 10985 1170 11076 1186
rect 10373 810 10443 1147
rect 10555 912 10613 918
rect 10555 878 10567 912
rect 10555 872 10613 878
rect 10831 859 10865 869
rect 11147 859 11181 869
rect 10831 851 11181 859
rect 10373 776 10444 810
rect 10795 789 11217 851
rect 10373 740 10426 776
rect 10004 634 10057 670
rect 9416 556 9425 560
rect 9437 556 9450 560
rect 9462 547 9518 560
rect 9525 556 9538 560
rect 9462 544 9528 547
rect 9357 445 9390 522
rect 9459 479 9528 544
rect 9553 534 9576 620
rect 9553 532 9572 534
rect 9559 522 9572 532
rect 9459 464 9517 479
rect 9584 465 9605 632
rect 9565 464 9605 465
rect 9618 464 9652 634
rect 9457 463 9510 464
rect 9517 463 9547 464
rect 9584 460 9593 464
rect 9357 411 9391 445
rect 9515 411 9549 445
rect 9618 426 9627 464
rect 9398 377 9425 411
rect 9488 400 9583 411
rect 9499 388 9583 400
rect 9639 388 9652 464
rect 9488 383 9583 388
rect 9488 377 9576 383
rect 9673 377 9706 634
rect 10186 619 10244 625
rect 10186 585 10198 619
rect 10186 579 10244 585
rect 11726 569 11772 580
rect 10140 493 10159 569
rect 11726 567 11744 569
rect 10168 542 10193 544
rect 10168 516 10196 542
rect 11727 510 11744 523
rect 10989 383 11023 417
rect 2021 348 2303 349
rect 3495 348 3777 349
rect 4969 348 5251 349
rect 6443 348 6725 349
rect 7917 348 8199 349
rect 9391 348 9673 349
rect 10865 348 11147 349
rect 2021 314 2303 315
rect 3495 314 3777 315
rect 4969 314 5251 315
rect 6443 314 6725 315
rect 7917 314 8199 315
rect 9391 314 9673 315
rect 10865 314 11147 315
rect 2083 255 2241 314
rect 3557 255 3715 314
rect 5031 255 5189 314
rect 6505 255 6663 314
rect 7979 255 8137 314
rect 9453 255 9611 314
rect 10927 255 11085 314
rect 9 141 21 168
rect -19 49 -7 77
rect 9 28 21 49
<< nwell >>
rect 10300 1147 10722 1823
rect 11303 1155 11816 1904
<< pwell >>
rect 10298 1904 10482 2452
rect 11528 1904 11816 2452
rect 10298 1877 10648 1904
rect 10318 1823 10648 1877
<< metal1 >>
rect 10332 2463 10476 2601
rect -54 2372 10476 2463
rect 11492 2452 11816 2601
rect -54 2280 -44 2372
rect 28 2326 10476 2372
rect 28 2280 38 2326
rect 9123 2320 10476 2326
rect -54 2186 4 2280
rect 10851 1913 10861 1976
rect 10949 1913 10959 1976
rect 11052 1794 11062 1877
rect 11150 1794 11160 1877
rect 547 1684 557 1756
rect 618 1684 628 1756
rect 1073 1684 1083 1756
rect 1144 1684 1154 1756
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 3495 1684 3505 1756
rect 3566 1684 3576 1756
rect 4021 1684 4031 1756
rect 4092 1684 4102 1756
rect 4969 1684 4979 1756
rect 5040 1684 5050 1756
rect 5495 1684 5505 1756
rect 5566 1684 5576 1756
rect 6443 1684 6453 1756
rect 6514 1684 6524 1756
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 7917 1684 7927 1756
rect 7988 1684 7998 1756
rect 8443 1684 8453 1756
rect 8514 1684 8524 1756
rect 9391 1684 9401 1756
rect 9462 1684 9472 1756
rect 9917 1684 9927 1756
rect 9988 1684 9998 1756
rect 328 1218 9266 1224
rect 0 1136 9266 1218
rect 10648 1136 11366 1190
rect 328 1130 9268 1136
rect -7 141 9 168
rect -7 49 3 141
rect 75 49 85 141
rect -7 28 9 49
<< via1 >>
rect -44 2280 28 2372
rect 10861 1913 10949 1976
rect 11062 1794 11150 1877
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
rect 3 49 75 141
<< metal2 >>
rect 62 2537 1547 2538
rect 62 2486 5975 2537
rect -44 2372 28 2382
rect -208 2280 -44 2365
rect -208 2278 28 2280
rect -208 124 -124 2278
rect -44 2270 28 2278
rect 15 1812 23 1838
rect 62 1826 114 2486
rect 1495 2485 5975 2486
rect 62 1812 79 1826
rect 1495 1811 1547 2485
rect 2972 2330 3043 2340
rect 2972 2246 3043 2256
rect 2981 1839 3033 2246
rect 2973 1813 3033 1839
rect 4451 1837 4503 2485
rect 2981 1812 3033 1813
rect 4436 1814 4503 1837
rect 5923 1817 5975 2485
rect 7396 2514 7467 2524
rect 7396 2420 7467 2430
rect 7404 1836 7456 2420
rect 4436 1811 4461 1814
rect 5923 1811 5948 1817
rect 7388 1813 7456 1836
rect 7388 1810 7413 1813
rect 8879 1810 8931 2443
rect 10861 1976 10949 1986
rect 10133 1970 10134 1973
rect 10087 1924 10861 1970
rect 10087 1804 10133 1924
rect 10861 1903 10949 1913
rect 11062 1877 11150 1887
rect 11062 1784 11150 1794
rect 557 1756 618 1766
rect 557 1674 618 1684
rect 1083 1756 1144 1766
rect 1083 1674 1144 1684
rect 2031 1756 2092 1766
rect 2031 1674 2092 1684
rect 2557 1756 2618 1766
rect 2557 1674 2618 1684
rect 3505 1756 3566 1766
rect 3505 1674 3566 1684
rect 4031 1756 4092 1766
rect 4031 1674 4092 1684
rect 4979 1756 5040 1766
rect 4979 1674 5040 1684
rect 5505 1756 5566 1766
rect 5505 1674 5566 1684
rect 6453 1756 6514 1766
rect 6453 1674 6514 1684
rect 6979 1756 7040 1766
rect 6979 1674 7040 1684
rect 7927 1756 7988 1766
rect 7927 1674 7988 1684
rect 8453 1756 8514 1766
rect 8453 1674 8514 1684
rect 9401 1756 9462 1766
rect 9401 1674 9462 1684
rect 9927 1756 9988 1766
rect 9927 1674 9988 1684
rect 11073 1409 11133 1784
rect 10952 1349 11133 1409
rect 10952 756 11012 1349
rect 10952 682 11012 692
rect 19 559 80 569
rect 19 493 80 503
rect 1671 559 1732 569
rect 3348 559 3409 569
rect 1732 518 1751 544
rect 1671 493 1732 503
rect 5035 559 5096 569
rect 3421 520 3446 546
rect 3348 493 3409 503
rect 6725 559 6786 569
rect 5106 519 5131 545
rect 5035 493 5096 503
rect 8413 559 8474 569
rect 6790 520 6815 546
rect 6725 493 6786 503
rect 10098 559 10159 569
rect 11744 567 11805 569
rect 8481 514 8506 540
rect 8413 493 8474 503
rect 11726 559 11805 567
rect 11726 552 11744 559
rect 10168 516 10193 542
rect 10098 493 10159 503
rect 11727 503 11744 510
rect 11727 495 11805 503
rect 11744 493 11805 495
rect 3 141 75 151
rect -208 49 3 124
rect -208 40 75 49
rect 3 39 75 40
<< via2 >>
rect 2972 2256 3043 2330
rect 7396 2430 7467 2514
rect 557 1684 618 1756
rect 1083 1684 1144 1756
rect 2031 1684 2092 1756
rect 2557 1684 2618 1756
rect 3505 1684 3566 1756
rect 4031 1684 4092 1756
rect 4979 1684 5040 1756
rect 5505 1684 5566 1756
rect 6453 1684 6514 1756
rect 6979 1684 7040 1756
rect 7927 1684 7988 1756
rect 8453 1684 8514 1756
rect 9401 1684 9462 1756
rect 9927 1684 9988 1756
rect 10952 692 11012 756
rect 19 503 80 559
rect 1671 503 1732 559
rect 3348 503 3409 559
rect 5035 503 5096 559
rect 6725 503 6786 559
rect 8413 503 8474 559
rect 10098 503 10159 559
rect 11744 503 11805 559
<< metal3 >>
rect 2981 2514 7477 2553
rect 2981 2493 7396 2514
rect 2981 2335 3041 2493
rect 7386 2430 7396 2493
rect 7467 2430 7477 2514
rect 7386 2425 7477 2430
rect 2962 2330 3053 2335
rect 2962 2256 2972 2330
rect 3043 2256 3053 2330
rect 2962 2251 3053 2256
rect 4497 2265 7957 2337
rect 1632 2014 3218 2086
rect 1632 1925 1704 2014
rect 1171 1853 1704 1925
rect 2753 1859 2903 1919
rect 2782 1848 2903 1859
rect 525 1756 628 1761
rect 525 1684 557 1756
rect 618 1684 628 1756
rect 525 1679 628 1684
rect 1054 1756 1154 1761
rect 1054 1684 1083 1756
rect 1144 1684 1154 1756
rect 1054 1679 1154 1684
rect 2021 1756 2102 1761
rect 2021 1684 2031 1756
rect 2092 1684 2102 1756
rect 2021 1679 2102 1684
rect 2547 1756 2628 1761
rect 2547 1684 2557 1756
rect 2618 1684 2628 1756
rect 2547 1679 2628 1684
rect 525 1183 585 1679
rect 26 1123 585 1183
rect 1054 1173 1114 1679
rect 26 564 86 1123
rect 1054 1113 1725 1173
rect 1665 564 1725 1113
rect 2031 699 2091 1679
rect 2564 867 2624 1679
rect 2843 1536 2903 1848
rect 3146 1769 3218 2014
rect 4497 1925 4569 2265
rect 6173 2039 7718 2111
rect 6173 1925 6245 2039
rect 4119 1853 4569 1925
rect 5593 1853 6245 1925
rect 7067 1853 7366 1925
rect 3146 1761 3560 1769
rect 3146 1756 3576 1761
rect 3146 1697 3505 1756
rect 3495 1684 3505 1697
rect 3566 1684 3576 1756
rect 4021 1756 4102 1761
rect 4021 1734 4031 1756
rect 3495 1679 3576 1684
rect 4020 1684 4031 1734
rect 4092 1684 4102 1756
rect 4020 1679 4102 1684
rect 4969 1756 5050 1761
rect 4969 1684 4979 1756
rect 5040 1748 5050 1756
rect 5495 1756 5576 1761
rect 5040 1684 5060 1748
rect 4969 1679 5060 1684
rect 5495 1684 5505 1756
rect 5566 1743 5576 1756
rect 6443 1756 6524 1761
rect 5566 1684 5585 1743
rect 5495 1679 5585 1684
rect 6443 1684 6453 1756
rect 6514 1734 6524 1756
rect 6969 1756 7050 1761
rect 6514 1684 6525 1734
rect 6443 1679 6525 1684
rect 6969 1684 6979 1756
rect 7040 1684 7050 1756
rect 6969 1679 7050 1684
rect 4020 1536 4080 1679
rect 2843 1476 4080 1536
rect 5000 1067 5060 1679
rect 5000 1007 5405 1067
rect 2564 807 5099 867
rect 2031 639 3414 699
rect 3354 564 3414 639
rect 5039 564 5099 807
rect 5345 809 5405 1007
rect 5525 950 5585 1679
rect 6465 1150 6525 1679
rect 6980 1335 7040 1679
rect 7294 1574 7366 1853
rect 7646 1774 7718 2039
rect 7885 2090 7957 2265
rect 7885 2018 9156 2090
rect 8541 1853 8845 1925
rect 7646 1761 7996 1774
rect 7646 1756 7998 1761
rect 7646 1702 7927 1756
rect 7917 1684 7927 1702
rect 7988 1684 7998 1756
rect 8443 1756 8524 1761
rect 8443 1742 8453 1756
rect 7917 1679 7998 1684
rect 8438 1684 8453 1742
rect 8514 1684 8524 1756
rect 8438 1679 8524 1684
rect 8438 1574 8510 1679
rect 7294 1502 8510 1574
rect 8773 1554 8845 1853
rect 9084 1769 9156 2018
rect 9084 1761 9446 1769
rect 9084 1756 9472 1761
rect 9084 1697 9401 1756
rect 9391 1684 9401 1697
rect 9462 1684 9472 1756
rect 9917 1756 9998 1761
rect 9917 1748 9927 1756
rect 9391 1679 9472 1684
rect 9902 1684 9927 1748
rect 9988 1684 9998 1756
rect 9902 1679 9998 1684
rect 9902 1554 9974 1679
rect 8773 1482 9974 1554
rect 6980 1275 10476 1335
rect 6465 1090 10166 1150
rect 5525 890 8474 950
rect 5345 749 6788 809
rect 6728 564 6788 749
rect 8414 564 8474 890
rect 10106 564 10166 1090
rect 10416 931 10476 1275
rect 10416 871 11810 931
rect 10942 756 11022 761
rect 10942 692 10952 756
rect 11012 692 11022 756
rect 10942 687 11022 692
rect 9 563 90 564
rect 9 559 145 563
rect 9 503 19 559
rect 80 503 145 559
rect 9 498 145 503
rect 1661 559 1742 564
rect 1661 503 1671 559
rect 1732 503 1742 559
rect 1661 498 1742 503
rect 3338 559 3419 564
rect 3338 503 3348 559
rect 3409 503 3419 559
rect 3338 498 3419 503
rect 5025 559 5106 564
rect 5025 503 5035 559
rect 5096 503 5106 559
rect 5025 498 5106 503
rect 6715 559 6796 564
rect 6715 503 6725 559
rect 6786 503 6796 559
rect 6715 498 6796 503
rect 8403 559 8484 564
rect 8403 503 8413 559
rect 8474 503 8484 559
rect 8403 498 8484 503
rect 10088 559 10169 564
rect 10088 503 10098 559
rect 10159 503 10169 559
rect 10088 498 10169 503
rect 85 112 145 498
rect 10952 112 11012 687
rect 11750 564 11810 871
rect 11734 559 11815 564
rect 11734 503 11744 559
rect 11805 503 11815 559
rect 11734 498 11815 503
rect 85 52 11012 112
use buffer_no_inv_x05  buffer_no_inv_x05_0
timestamp 1623938174
transform 1 0 -10 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_1
timestamp 1623938174
transform 1 0 834 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_2
timestamp 1623938174
transform 1 0 1678 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_0
timestamp 1624053917
transform 1 0 475 0 -1 1770
box -475 -2400 1898 1551
use mux_2to1_logic  mux_2to1_logic_1
timestamp 1624053917
transform 1 0 1949 0 -1 1770
box -475 -2400 1898 1551
use buffer_no_inv_x05  buffer_no_inv_x05_3
timestamp 1623938174
transform 1 0 2522 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_4
timestamp 1623938174
transform 1 0 3366 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_5
timestamp 1623938174
transform 1 0 4210 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_3
timestamp 1624053917
transform 1 0 4897 0 -1 1770
box -475 -2400 1898 1551
use mux_2to1_logic  mux_2to1_logic_2
timestamp 1624053917
transform 1 0 3423 0 -1 1770
box -475 -2400 1898 1551
use buffer_no_inv_x05  buffer_no_inv_x05_6
timestamp 1623938174
transform 1 0 5054 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_7
timestamp 1623938174
transform 1 0 5898 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_8
timestamp 1623938174
transform 1 0 6742 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_4
timestamp 1624053917
transform 1 0 6371 0 -1 1770
box -475 -2400 1898 1551
use buffer_no_inv_x05  buffer_no_inv_x05_9
timestamp 1623938174
transform 1 0 7586 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_10
timestamp 1623938174
transform 1 0 8430 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_11
timestamp 1623938174
transform 1 0 9274 0 1 -10
box 10 10 854 1173
use mux_2to1_logic  mux_2to1_logic_6
timestamp 1624053917
transform 1 0 9319 0 -1 1770
box -475 -2400 1898 1551
use mux_2to1_logic  mux_2to1_logic_5
timestamp 1624053917
transform 1 0 7845 0 -1 1770
box -475 -2400 1898 1551
use buffer_no_inv_x05  buffer_no_inv_x05_12
timestamp 1623938174
transform 1 0 10118 0 1 -10
box 10 10 854 1173
use buffer_no_inv_x05  buffer_no_inv_x05_13
timestamp 1623938174
transform 1 0 10962 0 1 -10
box 10 10 854 1173
use nand_logic  nand_logic_0
timestamp 1623952422
transform 1 0 10695 0 -1 1870
box -219 -731 833 707
<< labels >>
rlabel via2 30 516 55 542 1 clk
rlabel metal2 8893 2121 8918 2147 1 reg0
rlabel metal3 6059 2508 6084 2534 1 reg1
rlabel space 11254 1972 11279 1998 1 clk_out
rlabel metal2 80 2501 105 2527 1 reg2
rlabel space 32 1216 57 1242 1 avdd1p8
rlabel space 146 2318 171 2344 1 avss1p8
<< end >>
