magic
tech sky130A
timestamp 1616191796
<< error_s >>
rect 877 893 920 977
rect 961 891 1015 893
<< nwell >>
rect 1539 1212 1676 1213
rect 931 891 961 1211
rect 1533 893 2935 1212
<< pwell >>
rect 931 544 1786 836
rect 916 415 1786 544
rect 2776 -54 2804 -16
<< poly >>
rect 1571 1180 1590 1181
rect 2556 1180 2576 1181
rect 1571 1155 2576 1180
rect 1571 1093 1590 1155
rect 1277 1070 1590 1093
rect 931 846 982 876
rect 1114 867 1145 876
rect 1114 849 1122 867
rect 1139 849 1145 867
rect 1114 837 1145 849
rect 1567 869 1593 870
rect 1567 839 1598 869
rect 1567 384 1593 839
rect 2556 773 2576 1155
rect 2556 743 2612 773
rect 2597 708 2612 743
rect 2597 704 2637 708
rect 2597 679 2667 704
rect 1538 352 1618 384
rect 1538 314 1558 352
rect 1598 314 1618 352
rect 1538 289 1618 314
rect 2748 151 2774 157
rect 2719 119 2799 151
rect 2719 81 2739 119
rect 2779 81 2799 119
rect 2719 56 2799 81
rect 2484 -25 2507 56
rect 2752 -25 2775 56
rect 2484 -48 2776 -25
<< polycont >>
rect 1122 849 1139 867
rect 1558 314 1598 352
rect 2739 81 2779 119
<< locali >>
rect 1114 870 1145 877
rect 1114 843 1117 870
rect 1142 843 1145 870
rect 1114 837 1145 843
rect 1537 370 1618 371
rect 1537 302 1545 370
rect 1611 302 1618 370
rect 2718 137 2799 138
rect 2718 69 2726 137
rect 2792 69 2799 137
<< viali >>
rect 1117 867 1142 870
rect 1117 849 1122 867
rect 1122 849 1139 867
rect 1139 849 1142 867
rect 1117 843 1142 849
rect 1545 352 1611 370
rect 1545 314 1558 352
rect 1558 314 1598 352
rect 1598 314 1611 352
rect 1545 298 1611 314
rect 2726 119 2792 137
rect 2726 81 2739 119
rect 2739 81 2779 119
rect 2779 81 2792 119
rect 2726 65 2792 81
<< metal1 >>
rect 1114 875 1145 876
rect 1109 837 1114 875
rect 1146 837 1151 875
rect 1548 800 1566 820
rect 1536 742 1566 800
rect 1548 651 1566 742
rect 2529 655 2534 696
rect 2563 655 2568 696
rect 1548 610 1717 651
rect 1538 370 1618 384
rect 1538 298 1545 370
rect 1611 298 1618 370
rect 1538 289 1618 298
rect 2719 137 2799 151
rect 2719 65 2726 137
rect 2792 65 2799 137
rect 2719 56 2799 65
<< via1 >>
rect 1114 870 1146 875
rect 1114 843 1117 870
rect 1117 843 1142 870
rect 1142 843 1146 870
rect 1114 837 1146 843
rect 2534 655 2563 696
rect 1545 298 1611 370
rect 2726 65 2792 137
<< metal2 >>
rect 1109 875 1146 880
rect 1109 869 1114 875
rect 931 837 1114 869
rect 1146 837 1150 851
rect 931 835 1142 837
rect 2534 696 2563 701
rect 2534 650 2563 655
rect 1545 370 1611 375
rect 1545 293 1611 298
rect 2726 137 2792 142
rect 2726 60 2792 65
use xor2  xor2_0
timestamp 1616170071
transform -1 0 1538 0 1 893
box -26 -454 618 319
use dffc  dffc_0
timestamp 1616191617
transform 1 0 2027 0 1 396
box -433 -545 907 731
<< end >>
