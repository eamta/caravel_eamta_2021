magic
tech sky130A
magscale 1 2
timestamp 1615944125
<< pwell >>
rect -546 -1326 3146 174
<< metal1 >>
rect 370 207 2174 243
rect 370 127 1122 207
rect 1202 127 1231 207
rect 1311 127 1340 207
rect 1420 127 2174 207
rect 370 91 2174 127
rect 370 -237 522 91
rect 2022 -237 2174 91
rect -114 -283 2776 -237
rect -180 -903 -170 -327
rect -118 -903 -108 -327
rect -50 -1065 -3 -315
rect 56 -903 66 -327
rect 118 -903 128 -327
rect 186 -1065 233 -315
rect 292 -903 302 -327
rect 354 -903 364 -327
rect 422 -1065 469 -315
rect 528 -903 538 -327
rect 590 -903 600 -327
rect 658 -1065 705 -315
rect 764 -903 774 -327
rect 826 -903 836 -327
rect 894 -1065 941 -315
rect 1000 -903 1010 -327
rect 1062 -903 1072 -327
rect 1130 -1065 1177 -315
rect 1236 -903 1246 -327
rect 1298 -903 1308 -327
rect 1366 -1065 1413 -315
rect 1472 -903 1482 -327
rect 1534 -903 1544 -327
rect 1602 -1065 1649 -315
rect 1708 -903 1718 -327
rect 1770 -903 1780 -327
rect 1838 -1065 1885 -315
rect 1944 -903 1954 -327
rect 2006 -903 2016 -327
rect 2074 -1065 2121 -315
rect 2180 -903 2190 -327
rect 2242 -903 2252 -327
rect 2310 -1065 2357 -315
rect 2416 -903 2426 -327
rect 2478 -903 2488 -327
rect 2546 -1065 2593 -315
rect 2652 -903 2662 -327
rect 2714 -903 2724 -327
rect 2782 -1065 2829 -315
rect -50 -1075 2829 -1065
rect -50 -1135 1272 -1075
rect 1332 -1135 1360 -1075
rect 1420 -1135 1448 -1075
rect 1508 -1135 2829 -1075
rect -50 -1145 2829 -1135
<< via1 >>
rect 1122 127 1202 207
rect 1231 127 1311 207
rect 1340 127 1420 207
rect -170 -903 -118 -327
rect 66 -903 118 -327
rect 302 -903 354 -327
rect 538 -903 590 -327
rect 774 -903 826 -327
rect 1010 -903 1062 -327
rect 1246 -903 1298 -327
rect 1482 -903 1534 -327
rect 1718 -903 1770 -327
rect 1954 -903 2006 -327
rect 2190 -903 2242 -327
rect 2426 -903 2478 -327
rect 2662 -903 2714 -327
rect 1272 -1135 1332 -1075
rect 1360 -1135 1420 -1075
rect 1448 -1135 1508 -1075
<< metal2 >>
rect 1122 207 1202 217
rect 1122 117 1202 127
rect 1231 207 1311 217
rect 1231 117 1311 127
rect 1340 207 1420 217
rect 1340 117 1420 127
rect -170 -16 2714 -6
rect -170 -76 1161 -16
rect 1221 -76 1245 -16
rect 1305 -76 1329 -16
rect 1389 -76 2714 -16
rect -170 -86 2714 -76
rect -170 -327 -118 -86
rect -170 -913 -118 -903
rect 66 -327 118 -86
rect 66 -913 118 -903
rect 302 -327 354 -86
rect 302 -913 354 -903
rect 538 -327 590 -86
rect 538 -913 590 -903
rect 774 -327 826 -86
rect 774 -913 826 -903
rect 1010 -327 1062 -86
rect 1010 -913 1062 -903
rect 1246 -327 1298 -86
rect 1246 -913 1298 -903
rect 1482 -327 1534 -86
rect 1482 -913 1534 -903
rect 1718 -327 1770 -86
rect 1718 -913 1770 -903
rect 1954 -327 2006 -86
rect 1954 -913 2006 -903
rect 2190 -327 2242 -86
rect 2190 -913 2242 -903
rect 2426 -327 2478 -86
rect 2426 -913 2478 -903
rect 2662 -327 2714 -86
rect 2662 -913 2714 -903
rect 1272 -1075 1332 -1065
rect 1272 -1145 1332 -1135
rect 1360 -1075 1420 -1065
rect 1360 -1145 1420 -1135
rect 1448 -1075 1508 -1065
rect 1448 -1145 1508 -1135
<< via2 >>
rect 1161 -76 1221 -16
rect 1245 -76 1305 -16
rect 1329 -76 1389 -16
rect 1272 -1135 1332 -1075
rect 1360 -1135 1420 -1075
rect 1448 -1135 1508 -1075
<< metal3 >>
rect 1156 -16 1394 -6
rect 1156 -76 1161 -16
rect 1221 -76 1245 -16
rect 1305 -76 1329 -16
rect 1389 -76 1394 -16
rect 1156 -86 1394 -76
rect 1259 -1075 1526 -1063
rect 1259 -1135 1272 -1075
rect 1332 -1135 1360 -1075
rect 1420 -1135 1448 -1075
rect 1508 -1135 1526 -1075
rect 1259 -1146 1526 -1135
use sky130_fd_pr__nfet_01v8_QMU5EQ  sky130_fd_pr__nfet_01v8_QMU5EQ_0
timestamp 1615944125
transform 1 0 1331 0 1 -584
box -1642 -479 1642 479
<< end >>
