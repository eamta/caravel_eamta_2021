magic
tech sky130A
magscale 1 2
timestamp 1615898364
<< nwell >>
rect -1157 -884 1157 884
<< pmos >>
rect -961 -664 -821 736
rect -763 -664 -623 736
rect -565 -664 -425 736
rect -367 -664 -227 736
rect -169 -664 -29 736
rect 29 -664 169 736
rect 227 -664 367 736
rect 425 -664 565 736
rect 623 -664 763 736
rect 821 -664 961 736
<< pdiff >>
rect -1019 724 -961 736
rect -1019 -652 -1007 724
rect -973 -652 -961 724
rect -1019 -664 -961 -652
rect -821 724 -763 736
rect -821 -652 -809 724
rect -775 -652 -763 724
rect -821 -664 -763 -652
rect -623 724 -565 736
rect -623 -652 -611 724
rect -577 -652 -565 724
rect -623 -664 -565 -652
rect -425 724 -367 736
rect -425 -652 -413 724
rect -379 -652 -367 724
rect -425 -664 -367 -652
rect -227 724 -169 736
rect -227 -652 -215 724
rect -181 -652 -169 724
rect -227 -664 -169 -652
rect -29 724 29 736
rect -29 -652 -17 724
rect 17 -652 29 724
rect -29 -664 29 -652
rect 169 724 227 736
rect 169 -652 181 724
rect 215 -652 227 724
rect 169 -664 227 -652
rect 367 724 425 736
rect 367 -652 379 724
rect 413 -652 425 724
rect 367 -664 425 -652
rect 565 724 623 736
rect 565 -652 577 724
rect 611 -652 623 724
rect 565 -664 623 -652
rect 763 724 821 736
rect 763 -652 775 724
rect 809 -652 821 724
rect 763 -664 821 -652
rect 961 724 1019 736
rect 961 -652 973 724
rect 1007 -652 1019 724
rect 961 -664 1019 -652
<< pdiffc >>
rect -1007 -652 -973 724
rect -809 -652 -775 724
rect -611 -652 -577 724
rect -413 -652 -379 724
rect -215 -652 -181 724
rect -17 -652 17 724
rect 181 -652 215 724
rect 379 -652 413 724
rect 577 -652 611 724
rect 775 -652 809 724
rect 973 -652 1007 724
<< nsubdiff >>
rect -1121 814 -1025 848
rect 1025 814 1121 848
rect -1121 751 -1087 814
rect 1087 751 1121 814
rect -1121 -814 -1087 -751
rect 1087 -814 1121 -751
rect -1121 -848 -1025 -814
rect 1025 -848 1121 -814
<< nsubdiffcont >>
rect -1025 814 1025 848
rect -1121 -751 -1087 751
rect 1087 -751 1121 751
rect -1025 -848 1025 -814
<< poly >>
rect -961 736 -821 762
rect -763 736 -623 762
rect -565 736 -425 762
rect -367 736 -227 762
rect -169 736 -29 762
rect 29 736 169 762
rect 227 736 367 762
rect 425 736 565 762
rect 623 736 763 762
rect 821 736 961 762
rect -961 -711 -821 -664
rect -961 -745 -945 -711
rect -837 -745 -821 -711
rect -961 -761 -821 -745
rect -763 -711 -623 -664
rect -763 -745 -747 -711
rect -639 -745 -623 -711
rect -763 -761 -623 -745
rect -565 -711 -425 -664
rect -565 -745 -549 -711
rect -441 -745 -425 -711
rect -565 -761 -425 -745
rect -367 -711 -227 -664
rect -367 -745 -351 -711
rect -243 -745 -227 -711
rect -367 -761 -227 -745
rect -169 -711 -29 -664
rect -169 -745 -153 -711
rect -45 -745 -29 -711
rect -169 -761 -29 -745
rect 29 -711 169 -664
rect 29 -745 45 -711
rect 153 -745 169 -711
rect 29 -761 169 -745
rect 227 -711 367 -664
rect 227 -745 243 -711
rect 351 -745 367 -711
rect 227 -761 367 -745
rect 425 -711 565 -664
rect 425 -745 441 -711
rect 549 -745 565 -711
rect 425 -761 565 -745
rect 623 -711 763 -664
rect 623 -745 639 -711
rect 747 -745 763 -711
rect 623 -761 763 -745
rect 821 -711 961 -664
rect 821 -745 837 -711
rect 945 -745 961 -711
rect 821 -761 961 -745
<< polycont >>
rect -945 -745 -837 -711
rect -747 -745 -639 -711
rect -549 -745 -441 -711
rect -351 -745 -243 -711
rect -153 -745 -45 -711
rect 45 -745 153 -711
rect 243 -745 351 -711
rect 441 -745 549 -711
rect 639 -745 747 -711
rect 837 -745 945 -711
<< locali >>
rect -1121 814 -1025 848
rect 1025 814 1121 848
rect -1121 751 -1087 814
rect 1087 751 1121 814
rect -1007 724 -973 740
rect -1007 -668 -973 -652
rect -809 724 -775 740
rect -809 -668 -775 -652
rect -611 724 -577 740
rect -611 -668 -577 -652
rect -413 724 -379 740
rect -413 -668 -379 -652
rect -215 724 -181 740
rect -215 -668 -181 -652
rect -17 724 17 740
rect -17 -668 17 -652
rect 181 724 215 740
rect 181 -668 215 -652
rect 379 724 413 740
rect 379 -668 413 -652
rect 577 724 611 740
rect 577 -668 611 -652
rect 775 724 809 740
rect 775 -668 809 -652
rect 973 724 1007 740
rect 973 -668 1007 -652
rect -961 -745 -945 -711
rect -837 -745 -821 -711
rect -763 -745 -747 -711
rect -639 -745 -623 -711
rect -565 -745 -549 -711
rect -441 -745 -425 -711
rect -367 -745 -351 -711
rect -243 -745 -227 -711
rect -169 -745 -153 -711
rect -45 -745 -29 -711
rect 29 -745 45 -711
rect 153 -745 169 -711
rect 227 -745 243 -711
rect 351 -745 367 -711
rect 425 -745 441 -711
rect 549 -745 565 -711
rect 623 -745 639 -711
rect 747 -745 763 -711
rect 821 -745 837 -711
rect 945 -745 961 -711
rect -1121 -814 -1087 -751
rect 1087 -814 1121 -751
rect -1121 -848 -1025 -814
rect 1025 -848 1121 -814
<< viali >>
rect -1007 -652 -973 724
rect -809 -652 -775 724
rect -611 -652 -577 724
rect -413 -652 -379 724
rect -215 -652 -181 724
rect -17 -652 17 724
rect 181 -652 215 724
rect 379 -652 413 724
rect 577 -652 611 724
rect 775 -652 809 724
rect 973 -652 1007 724
rect -945 -745 -837 -711
rect -747 -745 -639 -711
rect -549 -745 -441 -711
rect -351 -745 -243 -711
rect -153 -745 -45 -711
rect 45 -745 153 -711
rect 243 -745 351 -711
rect 441 -745 549 -711
rect 639 -745 747 -711
rect 837 -745 945 -711
<< metal1 >>
rect -1013 724 -967 736
rect -1013 -652 -1007 724
rect -973 -652 -967 724
rect -1013 -664 -967 -652
rect -815 724 -769 736
rect -815 -652 -809 724
rect -775 -652 -769 724
rect -815 -664 -769 -652
rect -617 724 -571 736
rect -617 -652 -611 724
rect -577 -652 -571 724
rect -617 -664 -571 -652
rect -419 724 -373 736
rect -419 -652 -413 724
rect -379 -652 -373 724
rect -419 -664 -373 -652
rect -221 724 -175 736
rect -221 -652 -215 724
rect -181 -652 -175 724
rect -221 -664 -175 -652
rect -23 724 23 736
rect -23 -652 -17 724
rect 17 -652 23 724
rect -23 -664 23 -652
rect 175 724 221 736
rect 175 -652 181 724
rect 215 -652 221 724
rect 175 -664 221 -652
rect 373 724 419 736
rect 373 -652 379 724
rect 413 -652 419 724
rect 373 -664 419 -652
rect 571 724 617 736
rect 571 -652 577 724
rect 611 -652 617 724
rect 571 -664 617 -652
rect 769 724 815 736
rect 769 -652 775 724
rect 809 -652 815 724
rect 769 -664 815 -652
rect 967 724 1013 736
rect 967 -652 973 724
rect 1007 -652 1013 724
rect 967 -664 1013 -652
rect -957 -711 -825 -705
rect -957 -745 -945 -711
rect -837 -745 -825 -711
rect -957 -751 -825 -745
rect -759 -711 -627 -705
rect -759 -745 -747 -711
rect -639 -745 -627 -711
rect -759 -751 -627 -745
rect -561 -711 -429 -705
rect -561 -745 -549 -711
rect -441 -745 -429 -711
rect -561 -751 -429 -745
rect -363 -711 -231 -705
rect -363 -745 -351 -711
rect -243 -745 -231 -711
rect -363 -751 -231 -745
rect -165 -711 -33 -705
rect -165 -745 -153 -711
rect -45 -745 -33 -711
rect -165 -751 -33 -745
rect 33 -711 165 -705
rect 33 -745 45 -711
rect 153 -745 165 -711
rect 33 -751 165 -745
rect 231 -711 363 -705
rect 231 -745 243 -711
rect 351 -745 363 -711
rect 231 -751 363 -745
rect 429 -711 561 -705
rect 429 -745 441 -711
rect 549 -745 561 -711
rect 429 -751 561 -745
rect 627 -711 759 -705
rect 627 -745 639 -711
rect 747 -745 759 -711
rect 627 -751 759 -745
rect 825 -711 957 -705
rect 825 -745 837 -711
rect 945 -745 957 -711
rect 825 -751 957 -745
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1104 -831 1104 831
string parameters w 7 l 0.7 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
