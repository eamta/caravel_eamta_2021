magic
tech sky130A
magscale 1 2
timestamp 1619394249
<< viali >>
rect 800 9460 960 9480
rect 1740 9460 1880 9480
rect 2660 9460 2800 9480
rect 3600 9460 3740 9480
rect 4520 9460 4660 9480
rect 5460 9460 5600 9480
rect 6380 9460 6520 9480
rect -20 9420 7360 9460
rect -20 7660 20 9420
rect 800 7660 960 9420
rect 1740 7660 1880 9420
rect 2660 7660 2800 9420
rect 3600 7660 3740 9420
rect 4520 7660 4660 9420
rect 5460 7660 5600 9420
rect 6380 7660 6520 9420
rect 7320 7660 7360 9420
rect -20 7500 7360 7660
rect -20 5740 20 7500
rect 800 5740 960 7500
rect 1740 5740 1880 7500
rect 2660 5740 2800 7500
rect 3600 5740 3740 7500
rect 4520 5740 4660 7500
rect 5460 5740 5600 7500
rect 6380 5740 6520 7500
rect 7320 5740 7360 7500
rect -20 5600 7360 5740
rect -20 3840 20 5600
rect 800 3840 960 5600
rect 1740 3840 1880 5600
rect 2660 3840 2800 5600
rect 3600 3840 3740 5600
rect 4520 3840 4660 5600
rect 5460 3840 5600 5600
rect 6380 3840 6520 5600
rect 7320 3840 7360 5600
rect -20 3700 7360 3840
rect -20 1920 20 3700
rect 800 1920 960 3700
rect 1740 1920 1880 3700
rect 2660 1920 2800 3700
rect 3600 1920 3740 3700
rect 4520 1920 4660 3700
rect 5460 1920 5600 3700
rect 6380 1920 6520 3700
rect 7320 1920 7360 3700
rect -20 1780 7360 1920
rect -1600 1160 -140 1200
rect -1600 40 -1560 1160
rect -180 40 -140 1160
rect -1600 0 -140 40
rect -20 20 20 1780
rect 800 20 960 1780
rect 1740 20 1880 1780
rect 2660 20 2800 1780
rect 3600 20 3740 1780
rect 4520 20 4660 1780
rect 5460 20 5600 1780
rect 6380 20 6520 1780
rect 7320 20 7360 1780
rect -20 -20 7360 20
<< metal1 >>
rect -100 10400 -40 10500
rect 20 10400 900 10500
rect 960 10400 1840 10500
rect 1900 10400 2760 10500
rect 2820 10400 3700 10500
rect 3760 10400 4620 10500
rect 4680 10400 5560 10500
rect 5620 10400 6480 10500
rect 6540 10400 7400 10500
rect -100 10200 800 10300
rect 860 10200 1740 10300
rect 1800 10200 2660 10300
rect 2720 10200 3600 10300
rect 3660 10200 4520 10300
rect 4580 10200 5460 10300
rect 5520 10200 6380 10300
rect 6440 10200 7320 10300
rect 7380 10200 7400 10300
rect -100 10000 300 10100
rect 500 10000 1300 10100
rect 1400 10000 2200 10100
rect 2300 10000 3100 10100
rect 3300 10000 4100 10100
rect 4200 10000 5000 10100
rect 5100 10000 5900 10100
rect 6100 10000 6900 10100
rect 7000 10000 7400 10100
rect -340 9800 -180 9900
rect -80 9800 80 9900
rect 140 9800 1020 9900
rect 1080 9800 1940 9900
rect 2000 9800 2880 9900
rect 2940 9800 3800 9900
rect 3860 9800 4720 9900
rect 4780 9800 5660 9900
rect 5720 9800 6600 9900
rect 6660 9800 7400 9900
rect -340 9600 -320 9700
rect -220 9600 680 9700
rect 740 9600 1620 9700
rect 1680 9600 2540 9700
rect 2600 9600 3480 9700
rect 3540 9600 4400 9700
rect 4460 9600 5340 9700
rect 5400 9600 6260 9700
rect 6320 9600 7200 9700
rect 7260 9600 7400 9700
rect 794 9480 966 9492
rect 1734 9480 1886 9492
rect 2654 9480 2806 9492
rect 3594 9480 3746 9492
rect 4514 9480 4666 9492
rect 5454 9480 5606 9492
rect 6374 9480 6526 9492
rect 370 9466 380 9480
rect -32 9460 380 9466
rect 440 9466 450 9480
rect 794 9466 800 9480
rect 440 9460 800 9466
rect 960 9466 966 9480
rect 1310 9466 1320 9480
rect 960 9460 1320 9466
rect 1380 9466 1390 9480
rect 1734 9466 1740 9480
rect 1380 9460 1740 9466
rect 1880 9466 1886 9480
rect 2230 9466 2240 9480
rect 1880 9460 2240 9466
rect 2300 9466 2310 9480
rect 2654 9466 2660 9480
rect 2300 9460 2660 9466
rect 2800 9466 2806 9480
rect 3170 9466 3180 9480
rect 2800 9460 3180 9466
rect 3240 9466 3250 9480
rect 3594 9466 3600 9480
rect 3240 9460 3600 9466
rect 3740 9466 3746 9480
rect 4090 9466 4100 9480
rect 3740 9460 4100 9466
rect 4160 9466 4170 9480
rect 4514 9466 4520 9480
rect 4160 9460 4520 9466
rect 4660 9466 4666 9480
rect 5030 9466 5040 9480
rect 4660 9460 5040 9466
rect 5100 9466 5110 9480
rect 5454 9466 5460 9480
rect 5100 9460 5460 9466
rect 5600 9466 5606 9480
rect 5950 9466 5960 9480
rect 5600 9460 5960 9466
rect 6020 9466 6030 9480
rect 6374 9466 6380 9480
rect 6020 9460 6380 9466
rect 6520 9466 6526 9480
rect 6890 9466 6900 9480
rect 6520 9460 6900 9466
rect 6960 9466 6970 9480
rect 6960 9460 7372 9466
rect -32 9414 -20 9460
rect -26 7666 -20 9414
rect -32 7494 -20 7666
rect 20 9414 800 9420
rect 20 7666 26 9414
rect 190 9360 200 9380
rect 140 9320 200 9360
rect 190 9280 200 9320
rect 320 9360 330 9380
rect 490 9360 500 9380
rect 320 9320 380 9360
rect 440 9320 500 9360
rect 320 9280 330 9320
rect 490 9280 500 9320
rect 620 9360 630 9380
rect 620 9320 680 9360
rect 620 9280 630 9320
rect 70 7800 80 9260
rect 140 7800 150 9260
rect 370 7800 380 9260
rect 440 7800 450 9260
rect 670 7800 680 9260
rect 740 7800 750 9260
rect 190 7760 200 7800
rect 140 7720 200 7760
rect 190 7700 200 7720
rect 320 7760 330 7800
rect 490 7760 500 7800
rect 320 7720 380 7760
rect 440 7720 500 7760
rect 320 7700 330 7720
rect 490 7700 500 7720
rect 620 7760 630 7800
rect 620 7720 680 7760
rect 620 7700 630 7720
rect 794 7666 800 9414
rect 20 7660 800 7666
rect 960 9414 1740 9420
rect 960 7666 966 9414
rect 1130 9360 1140 9380
rect 1080 9320 1140 9360
rect 1130 9280 1140 9320
rect 1260 9360 1270 9380
rect 1410 9360 1420 9380
rect 1260 9320 1320 9360
rect 1380 9320 1420 9360
rect 1260 9280 1270 9320
rect 1410 9280 1420 9320
rect 1540 9360 1550 9380
rect 1540 9320 1620 9360
rect 1540 9280 1550 9320
rect 1010 7800 1020 9260
rect 1080 7800 1090 9260
rect 1310 7800 1320 9260
rect 1380 7800 1390 9260
rect 1610 7800 1620 9260
rect 1680 7800 1690 9260
rect 1130 7760 1140 7800
rect 1080 7720 1140 7760
rect 1130 7700 1140 7720
rect 1260 7760 1270 7800
rect 1430 7760 1440 7800
rect 1260 7720 1320 7760
rect 1380 7720 1440 7760
rect 1260 7700 1270 7720
rect 1430 7700 1440 7720
rect 1560 7760 1570 7800
rect 1560 7720 1620 7760
rect 1560 7700 1570 7720
rect 1734 7666 1740 9414
rect 960 7660 1740 7666
rect 1880 9414 2660 9420
rect 1880 7666 1886 9414
rect 2050 9360 2060 9380
rect 2000 9320 2060 9360
rect 2050 9280 2060 9320
rect 2180 9360 2190 9380
rect 2350 9360 2360 9380
rect 2180 9320 2240 9360
rect 2300 9320 2360 9360
rect 2180 9280 2190 9320
rect 2350 9280 2360 9320
rect 2480 9360 2490 9380
rect 2480 9320 2540 9360
rect 2480 9280 2490 9320
rect 1930 7800 1940 9260
rect 2000 7800 2010 9260
rect 2230 7800 2240 9260
rect 2300 7800 2310 9260
rect 2530 7800 2540 9260
rect 2600 7800 2610 9260
rect 2050 7760 2060 7800
rect 2000 7720 2060 7760
rect 2050 7700 2060 7720
rect 2180 7760 2190 7800
rect 2350 7760 2360 7800
rect 2180 7720 2240 7760
rect 2300 7720 2360 7760
rect 2180 7700 2190 7720
rect 2350 7700 2360 7720
rect 2480 7760 2490 7800
rect 2480 7720 2540 7760
rect 2480 7700 2490 7720
rect 2654 7666 2660 9414
rect 1880 7660 2660 7666
rect 2800 9414 3600 9420
rect 2800 7666 2806 9414
rect 2990 9360 3000 9380
rect 2920 9320 3000 9360
rect 2990 9280 3000 9320
rect 3120 9360 3130 9380
rect 3290 9360 3300 9380
rect 3120 9320 3180 9360
rect 3240 9320 3300 9360
rect 3120 9280 3130 9320
rect 3290 9280 3300 9320
rect 3420 9360 3430 9380
rect 3420 9320 3460 9360
rect 3420 9280 3430 9320
rect 2870 7800 2880 9260
rect 2940 7800 2950 9260
rect 3170 7800 3180 9260
rect 3240 7800 3250 9260
rect 3470 7800 3480 9260
rect 3540 7800 3550 9260
rect 2990 7700 3000 7800
rect 3120 7700 3130 7800
rect 3290 7700 3300 7800
rect 3420 7700 3430 7800
rect 3594 7666 3600 9414
rect 2800 7660 3600 7666
rect 3740 9414 4520 9420
rect 3740 7666 3746 9414
rect 3910 9360 3920 9380
rect 3860 9320 3920 9360
rect 3910 9280 3920 9320
rect 4040 9360 4050 9380
rect 4210 9360 4220 9380
rect 4040 9320 4100 9360
rect 4160 9320 4220 9360
rect 4040 9280 4050 9320
rect 4210 9280 4220 9320
rect 4340 9360 4350 9380
rect 4340 9320 4400 9360
rect 4340 9280 4350 9320
rect 3790 7800 3800 9260
rect 3860 7800 3870 9260
rect 4090 7800 4100 9260
rect 4160 7800 4170 9260
rect 4390 7800 4400 9260
rect 4460 7800 4470 9260
rect 3910 7700 3920 7800
rect 4040 7700 4050 7800
rect 4210 7700 4220 7800
rect 4340 7700 4350 7800
rect 4514 7666 4520 9414
rect 3740 7660 4520 7666
rect 4660 9414 5460 9420
rect 4660 7666 4666 9414
rect 4850 9360 4860 9380
rect 4800 9320 4860 9360
rect 4850 9280 4860 9320
rect 4980 9360 4990 9380
rect 5150 9360 5160 9380
rect 4980 9320 5040 9360
rect 5100 9320 5160 9360
rect 4980 9280 4990 9320
rect 5150 9280 5160 9320
rect 5280 9360 5290 9380
rect 5280 9320 5340 9360
rect 5280 9280 5290 9320
rect 4720 7790 4730 9250
rect 4790 7790 4800 9250
rect 4830 7700 4840 7800
rect 4960 7700 4970 7800
rect 5020 7790 5030 9250
rect 5090 7790 5100 9250
rect 5150 7700 5160 7800
rect 5280 7700 5290 7800
rect 5320 7790 5330 9250
rect 5390 7790 5400 9250
rect 5454 7666 5460 9414
rect 4660 7660 5460 7666
rect 5600 9414 6380 9420
rect 5600 7666 5606 9414
rect 5770 9360 5780 9380
rect 5720 9320 5780 9360
rect 5770 9280 5780 9320
rect 5900 9360 5910 9380
rect 6070 9360 6080 9380
rect 5900 9320 5960 9360
rect 6020 9320 6080 9360
rect 5900 9280 5910 9320
rect 6070 9280 6080 9320
rect 6200 9360 6210 9380
rect 6200 9320 6260 9360
rect 6200 9280 6210 9320
rect 5650 7800 5660 9260
rect 5720 7800 5730 9260
rect 5950 7800 5960 9260
rect 6020 7800 6030 9260
rect 6250 7800 6260 9260
rect 6320 7800 6330 9260
rect 5770 7700 5780 7800
rect 5900 7700 5910 7800
rect 6070 7700 6080 7800
rect 6200 7700 6210 7800
rect 6374 7666 6380 9414
rect 5600 7660 6380 7666
rect 6520 9414 7320 9420
rect 6520 7666 6526 9414
rect 6710 9360 6720 9380
rect 6660 9320 6720 9360
rect 6710 9280 6720 9320
rect 6840 9360 6850 9380
rect 7010 9360 7020 9380
rect 6840 9320 6900 9360
rect 6960 9320 7020 9360
rect 6840 9280 6850 9320
rect 7010 9280 7020 9320
rect 7140 9360 7150 9380
rect 7140 9320 7200 9360
rect 7140 9280 7150 9320
rect 6580 7800 6590 9260
rect 6650 7800 6660 9260
rect 6880 7800 6890 9260
rect 6950 7800 6960 9260
rect 7180 7800 7190 9260
rect 7250 7800 7260 9260
rect 6710 7700 6720 7800
rect 6840 7700 6850 7800
rect 7010 7700 7020 7800
rect 7140 7700 7150 7800
rect 7314 7666 7320 9414
rect 6520 7660 7320 7666
rect 7360 9414 7372 9460
rect 7360 7666 7366 9414
rect -26 5746 -20 7494
rect -32 5594 -20 5746
rect 20 7494 800 7500
rect 20 5746 26 7494
rect 190 7440 200 7460
rect 140 7400 200 7440
rect 190 7360 200 7400
rect 320 7440 330 7460
rect 490 7440 500 7460
rect 320 7400 380 7440
rect 440 7400 500 7440
rect 320 7360 330 7400
rect 490 7360 500 7400
rect 620 7440 630 7460
rect 620 7400 680 7440
rect 620 7360 630 7400
rect 70 5890 80 7350
rect 140 5890 150 7350
rect 370 5890 380 7350
rect 440 5890 450 7350
rect 670 5890 680 7350
rect 740 5890 750 7350
rect 190 5780 200 5880
rect 320 5780 330 5880
rect 490 5780 500 5880
rect 620 5780 630 5880
rect 794 5746 800 7494
rect 20 5740 800 5746
rect 960 7494 1740 7500
rect 960 5746 966 7494
rect 1130 7440 1140 7460
rect 1080 7400 1140 7440
rect 1130 7360 1140 7400
rect 1260 7440 1270 7460
rect 1430 7440 1440 7460
rect 1260 7400 1300 7440
rect 1360 7400 1440 7440
rect 1260 7360 1270 7400
rect 1430 7360 1440 7400
rect 1560 7440 1570 7460
rect 1560 7400 1620 7440
rect 1560 7360 1570 7400
rect 1000 5900 1010 7360
rect 1070 5900 1080 7360
rect 1300 5900 1310 7360
rect 1370 5900 1380 7360
rect 1600 5900 1610 7360
rect 1670 5900 1680 7360
rect 1130 5780 1140 5880
rect 1260 5780 1270 5880
rect 1430 5780 1440 5880
rect 1560 5780 1570 5880
rect 1734 5746 1740 7494
rect 960 5740 1740 5746
rect 1880 7494 2660 7500
rect 1880 5746 1886 7494
rect 2050 7440 2060 7460
rect 2000 7400 2060 7440
rect 2050 7360 2060 7400
rect 2180 7440 2190 7460
rect 2350 7440 2360 7460
rect 2180 7400 2240 7440
rect 2300 7400 2360 7440
rect 2180 7360 2190 7400
rect 2350 7360 2360 7400
rect 2480 7440 2490 7460
rect 2480 7400 2540 7440
rect 2480 7360 2490 7400
rect 1930 5900 1940 7360
rect 2000 5900 2010 7360
rect 2230 5900 2240 7360
rect 2300 5900 2310 7360
rect 2530 5900 2540 7360
rect 2600 5900 2610 7360
rect 2050 5780 2060 5880
rect 2180 5780 2190 5880
rect 2350 5780 2360 5880
rect 2480 5780 2490 5880
rect 2654 5746 2660 7494
rect 1880 5740 2660 5746
rect 2800 7494 3600 7500
rect 2800 5746 2806 7494
rect 2990 7360 3000 7460
rect 3120 7360 3130 7460
rect 3270 7360 3280 7460
rect 3400 7360 3410 7460
rect 2860 5890 2870 7350
rect 2930 5890 2940 7350
rect 3160 5890 3170 7350
rect 3230 5890 3240 7350
rect 3460 5890 3470 7350
rect 3530 5890 3540 7350
rect 2990 5780 3000 5880
rect 3120 5780 3130 5880
rect 3290 5780 3300 5880
rect 3420 5780 3430 5880
rect 3594 5746 3600 7494
rect 2800 5740 3600 5746
rect 3740 7494 4520 7500
rect 3740 5746 3746 7494
rect 3910 7360 3920 7460
rect 4040 7360 4050 7460
rect 4210 7360 4220 7460
rect 4340 7360 4350 7460
rect 3790 5890 3800 7350
rect 3860 5890 3870 7350
rect 4090 5890 4100 7350
rect 4160 5890 4170 7350
rect 4390 5890 4400 7350
rect 4460 5890 4470 7350
rect 3910 5780 3920 5880
rect 4040 5780 4050 5880
rect 4210 5780 4220 5880
rect 4340 5780 4350 5880
rect 4514 5746 4520 7494
rect 3740 5740 4520 5746
rect 4660 7494 5460 7500
rect 4660 5746 4666 7494
rect 4840 7360 4850 7460
rect 4970 7360 4980 7460
rect 5130 7360 5140 7460
rect 5260 7360 5270 7460
rect 4720 5890 4730 7350
rect 4790 5890 4800 7350
rect 5020 5890 5030 7350
rect 5090 5890 5100 7350
rect 5320 5890 5330 7350
rect 5390 5890 5400 7350
rect 4840 5780 4850 5880
rect 4970 5780 4980 5880
rect 5150 5780 5160 5880
rect 5280 5780 5290 5880
rect 5454 5746 5460 7494
rect 4660 5740 5460 5746
rect 5600 7494 6380 7500
rect 5600 5746 5606 7494
rect 5770 7360 5780 7460
rect 5900 7360 5910 7460
rect 6070 7360 6080 7460
rect 6200 7360 6210 7460
rect 5650 5890 5660 7350
rect 5720 5890 5730 7350
rect 5950 5890 5960 7350
rect 6020 5890 6030 7350
rect 6250 5890 6260 7350
rect 6320 5890 6330 7350
rect 5770 5780 5780 5880
rect 5900 5780 5910 5880
rect 6080 5780 6090 5880
rect 6210 5780 6220 5880
rect 6374 5746 6380 7494
rect 5600 5740 6380 5746
rect 6520 7494 7320 7500
rect 6520 5746 6526 7494
rect 6710 7360 6720 7460
rect 6840 7360 6850 7460
rect 7010 7360 7020 7460
rect 7140 7360 7150 7460
rect 6580 5890 6590 7350
rect 6650 5890 6660 7350
rect 6880 5890 6890 7350
rect 6950 5890 6960 7350
rect 7180 5890 7190 7350
rect 7250 5890 7260 7350
rect 6700 5780 6710 5880
rect 6830 5780 6840 5880
rect 7000 5780 7010 5880
rect 7130 5780 7140 5880
rect 7314 5746 7320 7494
rect 6520 5740 7320 5746
rect 7360 7494 7372 7666
rect 7360 5746 7366 7494
rect -26 3846 -20 5594
rect -32 3694 -20 3846
rect 20 5594 800 5600
rect 20 3846 26 5594
rect 190 5460 200 5560
rect 320 5460 330 5560
rect 500 5460 510 5560
rect 630 5460 640 5560
rect 70 3980 80 5440
rect 140 3980 150 5440
rect 180 3890 190 3990
rect 310 3890 320 3990
rect 370 3980 380 5440
rect 440 3980 450 5440
rect 500 3890 510 3990
rect 630 3890 640 3990
rect 670 3980 680 5440
rect 740 3980 750 5440
rect 794 3846 800 5594
rect 20 3840 800 3846
rect 960 5594 1740 5600
rect 960 3846 966 5594
rect 1120 5460 1130 5560
rect 1250 5460 1260 5560
rect 1430 5460 1440 5560
rect 1560 5460 1570 5560
rect 1000 3990 1010 5450
rect 1070 3990 1080 5450
rect 1300 3990 1310 5450
rect 1370 3990 1380 5450
rect 1600 3990 1610 5450
rect 1670 3990 1680 5450
rect 1120 3890 1130 3990
rect 1250 3890 1260 3990
rect 1420 3890 1430 3990
rect 1550 3890 1560 3990
rect 1734 3846 1740 5594
rect 960 3840 1740 3846
rect 1880 5594 2660 5600
rect 1880 3846 1886 5594
rect 2050 5460 2060 5560
rect 2180 5460 2190 5560
rect 2360 5460 2370 5560
rect 2490 5460 2500 5560
rect 1930 3990 1940 5450
rect 2000 3990 2010 5450
rect 2230 3990 2240 5450
rect 2300 3990 2310 5450
rect 2530 3990 2540 5450
rect 2600 3990 2610 5450
rect 2040 3890 2050 3990
rect 2170 3890 2180 3990
rect 2340 3890 2350 3990
rect 2470 3890 2480 3990
rect 2654 3846 2660 5594
rect 1880 3840 2660 3846
rect 2800 5594 3600 5600
rect 2800 3846 2806 5594
rect 2990 5460 3000 5560
rect 3120 5460 3130 5560
rect 3290 5460 3300 5560
rect 3420 5460 3430 5560
rect 2860 3980 2870 5440
rect 2930 3980 2940 5440
rect 2980 3890 2990 3990
rect 3110 3890 3120 3990
rect 3160 3980 3170 5440
rect 3230 3980 3240 5440
rect 3280 3890 3290 3990
rect 3410 3890 3420 3990
rect 3460 3980 3470 5440
rect 3530 3980 3540 5440
rect 3594 3846 3600 5594
rect 2800 3840 3600 3846
rect 3740 5594 4520 5600
rect 3740 3846 3746 5594
rect 3920 5460 3930 5560
rect 4050 5460 4060 5560
rect 4210 5460 4220 5560
rect 4340 5460 4350 5560
rect 3790 3970 3800 5430
rect 3860 3970 3870 5430
rect 3920 3890 3930 3990
rect 4050 3890 4060 3990
rect 4090 3970 4100 5430
rect 4160 3970 4170 5430
rect 4200 3890 4210 3990
rect 4330 3890 4340 3990
rect 4390 3970 4400 5430
rect 4460 3970 4470 5430
rect 4514 3846 4520 5594
rect 3740 3840 4520 3846
rect 4660 5594 5460 5600
rect 4660 3846 4666 5594
rect 4840 5460 4850 5560
rect 4970 5460 4980 5560
rect 5150 5460 5160 5560
rect 5280 5460 5290 5560
rect 4720 3970 4730 5430
rect 4790 3970 4800 5430
rect 4840 3890 4850 3990
rect 4970 3890 4980 3990
rect 5020 3970 5030 5430
rect 5090 3970 5100 5430
rect 5140 3890 5150 3990
rect 5270 3890 5280 3990
rect 5320 3970 5330 5430
rect 5390 3970 5400 5430
rect 5454 3846 5460 5594
rect 4660 3840 5460 3846
rect 5600 5594 6380 5600
rect 5600 3846 5606 5594
rect 5780 5460 5790 5560
rect 5910 5460 5920 5560
rect 6080 5460 6090 5560
rect 6210 5460 6220 5560
rect 5650 3970 5660 5430
rect 5720 3970 5730 5430
rect 5780 3890 5790 3990
rect 5910 3890 5920 3990
rect 5950 3970 5960 5430
rect 6020 3970 6030 5430
rect 6070 3880 6080 3980
rect 6200 3880 6210 3980
rect 6250 3970 6260 5430
rect 6320 3970 6330 5430
rect 6374 3846 6380 5594
rect 5600 3840 6380 3846
rect 6520 5594 7320 5600
rect 6520 3846 6526 5594
rect 6690 5460 6700 5560
rect 6820 5460 6830 5560
rect 7010 5460 7020 5560
rect 7140 5460 7150 5560
rect 6580 3980 6590 5440
rect 6650 3980 6660 5440
rect 6880 3980 6890 5440
rect 6950 3980 6960 5440
rect 7180 3980 7190 5440
rect 7250 3980 7260 5440
rect 6700 3880 6710 3980
rect 6830 3880 6840 3980
rect 7010 3880 7020 3980
rect 7140 3880 7150 3980
rect 7314 3846 7320 5594
rect 6520 3840 7320 3846
rect 7360 5594 7372 5746
rect 7360 3846 7366 5594
rect -26 1926 -20 3694
rect -32 1774 -20 1926
rect 20 3694 800 3700
rect 20 1926 26 3694
rect 200 3550 210 3650
rect 330 3550 340 3650
rect 500 3550 510 3650
rect 630 3550 640 3650
rect 70 2080 80 3540
rect 140 2080 150 3540
rect 370 2080 380 3540
rect 440 2080 450 3540
rect 670 2080 680 3540
rect 740 2080 750 3540
rect 180 1970 190 2070
rect 310 1970 320 2070
rect 500 1970 510 2070
rect 630 1970 640 2070
rect 794 1926 800 3694
rect 20 1920 800 1926
rect 960 3694 1740 3700
rect 960 1926 966 3694
rect 1120 3550 1130 3650
rect 1250 3550 1260 3650
rect 1420 3550 1430 3650
rect 1550 3550 1560 3650
rect 1000 2080 1010 3540
rect 1070 2080 1080 3540
rect 1300 2080 1310 3540
rect 1370 2080 1380 3540
rect 1600 2080 1610 3540
rect 1670 2080 1680 3540
rect 1120 1970 1130 2070
rect 1250 1970 1260 2070
rect 1420 1970 1430 2070
rect 1550 1970 1560 2070
rect 1734 1926 1740 3694
rect 960 1920 1740 1926
rect 1880 3694 2660 3700
rect 1880 1926 1886 3694
rect 2060 3550 2070 3650
rect 2190 3550 2200 3650
rect 2360 3550 2370 3650
rect 2490 3550 2500 3650
rect 1930 2080 1940 3540
rect 2000 2080 2010 3540
rect 2230 2080 2240 3540
rect 2300 2080 2310 3540
rect 2530 2080 2540 3540
rect 2600 2080 2610 3540
rect 2040 1970 2050 2070
rect 2170 1970 2180 2070
rect 2360 1970 2370 2070
rect 2490 1970 2500 2070
rect 2654 1926 2660 3694
rect 1880 1920 2660 1926
rect 2800 3694 3600 3700
rect 2800 1926 2806 3694
rect 2980 3550 2990 3650
rect 3110 3550 3120 3650
rect 3300 3550 3310 3650
rect 3430 3550 3440 3650
rect 2870 2110 2880 3470
rect 2940 2110 2950 3470
rect 3170 2110 3180 3470
rect 3240 2110 3250 3470
rect 3470 2110 3480 3470
rect 3540 2110 3550 3470
rect 2980 1970 2990 2070
rect 3110 1970 3120 2070
rect 3280 1970 3290 2070
rect 3410 1970 3420 2070
rect 3594 1926 3600 3694
rect 2800 1920 3600 1926
rect 3740 3694 4520 3700
rect 3740 1926 3746 3694
rect 3920 3550 3930 3650
rect 4050 3550 4060 3650
rect 4220 3550 4230 3650
rect 4350 3550 4360 3650
rect 3790 2070 3800 3530
rect 3860 2070 3870 3530
rect 4090 2070 4100 3530
rect 4160 2070 4170 3530
rect 4390 2070 4400 3530
rect 4460 2070 4470 3530
rect 3900 1970 3910 2070
rect 4030 1970 4040 2070
rect 4220 1970 4230 2070
rect 4350 1970 4360 2070
rect 4514 1926 4520 3694
rect 3740 1920 4520 1926
rect 4660 3694 5460 3700
rect 4660 1926 4666 3694
rect 4840 3550 4850 3650
rect 4970 3550 4980 3650
rect 5140 3550 5150 3650
rect 5270 3550 5280 3650
rect 4720 2070 4730 3530
rect 4790 2070 4800 3530
rect 5020 2070 5030 3530
rect 5090 2070 5100 3530
rect 5320 2070 5330 3530
rect 5390 2070 5400 3530
rect 4840 1970 4850 2070
rect 4970 1970 4980 2070
rect 5140 1970 5150 2070
rect 5270 1970 5280 2070
rect 5454 1926 5460 3694
rect 4660 1920 5460 1926
rect 5600 3694 6380 3700
rect 5600 1926 5606 3694
rect 5780 3550 5790 3650
rect 5910 3550 5920 3650
rect 6060 3550 6070 3650
rect 6190 3550 6200 3650
rect 5650 2080 5660 3540
rect 5720 2080 5730 3540
rect 5950 2080 5960 3540
rect 6020 2080 6030 3540
rect 6250 2080 6260 3540
rect 6320 2080 6330 3540
rect 5780 1970 5790 2070
rect 5910 1970 5920 2070
rect 6080 1970 6090 2070
rect 6210 1970 6220 2070
rect 6374 1926 6380 3694
rect 5600 1920 6380 1926
rect 6520 3694 7320 3700
rect 6520 1926 6526 3694
rect 6700 3550 6710 3650
rect 6830 3550 6840 3650
rect 7000 3550 7010 3650
rect 7130 3550 7140 3650
rect 6580 2080 6590 3540
rect 6650 2080 6660 3540
rect 6880 2080 6890 3540
rect 6950 2080 6960 3540
rect 7180 2080 7190 3540
rect 7250 2080 7260 3540
rect 6700 1970 6710 2070
rect 6830 1970 6840 2070
rect 7000 1970 7010 2070
rect 7130 1970 7140 2070
rect 7314 1926 7320 3694
rect 6520 1920 7320 1926
rect 7360 3694 7372 3846
rect 7360 1926 7366 3694
rect -1400 1500 -1340 1600
rect -1280 1500 -740 1600
rect -680 1500 -320 1600
rect -220 1500 -100 1600
rect -1400 1300 -1040 1400
rect -980 1300 -460 1400
rect -400 1300 -180 1400
rect -80 1300 -70 1400
rect -1606 1206 -1554 1212
rect -186 1206 -134 1212
rect -1612 1200 -128 1206
rect -1612 1154 -1600 1200
rect -1606 46 -1600 1154
rect -1612 0 -1600 46
rect -1560 1154 -180 1160
rect -1560 46 -1554 1154
rect -1440 1040 -300 1100
rect -1360 960 -1260 1040
rect -760 960 -680 1040
rect -1510 220 -1500 960
rect -1440 220 -1430 960
rect -1350 220 -1340 960
rect -1280 220 -1270 960
rect -1210 220 -1200 960
rect -1140 220 -1130 960
rect -1050 220 -1040 960
rect -980 220 -970 960
rect -910 220 -900 960
rect -840 220 -830 960
rect -750 220 -740 960
rect -680 220 -670 960
rect -610 220 -600 960
rect -540 220 -530 960
rect -470 220 -460 960
rect -400 220 -390 960
rect -310 220 -300 960
rect -240 220 -230 960
rect -1340 140 -1280 220
rect -760 140 -680 220
rect -1440 100 -300 140
rect -186 46 -180 1154
rect -1560 40 -180 46
rect -140 1154 -128 1200
rect -140 46 -134 1154
rect -140 0 -128 46
rect -26 26 -20 1774
rect -1612 -6 -128 0
rect -1606 -12 -134 -6
rect -1600 -40 -140 -12
rect -32 -20 -20 26
rect 20 1774 800 1780
rect 20 26 26 1774
rect 70 180 80 1640
rect 140 180 150 1640
rect 180 1630 190 1730
rect 310 1630 320 1730
rect 370 180 380 1640
rect 440 180 450 1640
rect 500 1630 510 1730
rect 630 1630 640 1730
rect 670 180 680 1640
rect 740 180 750 1640
rect 200 70 210 170
rect 330 70 340 170
rect 500 70 510 170
rect 630 70 640 170
rect 794 26 800 1774
rect 20 20 800 26
rect 960 1774 1740 1780
rect 960 26 966 1774
rect 1120 1630 1130 1730
rect 1250 1630 1260 1730
rect 1420 1630 1430 1730
rect 1550 1630 1560 1730
rect 1010 210 1020 1570
rect 1080 210 1090 1570
rect 1310 210 1320 1570
rect 1380 210 1390 1570
rect 1610 210 1620 1570
rect 1680 210 1690 1570
rect 1120 70 1130 170
rect 1250 70 1260 170
rect 1440 70 1450 170
rect 1570 70 1580 170
rect 1734 26 1740 1774
rect 960 20 1740 26
rect 1880 1774 2660 1780
rect 1880 26 1886 1774
rect 2060 1630 2070 1730
rect 2190 1630 2200 1730
rect 2360 1630 2370 1730
rect 2490 1630 2500 1730
rect 1930 170 1940 1630
rect 2000 170 2010 1630
rect 2230 170 2240 1630
rect 2300 170 2310 1630
rect 2530 170 2540 1630
rect 2600 170 2610 1630
rect 2060 70 2070 170
rect 2190 70 2200 170
rect 2340 70 2350 170
rect 2470 70 2480 170
rect 2654 26 2660 1774
rect 1880 20 2660 26
rect 2800 1774 3600 1780
rect 2800 26 2806 1774
rect 3000 1630 3010 1730
rect 3130 1630 3140 1730
rect 3300 1630 3310 1730
rect 3430 1630 3440 1730
rect 2860 210 2870 1570
rect 2930 210 2940 1570
rect 3160 210 3170 1570
rect 3230 210 3240 1570
rect 3460 210 3470 1570
rect 3530 210 3540 1570
rect 2980 70 2990 170
rect 3110 70 3120 170
rect 3280 70 3290 170
rect 3410 70 3420 170
rect 3594 26 3600 1774
rect 2800 20 3600 26
rect 3740 1774 4520 1780
rect 3740 26 3746 1774
rect 3920 1630 3930 1730
rect 4050 1630 4060 1730
rect 4220 1630 4230 1730
rect 4350 1630 4360 1730
rect 3800 210 3810 1570
rect 3870 210 3880 1570
rect 4100 210 4110 1570
rect 4170 210 4180 1570
rect 4400 210 4410 1570
rect 4470 210 4480 1570
rect 3920 70 3930 170
rect 4050 70 4060 170
rect 4220 70 4230 170
rect 4350 70 4360 170
rect 4514 26 4520 1774
rect 3740 20 4520 26
rect 4660 1774 5460 1780
rect 4660 26 4666 1774
rect 4840 1630 4850 1730
rect 4970 1630 4980 1730
rect 5140 1630 5150 1730
rect 5270 1630 5280 1730
rect 4720 210 4730 1570
rect 4790 210 4800 1570
rect 5020 210 5030 1570
rect 5090 210 5100 1570
rect 5320 210 5330 1570
rect 5390 210 5400 1570
rect 4840 70 4850 170
rect 4970 70 4980 170
rect 5140 70 5150 170
rect 5270 70 5280 170
rect 5454 26 5460 1774
rect 4660 20 5460 26
rect 5600 1774 6380 1780
rect 5600 26 5606 1774
rect 5760 1630 5770 1730
rect 5890 1630 5900 1730
rect 6080 1630 6090 1730
rect 6210 1630 6220 1730
rect 5650 210 5660 1570
rect 5720 210 5730 1570
rect 5950 210 5960 1570
rect 6020 210 6030 1570
rect 6250 210 6260 1570
rect 6320 210 6330 1570
rect 5760 70 5770 170
rect 5890 70 5900 170
rect 6060 70 6070 170
rect 6190 70 6200 170
rect 6374 26 6380 1774
rect 5600 20 6380 26
rect 6520 1774 7320 1780
rect 6520 26 6526 1774
rect 6700 1630 6710 1730
rect 6830 1630 6840 1730
rect 7000 1630 7010 1730
rect 7130 1630 7140 1730
rect 6590 210 6600 1570
rect 6660 210 6670 1570
rect 6890 210 6900 1570
rect 6960 210 6970 1570
rect 7190 210 7200 1570
rect 7260 210 7270 1570
rect 6700 70 6710 170
rect 6830 70 6840 170
rect 7000 70 7010 170
rect 7130 70 7140 170
rect 7314 26 7320 1774
rect 6520 20 7320 26
rect 7360 1774 7372 1926
rect 7360 26 7366 1774
rect 7360 -20 7372 26
rect -32 -26 7372 -20
rect -26 -32 26 -26
rect 794 -32 966 -26
rect 1734 -32 1886 -26
rect 2654 -32 2806 -26
rect 3594 -32 3746 -26
rect 4514 -32 4666 -26
rect 5454 -32 5606 -26
rect 6374 -32 6526 -26
rect 7314 -32 7366 -26
rect -1600 -400 -1500 -40
rect -1440 -400 -1200 -40
rect -1140 -400 -900 -40
rect -840 -400 -600 -40
rect -540 -400 -300 -40
rect -240 -140 -140 -40
rect -240 -400 7360 -140
<< via1 >>
rect -40 10400 20 10500
rect 900 10400 960 10500
rect 1840 10400 1900 10500
rect 2760 10400 2820 10500
rect 3700 10400 3760 10500
rect 4620 10400 4680 10500
rect 5560 10400 5620 10500
rect 6480 10400 6540 10500
rect 800 10200 860 10300
rect 1740 10200 1800 10300
rect 2660 10200 2720 10300
rect 3600 10200 3660 10300
rect 4520 10200 4580 10300
rect 5460 10200 5520 10300
rect 6380 10200 6440 10300
rect 7320 10200 7380 10300
rect 300 10000 500 10100
rect 1300 10000 1400 10100
rect 2200 10000 2300 10100
rect 3100 10000 3300 10100
rect 4100 10000 4200 10100
rect 5000 10000 5100 10100
rect 5900 10000 6100 10100
rect 6900 10000 7000 10100
rect -180 9800 -80 9900
rect 80 9800 140 9900
rect 1020 9800 1080 9900
rect 1940 9800 2000 9900
rect 2880 9800 2940 9900
rect 3800 9800 3860 9900
rect 4720 9800 4780 9900
rect 5660 9800 5720 9900
rect 6600 9800 6660 9900
rect -320 9600 -220 9700
rect 680 9600 740 9700
rect 1620 9600 1680 9700
rect 2540 9600 2600 9700
rect 3480 9600 3540 9700
rect 4400 9600 4460 9700
rect 5340 9600 5400 9700
rect 6260 9600 6320 9700
rect 7200 9600 7260 9700
rect 380 9460 440 9480
rect 1320 9460 1380 9480
rect 2240 9460 2300 9480
rect 3180 9460 3240 9480
rect 4100 9460 4160 9480
rect 5040 9460 5100 9480
rect 5960 9460 6020 9480
rect 6900 9460 6960 9480
rect 380 9420 440 9460
rect 1320 9420 1380 9460
rect 2240 9420 2300 9460
rect 3180 9420 3240 9460
rect 4100 9420 4160 9460
rect 5040 9420 5100 9460
rect 5960 9420 6020 9460
rect 6900 9420 6960 9460
rect 200 9280 320 9380
rect 500 9280 620 9380
rect 80 7800 140 9260
rect 380 7800 440 9260
rect 680 7800 740 9260
rect 200 7700 320 7800
rect 500 7700 620 7800
rect 1140 9280 1260 9380
rect 1420 9280 1540 9380
rect 1020 7800 1080 9260
rect 1320 7800 1380 9260
rect 1620 7800 1680 9260
rect 1140 7700 1260 7800
rect 1440 7700 1560 7800
rect 2060 9280 2180 9380
rect 2360 9280 2480 9380
rect 1940 7800 2000 9260
rect 2240 7800 2300 9260
rect 2540 7800 2600 9260
rect 2060 7700 2180 7800
rect 2360 7700 2480 7800
rect 3000 9280 3120 9380
rect 3300 9280 3420 9380
rect 2880 7800 2940 9260
rect 3180 7800 3240 9260
rect 3480 7800 3540 9260
rect 3000 7700 3120 7800
rect 3300 7700 3420 7800
rect 3920 9280 4040 9380
rect 4220 9280 4340 9380
rect 3800 7800 3860 9260
rect 4100 7800 4160 9260
rect 4400 7800 4460 9260
rect 3920 7700 4040 7800
rect 4220 7700 4340 7800
rect 4860 9280 4980 9380
rect 5160 9280 5280 9380
rect 4730 7790 4790 9250
rect 4840 7700 4960 7800
rect 5030 7790 5090 9250
rect 5160 7700 5280 7800
rect 5330 7790 5390 9250
rect 5780 9280 5900 9380
rect 6080 9280 6200 9380
rect 5660 7800 5720 9260
rect 5960 7800 6020 9260
rect 6260 7800 6320 9260
rect 5780 7700 5900 7800
rect 6080 7700 6200 7800
rect 6720 9280 6840 9380
rect 7020 9280 7140 9380
rect 6590 7800 6650 9260
rect 6890 7800 6950 9260
rect 7190 7800 7250 9260
rect 6720 7700 6840 7800
rect 7020 7700 7140 7800
rect 200 7360 320 7460
rect 500 7360 620 7460
rect 80 5890 140 7350
rect 380 5890 440 7350
rect 680 5890 740 7350
rect 200 5780 320 5880
rect 500 5780 620 5880
rect 1140 7360 1260 7460
rect 1440 7360 1560 7460
rect 1010 5900 1070 7360
rect 1310 5900 1370 7360
rect 1610 5900 1670 7360
rect 1140 5780 1260 5880
rect 1440 5780 1560 5880
rect 2060 7360 2180 7460
rect 2360 7360 2480 7460
rect 1940 5900 2000 7360
rect 2240 5900 2300 7360
rect 2540 5900 2600 7360
rect 2060 5780 2180 5880
rect 2360 5780 2480 5880
rect 3000 7360 3120 7460
rect 3280 7360 3400 7460
rect 2870 5890 2930 7350
rect 3170 5890 3230 7350
rect 3470 5890 3530 7350
rect 3000 5780 3120 5880
rect 3300 5780 3420 5880
rect 3920 7360 4040 7460
rect 4220 7360 4340 7460
rect 3800 5890 3860 7350
rect 4100 5890 4160 7350
rect 4400 5890 4460 7350
rect 3920 5780 4040 5880
rect 4220 5780 4340 5880
rect 4850 7360 4970 7460
rect 5140 7360 5260 7460
rect 4730 5890 4790 7350
rect 5030 5890 5090 7350
rect 5330 5890 5390 7350
rect 4850 5780 4970 5880
rect 5160 5780 5280 5880
rect 5780 7360 5900 7460
rect 6080 7360 6200 7460
rect 5660 5890 5720 7350
rect 5960 5890 6020 7350
rect 6260 5890 6320 7350
rect 5780 5780 5900 5880
rect 6090 5780 6210 5880
rect 6720 7360 6840 7460
rect 7020 7360 7140 7460
rect 6590 5890 6650 7350
rect 6890 5890 6950 7350
rect 7190 5890 7250 7350
rect 6710 5780 6830 5880
rect 7010 5780 7130 5880
rect 200 5460 320 5560
rect 510 5460 630 5560
rect 80 3980 140 5440
rect 190 3890 310 3990
rect 380 3980 440 5440
rect 510 3890 630 3990
rect 680 3980 740 5440
rect 1130 5460 1250 5560
rect 1440 5460 1560 5560
rect 1010 3990 1070 5450
rect 1310 3990 1370 5450
rect 1610 3990 1670 5450
rect 1130 3890 1250 3990
rect 1430 3890 1550 3990
rect 2060 5460 2180 5560
rect 2370 5460 2490 5560
rect 1940 3990 2000 5450
rect 2240 3990 2300 5450
rect 2540 3990 2600 5450
rect 2050 3890 2170 3990
rect 2350 3890 2470 3990
rect 3000 5460 3120 5560
rect 3300 5460 3420 5560
rect 2870 3980 2930 5440
rect 2990 3890 3110 3990
rect 3170 3980 3230 5440
rect 3290 3890 3410 3990
rect 3470 3980 3530 5440
rect 3930 5460 4050 5560
rect 4220 5460 4340 5560
rect 3800 3970 3860 5430
rect 3930 3890 4050 3990
rect 4100 3970 4160 5430
rect 4210 3890 4330 3990
rect 4400 3970 4460 5430
rect 4850 5460 4970 5560
rect 5160 5460 5280 5560
rect 4730 3970 4790 5430
rect 4850 3890 4970 3990
rect 5030 3970 5090 5430
rect 5150 3890 5270 3990
rect 5330 3970 5390 5430
rect 5790 5460 5910 5560
rect 6090 5460 6210 5560
rect 5660 3970 5720 5430
rect 5790 3890 5910 3990
rect 5960 3970 6020 5430
rect 6080 3880 6200 3980
rect 6260 3970 6320 5430
rect 6700 5460 6820 5560
rect 7020 5460 7140 5560
rect 6590 3980 6650 5440
rect 6890 3980 6950 5440
rect 7190 3980 7250 5440
rect 6710 3880 6830 3980
rect 7020 3880 7140 3980
rect 210 3550 330 3650
rect 510 3550 630 3650
rect 80 2080 140 3540
rect 380 2080 440 3540
rect 680 2080 740 3540
rect 190 1970 310 2070
rect 510 1970 630 2070
rect 1130 3550 1250 3650
rect 1430 3550 1550 3650
rect 1010 2080 1070 3540
rect 1310 2080 1370 3540
rect 1610 2080 1670 3540
rect 1130 1970 1250 2070
rect 1430 1970 1550 2070
rect 2070 3550 2190 3650
rect 2370 3550 2490 3650
rect 1940 2080 2000 3540
rect 2240 2080 2300 3540
rect 2540 2080 2600 3540
rect 2050 1970 2170 2070
rect 2370 1970 2490 2070
rect 2990 3550 3110 3650
rect 3310 3550 3430 3650
rect 2880 2110 2940 3470
rect 3180 2110 3240 3470
rect 3480 2110 3540 3470
rect 2990 1970 3110 2070
rect 3290 1970 3410 2070
rect 3930 3550 4050 3650
rect 4230 3550 4350 3650
rect 3800 2070 3860 3530
rect 4100 2070 4160 3530
rect 4400 2070 4460 3530
rect 3910 1970 4030 2070
rect 4230 1970 4350 2070
rect 4850 3550 4970 3650
rect 5150 3550 5270 3650
rect 4730 2070 4790 3530
rect 5030 2070 5090 3530
rect 5330 2070 5390 3530
rect 4850 1970 4970 2070
rect 5150 1970 5270 2070
rect 5790 3550 5910 3650
rect 6070 3550 6190 3650
rect 5660 2080 5720 3540
rect 5960 2080 6020 3540
rect 6260 2080 6320 3540
rect 5790 1970 5910 2070
rect 6090 1970 6210 2070
rect 6710 3550 6830 3650
rect 7010 3550 7130 3650
rect 6590 2080 6650 3540
rect 6890 2080 6950 3540
rect 7190 2080 7250 3540
rect 6710 1970 6830 2070
rect 7010 1970 7130 2070
rect -1340 1500 -1280 1600
rect -740 1500 -680 1600
rect -320 1500 -220 1600
rect -1040 1300 -980 1400
rect -460 1300 -400 1400
rect -180 1300 -80 1400
rect -1500 220 -1440 960
rect -1340 220 -1280 960
rect -1200 220 -1140 960
rect -1040 220 -980 960
rect -900 220 -840 960
rect -740 220 -680 960
rect -600 220 -540 960
rect -460 220 -400 960
rect -300 220 -240 960
rect 80 180 140 1640
rect 190 1630 310 1730
rect 380 180 440 1640
rect 510 1630 630 1730
rect 680 180 740 1640
rect 210 70 330 170
rect 510 70 630 170
rect 1130 1630 1250 1730
rect 1430 1630 1550 1730
rect 1020 210 1080 1570
rect 1320 210 1380 1570
rect 1620 210 1680 1570
rect 1130 70 1250 170
rect 1450 70 1570 170
rect 2070 1630 2190 1730
rect 2370 1630 2490 1730
rect 1940 170 2000 1630
rect 2240 170 2300 1630
rect 2540 170 2600 1630
rect 2070 70 2190 170
rect 2350 70 2470 170
rect 3010 1630 3130 1730
rect 3310 1630 3430 1730
rect 2870 210 2930 1570
rect 3170 210 3230 1570
rect 3470 210 3530 1570
rect 2990 70 3110 170
rect 3290 70 3410 170
rect 3930 1630 4050 1730
rect 4230 1630 4350 1730
rect 3810 210 3870 1570
rect 4110 210 4170 1570
rect 4410 210 4470 1570
rect 3930 70 4050 170
rect 4230 70 4350 170
rect 4850 1630 4970 1730
rect 5150 1630 5270 1730
rect 4730 210 4790 1570
rect 5030 210 5090 1570
rect 5330 210 5390 1570
rect 4850 70 4970 170
rect 5150 70 5270 170
rect 5770 1630 5890 1730
rect 6090 1630 6210 1730
rect 5660 210 5720 1570
rect 5960 210 6020 1570
rect 6260 210 6320 1570
rect 5770 70 5890 170
rect 6070 70 6190 170
rect 6710 1630 6830 1730
rect 7010 1630 7130 1730
rect 6600 210 6660 1570
rect 6900 210 6960 1570
rect 7200 210 7260 1570
rect 6710 70 6830 170
rect 7010 70 7130 170
rect -1500 -400 -1440 -40
rect -1200 -400 -1140 -40
rect -900 -400 -840 -40
rect -600 -400 -540 -40
rect -300 -400 -240 -40
<< metal2 >>
rect -40 10500 20 10510
rect 900 10500 960 10510
rect 1840 10500 1900 10510
rect 2760 10500 2820 10510
rect 3700 10500 3760 10510
rect 4620 10500 4680 10510
rect 5560 10500 5620 10510
rect 6480 10500 6540 10510
rect -180 9900 -80 9910
rect -320 9700 -220 9900
rect -1340 1600 -1280 1610
rect -740 1600 -680 1610
rect -320 1600 -220 9600
rect -1500 960 -1440 1020
rect -1500 -40 -1440 220
rect -1340 960 -1280 1500
rect -1040 1400 -980 1600
rect -1340 180 -1280 220
rect -1200 960 -1140 1020
rect -1500 -410 -1440 -400
rect -1200 -40 -1140 220
rect -1040 960 -980 1300
rect -1040 180 -980 220
rect -900 960 -840 1020
rect -1200 -410 -1140 -400
rect -900 -40 -840 220
rect -740 960 -680 1500
rect -460 1400 -400 1600
rect -320 1300 -220 1500
rect -180 1400 -80 9800
rect -740 180 -680 220
rect -600 960 -540 1020
rect -900 -410 -840 -400
rect -600 -40 -540 220
rect -460 960 -400 1300
rect -180 1290 -80 1300
rect -40 9440 20 10400
rect -40 7860 20 9380
rect -40 7520 20 7800
rect -40 5940 20 7460
rect -40 5620 20 5880
rect -40 4040 20 5560
rect -40 3700 20 3980
rect -40 2120 20 3640
rect -40 1780 20 2060
rect -460 180 -400 220
rect -300 960 -240 1020
rect -600 -410 -540 -400
rect -300 -40 -240 220
rect -40 220 20 1720
rect -40 -60 20 160
rect 80 9900 140 10500
rect 380 10110 440 10500
rect 300 10100 500 10110
rect 300 9990 500 10000
rect 80 9260 140 9800
rect 380 9480 440 9990
rect 200 9380 320 9390
rect 200 9270 320 9280
rect 380 9260 440 9420
rect 680 9700 740 10500
rect 500 9380 620 9390
rect 500 9270 620 9280
rect 80 7350 140 7800
rect 200 7800 320 7810
rect 200 7690 320 7700
rect 680 9260 740 9600
rect 200 7460 320 7470
rect 200 7350 320 7360
rect 380 7350 440 7800
rect 500 7800 620 7810
rect 500 7690 620 7700
rect 500 7460 620 7470
rect 500 7350 620 7360
rect 680 7350 740 7800
rect 80 5440 140 5890
rect 200 5880 320 5890
rect 200 5770 320 5780
rect 200 5560 320 5570
rect 200 5450 320 5460
rect 380 5440 440 5890
rect 500 5880 620 5890
rect 500 5770 620 5780
rect 510 5560 630 5570
rect 510 5450 630 5460
rect 80 3540 140 3980
rect 190 3990 310 4000
rect 190 3880 310 3890
rect 680 5440 740 5890
rect 210 3650 330 3660
rect 210 3540 330 3550
rect 380 3540 440 3980
rect 510 3990 630 4000
rect 510 3880 630 3890
rect 510 3650 630 3660
rect 510 3540 630 3550
rect 680 3540 740 3980
rect 80 1640 140 2080
rect 190 2070 310 2080
rect 190 1960 310 1970
rect 190 1730 310 1740
rect 190 1620 310 1630
rect 380 1640 440 2080
rect 510 2070 630 2080
rect 510 1960 630 1970
rect 510 1730 630 1740
rect 510 1620 630 1630
rect 680 1640 740 2080
rect 80 -60 140 180
rect 210 170 330 180
rect 210 60 330 70
rect 380 -60 440 180
rect 510 170 630 180
rect 510 60 630 70
rect 680 -60 740 180
rect 800 10300 860 10500
rect 800 9280 860 10200
rect 800 7700 860 9220
rect 800 7360 860 7640
rect 800 5780 860 7300
rect 800 5460 860 5720
rect 800 3880 860 5400
rect 800 3560 860 3820
rect 800 1980 860 3500
rect 800 1640 860 1920
rect 800 60 860 1580
rect 800 -60 860 0
rect 900 9440 960 10400
rect 900 7860 960 9380
rect 900 7520 960 7800
rect 900 5940 960 7460
rect 1020 9900 1080 10500
rect 1320 10110 1380 10500
rect 1300 10100 1400 10110
rect 1300 9990 1400 10000
rect 1020 9260 1080 9800
rect 1320 9480 1380 9990
rect 1140 9380 1260 9390
rect 1140 9270 1260 9280
rect 1320 9260 1380 9420
rect 1620 9700 1680 10500
rect 1420 9380 1540 9390
rect 1420 9270 1540 9280
rect 1020 7370 1080 7800
rect 1140 7800 1260 7810
rect 1140 7690 1260 7700
rect 1620 9260 1680 9600
rect 1010 7360 1080 7370
rect 1070 5900 1080 7360
rect 1140 7460 1260 7470
rect 1320 7370 1380 7800
rect 1440 7800 1560 7810
rect 1440 7690 1560 7700
rect 1140 7350 1260 7360
rect 1310 7360 1380 7370
rect 1010 5890 1080 5900
rect 1370 5900 1380 7360
rect 1440 7460 1560 7470
rect 1620 7370 1680 7800
rect 1440 7350 1560 7360
rect 1610 7360 1680 7370
rect 1310 5890 1380 5900
rect 1670 5900 1680 7360
rect 1610 5890 1680 5900
rect 900 5620 960 5880
rect 900 4040 960 5560
rect 1020 5460 1080 5890
rect 1140 5880 1260 5890
rect 1140 5770 1260 5780
rect 1010 5450 1080 5460
rect 1130 5560 1250 5570
rect 1320 5460 1380 5890
rect 1440 5880 1560 5890
rect 1440 5770 1560 5780
rect 1130 5450 1250 5460
rect 1310 5450 1380 5460
rect 1440 5560 1560 5570
rect 1620 5460 1680 5890
rect 1440 5450 1560 5460
rect 1610 5450 1680 5460
rect 1070 3990 1080 5450
rect 1010 3980 1080 3990
rect 900 3720 960 3980
rect 900 2140 960 3660
rect 1020 3550 1080 3980
rect 1130 3990 1250 4000
rect 1370 3990 1380 5450
rect 1310 3980 1380 3990
rect 1130 3880 1250 3890
rect 900 1800 960 2080
rect 1010 3540 1080 3550
rect 1130 3650 1250 3660
rect 1320 3550 1380 3980
rect 1430 3990 1550 4000
rect 1670 3990 1680 5450
rect 1610 3980 1680 3990
rect 1430 3880 1550 3890
rect 1130 3540 1250 3550
rect 1310 3540 1380 3550
rect 1430 3650 1550 3660
rect 1620 3550 1680 3980
rect 1430 3540 1550 3550
rect 1610 3540 1680 3550
rect 1070 2080 1080 3540
rect 1370 2080 1380 3540
rect 1670 2080 1680 3540
rect 1010 2070 1080 2080
rect 900 220 960 1740
rect 900 -60 960 160
rect 1020 1570 1080 2070
rect 1130 2070 1250 2080
rect 1310 2070 1380 2080
rect 1130 1960 1250 1970
rect 1130 1730 1250 1740
rect 1130 1620 1250 1630
rect 1020 -60 1080 210
rect 1320 1570 1380 2070
rect 1430 2070 1550 2080
rect 1610 2070 1680 2080
rect 1430 1960 1550 1970
rect 1430 1730 1550 1740
rect 1430 1620 1550 1630
rect 1130 170 1250 180
rect 1130 60 1250 70
rect 1320 -60 1380 210
rect 1620 1570 1680 2070
rect 1450 170 1570 180
rect 1450 60 1570 70
rect 1620 -60 1680 210
rect 1740 10300 1800 10500
rect 1740 9280 1800 10200
rect 1740 7700 1800 9220
rect 1740 7360 1800 7640
rect 1740 5780 1800 7300
rect 1740 5460 1800 5720
rect 1740 3880 1800 5400
rect 1740 3560 1800 3820
rect 1740 1980 1800 3500
rect 1740 1640 1800 1920
rect 1740 60 1800 1580
rect 1740 -60 1800 0
rect 1840 9440 1900 10400
rect 1840 7860 1900 9380
rect 1840 7520 1900 7800
rect 1840 5940 1900 7460
rect 1840 5620 1900 5880
rect 1840 4040 1900 5560
rect 1840 3720 1900 3980
rect 1840 2140 1900 3660
rect 1840 1800 1900 2080
rect 1840 220 1900 1740
rect 1840 -60 1900 160
rect 1940 9900 2000 10500
rect 2240 10110 2300 10500
rect 2200 10100 2300 10110
rect 2200 9990 2300 10000
rect 1940 9260 2000 9800
rect 2240 9480 2300 9990
rect 2060 9380 2180 9390
rect 2060 9270 2180 9280
rect 2240 9260 2300 9420
rect 2540 9700 2600 10500
rect 2360 9380 2480 9390
rect 2360 9270 2480 9280
rect 1940 7360 2000 7800
rect 2060 7800 2180 7810
rect 2060 7690 2180 7700
rect 2540 9260 2600 9600
rect 2060 7460 2180 7470
rect 2060 7350 2180 7360
rect 2240 7360 2300 7800
rect 2360 7800 2480 7810
rect 2360 7690 2480 7700
rect 1940 5450 2000 5900
rect 2360 7460 2480 7470
rect 2360 7350 2480 7360
rect 2540 7360 2600 7800
rect 2060 5880 2180 5890
rect 2060 5770 2180 5780
rect 2060 5560 2180 5570
rect 2060 5450 2180 5460
rect 2240 5450 2300 5900
rect 2360 5880 2480 5890
rect 2360 5770 2480 5780
rect 2370 5560 2490 5570
rect 2370 5450 2490 5460
rect 2540 5450 2600 5900
rect 1940 3540 2000 3990
rect 2050 3990 2170 4000
rect 2050 3880 2170 3890
rect 2070 3650 2190 3660
rect 2070 3540 2190 3550
rect 2240 3540 2300 3990
rect 2350 3990 2470 4000
rect 2350 3880 2470 3890
rect 2370 3650 2490 3660
rect 2370 3540 2490 3550
rect 2540 3540 2600 3990
rect 1940 1630 2000 2080
rect 2050 2070 2170 2080
rect 2050 1960 2170 1970
rect 2070 1730 2190 1740
rect 2070 1620 2190 1630
rect 2240 1630 2300 2080
rect 2370 2070 2490 2080
rect 2370 1960 2490 1970
rect 1940 -60 2000 170
rect 2070 170 2190 180
rect 2070 60 2190 70
rect 2370 1730 2490 1740
rect 2370 1620 2490 1630
rect 2540 1630 2600 2080
rect 2240 -60 2300 170
rect 2350 170 2470 180
rect 2350 60 2470 70
rect 2540 -60 2600 170
rect 2660 10300 2720 10500
rect 2660 9280 2720 10200
rect 2660 7700 2720 9220
rect 2660 7360 2720 7640
rect 2660 5780 2720 7300
rect 2660 5460 2720 5720
rect 2660 3900 2720 5400
rect 2660 3560 2720 3840
rect 2660 1980 2720 3500
rect 2660 1640 2720 1920
rect 2660 80 2720 1580
rect 2660 -60 2720 20
rect 2760 9440 2820 10400
rect 2760 7860 2820 9380
rect 2760 7520 2820 7800
rect 2760 5940 2820 7460
rect 2880 9900 2940 10500
rect 3180 10110 3240 10500
rect 3100 10100 3300 10110
rect 3100 9990 3300 10000
rect 2880 9260 2940 9800
rect 3180 9480 3240 9990
rect 3000 9380 3120 9390
rect 3000 9270 3120 9280
rect 3180 9260 3240 9420
rect 3480 9700 3540 10500
rect 3300 9380 3420 9390
rect 3300 9270 3420 9280
rect 2880 7360 2940 7800
rect 3000 7800 3120 7810
rect 3000 7690 3120 7700
rect 3480 9260 3540 9600
rect 2870 7350 2940 7360
rect 3000 7460 3120 7470
rect 3180 7360 3240 7800
rect 3300 7800 3420 7810
rect 3300 7690 3420 7700
rect 3000 7350 3120 7360
rect 3170 7350 3240 7360
rect 3280 7460 3400 7470
rect 3480 7360 3540 7800
rect 3280 7350 3400 7360
rect 3470 7350 3540 7360
rect 2930 5890 2940 7350
rect 3230 5890 3240 7350
rect 3530 5890 3540 7350
rect 2870 5880 2940 5890
rect 2760 5620 2820 5880
rect 2760 4060 2820 5560
rect 2880 5450 2940 5880
rect 3000 5880 3120 5890
rect 3170 5880 3240 5890
rect 3000 5770 3120 5780
rect 3000 5560 3120 5570
rect 3000 5450 3120 5460
rect 3180 5450 3240 5880
rect 3300 5880 3420 5890
rect 3470 5880 3540 5890
rect 3300 5770 3420 5780
rect 3300 5560 3420 5570
rect 3300 5450 3420 5460
rect 3480 5450 3540 5880
rect 2760 3720 2820 4000
rect 2870 5440 2940 5450
rect 2930 3980 2940 5440
rect 3170 5440 3240 5450
rect 2870 3970 2940 3980
rect 2760 2140 2820 3660
rect 2760 1800 2820 2080
rect 2760 240 2820 1740
rect 2880 3470 2940 3970
rect 2990 3990 3110 4000
rect 3230 3980 3240 5440
rect 3470 5440 3540 5450
rect 3170 3970 3240 3980
rect 2990 3880 3110 3890
rect 2990 3650 3110 3660
rect 2990 3540 3110 3550
rect 2880 1580 2940 2110
rect 3180 3470 3240 3970
rect 3290 3990 3410 4000
rect 3530 3980 3540 5440
rect 3470 3970 3540 3980
rect 3290 3880 3410 3890
rect 3310 3650 3430 3660
rect 3310 3540 3430 3550
rect 2990 2070 3110 2080
rect 2990 1960 3110 1970
rect 3010 1730 3130 1740
rect 3010 1620 3130 1630
rect 3180 1580 3240 2110
rect 3480 3470 3540 3970
rect 3290 2070 3410 2080
rect 3290 1960 3410 1970
rect 3310 1730 3430 1740
rect 3310 1620 3430 1630
rect 3480 1580 3540 2110
rect 2870 1570 2940 1580
rect 2930 210 2940 1570
rect 2870 200 2940 210
rect 3170 1570 3240 1580
rect 3230 210 3240 1570
rect 3170 200 3240 210
rect 3470 1570 3540 1580
rect 3530 210 3540 1570
rect 3470 200 3540 210
rect 2760 -60 2820 180
rect 2880 -60 2940 200
rect 2990 170 3110 180
rect 2990 60 3110 70
rect 3180 -40 3240 200
rect 3290 170 3410 180
rect 3290 60 3410 70
rect 3480 -60 3540 200
rect 3600 10300 3660 10500
rect 3600 9280 3660 10200
rect 3600 7700 3660 9220
rect 3600 7360 3660 7640
rect 3600 5780 3660 7300
rect 3600 5460 3660 5720
rect 3600 3900 3660 5400
rect 3600 3560 3660 3840
rect 3600 1980 3660 3500
rect 3600 1640 3660 1920
rect 3600 80 3660 1580
rect 3600 -60 3660 20
rect 3700 9440 3760 10400
rect 3700 7860 3760 9380
rect 3700 7520 3760 7800
rect 3700 5940 3760 7460
rect 3700 5620 3760 5880
rect 3700 4060 3760 5560
rect 3700 3720 3760 4000
rect 3700 2140 3760 3660
rect 3700 1800 3760 2080
rect 3700 240 3760 1740
rect 3700 -60 3760 180
rect 3800 9900 3860 10500
rect 3800 9260 3860 9800
rect 4100 10110 4160 10500
rect 4100 10100 4200 10110
rect 4100 9990 4200 10000
rect 4100 9480 4160 9990
rect 3920 9380 4040 9390
rect 3920 9270 4040 9280
rect 4100 9260 4160 9420
rect 4400 9700 4460 10500
rect 4220 9380 4340 9390
rect 4220 9270 4340 9280
rect 3800 7350 3860 7800
rect 3920 7800 4040 7810
rect 3920 7690 4040 7700
rect 4400 9260 4460 9600
rect 3920 7460 4040 7470
rect 3920 7350 4040 7360
rect 4100 7350 4160 7800
rect 4220 7800 4340 7810
rect 4220 7690 4340 7700
rect 4220 7460 4340 7470
rect 4220 7350 4340 7360
rect 4400 7350 4460 7800
rect 3800 5430 3860 5890
rect 3920 5880 4040 5890
rect 3920 5770 4040 5780
rect 3930 5560 4050 5570
rect 3930 5450 4050 5460
rect 4100 5430 4160 5890
rect 4220 5880 4340 5890
rect 4220 5770 4340 5780
rect 4220 5560 4340 5570
rect 4220 5450 4340 5460
rect 3800 3530 3860 3970
rect 3930 3990 4050 4000
rect 3930 3880 4050 3890
rect 4400 5430 4460 5890
rect 3930 3650 4050 3660
rect 3930 3540 4050 3550
rect 4100 3530 4160 3970
rect 4210 3990 4330 4000
rect 4210 3880 4330 3890
rect 4230 3650 4350 3660
rect 4230 3540 4350 3550
rect 3800 1580 3860 2070
rect 3910 2070 4030 2080
rect 3910 1960 4030 1970
rect 4400 3530 4460 3970
rect 3930 1730 4050 1740
rect 3930 1620 4050 1630
rect 4100 1580 4160 2070
rect 4230 2070 4350 2080
rect 4230 1960 4350 1970
rect 4230 1730 4350 1740
rect 4230 1620 4350 1630
rect 4400 1580 4460 2070
rect 4520 10300 4580 10500
rect 4520 9300 4580 10200
rect 4520 7700 4580 9240
rect 4520 7360 4580 7640
rect 4520 5780 4580 7300
rect 4520 5480 4580 5720
rect 4520 3900 4580 5420
rect 4520 3560 4580 3840
rect 4520 1980 4580 3500
rect 4520 1640 4580 1920
rect 3800 1570 3870 1580
rect 3800 210 3810 1570
rect 3800 200 3870 210
rect 4100 1570 4170 1580
rect 4100 210 4110 1570
rect 4100 200 4170 210
rect 4400 1570 4470 1580
rect 4400 210 4410 1570
rect 4400 200 4470 210
rect 3800 -60 3860 200
rect 3930 170 4050 180
rect 3930 60 4050 70
rect 4100 -60 4160 200
rect 4230 170 4350 180
rect 4230 60 4350 70
rect 4400 -60 4460 200
rect 4520 80 4580 1580
rect 4520 -60 4580 20
rect 4620 9460 4680 10400
rect 4620 7860 4680 9400
rect 4620 7520 4680 7800
rect 4620 5940 4680 7460
rect 4620 5640 4680 5880
rect 4620 4060 4680 5580
rect 4620 3720 4680 4000
rect 4620 2140 4680 3660
rect 4620 1800 4680 2080
rect 4620 240 4680 1740
rect 4620 -60 4680 180
rect 4720 9900 4780 10500
rect 5040 10110 5100 10500
rect 5000 10100 5100 10110
rect 5000 9990 5100 10000
rect 4720 9260 4780 9800
rect 5040 9480 5100 9990
rect 4860 9380 4980 9390
rect 4860 9270 4980 9280
rect 5040 9260 5100 9420
rect 5340 9700 5400 10500
rect 5160 9380 5280 9390
rect 5160 9270 5280 9280
rect 5340 9260 5400 9600
rect 4720 9250 4790 9260
rect 4720 7790 4730 9250
rect 5030 9250 5100 9260
rect 4720 7780 4790 7790
rect 4840 7800 4960 7810
rect 4720 7360 4780 7780
rect 5090 7790 5100 9250
rect 5330 9250 5400 9260
rect 5030 7780 5100 7790
rect 4840 7690 4960 7700
rect 4850 7460 4970 7470
rect 5040 7360 5100 7780
rect 5160 7800 5280 7810
rect 5390 7790 5400 9250
rect 5330 7780 5400 7790
rect 5160 7690 5280 7700
rect 4720 7350 4790 7360
rect 4850 7350 4970 7360
rect 5030 7350 5100 7360
rect 5140 7460 5260 7470
rect 5340 7360 5400 7780
rect 5140 7350 5260 7360
rect 5330 7350 5400 7360
rect 4720 5890 4730 7350
rect 5090 5890 5100 7350
rect 5390 5890 5400 7350
rect 4720 5880 4790 5890
rect 4850 5880 4970 5890
rect 5030 5880 5100 5890
rect 4720 5440 4780 5880
rect 4850 5770 4970 5780
rect 4850 5560 4970 5570
rect 4850 5450 4970 5460
rect 5040 5440 5100 5880
rect 5160 5880 5280 5890
rect 5330 5880 5400 5890
rect 5160 5770 5280 5780
rect 5160 5560 5280 5570
rect 5160 5450 5280 5460
rect 5340 5440 5400 5880
rect 4720 5430 4790 5440
rect 4720 3970 4730 5430
rect 5030 5430 5100 5440
rect 4720 3960 4790 3970
rect 4850 3990 4970 4000
rect 4720 3540 4780 3960
rect 5090 3970 5100 5430
rect 5330 5430 5400 5440
rect 5030 3960 5100 3970
rect 4850 3880 4970 3890
rect 4850 3650 4970 3660
rect 4850 3540 4970 3550
rect 5040 3540 5100 3960
rect 5150 3990 5270 4000
rect 5390 3970 5400 5430
rect 5330 3960 5400 3970
rect 5150 3880 5270 3890
rect 5150 3650 5270 3660
rect 5150 3540 5270 3550
rect 5340 3540 5400 3960
rect 4720 3530 4790 3540
rect 4720 2070 4730 3530
rect 5030 3530 5100 3540
rect 4720 2060 4790 2070
rect 4850 2070 4970 2080
rect 4720 1580 4780 2060
rect 5090 2070 5100 3530
rect 5330 3530 5400 3540
rect 5030 2060 5100 2070
rect 4850 1960 4970 1970
rect 4850 1730 4970 1740
rect 4850 1620 4970 1630
rect 5040 1580 5100 2060
rect 5150 2070 5270 2080
rect 5390 2070 5400 3530
rect 5330 2060 5400 2070
rect 5150 1960 5270 1970
rect 5150 1730 5270 1740
rect 5150 1620 5270 1630
rect 5340 1580 5400 2060
rect 4720 1570 4790 1580
rect 4720 210 4730 1570
rect 4720 200 4790 210
rect 5030 1570 5100 1580
rect 5090 210 5100 1570
rect 5030 200 5100 210
rect 5330 1570 5400 1580
rect 5390 210 5400 1570
rect 5330 200 5400 210
rect 4720 -60 4780 200
rect 4850 170 4970 180
rect 4850 60 4970 70
rect 5040 -60 5100 200
rect 5150 170 5270 180
rect 5150 60 5270 70
rect 5340 -60 5400 200
rect 5460 10300 5520 10500
rect 5460 9280 5520 10200
rect 5460 7700 5520 9220
rect 5460 7360 5520 7640
rect 5460 5780 5520 7300
rect 5460 5460 5520 5720
rect 5460 3900 5520 5400
rect 5460 3560 5520 3840
rect 5460 1980 5520 3500
rect 5460 1640 5520 1920
rect 5460 80 5520 1580
rect 5460 -60 5520 20
rect 5560 9440 5620 10400
rect 5560 7860 5620 9380
rect 5560 7520 5620 7800
rect 5560 5940 5620 7460
rect 5560 5620 5620 5880
rect 5560 4060 5620 5560
rect 5560 3720 5620 4000
rect 5560 2140 5620 3660
rect 5560 1800 5620 2080
rect 5560 240 5620 1740
rect 5560 -60 5620 180
rect 5660 9900 5720 10500
rect 5960 10110 6020 10500
rect 5900 10100 6100 10110
rect 5900 9990 6100 10000
rect 5660 9260 5720 9800
rect 5960 9480 6020 9990
rect 5780 9380 5900 9390
rect 5780 9270 5900 9280
rect 5960 9260 6020 9420
rect 6260 9700 6320 10500
rect 6080 9380 6200 9390
rect 6080 9270 6200 9280
rect 5660 7350 5720 7800
rect 5780 7800 5900 7810
rect 5780 7690 5900 7700
rect 6260 9260 6320 9600
rect 5780 7460 5900 7470
rect 5780 7350 5900 7360
rect 5960 7350 6020 7800
rect 6080 7800 6200 7810
rect 6080 7690 6200 7700
rect 6080 7460 6200 7470
rect 6080 7350 6200 7360
rect 6260 7350 6320 7800
rect 5660 5430 5720 5890
rect 5780 5880 5900 5890
rect 5780 5770 5900 5780
rect 5790 5560 5910 5570
rect 5790 5450 5910 5460
rect 5960 5430 6020 5890
rect 6090 5880 6210 5890
rect 6090 5770 6210 5780
rect 6090 5560 6210 5570
rect 6090 5450 6210 5460
rect 5660 3540 5720 3970
rect 5790 3990 5910 4000
rect 5790 3880 5910 3890
rect 6260 5430 6320 5890
rect 5790 3650 5910 3660
rect 5790 3540 5910 3550
rect 5960 3540 6020 3970
rect 6080 3980 6200 3990
rect 6080 3870 6200 3880
rect 6070 3650 6190 3660
rect 6070 3540 6190 3550
rect 6260 3540 6320 3970
rect 5660 1570 5720 2080
rect 5790 2070 5910 2080
rect 5790 1960 5910 1970
rect 5770 1730 5890 1740
rect 5770 1620 5890 1630
rect 5660 -60 5720 210
rect 5960 1570 6020 2080
rect 6090 2070 6210 2080
rect 6090 1960 6210 1970
rect 6090 1730 6210 1740
rect 6090 1620 6210 1630
rect 5770 170 5890 180
rect 5770 60 5890 70
rect 5960 -80 6020 210
rect 6260 1570 6320 2080
rect 6070 170 6190 180
rect 6070 60 6190 70
rect 6260 -60 6320 210
rect 6380 10300 6440 10500
rect 6380 9280 6440 10200
rect 6380 7700 6440 9220
rect 6380 7360 6440 7640
rect 6380 5780 6440 7300
rect 6380 5460 6440 5720
rect 6380 3880 6440 5400
rect 6380 3560 6440 3820
rect 6380 1980 6440 3500
rect 6380 1640 6440 1920
rect 6380 80 6440 1580
rect 6380 -60 6440 20
rect 6480 9440 6540 10400
rect 6480 7860 6540 9380
rect 6600 9900 6660 10500
rect 6600 9270 6660 9800
rect 6900 10110 6960 10500
rect 6900 10100 7000 10110
rect 6900 9990 7000 10000
rect 6900 9480 6960 9990
rect 6720 9380 6840 9390
rect 6720 9270 6840 9280
rect 6900 9270 6960 9420
rect 7200 9700 7260 10500
rect 7020 9380 7140 9390
rect 7020 9270 7140 9280
rect 7200 9270 7260 9600
rect 6480 7520 6540 7800
rect 6590 9260 6660 9270
rect 6650 7800 6660 9260
rect 6890 9260 6960 9270
rect 6590 7790 6660 7800
rect 6480 5940 6540 7460
rect 6600 7360 6660 7790
rect 6720 7800 6840 7810
rect 6950 7800 6960 9260
rect 7190 9260 7260 9270
rect 6890 7790 6960 7800
rect 6720 7690 6840 7700
rect 6590 7350 6660 7360
rect 6720 7460 6840 7470
rect 6900 7360 6960 7790
rect 7020 7800 7140 7810
rect 7250 7800 7260 9260
rect 7190 7790 7260 7800
rect 7020 7690 7140 7700
rect 6720 7350 6840 7360
rect 6890 7350 6960 7360
rect 7020 7460 7140 7470
rect 7200 7360 7260 7790
rect 7020 7350 7140 7360
rect 7190 7350 7260 7360
rect 6650 5890 6660 7350
rect 6950 5890 6960 7350
rect 7250 5890 7260 7350
rect 6590 5880 6660 5890
rect 6480 5620 6540 5880
rect 6480 4040 6540 5560
rect 6600 5450 6660 5880
rect 6710 5880 6830 5890
rect 6890 5880 6960 5890
rect 6710 5770 6830 5780
rect 6700 5560 6820 5570
rect 6700 5450 6820 5460
rect 6900 5450 6960 5880
rect 7010 5880 7130 5890
rect 7190 5880 7260 5890
rect 7010 5770 7130 5780
rect 7020 5560 7140 5570
rect 7020 5450 7140 5460
rect 7200 5450 7260 5880
rect 6480 3720 6540 3980
rect 6590 5440 6660 5450
rect 6650 3980 6660 5440
rect 6890 5440 6960 5450
rect 6590 3970 6660 3980
rect 6480 2140 6540 3660
rect 6600 3550 6660 3970
rect 6710 3980 6830 3990
rect 6950 3980 6960 5440
rect 7190 5440 7260 5450
rect 6890 3970 6960 3980
rect 6710 3870 6830 3880
rect 6480 1800 6540 2080
rect 6590 3540 6660 3550
rect 6710 3650 6830 3660
rect 6900 3550 6960 3970
rect 7020 3980 7140 3990
rect 7250 3980 7260 5440
rect 7190 3970 7260 3980
rect 7020 3870 7140 3880
rect 6710 3540 6830 3550
rect 6890 3540 6960 3550
rect 7010 3650 7130 3660
rect 7200 3550 7260 3970
rect 7010 3540 7130 3550
rect 7190 3540 7260 3550
rect 6650 2080 6660 3540
rect 6950 2080 6960 3540
rect 7250 2080 7260 3540
rect 6590 2070 6660 2080
rect 6480 240 6540 1740
rect 6480 -60 6540 180
rect 6600 1570 6660 2070
rect 6710 2070 6830 2080
rect 6890 2070 6960 2080
rect 6710 1960 6830 1970
rect 6710 1730 6830 1740
rect 6710 1620 6830 1630
rect 6600 -60 6660 210
rect 6900 1570 6960 2070
rect 7010 2070 7130 2080
rect 7190 2070 7260 2080
rect 7010 1960 7130 1970
rect 7010 1730 7130 1740
rect 7010 1620 7130 1630
rect 6710 170 6830 180
rect 6710 60 6830 70
rect 6900 -60 6960 210
rect 7200 1570 7260 2070
rect 7010 170 7130 180
rect 7010 60 7130 70
rect 7200 -60 7260 210
rect 7320 10300 7380 10500
rect 7320 9280 7380 10200
rect 7320 7700 7380 9220
rect 7320 7360 7380 7640
rect 7320 5780 7380 7300
rect 7320 5460 7380 5720
rect 7320 3880 7380 5400
rect 7320 3560 7380 3820
rect 7320 1980 7380 3500
rect 7320 1640 7380 1920
rect 7320 80 7380 1580
rect 7320 -60 7380 20
rect -300 -410 -240 -400
<< via2 >>
rect -40 9380 20 9440
rect -40 7800 20 7860
rect -40 7460 20 7520
rect -40 5880 20 5940
rect -40 5560 20 5620
rect -40 3980 20 4040
rect -40 3640 20 3700
rect -40 2060 20 2120
rect -40 1720 20 1780
rect -40 160 20 220
rect 200 9280 320 9380
rect 500 9280 620 9380
rect 200 7700 320 7800
rect 200 7360 320 7460
rect 500 7700 620 7800
rect 500 7360 620 7460
rect 200 5780 320 5880
rect 200 5460 320 5560
rect 500 5780 620 5880
rect 510 5460 630 5560
rect 190 3890 310 3990
rect 210 3550 330 3650
rect 510 3890 630 3990
rect 510 3550 630 3650
rect 190 1970 310 2070
rect 190 1630 310 1730
rect 510 1970 630 2070
rect 510 1630 630 1730
rect 210 70 330 170
rect 510 70 630 170
rect 800 9220 860 9280
rect 800 7640 860 7700
rect 800 7300 860 7360
rect 800 5720 860 5780
rect 800 5400 860 5460
rect 800 3820 860 3880
rect 800 3500 860 3560
rect 800 1920 860 1980
rect 800 1580 860 1640
rect 800 0 860 60
rect 900 9380 960 9440
rect 900 7800 960 7860
rect 900 7460 960 7520
rect 1140 9280 1260 9380
rect 1420 9280 1540 9380
rect 1140 7700 1260 7800
rect 900 5880 960 5940
rect 1140 7360 1260 7460
rect 1440 7700 1560 7800
rect 1440 7360 1560 7460
rect 900 5560 960 5620
rect 1140 5780 1260 5880
rect 900 3980 960 4040
rect 1130 5460 1250 5560
rect 1440 5780 1560 5880
rect 1440 5460 1560 5560
rect 900 3660 960 3720
rect 1130 3890 1250 3990
rect 900 2080 960 2140
rect 1130 3550 1250 3650
rect 1430 3890 1550 3990
rect 1430 3550 1550 3650
rect 900 1740 960 1800
rect 900 160 960 220
rect 1130 1970 1250 2070
rect 1130 1630 1250 1730
rect 1430 1970 1550 2070
rect 1430 1630 1550 1730
rect 1130 70 1250 170
rect 1450 70 1570 170
rect 1740 9220 1800 9280
rect 1740 7640 1800 7700
rect 1740 7300 1800 7360
rect 1740 5720 1800 5780
rect 1740 5400 1800 5460
rect 1740 3820 1800 3880
rect 1740 3500 1800 3560
rect 1740 1920 1800 1980
rect 1740 1580 1800 1640
rect 1740 0 1800 60
rect 1840 9380 1900 9440
rect 1840 7800 1900 7860
rect 1840 7460 1900 7520
rect 1840 5880 1900 5940
rect 1840 5560 1900 5620
rect 1840 3980 1900 4040
rect 1840 3660 1900 3720
rect 1840 2080 1900 2140
rect 1840 1740 1900 1800
rect 1840 160 1900 220
rect 2060 9280 2180 9380
rect 2360 9280 2480 9380
rect 2060 7700 2180 7800
rect 2060 7360 2180 7460
rect 2360 7700 2480 7800
rect 2360 7360 2480 7460
rect 2060 5780 2180 5880
rect 2060 5460 2180 5560
rect 2360 5780 2480 5880
rect 2370 5460 2490 5560
rect 2050 3890 2170 3990
rect 2070 3550 2190 3650
rect 2350 3890 2470 3990
rect 2370 3550 2490 3650
rect 2050 1970 2170 2070
rect 2070 1630 2190 1730
rect 2370 1970 2490 2070
rect 2070 70 2190 170
rect 2370 1630 2490 1730
rect 2350 70 2470 170
rect 2660 9220 2720 9280
rect 2660 7640 2720 7700
rect 2660 7300 2720 7360
rect 2660 5720 2720 5780
rect 2660 5400 2720 5460
rect 2660 3840 2720 3900
rect 2660 3500 2720 3560
rect 2660 1920 2720 1980
rect 2660 1580 2720 1640
rect 2660 20 2720 80
rect 2760 9380 2820 9440
rect 2760 7800 2820 7860
rect 2760 7460 2820 7520
rect 3000 9280 3120 9380
rect 3300 9280 3420 9380
rect 3000 7700 3120 7800
rect 2760 5880 2820 5940
rect 3000 7360 3120 7460
rect 3300 7700 3420 7800
rect 3280 7360 3400 7460
rect 2760 5560 2820 5620
rect 3000 5780 3120 5880
rect 3000 5460 3120 5560
rect 3300 5780 3420 5880
rect 3300 5460 3420 5560
rect 2760 4000 2820 4060
rect 2760 3660 2820 3720
rect 2760 2080 2820 2140
rect 2760 1740 2820 1800
rect 2990 3890 3110 3990
rect 2990 3550 3110 3650
rect 3290 3890 3410 3990
rect 3310 3550 3430 3650
rect 2990 1970 3110 2070
rect 3010 1630 3130 1730
rect 3290 1970 3410 2070
rect 3310 1630 3430 1730
rect 2760 180 2820 240
rect 2990 70 3110 170
rect 3290 70 3410 170
rect 3600 9220 3660 9280
rect 3600 7640 3660 7700
rect 3600 7300 3660 7360
rect 3600 5720 3660 5780
rect 3600 5400 3660 5460
rect 3600 3840 3660 3900
rect 3600 3500 3660 3560
rect 3600 1920 3660 1980
rect 3600 1580 3660 1640
rect 3600 20 3660 80
rect 3700 9380 3760 9440
rect 3700 7800 3760 7860
rect 3700 7460 3760 7520
rect 3700 5880 3760 5940
rect 3700 5560 3760 5620
rect 3700 4000 3760 4060
rect 3700 3660 3760 3720
rect 3700 2080 3760 2140
rect 3700 1740 3760 1800
rect 3700 180 3760 240
rect 3920 9280 4040 9380
rect 4220 9280 4340 9380
rect 3920 7700 4040 7800
rect 3920 7360 4040 7460
rect 4220 7700 4340 7800
rect 4220 7360 4340 7460
rect 3920 5780 4040 5880
rect 3930 5460 4050 5560
rect 4220 5780 4340 5880
rect 4220 5460 4340 5560
rect 3930 3890 4050 3990
rect 3930 3550 4050 3650
rect 4210 3890 4330 3990
rect 4230 3550 4350 3650
rect 3910 1970 4030 2070
rect 3930 1630 4050 1730
rect 4230 1970 4350 2070
rect 4230 1630 4350 1730
rect 4520 9240 4580 9300
rect 4520 7640 4580 7700
rect 4520 7300 4580 7360
rect 4520 5720 4580 5780
rect 4520 5420 4580 5480
rect 4520 3840 4580 3900
rect 4520 3500 4580 3560
rect 4520 1920 4580 1980
rect 4520 1580 4580 1640
rect 3930 70 4050 170
rect 4230 70 4350 170
rect 4520 20 4580 80
rect 4620 9400 4680 9460
rect 4620 7800 4680 7860
rect 4620 7460 4680 7520
rect 4620 5880 4680 5940
rect 4620 5580 4680 5640
rect 4620 4000 4680 4060
rect 4620 3660 4680 3720
rect 4620 2080 4680 2140
rect 4620 1740 4680 1800
rect 4620 180 4680 240
rect 4860 9280 4980 9380
rect 5160 9280 5280 9380
rect 4840 7700 4960 7800
rect 4850 7360 4970 7460
rect 5160 7700 5280 7800
rect 5140 7360 5260 7460
rect 4850 5780 4970 5880
rect 4850 5460 4970 5560
rect 5160 5780 5280 5880
rect 5160 5460 5280 5560
rect 4850 3890 4970 3990
rect 4850 3550 4970 3650
rect 5150 3890 5270 3990
rect 5150 3550 5270 3650
rect 4850 1970 4970 2070
rect 4850 1630 4970 1730
rect 5150 1970 5270 2070
rect 5150 1630 5270 1730
rect 4850 70 4970 170
rect 5150 70 5270 170
rect 5460 9220 5520 9280
rect 5460 7640 5520 7700
rect 5460 7300 5520 7360
rect 5460 5720 5520 5780
rect 5460 5400 5520 5460
rect 5460 3840 5520 3900
rect 5460 3500 5520 3560
rect 5460 1920 5520 1980
rect 5460 1580 5520 1640
rect 5460 20 5520 80
rect 5560 9380 5620 9440
rect 5560 7800 5620 7860
rect 5560 7460 5620 7520
rect 5560 5880 5620 5940
rect 5560 5560 5620 5620
rect 5560 4000 5620 4060
rect 5560 3660 5620 3720
rect 5560 2080 5620 2140
rect 5560 1740 5620 1800
rect 5560 180 5620 240
rect 5780 9280 5900 9380
rect 6080 9280 6200 9380
rect 5780 7700 5900 7800
rect 5780 7360 5900 7460
rect 6080 7700 6200 7800
rect 6080 7360 6200 7460
rect 5780 5780 5900 5880
rect 5790 5460 5910 5560
rect 6090 5780 6210 5880
rect 6090 5460 6210 5560
rect 5790 3890 5910 3990
rect 5790 3550 5910 3650
rect 6080 3880 6200 3980
rect 6070 3550 6190 3650
rect 5790 1970 5910 2070
rect 5770 1630 5890 1730
rect 6090 1970 6210 2070
rect 6090 1630 6210 1730
rect 5770 70 5890 170
rect 6070 70 6190 170
rect 6380 9220 6440 9280
rect 6380 7640 6440 7700
rect 6380 7300 6440 7360
rect 6380 5720 6440 5780
rect 6380 5400 6440 5460
rect 6380 3820 6440 3880
rect 6380 3500 6440 3560
rect 6380 1920 6440 1980
rect 6380 1580 6440 1640
rect 6380 20 6440 80
rect 6480 9380 6540 9440
rect 6720 9280 6840 9380
rect 7020 9280 7140 9380
rect 6480 7800 6540 7860
rect 6480 7460 6540 7520
rect 6720 7700 6840 7800
rect 6480 5880 6540 5940
rect 6720 7360 6840 7460
rect 7020 7700 7140 7800
rect 7020 7360 7140 7460
rect 6480 5560 6540 5620
rect 6710 5780 6830 5880
rect 6700 5460 6820 5560
rect 7010 5780 7130 5880
rect 7020 5460 7140 5560
rect 6480 3980 6540 4040
rect 6480 3660 6540 3720
rect 6710 3880 6830 3980
rect 6480 2080 6540 2140
rect 6710 3550 6830 3650
rect 7020 3880 7140 3980
rect 7010 3550 7130 3650
rect 6480 1740 6540 1800
rect 6480 180 6540 240
rect 6710 1970 6830 2070
rect 6710 1630 6830 1730
rect 7010 1970 7130 2070
rect 7010 1630 7130 1730
rect 6710 70 6830 170
rect 7010 70 7130 170
rect 7320 9220 7380 9280
rect 7320 7640 7380 7700
rect 7320 7300 7380 7360
rect 7320 5720 7380 5780
rect 7320 5400 7380 5460
rect 7320 3820 7380 3880
rect 7320 3500 7380 3560
rect 7320 1920 7380 1980
rect 7320 1580 7380 1640
rect 7320 20 7380 80
<< metal3 >>
rect 4610 9460 4690 9465
rect -50 9440 30 9445
rect 890 9440 970 9445
rect 1830 9440 1910 9445
rect 2750 9440 2830 9445
rect 3690 9440 3770 9445
rect -50 9380 -40 9440
rect 20 9380 340 9440
rect -50 9375 30 9380
rect 140 9320 200 9380
rect 190 9280 200 9320
rect 320 9320 340 9380
rect 490 9380 630 9385
rect 490 9340 500 9380
rect 320 9280 330 9320
rect 190 9275 330 9280
rect 480 9280 500 9340
rect 620 9340 630 9380
rect 890 9380 900 9440
rect 960 9380 1280 9440
rect 890 9375 970 9380
rect 620 9280 640 9340
rect 1120 9320 1140 9380
rect 790 9280 870 9285
rect 480 9220 800 9280
rect 860 9220 870 9280
rect 1130 9280 1140 9320
rect 1260 9320 1280 9380
rect 1410 9380 1550 9385
rect 1260 9280 1270 9320
rect 1130 9275 1270 9280
rect 1410 9280 1420 9380
rect 1540 9340 1550 9380
rect 1830 9380 1840 9440
rect 1900 9380 2220 9440
rect 1830 9375 1910 9380
rect 1540 9280 1620 9340
rect 2020 9320 2060 9380
rect 1730 9280 1810 9285
rect 1410 9275 1740 9280
rect 1420 9220 1740 9275
rect 1800 9220 1810 9280
rect 2050 9280 2060 9320
rect 2180 9320 2220 9380
rect 2350 9380 2490 9385
rect 2350 9340 2360 9380
rect 2180 9280 2190 9320
rect 2050 9275 2190 9280
rect 2340 9280 2360 9340
rect 2480 9340 2490 9380
rect 2750 9380 2760 9440
rect 2820 9380 3140 9440
rect 2750 9375 2830 9380
rect 2480 9280 2540 9340
rect 2940 9320 3000 9380
rect 2650 9280 2730 9285
rect 2340 9220 2660 9280
rect 2720 9220 2730 9280
rect 2990 9280 3000 9320
rect 3120 9320 3140 9380
rect 3290 9380 3430 9385
rect 3290 9340 3300 9380
rect 3120 9280 3130 9320
rect 2990 9275 3130 9280
rect 3280 9280 3300 9340
rect 3420 9340 3430 9380
rect 3690 9380 3700 9440
rect 3760 9380 4080 9440
rect 4610 9400 4620 9460
rect 4680 9400 5000 9460
rect 4610 9395 4690 9400
rect 3690 9375 3770 9380
rect 3420 9280 3480 9340
rect 3880 9320 3920 9380
rect 3590 9280 3670 9285
rect 3280 9220 3600 9280
rect 3660 9220 3670 9280
rect 3910 9280 3920 9320
rect 4040 9320 4080 9380
rect 4210 9380 4350 9385
rect 4210 9360 4220 9380
rect 4040 9280 4050 9320
rect 3910 9275 4050 9280
rect 4200 9280 4220 9360
rect 4340 9360 4350 9380
rect 4800 9380 5000 9400
rect 5550 9440 5630 9445
rect 6470 9440 6550 9445
rect 4340 9300 4400 9360
rect 4800 9340 4860 9380
rect 4510 9300 4590 9305
rect 4340 9280 4520 9300
rect 4200 9240 4520 9280
rect 4580 9240 4590 9300
rect 4850 9280 4860 9340
rect 4980 9340 5000 9380
rect 5150 9380 5290 9385
rect 5150 9340 5160 9380
rect 4980 9280 4990 9340
rect 4850 9275 4990 9280
rect 5140 9280 5160 9340
rect 5280 9340 5290 9380
rect 5550 9380 5560 9440
rect 5620 9380 5940 9440
rect 5550 9375 5630 9380
rect 5280 9280 5340 9340
rect 5740 9320 5780 9380
rect 5450 9280 5530 9285
rect 4510 9235 4590 9240
rect 5140 9220 5460 9280
rect 5520 9220 5530 9280
rect 5770 9280 5780 9320
rect 5900 9320 5940 9380
rect 6070 9380 6210 9385
rect 6070 9340 6080 9380
rect 5900 9280 5910 9320
rect 5770 9275 5910 9280
rect 6060 9280 6080 9340
rect 6200 9340 6210 9380
rect 6470 9380 6480 9440
rect 6540 9380 6860 9440
rect 6470 9375 6550 9380
rect 6200 9280 6260 9340
rect 6660 9320 6720 9380
rect 6370 9280 6450 9285
rect 6060 9220 6380 9280
rect 6440 9220 6450 9280
rect 6710 9280 6720 9320
rect 6840 9320 6860 9380
rect 7010 9380 7150 9385
rect 7010 9340 7020 9380
rect 6840 9280 6850 9320
rect 6710 9275 6850 9280
rect 7000 9280 7020 9340
rect 7140 9340 7150 9380
rect 7140 9280 7200 9340
rect 7310 9280 7390 9285
rect 7000 9220 7320 9280
rect 7380 9220 7390 9280
rect 790 9215 870 9220
rect 1730 9215 1810 9220
rect 2650 9215 2730 9220
rect 3590 9215 3670 9220
rect 5450 9215 5530 9220
rect 6370 9215 6450 9220
rect 7310 9215 7390 9220
rect -50 7860 30 7865
rect 890 7860 970 7865
rect 1830 7860 1910 7865
rect 2750 7860 2830 7865
rect 3690 7860 3770 7865
rect 4610 7860 4690 7865
rect 5550 7860 5630 7865
rect 6470 7860 6550 7865
rect -50 7800 -40 7860
rect 20 7800 340 7860
rect -50 7795 30 7800
rect 140 7740 200 7800
rect 190 7700 200 7740
rect 320 7740 340 7800
rect 490 7800 630 7805
rect 490 7760 500 7800
rect 320 7700 330 7740
rect 190 7695 330 7700
rect 480 7700 500 7760
rect 620 7760 630 7800
rect 890 7800 900 7860
rect 960 7800 1280 7860
rect 890 7795 970 7800
rect 620 7700 640 7760
rect 1120 7740 1140 7800
rect 790 7700 870 7705
rect 480 7640 800 7700
rect 860 7640 870 7700
rect 1130 7700 1140 7740
rect 1260 7740 1280 7800
rect 1430 7800 1570 7805
rect 1430 7760 1440 7800
rect 1260 7700 1270 7740
rect 1130 7695 1270 7700
rect 1420 7700 1440 7760
rect 1560 7760 1570 7800
rect 1830 7800 1840 7860
rect 1900 7800 2220 7860
rect 1830 7795 1910 7800
rect 1560 7700 1620 7760
rect 2020 7740 2060 7800
rect 1730 7700 1810 7705
rect 1420 7640 1740 7700
rect 1800 7640 1810 7700
rect 2050 7700 2060 7740
rect 2180 7740 2220 7800
rect 2350 7800 2490 7805
rect 2350 7760 2360 7800
rect 2180 7700 2190 7740
rect 2050 7695 2190 7700
rect 2340 7700 2360 7760
rect 2480 7760 2490 7800
rect 2750 7800 2760 7860
rect 2820 7800 3140 7860
rect 2750 7795 2830 7800
rect 2480 7700 2540 7760
rect 2940 7740 3000 7800
rect 2650 7700 2730 7705
rect 2340 7640 2660 7700
rect 2720 7640 2730 7700
rect 2990 7700 3000 7740
rect 3120 7740 3140 7800
rect 3290 7800 3430 7805
rect 3290 7760 3300 7800
rect 3120 7700 3130 7740
rect 2990 7695 3130 7700
rect 3280 7700 3300 7760
rect 3420 7760 3430 7800
rect 3690 7800 3700 7860
rect 3760 7800 4080 7860
rect 3690 7795 3770 7800
rect 3420 7700 3480 7760
rect 3880 7740 3920 7800
rect 3590 7700 3670 7705
rect 3280 7640 3600 7700
rect 3660 7640 3670 7700
rect 3910 7700 3920 7740
rect 4040 7740 4080 7800
rect 4210 7800 4350 7805
rect 4210 7760 4220 7800
rect 4040 7700 4050 7740
rect 3910 7695 4050 7700
rect 4200 7700 4220 7760
rect 4340 7760 4350 7800
rect 4610 7800 4620 7860
rect 4680 7800 5000 7860
rect 4610 7795 4690 7800
rect 4340 7700 4400 7760
rect 4800 7740 4840 7800
rect 4510 7700 4590 7705
rect 4200 7640 4520 7700
rect 4580 7640 4590 7700
rect 4830 7700 4840 7740
rect 4960 7740 5000 7800
rect 5150 7800 5290 7805
rect 5150 7760 5160 7800
rect 4960 7700 4970 7740
rect 4830 7695 4970 7700
rect 5140 7700 5160 7760
rect 5280 7760 5290 7800
rect 5550 7800 5560 7860
rect 5620 7800 5940 7860
rect 5550 7795 5630 7800
rect 5280 7700 5340 7760
rect 5740 7740 5780 7800
rect 5450 7700 5530 7705
rect 5140 7640 5460 7700
rect 5520 7640 5530 7700
rect 5770 7700 5780 7740
rect 5900 7740 5940 7800
rect 6070 7800 6210 7805
rect 6070 7760 6080 7800
rect 5900 7700 5910 7740
rect 5770 7695 5910 7700
rect 6060 7700 6080 7760
rect 6200 7760 6210 7800
rect 6470 7800 6480 7860
rect 6540 7800 6860 7860
rect 6470 7795 6550 7800
rect 6200 7700 6260 7760
rect 6660 7740 6720 7800
rect 6370 7700 6450 7705
rect 6060 7640 6380 7700
rect 6440 7640 6450 7700
rect 6710 7700 6720 7740
rect 6840 7740 6860 7800
rect 7010 7800 7150 7805
rect 7010 7760 7020 7800
rect 6840 7700 6850 7740
rect 6710 7695 6850 7700
rect 7000 7700 7020 7760
rect 7140 7760 7150 7800
rect 7140 7700 7200 7760
rect 7310 7700 7390 7705
rect 7000 7640 7320 7700
rect 7380 7640 7390 7700
rect 790 7635 870 7640
rect 1730 7635 1810 7640
rect 2650 7635 2730 7640
rect 3590 7635 3670 7640
rect 4510 7635 4590 7640
rect 5450 7635 5530 7640
rect 6370 7635 6450 7640
rect 7310 7635 7390 7640
rect -50 7520 30 7525
rect 890 7520 970 7525
rect 1830 7520 1910 7525
rect 2750 7520 2830 7525
rect 3690 7520 3770 7525
rect 4610 7520 4690 7525
rect 5550 7520 5630 7525
rect 6470 7520 6550 7525
rect -50 7460 -40 7520
rect 20 7460 340 7520
rect -50 7455 30 7460
rect 140 7400 200 7460
rect 190 7360 200 7400
rect 320 7400 340 7460
rect 490 7460 630 7465
rect 490 7420 500 7460
rect 320 7360 330 7400
rect 190 7355 330 7360
rect 480 7360 500 7420
rect 620 7420 630 7460
rect 890 7460 900 7520
rect 960 7460 1280 7520
rect 890 7455 970 7460
rect 620 7360 640 7420
rect 1120 7400 1140 7460
rect 790 7360 870 7365
rect 480 7300 800 7360
rect 860 7300 870 7360
rect 1130 7360 1140 7400
rect 1260 7400 1280 7460
rect 1430 7460 1570 7465
rect 1430 7420 1440 7460
rect 1260 7360 1270 7400
rect 1130 7355 1270 7360
rect 1420 7360 1440 7420
rect 1560 7420 1570 7460
rect 1830 7460 1840 7520
rect 1900 7460 2220 7520
rect 1830 7455 1910 7460
rect 1560 7360 1620 7420
rect 2020 7400 2060 7460
rect 1730 7360 1810 7365
rect 1420 7300 1740 7360
rect 1800 7300 1810 7360
rect 2050 7360 2060 7400
rect 2180 7400 2220 7460
rect 2350 7460 2490 7465
rect 2350 7420 2360 7460
rect 2180 7360 2190 7400
rect 2050 7355 2190 7360
rect 2340 7360 2360 7420
rect 2480 7420 2490 7460
rect 2750 7460 2760 7520
rect 2820 7460 3140 7520
rect 2750 7455 2830 7460
rect 2480 7360 2540 7420
rect 2940 7400 3000 7460
rect 2650 7360 2730 7365
rect 2340 7300 2660 7360
rect 2720 7300 2730 7360
rect 2990 7360 3000 7400
rect 3120 7400 3140 7460
rect 3270 7460 3410 7465
rect 3120 7360 3130 7400
rect 2990 7355 3130 7360
rect 3270 7360 3280 7460
rect 3400 7420 3410 7460
rect 3690 7460 3700 7520
rect 3760 7460 4080 7520
rect 3690 7455 3770 7460
rect 3400 7360 3480 7420
rect 3880 7400 3920 7460
rect 3590 7360 3670 7365
rect 3270 7355 3600 7360
rect 3280 7300 3600 7355
rect 3660 7300 3670 7360
rect 3910 7360 3920 7400
rect 4040 7400 4080 7460
rect 4210 7460 4350 7465
rect 4210 7420 4220 7460
rect 4040 7360 4050 7400
rect 3910 7355 4050 7360
rect 4200 7360 4220 7420
rect 4340 7420 4350 7460
rect 4610 7460 4620 7520
rect 4680 7460 5000 7520
rect 4610 7455 4690 7460
rect 4340 7360 4400 7420
rect 4800 7400 4850 7460
rect 4510 7360 4590 7365
rect 4200 7300 4520 7360
rect 4580 7300 4590 7360
rect 4840 7360 4850 7400
rect 4970 7400 5000 7460
rect 5130 7460 5270 7465
rect 4970 7360 4980 7400
rect 4840 7355 4980 7360
rect 5130 7360 5140 7460
rect 5260 7420 5270 7460
rect 5550 7460 5560 7520
rect 5620 7460 5940 7520
rect 5550 7455 5630 7460
rect 5260 7360 5340 7420
rect 5740 7400 5780 7460
rect 5450 7360 5530 7365
rect 5130 7355 5460 7360
rect 5140 7300 5460 7355
rect 5520 7300 5530 7360
rect 5770 7360 5780 7400
rect 5900 7400 5940 7460
rect 6070 7460 6210 7465
rect 6070 7420 6080 7460
rect 5900 7360 5910 7400
rect 5770 7355 5910 7360
rect 6060 7360 6080 7420
rect 6200 7420 6210 7460
rect 6470 7460 6480 7520
rect 6540 7460 6860 7520
rect 6470 7455 6550 7460
rect 6200 7360 6260 7420
rect 6660 7400 6720 7460
rect 6370 7360 6450 7365
rect 6060 7300 6380 7360
rect 6440 7300 6450 7360
rect 6710 7360 6720 7400
rect 6840 7400 6860 7460
rect 7010 7460 7150 7465
rect 7010 7420 7020 7460
rect 6840 7360 6850 7400
rect 6710 7355 6850 7360
rect 7000 7360 7020 7420
rect 7140 7420 7150 7460
rect 7140 7360 7200 7420
rect 7310 7360 7390 7365
rect 7000 7300 7320 7360
rect 7380 7300 7390 7360
rect 790 7295 870 7300
rect 1730 7295 1810 7300
rect 2650 7295 2730 7300
rect 3590 7295 3670 7300
rect 4510 7295 4590 7300
rect 5450 7295 5530 7300
rect 6370 7295 6450 7300
rect 7310 7295 7390 7300
rect -50 5940 30 5945
rect 890 5940 970 5945
rect 1830 5940 1910 5945
rect 2750 5940 2830 5945
rect 3690 5940 3770 5945
rect 4610 5940 4690 5945
rect 5550 5940 5630 5945
rect 6470 5940 6550 5945
rect -50 5880 -40 5940
rect 20 5880 340 5940
rect -50 5875 30 5880
rect 140 5820 200 5880
rect 190 5780 200 5820
rect 320 5820 340 5880
rect 490 5880 630 5885
rect 490 5840 500 5880
rect 320 5780 330 5820
rect 190 5775 330 5780
rect 480 5780 500 5840
rect 620 5840 630 5880
rect 890 5880 900 5940
rect 960 5880 1280 5940
rect 890 5875 970 5880
rect 620 5780 640 5840
rect 1120 5820 1140 5880
rect 790 5780 870 5785
rect 480 5720 800 5780
rect 860 5720 870 5780
rect 1130 5780 1140 5820
rect 1260 5820 1280 5880
rect 1430 5880 1570 5885
rect 1430 5840 1440 5880
rect 1260 5780 1270 5820
rect 1130 5775 1270 5780
rect 1420 5780 1440 5840
rect 1560 5840 1570 5880
rect 1830 5880 1840 5940
rect 1900 5880 2220 5940
rect 1830 5875 1910 5880
rect 1560 5780 1620 5840
rect 2020 5820 2060 5880
rect 1730 5780 1810 5785
rect 1420 5720 1740 5780
rect 1800 5720 1810 5780
rect 2050 5780 2060 5820
rect 2180 5820 2220 5880
rect 2350 5880 2490 5885
rect 2350 5840 2360 5880
rect 2180 5780 2190 5820
rect 2050 5775 2190 5780
rect 2340 5780 2360 5840
rect 2480 5840 2490 5880
rect 2750 5880 2760 5940
rect 2820 5880 3140 5940
rect 2750 5875 2830 5880
rect 2480 5780 2540 5840
rect 2940 5820 3000 5880
rect 2650 5780 2730 5785
rect 2340 5720 2660 5780
rect 2720 5720 2730 5780
rect 2990 5780 3000 5820
rect 3120 5820 3140 5880
rect 3290 5880 3430 5885
rect 3290 5840 3300 5880
rect 3120 5780 3130 5820
rect 2990 5775 3130 5780
rect 3280 5780 3300 5840
rect 3420 5840 3430 5880
rect 3690 5880 3700 5940
rect 3760 5880 4080 5940
rect 3690 5875 3770 5880
rect 3420 5780 3480 5840
rect 3880 5820 3920 5880
rect 3590 5780 3670 5785
rect 3280 5720 3600 5780
rect 3660 5720 3670 5780
rect 3910 5780 3920 5820
rect 4040 5820 4080 5880
rect 4210 5880 4350 5885
rect 4210 5840 4220 5880
rect 4040 5780 4050 5820
rect 3910 5775 4050 5780
rect 4200 5780 4220 5840
rect 4340 5840 4350 5880
rect 4610 5880 4620 5940
rect 4680 5880 5000 5940
rect 4610 5875 4690 5880
rect 4340 5780 4400 5840
rect 4800 5820 4850 5880
rect 4510 5780 4590 5785
rect 4200 5720 4520 5780
rect 4580 5720 4590 5780
rect 4840 5780 4850 5820
rect 4970 5820 5000 5880
rect 5150 5880 5290 5885
rect 5150 5840 5160 5880
rect 4970 5780 4980 5820
rect 4840 5775 4980 5780
rect 5140 5780 5160 5840
rect 5280 5840 5290 5880
rect 5550 5880 5560 5940
rect 5620 5880 5940 5940
rect 5550 5875 5630 5880
rect 5280 5780 5340 5840
rect 5740 5820 5780 5880
rect 5450 5780 5530 5785
rect 5140 5720 5460 5780
rect 5520 5720 5530 5780
rect 5770 5780 5780 5820
rect 5900 5820 5940 5880
rect 6080 5880 6220 5885
rect 6080 5840 6090 5880
rect 5900 5780 5910 5820
rect 5770 5775 5910 5780
rect 6060 5780 6090 5840
rect 6210 5840 6220 5880
rect 6470 5880 6480 5940
rect 6540 5880 6860 5940
rect 6470 5875 6550 5880
rect 6210 5780 6260 5840
rect 6660 5820 6710 5880
rect 6370 5780 6450 5785
rect 6060 5720 6380 5780
rect 6440 5720 6450 5780
rect 6700 5780 6710 5820
rect 6830 5820 6860 5880
rect 7000 5880 7140 5885
rect 6830 5780 6840 5820
rect 6700 5775 6840 5780
rect 7000 5780 7010 5880
rect 7130 5840 7140 5880
rect 7130 5780 7200 5840
rect 7310 5780 7390 5785
rect 7000 5720 7320 5780
rect 7380 5720 7390 5780
rect 790 5715 870 5720
rect 1730 5715 1810 5720
rect 2650 5715 2730 5720
rect 3590 5715 3670 5720
rect 4510 5715 4590 5720
rect 5450 5715 5530 5720
rect 6370 5715 6450 5720
rect 7310 5715 7390 5720
rect 4610 5640 4690 5645
rect -50 5620 30 5625
rect 890 5620 970 5625
rect 1830 5620 1910 5625
rect 2750 5620 2830 5625
rect 3690 5620 3770 5625
rect -50 5560 -40 5620
rect 20 5560 340 5620
rect -50 5555 30 5560
rect 140 5500 200 5560
rect 190 5460 200 5500
rect 320 5500 340 5560
rect 500 5560 640 5565
rect 500 5520 510 5560
rect 320 5460 330 5500
rect 190 5455 330 5460
rect 480 5460 510 5520
rect 630 5460 640 5560
rect 890 5560 900 5620
rect 960 5560 1280 5620
rect 890 5555 970 5560
rect 790 5460 870 5465
rect 480 5400 800 5460
rect 860 5400 870 5460
rect 1120 5460 1130 5560
rect 1250 5500 1280 5560
rect 1430 5560 1570 5565
rect 1430 5520 1440 5560
rect 1250 5460 1260 5500
rect 1120 5455 1260 5460
rect 1420 5460 1440 5520
rect 1560 5520 1570 5560
rect 1830 5560 1840 5620
rect 1900 5560 2220 5620
rect 1830 5555 1910 5560
rect 1560 5460 1620 5520
rect 2020 5500 2060 5560
rect 1730 5460 1810 5465
rect 1420 5400 1740 5460
rect 1800 5400 1810 5460
rect 2050 5460 2060 5500
rect 2180 5500 2220 5560
rect 2360 5560 2500 5565
rect 2360 5520 2370 5560
rect 2180 5460 2190 5500
rect 2050 5455 2190 5460
rect 2340 5460 2370 5520
rect 2490 5520 2500 5560
rect 2750 5560 2760 5620
rect 2820 5560 3140 5620
rect 2750 5555 2830 5560
rect 2490 5460 2540 5520
rect 2940 5500 3000 5560
rect 2650 5460 2730 5465
rect 2340 5400 2660 5460
rect 2720 5400 2730 5460
rect 2990 5460 3000 5500
rect 3120 5500 3140 5560
rect 3290 5560 3430 5565
rect 3290 5520 3300 5560
rect 3120 5460 3130 5500
rect 2990 5455 3130 5460
rect 3280 5460 3300 5520
rect 3420 5520 3430 5560
rect 3690 5560 3700 5620
rect 3760 5560 4080 5620
rect 4610 5580 4620 5640
rect 4680 5580 5000 5640
rect 4610 5575 4690 5580
rect 3690 5555 3770 5560
rect 3420 5460 3480 5520
rect 3880 5500 3930 5560
rect 3590 5460 3670 5465
rect 3280 5400 3600 5460
rect 3660 5400 3670 5460
rect 3920 5460 3930 5500
rect 4050 5500 4080 5560
rect 4210 5560 4350 5565
rect 4210 5540 4220 5560
rect 4050 5460 4060 5500
rect 3920 5455 4060 5460
rect 4200 5460 4220 5540
rect 4340 5540 4350 5560
rect 4800 5560 5000 5580
rect 5550 5620 5630 5625
rect 6470 5620 6550 5625
rect 4340 5480 4400 5540
rect 4800 5520 4850 5560
rect 4510 5480 4590 5485
rect 4340 5460 4520 5480
rect 4200 5420 4520 5460
rect 4580 5420 4590 5480
rect 4840 5460 4850 5520
rect 4970 5520 5000 5560
rect 5150 5560 5290 5565
rect 5150 5520 5160 5560
rect 4970 5460 4980 5520
rect 4840 5455 4980 5460
rect 5140 5460 5160 5520
rect 5280 5520 5290 5560
rect 5550 5560 5560 5620
rect 5620 5560 5940 5620
rect 5550 5555 5630 5560
rect 5280 5460 5340 5520
rect 5740 5500 5790 5560
rect 5450 5460 5530 5465
rect 4510 5415 4590 5420
rect 5140 5400 5460 5460
rect 5520 5400 5530 5460
rect 5780 5460 5790 5500
rect 5910 5500 5940 5560
rect 6080 5560 6220 5565
rect 6080 5520 6090 5560
rect 5910 5460 5920 5500
rect 5780 5455 5920 5460
rect 6060 5460 6090 5520
rect 6210 5520 6220 5560
rect 6470 5560 6480 5620
rect 6540 5560 6860 5620
rect 6470 5555 6550 5560
rect 6210 5460 6260 5520
rect 6660 5500 6700 5560
rect 6370 5460 6450 5465
rect 6060 5400 6380 5460
rect 6440 5400 6450 5460
rect 6690 5460 6700 5500
rect 6820 5500 6860 5560
rect 7010 5560 7150 5565
rect 7010 5520 7020 5560
rect 6820 5460 6830 5500
rect 6690 5455 6830 5460
rect 7000 5460 7020 5520
rect 7140 5520 7150 5560
rect 7140 5460 7200 5520
rect 7310 5460 7390 5465
rect 7000 5400 7320 5460
rect 7380 5400 7390 5460
rect 790 5395 870 5400
rect 1730 5395 1810 5400
rect 2650 5395 2730 5400
rect 3590 5395 3670 5400
rect 5450 5395 5530 5400
rect 6370 5395 6450 5400
rect 7310 5395 7390 5400
rect 2750 4060 2830 4065
rect 3690 4060 3770 4065
rect 4610 4060 4690 4065
rect 5550 4060 5630 4065
rect -50 4040 30 4045
rect 890 4040 970 4045
rect 1830 4040 1910 4045
rect -50 3980 -40 4040
rect 20 3990 340 4040
rect 20 3980 190 3990
rect -50 3975 30 3980
rect 140 3920 190 3980
rect 180 3890 190 3920
rect 310 3920 340 3990
rect 500 3990 640 3995
rect 500 3940 510 3990
rect 310 3890 320 3920
rect 180 3885 320 3890
rect 480 3890 510 3940
rect 630 3890 640 3990
rect 890 3980 900 4040
rect 960 3990 1280 4040
rect 960 3980 1130 3990
rect 890 3975 970 3980
rect 480 3880 640 3890
rect 1120 3890 1130 3980
rect 1250 3920 1280 3990
rect 1420 3990 1560 3995
rect 1250 3890 1260 3920
rect 1120 3885 1260 3890
rect 1420 3890 1430 3990
rect 1550 3940 1560 3990
rect 1830 3980 1840 4040
rect 1900 3990 2220 4040
rect 2750 4000 2760 4060
rect 2820 4000 3140 4060
rect 2750 3995 2830 4000
rect 1900 3980 2050 3990
rect 1830 3975 1910 3980
rect 1550 3890 1620 3940
rect 2020 3920 2050 3980
rect 790 3880 870 3885
rect 480 3820 800 3880
rect 860 3820 870 3880
rect 1420 3880 1620 3890
rect 2040 3890 2050 3920
rect 2170 3920 2220 3990
rect 2340 3990 2480 3995
rect 2170 3890 2180 3920
rect 2040 3885 2180 3890
rect 2340 3890 2350 3990
rect 2470 3960 2480 3990
rect 2940 3990 3140 4000
rect 3690 4000 3700 4060
rect 3760 4000 4080 4060
rect 3690 3995 3770 4000
rect 2470 3900 2540 3960
rect 2940 3940 2990 3990
rect 2650 3900 2730 3905
rect 2470 3890 2660 3900
rect 1730 3880 1810 3885
rect 1420 3820 1740 3880
rect 1800 3820 1810 3880
rect 2340 3840 2660 3890
rect 2720 3840 2730 3900
rect 2980 3890 2990 3940
rect 3110 3940 3140 3990
rect 3280 3990 3420 3995
rect 3110 3890 3120 3940
rect 2980 3885 3120 3890
rect 3280 3890 3290 3990
rect 3410 3960 3420 3990
rect 3880 3990 4080 4000
rect 4610 4000 4620 4060
rect 4680 4000 5000 4060
rect 4610 3995 4690 4000
rect 3410 3900 3480 3960
rect 3880 3940 3930 3990
rect 3590 3900 3670 3905
rect 3410 3890 3600 3900
rect 3280 3840 3600 3890
rect 3660 3840 3670 3900
rect 3920 3890 3930 3940
rect 4050 3940 4080 3990
rect 4200 3990 4340 3995
rect 4050 3890 4060 3940
rect 3920 3885 4060 3890
rect 4200 3890 4210 3990
rect 4330 3960 4340 3990
rect 4800 3990 5000 4000
rect 5550 4000 5560 4060
rect 5620 4000 5940 4060
rect 5550 3995 5630 4000
rect 4330 3900 4400 3960
rect 4800 3940 4850 3990
rect 4510 3900 4590 3905
rect 4330 3890 4520 3900
rect 4200 3840 4520 3890
rect 4580 3840 4590 3900
rect 4840 3890 4850 3940
rect 4970 3940 5000 3990
rect 5140 3990 5280 3995
rect 4970 3890 4980 3940
rect 4840 3885 4980 3890
rect 5140 3890 5150 3990
rect 5270 3960 5280 3990
rect 5740 3990 5940 4000
rect 5270 3900 5340 3960
rect 5740 3940 5790 3990
rect 5450 3900 5530 3905
rect 5270 3890 5460 3900
rect 5140 3840 5460 3890
rect 5520 3840 5530 3900
rect 5780 3890 5790 3940
rect 5910 3940 5940 3990
rect 6470 4040 6550 4045
rect 6070 3980 6210 3985
rect 6070 3940 6080 3980
rect 5910 3890 5920 3940
rect 5780 3885 5920 3890
rect 2650 3835 2730 3840
rect 3590 3835 3670 3840
rect 4510 3835 4590 3840
rect 5450 3835 5530 3840
rect 6060 3880 6080 3940
rect 6200 3940 6210 3980
rect 6470 3980 6480 4040
rect 6540 3980 6860 4040
rect 6470 3975 6550 3980
rect 6200 3880 6260 3940
rect 6660 3920 6710 3980
rect 6370 3880 6450 3885
rect 6060 3820 6380 3880
rect 6440 3820 6450 3880
rect 6700 3880 6710 3920
rect 6830 3920 6860 3980
rect 7010 3980 7150 3985
rect 7010 3940 7020 3980
rect 6830 3880 6840 3920
rect 6700 3875 6840 3880
rect 7000 3880 7020 3940
rect 7140 3940 7150 3980
rect 7140 3880 7200 3940
rect 7310 3880 7390 3885
rect 7000 3820 7320 3880
rect 7380 3820 7390 3880
rect 790 3815 870 3820
rect 1730 3815 1810 3820
rect 6370 3815 6450 3820
rect 7310 3815 7390 3820
rect 890 3720 970 3725
rect 1830 3720 1910 3725
rect 2750 3720 2830 3725
rect 3690 3720 3770 3725
rect 4610 3720 4690 3725
rect 5550 3720 5630 3725
rect 6470 3720 6550 3725
rect -50 3700 30 3705
rect -50 3640 -40 3700
rect 20 3650 340 3700
rect 890 3660 900 3720
rect 960 3660 1280 3720
rect 890 3655 970 3660
rect 20 3640 210 3650
rect -50 3635 30 3640
rect 140 3580 210 3640
rect 200 3550 210 3580
rect 330 3550 340 3650
rect 500 3650 640 3655
rect 500 3620 510 3650
rect 200 3545 340 3550
rect 480 3550 510 3620
rect 630 3560 640 3650
rect 1120 3650 1280 3660
rect 1830 3660 1840 3720
rect 1900 3660 2220 3720
rect 1830 3655 1910 3660
rect 790 3560 870 3565
rect 630 3550 800 3560
rect 480 3500 800 3550
rect 860 3500 870 3560
rect 1120 3550 1130 3650
rect 1250 3600 1280 3650
rect 1420 3650 1560 3655
rect 1250 3550 1260 3600
rect 1120 3545 1260 3550
rect 1420 3550 1430 3650
rect 1550 3620 1560 3650
rect 2020 3650 2220 3660
rect 2750 3660 2760 3720
rect 2820 3660 3140 3720
rect 2750 3655 2830 3660
rect 1550 3560 1620 3620
rect 2020 3600 2070 3650
rect 1730 3560 1810 3565
rect 1550 3550 1740 3560
rect 1420 3500 1740 3550
rect 1800 3500 1810 3560
rect 2060 3550 2070 3600
rect 2190 3600 2220 3650
rect 2360 3650 2500 3655
rect 2360 3620 2370 3650
rect 2190 3550 2200 3600
rect 2060 3545 2200 3550
rect 2340 3550 2370 3620
rect 2490 3620 2500 3650
rect 2940 3650 3140 3660
rect 3690 3660 3700 3720
rect 3760 3660 4080 3720
rect 3690 3655 3770 3660
rect 2490 3560 2540 3620
rect 2940 3600 2990 3650
rect 2650 3560 2730 3565
rect 2490 3550 2660 3560
rect 2340 3500 2660 3550
rect 2720 3500 2730 3560
rect 2980 3550 2990 3600
rect 3110 3600 3140 3650
rect 3300 3650 3440 3655
rect 3300 3620 3310 3650
rect 3110 3550 3120 3600
rect 2980 3545 3120 3550
rect 3280 3550 3310 3620
rect 3430 3620 3440 3650
rect 3880 3650 4080 3660
rect 4610 3660 4620 3720
rect 4680 3660 5000 3720
rect 4610 3655 4690 3660
rect 3430 3560 3480 3620
rect 3880 3600 3930 3650
rect 3590 3560 3670 3565
rect 3430 3550 3600 3560
rect 3280 3500 3600 3550
rect 3660 3500 3670 3560
rect 3920 3550 3930 3600
rect 4050 3600 4080 3650
rect 4220 3650 4360 3655
rect 4220 3620 4230 3650
rect 4050 3550 4060 3600
rect 3920 3545 4060 3550
rect 4200 3550 4230 3620
rect 4350 3620 4360 3650
rect 4800 3650 5000 3660
rect 5550 3660 5560 3720
rect 5620 3660 5940 3720
rect 5550 3655 5630 3660
rect 4350 3560 4400 3620
rect 4800 3600 4850 3650
rect 4510 3560 4590 3565
rect 4350 3550 4520 3560
rect 4200 3500 4520 3550
rect 4580 3500 4590 3560
rect 4840 3550 4850 3600
rect 4970 3600 5000 3650
rect 5140 3650 5280 3655
rect 4970 3550 4980 3600
rect 4840 3545 4980 3550
rect 5140 3550 5150 3650
rect 5270 3620 5280 3650
rect 5740 3650 5940 3660
rect 6470 3660 6480 3720
rect 6540 3660 6860 3720
rect 6470 3655 6550 3660
rect 5270 3560 5340 3620
rect 5740 3600 5790 3650
rect 5450 3560 5530 3565
rect 5270 3550 5460 3560
rect 5140 3500 5460 3550
rect 5520 3500 5530 3560
rect 5780 3550 5790 3600
rect 5910 3600 5940 3650
rect 6060 3650 6200 3655
rect 5910 3550 5920 3600
rect 5780 3545 5920 3550
rect 6060 3550 6070 3650
rect 6190 3620 6200 3650
rect 6660 3650 6860 3660
rect 6190 3560 6260 3620
rect 6660 3600 6710 3650
rect 6370 3560 6450 3565
rect 6190 3550 6380 3560
rect 6060 3500 6380 3550
rect 6440 3500 6450 3560
rect 6700 3550 6710 3600
rect 6830 3600 6860 3650
rect 7000 3650 7140 3655
rect 6830 3550 6840 3600
rect 6700 3545 6840 3550
rect 7000 3550 7010 3650
rect 7130 3620 7140 3650
rect 7130 3560 7200 3620
rect 7310 3560 7390 3565
rect 7130 3550 7320 3560
rect 7000 3500 7320 3550
rect 7380 3500 7390 3560
rect 790 3495 870 3500
rect 1730 3495 1810 3500
rect 2650 3495 2730 3500
rect 3590 3495 3670 3500
rect 4510 3495 4590 3500
rect 5450 3495 5530 3500
rect 6370 3495 6450 3500
rect 7310 3495 7390 3500
rect 890 2140 970 2145
rect 1830 2140 1910 2145
rect 2750 2140 2830 2145
rect 3690 2140 3770 2145
rect 4610 2140 4690 2145
rect 5550 2140 5630 2145
rect 6470 2140 6550 2145
rect -50 2120 30 2125
rect -50 2060 -40 2120
rect 20 2070 340 2120
rect 890 2080 900 2140
rect 960 2080 1280 2140
rect 890 2075 970 2080
rect 20 2060 190 2070
rect -50 2055 30 2060
rect 140 2000 190 2060
rect 180 1970 190 2000
rect 310 2000 340 2070
rect 500 2070 640 2075
rect 500 2040 510 2070
rect 310 1970 320 2000
rect 180 1965 320 1970
rect 480 1970 510 2040
rect 630 1980 640 2070
rect 1120 2070 1280 2080
rect 1830 2080 1840 2140
rect 1900 2080 2220 2140
rect 1830 2075 1910 2080
rect 790 1980 870 1985
rect 630 1970 800 1980
rect 480 1920 800 1970
rect 860 1920 870 1980
rect 1120 1970 1130 2070
rect 1250 2020 1280 2070
rect 1420 2070 1560 2075
rect 1250 1970 1260 2020
rect 1120 1965 1260 1970
rect 1420 1970 1430 2070
rect 1550 2040 1560 2070
rect 2020 2070 2220 2080
rect 2750 2080 2760 2140
rect 2820 2080 3140 2140
rect 2750 2075 2830 2080
rect 1550 1980 1620 2040
rect 2020 2020 2050 2070
rect 1730 1980 1810 1985
rect 1550 1970 1740 1980
rect 1420 1920 1740 1970
rect 1800 1920 1810 1980
rect 2040 1970 2050 2020
rect 2170 2020 2220 2070
rect 2360 2070 2500 2075
rect 2360 2040 2370 2070
rect 2170 1970 2180 2020
rect 2040 1965 2180 1970
rect 2340 1970 2370 2040
rect 2490 2040 2500 2070
rect 2940 2070 3140 2080
rect 3690 2080 3700 2140
rect 3760 2080 4080 2140
rect 3690 2075 3770 2080
rect 2490 1980 2540 2040
rect 2940 2020 2990 2070
rect 2650 1980 2730 1985
rect 2490 1970 2660 1980
rect 2340 1920 2660 1970
rect 2720 1920 2730 1980
rect 2980 1970 2990 2020
rect 3110 2020 3140 2070
rect 3280 2070 3420 2075
rect 3110 1970 3120 2020
rect 2980 1965 3120 1970
rect 3280 1970 3290 2070
rect 3410 2040 3420 2070
rect 3880 2070 4080 2080
rect 4610 2080 4620 2140
rect 4680 2080 5000 2140
rect 4610 2075 4690 2080
rect 3410 1980 3480 2040
rect 3880 2020 3910 2070
rect 3590 1980 3670 1985
rect 3410 1970 3600 1980
rect 3280 1920 3600 1970
rect 3660 1920 3670 1980
rect 3900 1970 3910 2020
rect 4030 2020 4080 2070
rect 4220 2070 4360 2075
rect 4220 2040 4230 2070
rect 4030 1970 4040 2020
rect 3900 1965 4040 1970
rect 4200 1970 4230 2040
rect 4350 2040 4360 2070
rect 4800 2070 5000 2080
rect 5550 2080 5560 2140
rect 5620 2080 5940 2140
rect 5550 2075 5630 2080
rect 4350 1980 4400 2040
rect 4800 2020 4850 2070
rect 4510 1980 4590 1985
rect 4350 1970 4520 1980
rect 4200 1920 4520 1970
rect 4580 1920 4590 1980
rect 4840 1970 4850 2020
rect 4970 2020 5000 2070
rect 5140 2070 5280 2075
rect 4970 1970 4980 2020
rect 4840 1965 4980 1970
rect 5140 1970 5150 2070
rect 5270 2040 5280 2070
rect 5740 2070 5940 2080
rect 6470 2080 6480 2140
rect 6540 2080 6860 2140
rect 6470 2075 6550 2080
rect 5270 1980 5340 2040
rect 5740 2020 5790 2070
rect 5450 1980 5530 1985
rect 5270 1970 5460 1980
rect 5140 1920 5460 1970
rect 5520 1920 5530 1980
rect 5780 1970 5790 2020
rect 5910 2020 5940 2070
rect 6080 2070 6220 2075
rect 6080 2040 6090 2070
rect 5910 1970 5920 2020
rect 5780 1965 5920 1970
rect 6060 1970 6090 2040
rect 6210 2040 6220 2070
rect 6660 2070 6860 2080
rect 6210 1980 6260 2040
rect 6660 2020 6710 2070
rect 6370 1980 6450 1985
rect 6210 1970 6380 1980
rect 6060 1920 6380 1970
rect 6440 1920 6450 1980
rect 6700 1970 6710 2020
rect 6830 2020 6860 2070
rect 7000 2070 7140 2075
rect 6830 1970 6840 2020
rect 6700 1965 6840 1970
rect 7000 1970 7010 2070
rect 7130 2040 7140 2070
rect 7130 1980 7200 2040
rect 7310 1980 7390 1985
rect 7130 1970 7320 1980
rect 7000 1920 7320 1970
rect 7380 1920 7390 1980
rect 790 1915 870 1920
rect 1730 1915 1810 1920
rect 2650 1915 2730 1920
rect 3590 1915 3670 1920
rect 4510 1915 4590 1920
rect 5450 1915 5530 1920
rect 6370 1915 6450 1920
rect 7310 1915 7390 1920
rect 890 1800 970 1805
rect 1830 1800 1910 1805
rect 2750 1800 2830 1805
rect 3690 1800 3770 1805
rect 4610 1800 4690 1805
rect 5550 1800 5630 1805
rect 6470 1800 6550 1805
rect -50 1780 30 1785
rect -50 1720 -40 1780
rect 20 1730 340 1780
rect 890 1740 900 1800
rect 960 1740 1280 1800
rect 890 1735 970 1740
rect 20 1720 190 1730
rect -50 1715 30 1720
rect 140 1660 190 1720
rect 180 1630 190 1660
rect 310 1660 340 1730
rect 500 1730 640 1735
rect 500 1700 510 1730
rect 310 1630 320 1660
rect 180 1625 320 1630
rect 480 1630 510 1700
rect 630 1640 640 1730
rect 1120 1730 1280 1740
rect 1830 1740 1840 1800
rect 1900 1740 2220 1800
rect 1830 1735 1910 1740
rect 790 1640 870 1645
rect 630 1630 800 1640
rect 480 1580 800 1630
rect 860 1580 870 1640
rect 1120 1630 1130 1730
rect 1250 1680 1280 1730
rect 1420 1730 1560 1735
rect 1250 1630 1260 1680
rect 1120 1625 1260 1630
rect 1420 1630 1430 1730
rect 1550 1700 1560 1730
rect 2060 1730 2220 1740
rect 2750 1740 2760 1800
rect 2820 1740 3140 1800
rect 2750 1735 2830 1740
rect 1550 1640 1580 1700
rect 1730 1640 1810 1645
rect 1550 1630 1740 1640
rect 1420 1580 1740 1630
rect 1800 1580 1810 1640
rect 2060 1630 2070 1730
rect 2190 1680 2220 1730
rect 2360 1730 2500 1735
rect 2360 1700 2370 1730
rect 2190 1630 2200 1680
rect 2060 1625 2200 1630
rect 2340 1630 2370 1700
rect 2490 1700 2500 1730
rect 2940 1730 3140 1740
rect 3690 1740 3700 1800
rect 3760 1740 4080 1800
rect 3690 1735 3770 1740
rect 2490 1640 2540 1700
rect 2940 1680 3010 1730
rect 2650 1640 2730 1645
rect 2490 1630 2660 1640
rect 2340 1580 2660 1630
rect 2720 1580 2730 1640
rect 3000 1630 3010 1680
rect 3130 1630 3140 1730
rect 3300 1730 3440 1735
rect 3300 1700 3310 1730
rect 3000 1625 3140 1630
rect 3280 1630 3310 1700
rect 3430 1700 3440 1730
rect 3880 1730 4080 1740
rect 4610 1740 4620 1800
rect 4680 1740 5000 1800
rect 4610 1735 4690 1740
rect 3430 1640 3480 1700
rect 3880 1680 3930 1730
rect 3590 1640 3670 1645
rect 3430 1630 3600 1640
rect 3280 1580 3600 1630
rect 3660 1580 3670 1640
rect 3920 1630 3930 1680
rect 4050 1680 4080 1730
rect 4220 1730 4360 1735
rect 4220 1700 4230 1730
rect 4050 1630 4060 1680
rect 3920 1625 4060 1630
rect 4200 1630 4230 1700
rect 4350 1700 4360 1730
rect 4800 1730 5000 1740
rect 5550 1740 5560 1800
rect 5620 1740 5940 1800
rect 5550 1735 5630 1740
rect 4350 1640 4400 1700
rect 4800 1680 4850 1730
rect 4510 1640 4590 1645
rect 4350 1630 4520 1640
rect 4200 1580 4520 1630
rect 4580 1580 4590 1640
rect 4840 1630 4850 1680
rect 4970 1680 5000 1730
rect 5140 1730 5280 1735
rect 4970 1630 4980 1680
rect 4840 1625 4980 1630
rect 5140 1630 5150 1730
rect 5270 1700 5280 1730
rect 5740 1730 5940 1740
rect 6470 1740 6480 1800
rect 6540 1740 6860 1800
rect 6470 1735 6550 1740
rect 5270 1640 5340 1700
rect 5740 1680 5770 1730
rect 5450 1640 5530 1645
rect 5270 1630 5460 1640
rect 5140 1580 5460 1630
rect 5520 1580 5530 1640
rect 5760 1630 5770 1680
rect 5890 1680 5940 1730
rect 6080 1730 6220 1735
rect 6080 1700 6090 1730
rect 5890 1630 5900 1680
rect 5760 1625 5900 1630
rect 6060 1630 6090 1700
rect 6210 1700 6220 1730
rect 6660 1730 6860 1740
rect 6210 1640 6260 1700
rect 6660 1680 6710 1730
rect 6370 1640 6450 1645
rect 6210 1630 6380 1640
rect 6060 1580 6380 1630
rect 6440 1580 6450 1640
rect 6700 1630 6710 1680
rect 6830 1680 6860 1730
rect 7000 1730 7140 1735
rect 6830 1630 6840 1680
rect 6700 1625 6840 1630
rect 7000 1630 7010 1730
rect 7130 1700 7140 1730
rect 7130 1640 7200 1700
rect 7310 1640 7390 1645
rect 7130 1630 7320 1640
rect 7000 1580 7320 1630
rect 7380 1580 7390 1640
rect 790 1575 870 1580
rect 1730 1575 1810 1580
rect 2650 1575 2730 1580
rect 3590 1575 3670 1580
rect 4510 1575 4590 1580
rect 5450 1575 5530 1580
rect 6370 1575 6450 1580
rect 7310 1575 7390 1580
rect 2750 240 2830 245
rect 3690 240 3770 245
rect 4610 240 4690 245
rect 5550 240 5630 245
rect 6470 240 6550 245
rect -50 220 30 225
rect 890 220 970 225
rect 1830 220 1910 225
rect -50 160 -40 220
rect 20 170 340 220
rect 20 160 210 170
rect -50 155 30 160
rect 140 100 210 160
rect 200 70 210 100
rect 330 70 340 170
rect 500 170 640 175
rect 500 120 510 170
rect 200 65 340 70
rect 480 70 510 120
rect 630 70 640 170
rect 890 160 900 220
rect 960 170 1280 220
rect 960 160 1130 170
rect 890 155 970 160
rect 480 60 640 70
rect 1120 70 1130 160
rect 1250 100 1280 170
rect 1440 170 1580 175
rect 1440 120 1450 170
rect 1250 70 1260 100
rect 1120 65 1260 70
rect 1420 70 1450 120
rect 1570 70 1580 170
rect 1830 160 1840 220
rect 1900 170 2220 220
rect 2750 180 2760 240
rect 2820 180 3140 240
rect 2750 175 2830 180
rect 1900 160 2070 170
rect 1830 155 1910 160
rect 790 60 870 65
rect 480 0 800 60
rect 860 0 870 60
rect 1420 60 1580 70
rect 2060 70 2070 160
rect 2190 100 2220 170
rect 2340 170 2480 175
rect 2190 70 2200 100
rect 2060 65 2200 70
rect 2340 70 2350 170
rect 2470 140 2480 170
rect 2940 170 3140 180
rect 3690 180 3700 240
rect 3760 180 4080 240
rect 3690 175 3770 180
rect 2470 80 2540 140
rect 2940 120 2990 170
rect 2650 80 2730 85
rect 2470 70 2660 80
rect 1730 60 1810 65
rect 1420 0 1740 60
rect 1800 0 1810 60
rect 2340 20 2660 70
rect 2720 20 2730 80
rect 2980 70 2990 120
rect 3110 120 3140 170
rect 3280 170 3420 175
rect 3110 70 3120 120
rect 2980 65 3120 70
rect 3280 70 3290 170
rect 3410 140 3420 170
rect 3880 170 4080 180
rect 4610 180 4620 240
rect 4680 180 5000 240
rect 4610 175 4690 180
rect 3410 80 3480 140
rect 3880 120 3930 170
rect 3590 80 3670 85
rect 3410 70 3600 80
rect 3280 20 3600 70
rect 3660 20 3670 80
rect 3920 70 3930 120
rect 4050 120 4080 170
rect 4220 170 4360 175
rect 4220 140 4230 170
rect 4050 70 4060 120
rect 3920 65 4060 70
rect 4200 70 4230 140
rect 4350 140 4360 170
rect 4800 170 5000 180
rect 5550 180 5560 240
rect 5620 180 5940 240
rect 5550 175 5630 180
rect 4350 80 4400 140
rect 4800 120 4850 170
rect 4510 80 4590 85
rect 4350 70 4520 80
rect 4200 20 4520 70
rect 4580 20 4590 80
rect 4840 70 4850 120
rect 4970 120 5000 170
rect 5140 170 5280 175
rect 4970 70 4980 120
rect 4840 65 4980 70
rect 5140 70 5150 170
rect 5270 140 5280 170
rect 5740 170 5940 180
rect 6470 180 6480 240
rect 6540 180 6860 240
rect 6470 175 6550 180
rect 5270 80 5340 140
rect 5740 120 5770 170
rect 5450 80 5530 85
rect 5270 70 5460 80
rect 5140 20 5460 70
rect 5520 20 5530 80
rect 5760 70 5770 120
rect 5890 120 5940 170
rect 6060 170 6200 175
rect 5890 70 5900 120
rect 5760 65 5900 70
rect 6060 70 6070 170
rect 6190 140 6200 170
rect 6660 170 6860 180
rect 6190 80 6260 140
rect 6660 120 6710 170
rect 6370 80 6450 85
rect 6190 70 6380 80
rect 6060 20 6380 70
rect 6440 20 6450 80
rect 6700 70 6710 120
rect 6830 120 6860 170
rect 7000 170 7140 175
rect 6830 70 6840 120
rect 6700 65 6840 70
rect 7000 70 7010 170
rect 7130 140 7140 170
rect 7130 80 7200 140
rect 7310 80 7390 85
rect 7130 70 7320 80
rect 7000 20 7320 70
rect 7380 20 7390 80
rect 2650 15 2730 20
rect 3590 15 3670 20
rect 4510 15 4590 20
rect 5450 15 5530 20
rect 6370 15 6450 20
rect 7310 15 7390 20
rect 790 -5 870 0
rect 1730 -5 1810 0
use sky130_fd_pr__nfet_01v8_ZWZ6GW  sky130_fd_pr__nfet_01v8_ZWZ6GW_0
timestamp 1619111721
transform 1 0 -867 0 1 592
box -759 -630 759 630
use sky130_fd_pr__pfet_01v8_lvt_CWLY9J  sky130_fd_pr__pfet_01v8_lvt_CWLY9J_0
array 0 7 930 0 4 1908
timestamp 1619111470
transform 1 0 412 0 1 901
box -465 -954 465 954
<< labels >>
rlabel metal1 -100 10400 7400 10500 1 vin_p
rlabel metal1 -100 10200 7400 10300 1 vin_n
rlabel metal1 -100 10000 7400 10100 1 iref
rlabel metal1 -100 9800 7400 9900 1 vout
rlabel metal1 -100 9600 7400 9700 1 vout_n
rlabel metal1 -1600 -400 7360 -140 1 vss
<< end >>
