magic
tech sky130A
magscale 1 2
timestamp 1615909117
<< error_p >>
rect -1445 -311 -1387 -305
rect -1327 -311 -1269 -305
rect -1209 -311 -1151 -305
rect -1091 -311 -1033 -305
rect -973 -311 -915 -305
rect -855 -311 -797 -305
rect -737 -311 -679 -305
rect -619 -311 -561 -305
rect -501 -311 -443 -305
rect -383 -311 -325 -305
rect -265 -311 -207 -305
rect -147 -311 -89 -305
rect -29 -311 29 -305
rect 89 -311 147 -305
rect 207 -311 265 -305
rect 325 -311 383 -305
rect 443 -311 501 -305
rect 561 -311 619 -305
rect 679 -311 737 -305
rect 797 -311 855 -305
rect 915 -311 973 -305
rect 1033 -311 1091 -305
rect 1151 -311 1209 -305
rect 1269 -311 1327 -305
rect 1387 -311 1445 -305
rect -1445 -345 -1433 -311
rect -1327 -345 -1315 -311
rect -1209 -345 -1197 -311
rect -1091 -345 -1079 -311
rect -973 -345 -961 -311
rect -855 -345 -843 -311
rect -737 -345 -725 -311
rect -619 -345 -607 -311
rect -501 -345 -489 -311
rect -383 -345 -371 -311
rect -265 -345 -253 -311
rect -147 -345 -135 -311
rect -29 -345 -17 -311
rect 89 -345 101 -311
rect 207 -345 219 -311
rect 325 -345 337 -311
rect 443 -345 455 -311
rect 561 -345 573 -311
rect 679 -345 691 -311
rect 797 -345 809 -311
rect 915 -345 927 -311
rect 1033 -345 1045 -311
rect 1151 -345 1163 -311
rect 1269 -345 1281 -311
rect 1387 -345 1399 -311
rect -1445 -351 -1387 -345
rect -1327 -351 -1269 -345
rect -1209 -351 -1151 -345
rect -1091 -351 -1033 -345
rect -973 -351 -915 -345
rect -855 -351 -797 -345
rect -737 -351 -679 -345
rect -619 -351 -561 -345
rect -501 -351 -443 -345
rect -383 -351 -325 -345
rect -265 -351 -207 -345
rect -147 -351 -89 -345
rect -29 -351 29 -345
rect 89 -351 147 -345
rect 207 -351 265 -345
rect 325 -351 383 -345
rect 443 -351 501 -345
rect 561 -351 619 -345
rect 679 -351 737 -345
rect 797 -351 855 -345
rect 915 -351 973 -345
rect 1033 -351 1091 -345
rect 1151 -351 1209 -345
rect 1269 -351 1327 -345
rect 1387 -351 1445 -345
<< nwell >>
rect -1642 -484 1642 484
<< pmos >>
rect -1446 -264 -1386 336
rect -1328 -264 -1268 336
rect -1210 -264 -1150 336
rect -1092 -264 -1032 336
rect -974 -264 -914 336
rect -856 -264 -796 336
rect -738 -264 -678 336
rect -620 -264 -560 336
rect -502 -264 -442 336
rect -384 -264 -324 336
rect -266 -264 -206 336
rect -148 -264 -88 336
rect -30 -264 30 336
rect 88 -264 148 336
rect 206 -264 266 336
rect 324 -264 384 336
rect 442 -264 502 336
rect 560 -264 620 336
rect 678 -264 738 336
rect 796 -264 856 336
rect 914 -264 974 336
rect 1032 -264 1092 336
rect 1150 -264 1210 336
rect 1268 -264 1328 336
rect 1386 -264 1446 336
<< pdiff >>
rect -1504 324 -1446 336
rect -1504 -252 -1492 324
rect -1458 -252 -1446 324
rect -1504 -264 -1446 -252
rect -1386 324 -1328 336
rect -1386 -252 -1374 324
rect -1340 -252 -1328 324
rect -1386 -264 -1328 -252
rect -1268 324 -1210 336
rect -1268 -252 -1256 324
rect -1222 -252 -1210 324
rect -1268 -264 -1210 -252
rect -1150 324 -1092 336
rect -1150 -252 -1138 324
rect -1104 -252 -1092 324
rect -1150 -264 -1092 -252
rect -1032 324 -974 336
rect -1032 -252 -1020 324
rect -986 -252 -974 324
rect -1032 -264 -974 -252
rect -914 324 -856 336
rect -914 -252 -902 324
rect -868 -252 -856 324
rect -914 -264 -856 -252
rect -796 324 -738 336
rect -796 -252 -784 324
rect -750 -252 -738 324
rect -796 -264 -738 -252
rect -678 324 -620 336
rect -678 -252 -666 324
rect -632 -252 -620 324
rect -678 -264 -620 -252
rect -560 324 -502 336
rect -560 -252 -548 324
rect -514 -252 -502 324
rect -560 -264 -502 -252
rect -442 324 -384 336
rect -442 -252 -430 324
rect -396 -252 -384 324
rect -442 -264 -384 -252
rect -324 324 -266 336
rect -324 -252 -312 324
rect -278 -252 -266 324
rect -324 -264 -266 -252
rect -206 324 -148 336
rect -206 -252 -194 324
rect -160 -252 -148 324
rect -206 -264 -148 -252
rect -88 324 -30 336
rect -88 -252 -76 324
rect -42 -252 -30 324
rect -88 -264 -30 -252
rect 30 324 88 336
rect 30 -252 42 324
rect 76 -252 88 324
rect 30 -264 88 -252
rect 148 324 206 336
rect 148 -252 160 324
rect 194 -252 206 324
rect 148 -264 206 -252
rect 266 324 324 336
rect 266 -252 278 324
rect 312 -252 324 324
rect 266 -264 324 -252
rect 384 324 442 336
rect 384 -252 396 324
rect 430 -252 442 324
rect 384 -264 442 -252
rect 502 324 560 336
rect 502 -252 514 324
rect 548 -252 560 324
rect 502 -264 560 -252
rect 620 324 678 336
rect 620 -252 632 324
rect 666 -252 678 324
rect 620 -264 678 -252
rect 738 324 796 336
rect 738 -252 750 324
rect 784 -252 796 324
rect 738 -264 796 -252
rect 856 324 914 336
rect 856 -252 868 324
rect 902 -252 914 324
rect 856 -264 914 -252
rect 974 324 1032 336
rect 974 -252 986 324
rect 1020 -252 1032 324
rect 974 -264 1032 -252
rect 1092 324 1150 336
rect 1092 -252 1104 324
rect 1138 -252 1150 324
rect 1092 -264 1150 -252
rect 1210 324 1268 336
rect 1210 -252 1222 324
rect 1256 -252 1268 324
rect 1210 -264 1268 -252
rect 1328 324 1386 336
rect 1328 -252 1340 324
rect 1374 -252 1386 324
rect 1328 -264 1386 -252
rect 1446 324 1504 336
rect 1446 -252 1458 324
rect 1492 -252 1504 324
rect 1446 -264 1504 -252
<< pdiffc >>
rect -1492 -252 -1458 324
rect -1374 -252 -1340 324
rect -1256 -252 -1222 324
rect -1138 -252 -1104 324
rect -1020 -252 -986 324
rect -902 -252 -868 324
rect -784 -252 -750 324
rect -666 -252 -632 324
rect -548 -252 -514 324
rect -430 -252 -396 324
rect -312 -252 -278 324
rect -194 -252 -160 324
rect -76 -252 -42 324
rect 42 -252 76 324
rect 160 -252 194 324
rect 278 -252 312 324
rect 396 -252 430 324
rect 514 -252 548 324
rect 632 -252 666 324
rect 750 -252 784 324
rect 868 -252 902 324
rect 986 -252 1020 324
rect 1104 -252 1138 324
rect 1222 -252 1256 324
rect 1340 -252 1374 324
rect 1458 -252 1492 324
<< nsubdiff >>
rect -1606 414 -1510 448
rect 1510 414 1606 448
rect -1606 351 -1572 414
rect 1572 351 1606 414
rect -1606 -414 -1572 -351
rect 1572 -414 1606 -351
rect -1606 -448 -1510 -414
rect 1510 -448 1606 -414
<< nsubdiffcont >>
rect -1510 414 1510 448
rect -1606 -351 -1572 351
rect 1572 -351 1606 351
rect -1510 -448 1510 -414
<< poly >>
rect -1446 336 -1386 362
rect -1328 336 -1268 362
rect -1210 336 -1150 362
rect -1092 336 -1032 362
rect -974 336 -914 362
rect -856 336 -796 362
rect -738 336 -678 362
rect -620 336 -560 362
rect -502 336 -442 362
rect -384 336 -324 362
rect -266 336 -206 362
rect -148 336 -88 362
rect -30 336 30 362
rect 88 336 148 362
rect 206 336 266 362
rect 324 336 384 362
rect 442 336 502 362
rect 560 336 620 362
rect 678 336 738 362
rect 796 336 856 362
rect 914 336 974 362
rect 1032 336 1092 362
rect 1150 336 1210 362
rect 1268 336 1328 362
rect 1386 336 1446 362
rect -1446 -295 -1386 -264
rect -1328 -295 -1268 -264
rect -1210 -295 -1150 -264
rect -1092 -295 -1032 -264
rect -974 -295 -914 -264
rect -856 -295 -796 -264
rect -738 -295 -678 -264
rect -620 -295 -560 -264
rect -502 -295 -442 -264
rect -384 -295 -324 -264
rect -266 -295 -206 -264
rect -148 -295 -88 -264
rect -30 -295 30 -264
rect 88 -295 148 -264
rect 206 -295 266 -264
rect 324 -295 384 -264
rect 442 -295 502 -264
rect 560 -295 620 -264
rect 678 -295 738 -264
rect 796 -295 856 -264
rect 914 -295 974 -264
rect 1032 -295 1092 -264
rect 1150 -295 1210 -264
rect 1268 -295 1328 -264
rect 1386 -295 1446 -264
rect -1449 -311 -1383 -295
rect -1449 -345 -1433 -311
rect -1399 -345 -1383 -311
rect -1449 -361 -1383 -345
rect -1331 -311 -1265 -295
rect -1331 -345 -1315 -311
rect -1281 -345 -1265 -311
rect -1331 -361 -1265 -345
rect -1213 -311 -1147 -295
rect -1213 -345 -1197 -311
rect -1163 -345 -1147 -311
rect -1213 -361 -1147 -345
rect -1095 -311 -1029 -295
rect -1095 -345 -1079 -311
rect -1045 -345 -1029 -311
rect -1095 -361 -1029 -345
rect -977 -311 -911 -295
rect -977 -345 -961 -311
rect -927 -345 -911 -311
rect -977 -361 -911 -345
rect -859 -311 -793 -295
rect -859 -345 -843 -311
rect -809 -345 -793 -311
rect -859 -361 -793 -345
rect -741 -311 -675 -295
rect -741 -345 -725 -311
rect -691 -345 -675 -311
rect -741 -361 -675 -345
rect -623 -311 -557 -295
rect -623 -345 -607 -311
rect -573 -345 -557 -311
rect -623 -361 -557 -345
rect -505 -311 -439 -295
rect -505 -345 -489 -311
rect -455 -345 -439 -311
rect -505 -361 -439 -345
rect -387 -311 -321 -295
rect -387 -345 -371 -311
rect -337 -345 -321 -311
rect -387 -361 -321 -345
rect -269 -311 -203 -295
rect -269 -345 -253 -311
rect -219 -345 -203 -311
rect -269 -361 -203 -345
rect -151 -311 -85 -295
rect -151 -345 -135 -311
rect -101 -345 -85 -311
rect -151 -361 -85 -345
rect -33 -311 33 -295
rect -33 -345 -17 -311
rect 17 -345 33 -311
rect -33 -361 33 -345
rect 85 -311 151 -295
rect 85 -345 101 -311
rect 135 -345 151 -311
rect 85 -361 151 -345
rect 203 -311 269 -295
rect 203 -345 219 -311
rect 253 -345 269 -311
rect 203 -361 269 -345
rect 321 -311 387 -295
rect 321 -345 337 -311
rect 371 -345 387 -311
rect 321 -361 387 -345
rect 439 -311 505 -295
rect 439 -345 455 -311
rect 489 -345 505 -311
rect 439 -361 505 -345
rect 557 -311 623 -295
rect 557 -345 573 -311
rect 607 -345 623 -311
rect 557 -361 623 -345
rect 675 -311 741 -295
rect 675 -345 691 -311
rect 725 -345 741 -311
rect 675 -361 741 -345
rect 793 -311 859 -295
rect 793 -345 809 -311
rect 843 -345 859 -311
rect 793 -361 859 -345
rect 911 -311 977 -295
rect 911 -345 927 -311
rect 961 -345 977 -311
rect 911 -361 977 -345
rect 1029 -311 1095 -295
rect 1029 -345 1045 -311
rect 1079 -345 1095 -311
rect 1029 -361 1095 -345
rect 1147 -311 1213 -295
rect 1147 -345 1163 -311
rect 1197 -345 1213 -311
rect 1147 -361 1213 -345
rect 1265 -311 1331 -295
rect 1265 -345 1281 -311
rect 1315 -345 1331 -311
rect 1265 -361 1331 -345
rect 1383 -311 1449 -295
rect 1383 -345 1399 -311
rect 1433 -345 1449 -311
rect 1383 -361 1449 -345
<< polycont >>
rect -1433 -345 -1399 -311
rect -1315 -345 -1281 -311
rect -1197 -345 -1163 -311
rect -1079 -345 -1045 -311
rect -961 -345 -927 -311
rect -843 -345 -809 -311
rect -725 -345 -691 -311
rect -607 -345 -573 -311
rect -489 -345 -455 -311
rect -371 -345 -337 -311
rect -253 -345 -219 -311
rect -135 -345 -101 -311
rect -17 -345 17 -311
rect 101 -345 135 -311
rect 219 -345 253 -311
rect 337 -345 371 -311
rect 455 -345 489 -311
rect 573 -345 607 -311
rect 691 -345 725 -311
rect 809 -345 843 -311
rect 927 -345 961 -311
rect 1045 -345 1079 -311
rect 1163 -345 1197 -311
rect 1281 -345 1315 -311
rect 1399 -345 1433 -311
<< locali >>
rect -1606 414 -1510 448
rect 1510 414 1606 448
rect -1606 351 -1572 414
rect 1572 351 1606 414
rect -1492 324 -1458 340
rect -1492 -268 -1458 -252
rect -1374 324 -1340 340
rect -1374 -268 -1340 -252
rect -1256 324 -1222 340
rect -1256 -268 -1222 -252
rect -1138 324 -1104 340
rect -1138 -268 -1104 -252
rect -1020 324 -986 340
rect -1020 -268 -986 -252
rect -902 324 -868 340
rect -902 -268 -868 -252
rect -784 324 -750 340
rect -784 -268 -750 -252
rect -666 324 -632 340
rect -666 -268 -632 -252
rect -548 324 -514 340
rect -548 -268 -514 -252
rect -430 324 -396 340
rect -430 -268 -396 -252
rect -312 324 -278 340
rect -312 -268 -278 -252
rect -194 324 -160 340
rect -194 -268 -160 -252
rect -76 324 -42 340
rect -76 -268 -42 -252
rect 42 324 76 340
rect 42 -268 76 -252
rect 160 324 194 340
rect 160 -268 194 -252
rect 278 324 312 340
rect 278 -268 312 -252
rect 396 324 430 340
rect 396 -268 430 -252
rect 514 324 548 340
rect 514 -268 548 -252
rect 632 324 666 340
rect 632 -268 666 -252
rect 750 324 784 340
rect 750 -268 784 -252
rect 868 324 902 340
rect 868 -268 902 -252
rect 986 324 1020 340
rect 986 -268 1020 -252
rect 1104 324 1138 340
rect 1104 -268 1138 -252
rect 1222 324 1256 340
rect 1222 -268 1256 -252
rect 1340 324 1374 340
rect 1340 -268 1374 -252
rect 1458 324 1492 340
rect 1458 -268 1492 -252
rect -1449 -345 -1433 -311
rect -1399 -345 -1383 -311
rect -1331 -345 -1315 -311
rect -1281 -345 -1265 -311
rect -1213 -345 -1197 -311
rect -1163 -345 -1147 -311
rect -1095 -345 -1079 -311
rect -1045 -345 -1029 -311
rect -977 -345 -961 -311
rect -927 -345 -911 -311
rect -859 -345 -843 -311
rect -809 -345 -793 -311
rect -741 -345 -725 -311
rect -691 -345 -675 -311
rect -623 -345 -607 -311
rect -573 -345 -557 -311
rect -505 -345 -489 -311
rect -455 -345 -439 -311
rect -387 -345 -371 -311
rect -337 -345 -321 -311
rect -269 -345 -253 -311
rect -219 -345 -203 -311
rect -151 -345 -135 -311
rect -101 -345 -85 -311
rect -33 -345 -17 -311
rect 17 -345 33 -311
rect 85 -345 101 -311
rect 135 -345 151 -311
rect 203 -345 219 -311
rect 253 -345 269 -311
rect 321 -345 337 -311
rect 371 -345 387 -311
rect 439 -345 455 -311
rect 489 -345 505 -311
rect 557 -345 573 -311
rect 607 -345 623 -311
rect 675 -345 691 -311
rect 725 -345 741 -311
rect 793 -345 809 -311
rect 843 -345 859 -311
rect 911 -345 927 -311
rect 961 -345 977 -311
rect 1029 -345 1045 -311
rect 1079 -345 1095 -311
rect 1147 -345 1163 -311
rect 1197 -345 1213 -311
rect 1265 -345 1281 -311
rect 1315 -345 1331 -311
rect 1383 -345 1399 -311
rect 1433 -345 1449 -311
rect -1606 -414 -1572 -351
rect 1572 -414 1606 -351
rect -1606 -448 -1510 -414
rect 1510 -448 1606 -414
<< viali >>
rect -1492 -252 -1458 324
rect -1374 -252 -1340 324
rect -1256 -252 -1222 324
rect -1138 -252 -1104 324
rect -1020 -252 -986 324
rect -902 -252 -868 324
rect -784 -252 -750 324
rect -666 -252 -632 324
rect -548 -252 -514 324
rect -430 -252 -396 324
rect -312 -252 -278 324
rect -194 -252 -160 324
rect -76 -252 -42 324
rect 42 -252 76 324
rect 160 -252 194 324
rect 278 -252 312 324
rect 396 -252 430 324
rect 514 -252 548 324
rect 632 -252 666 324
rect 750 -252 784 324
rect 868 -252 902 324
rect 986 -252 1020 324
rect 1104 -252 1138 324
rect 1222 -252 1256 324
rect 1340 -252 1374 324
rect 1458 -252 1492 324
rect -1433 -345 -1399 -311
rect -1315 -345 -1281 -311
rect -1197 -345 -1163 -311
rect -1079 -345 -1045 -311
rect -961 -345 -927 -311
rect -843 -345 -809 -311
rect -725 -345 -691 -311
rect -607 -345 -573 -311
rect -489 -345 -455 -311
rect -371 -345 -337 -311
rect -253 -345 -219 -311
rect -135 -345 -101 -311
rect -17 -345 17 -311
rect 101 -345 135 -311
rect 219 -345 253 -311
rect 337 -345 371 -311
rect 455 -345 489 -311
rect 573 -345 607 -311
rect 691 -345 725 -311
rect 809 -345 843 -311
rect 927 -345 961 -311
rect 1045 -345 1079 -311
rect 1163 -345 1197 -311
rect 1281 -345 1315 -311
rect 1399 -345 1433 -311
<< metal1 >>
rect -1498 324 -1452 336
rect -1498 -252 -1492 324
rect -1458 -252 -1452 324
rect -1498 -264 -1452 -252
rect -1380 324 -1334 336
rect -1380 -252 -1374 324
rect -1340 -252 -1334 324
rect -1380 -264 -1334 -252
rect -1262 324 -1216 336
rect -1262 -252 -1256 324
rect -1222 -252 -1216 324
rect -1262 -264 -1216 -252
rect -1144 324 -1098 336
rect -1144 -252 -1138 324
rect -1104 -252 -1098 324
rect -1144 -264 -1098 -252
rect -1026 324 -980 336
rect -1026 -252 -1020 324
rect -986 -252 -980 324
rect -1026 -264 -980 -252
rect -908 324 -862 336
rect -908 -252 -902 324
rect -868 -252 -862 324
rect -908 -264 -862 -252
rect -790 324 -744 336
rect -790 -252 -784 324
rect -750 -252 -744 324
rect -790 -264 -744 -252
rect -672 324 -626 336
rect -672 -252 -666 324
rect -632 -252 -626 324
rect -672 -264 -626 -252
rect -554 324 -508 336
rect -554 -252 -548 324
rect -514 -252 -508 324
rect -554 -264 -508 -252
rect -436 324 -390 336
rect -436 -252 -430 324
rect -396 -252 -390 324
rect -436 -264 -390 -252
rect -318 324 -272 336
rect -318 -252 -312 324
rect -278 -252 -272 324
rect -318 -264 -272 -252
rect -200 324 -154 336
rect -200 -252 -194 324
rect -160 -252 -154 324
rect -200 -264 -154 -252
rect -82 324 -36 336
rect -82 -252 -76 324
rect -42 -252 -36 324
rect -82 -264 -36 -252
rect 36 324 82 336
rect 36 -252 42 324
rect 76 -252 82 324
rect 36 -264 82 -252
rect 154 324 200 336
rect 154 -252 160 324
rect 194 -252 200 324
rect 154 -264 200 -252
rect 272 324 318 336
rect 272 -252 278 324
rect 312 -252 318 324
rect 272 -264 318 -252
rect 390 324 436 336
rect 390 -252 396 324
rect 430 -252 436 324
rect 390 -264 436 -252
rect 508 324 554 336
rect 508 -252 514 324
rect 548 -252 554 324
rect 508 -264 554 -252
rect 626 324 672 336
rect 626 -252 632 324
rect 666 -252 672 324
rect 626 -264 672 -252
rect 744 324 790 336
rect 744 -252 750 324
rect 784 -252 790 324
rect 744 -264 790 -252
rect 862 324 908 336
rect 862 -252 868 324
rect 902 -252 908 324
rect 862 -264 908 -252
rect 980 324 1026 336
rect 980 -252 986 324
rect 1020 -252 1026 324
rect 980 -264 1026 -252
rect 1098 324 1144 336
rect 1098 -252 1104 324
rect 1138 -252 1144 324
rect 1098 -264 1144 -252
rect 1216 324 1262 336
rect 1216 -252 1222 324
rect 1256 -252 1262 324
rect 1216 -264 1262 -252
rect 1334 324 1380 336
rect 1334 -252 1340 324
rect 1374 -252 1380 324
rect 1334 -264 1380 -252
rect 1452 324 1498 336
rect 1452 -252 1458 324
rect 1492 -252 1498 324
rect 1452 -264 1498 -252
rect -1445 -311 -1387 -305
rect -1445 -345 -1433 -311
rect -1399 -345 -1387 -311
rect -1445 -351 -1387 -345
rect -1327 -311 -1269 -305
rect -1327 -345 -1315 -311
rect -1281 -345 -1269 -311
rect -1327 -351 -1269 -345
rect -1209 -311 -1151 -305
rect -1209 -345 -1197 -311
rect -1163 -345 -1151 -311
rect -1209 -351 -1151 -345
rect -1091 -311 -1033 -305
rect -1091 -345 -1079 -311
rect -1045 -345 -1033 -311
rect -1091 -351 -1033 -345
rect -973 -311 -915 -305
rect -973 -345 -961 -311
rect -927 -345 -915 -311
rect -973 -351 -915 -345
rect -855 -311 -797 -305
rect -855 -345 -843 -311
rect -809 -345 -797 -311
rect -855 -351 -797 -345
rect -737 -311 -679 -305
rect -737 -345 -725 -311
rect -691 -345 -679 -311
rect -737 -351 -679 -345
rect -619 -311 -561 -305
rect -619 -345 -607 -311
rect -573 -345 -561 -311
rect -619 -351 -561 -345
rect -501 -311 -443 -305
rect -501 -345 -489 -311
rect -455 -345 -443 -311
rect -501 -351 -443 -345
rect -383 -311 -325 -305
rect -383 -345 -371 -311
rect -337 -345 -325 -311
rect -383 -351 -325 -345
rect -265 -311 -207 -305
rect -265 -345 -253 -311
rect -219 -345 -207 -311
rect -265 -351 -207 -345
rect -147 -311 -89 -305
rect -147 -345 -135 -311
rect -101 -345 -89 -311
rect -147 -351 -89 -345
rect -29 -311 29 -305
rect -29 -345 -17 -311
rect 17 -345 29 -311
rect -29 -351 29 -345
rect 89 -311 147 -305
rect 89 -345 101 -311
rect 135 -345 147 -311
rect 89 -351 147 -345
rect 207 -311 265 -305
rect 207 -345 219 -311
rect 253 -345 265 -311
rect 207 -351 265 -345
rect 325 -311 383 -305
rect 325 -345 337 -311
rect 371 -345 383 -311
rect 325 -351 383 -345
rect 443 -311 501 -305
rect 443 -345 455 -311
rect 489 -345 501 -311
rect 443 -351 501 -345
rect 561 -311 619 -305
rect 561 -345 573 -311
rect 607 -345 619 -311
rect 561 -351 619 -345
rect 679 -311 737 -305
rect 679 -345 691 -311
rect 725 -345 737 -311
rect 679 -351 737 -345
rect 797 -311 855 -305
rect 797 -345 809 -311
rect 843 -345 855 -311
rect 797 -351 855 -345
rect 915 -311 973 -305
rect 915 -345 927 -311
rect 961 -345 973 -311
rect 915 -351 973 -345
rect 1033 -311 1091 -305
rect 1033 -345 1045 -311
rect 1079 -345 1091 -311
rect 1033 -351 1091 -345
rect 1151 -311 1209 -305
rect 1151 -345 1163 -311
rect 1197 -345 1209 -311
rect 1151 -351 1209 -345
rect 1269 -311 1327 -305
rect 1269 -345 1281 -311
rect 1315 -345 1327 -311
rect 1269 -351 1327 -345
rect 1387 -311 1445 -305
rect 1387 -345 1399 -311
rect 1433 -345 1445 -311
rect 1387 -351 1445 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1589 -431 1589 431
string parameters w 3 l 0.3 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
