magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_p >>
rect -29 261 29 267
rect -29 227 -17 261
rect -29 221 29 227
rect -29 -227 29 -221
rect -29 -261 -17 -227
rect -29 -267 29 -261
<< nwell >>
rect -211 -399 211 399
<< pmos >>
rect -15 -180 15 180
<< pdiff >>
rect -73 168 -15 180
rect -73 -168 -61 168
rect -27 -168 -15 168
rect -73 -180 -15 -168
rect 15 168 73 180
rect 15 -168 27 168
rect 61 -168 73 168
rect 15 -180 73 -168
<< pdiffc >>
rect -61 -168 -27 168
rect 27 -168 61 168
<< nsubdiff >>
rect -175 329 -79 363
rect 79 329 175 363
rect -175 267 -141 329
rect 141 267 175 329
rect -175 -329 -141 -267
rect 141 -329 175 -267
rect -175 -363 -79 -329
rect 79 -363 175 -329
<< nsubdiffcont >>
rect -79 329 79 363
rect -175 -267 -141 267
rect 141 -267 175 267
rect -79 -363 79 -329
<< poly >>
rect -33 261 33 277
rect -33 227 -17 261
rect 17 227 33 261
rect -33 211 33 227
rect -15 180 15 211
rect -15 -211 15 -180
rect -33 -227 33 -211
rect -33 -261 -17 -227
rect 17 -261 33 -227
rect -33 -277 33 -261
<< polycont >>
rect -17 227 17 261
rect -17 -261 17 -227
<< locali >>
rect -175 329 -79 363
rect 79 329 175 363
rect -175 267 -141 329
rect 141 267 175 329
rect -33 227 -17 261
rect 17 227 33 261
rect -61 168 -27 184
rect -61 -184 -27 -168
rect 27 168 61 184
rect 27 -184 61 -168
rect -33 -261 -17 -227
rect 17 -261 33 -227
rect -175 -329 -141 -267
rect 141 -329 175 -267
rect -175 -363 -79 -329
rect 79 -363 175 -329
<< viali >>
rect -17 227 17 261
rect -61 -168 -27 168
rect 27 -168 61 168
rect -17 -261 17 -227
<< metal1 >>
rect -29 261 29 267
rect -29 227 -17 261
rect 17 227 29 261
rect -29 221 29 227
rect -67 168 -21 180
rect -67 -168 -61 168
rect -27 -168 -21 168
rect -67 -180 -21 -168
rect 21 168 67 180
rect 21 -168 27 168
rect 61 -168 67 168
rect 21 -180 67 -168
rect -29 -227 29 -221
rect -29 -261 -17 -227
rect 17 -261 29 -227
rect -29 -267 29 -261
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -346 158 346
string parameters w 1.8 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
