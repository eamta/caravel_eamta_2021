magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 352 1057 387 1075
rect 316 1042 387 1057
rect 667 1042 702 1076
rect 129 919 187 925
rect 129 908 141 919
rect 129 906 175 908
rect 316 906 386 1042
rect 668 1023 702 1042
rect 687 980 702 1023
rect 498 974 556 980
rect 498 940 510 974
rect 498 934 556 940
rect -53 870 386 906
rect 466 870 500 904
rect 554 870 588 904
rect 668 870 702 980
rect 721 989 756 1023
rect 721 870 755 989
rect 2512 957 2547 991
rect 867 921 925 927
rect 867 908 879 921
rect 867 906 913 908
rect 867 904 925 906
rect 863 887 929 904
rect 1037 898 1071 927
rect 1423 898 1634 953
rect 2513 938 2547 957
rect 867 881 925 887
rect 839 870 953 878
rect 1037 870 1380 898
rect -53 836 1380 870
rect -53 564 386 836
rect 454 818 469 833
rect 585 818 600 833
rect 454 788 512 818
rect 542 788 600 818
rect 454 772 480 788
rect 585 773 600 788
rect 454 728 488 772
rect 388 598 420 722
rect 454 713 495 728
rect 512 713 600 744
rect 452 682 480 713
rect 512 682 522 713
rect 554 709 588 713
rect 576 690 610 694
rect 494 616 522 682
rect 564 685 616 690
rect 564 675 610 685
rect 538 632 560 666
rect 542 626 556 632
rect 564 601 594 675
rect 570 598 594 601
rect 388 564 422 598
rect 576 594 582 598
rect 668 564 702 836
rect -53 547 434 564
rect 439 553 491 564
rect 448 550 480 553
rect 318 534 334 547
rect 352 538 434 547
rect 450 541 480 550
rect 352 530 387 538
rect 439 530 491 541
rect 564 530 702 564
rect 687 506 698 530
rect 721 511 755 836
rect 835 731 869 828
rect 923 798 957 828
rect 908 738 923 772
rect 954 754 969 769
rect 823 694 869 731
rect 823 690 874 694
rect 835 672 874 690
rect 840 660 874 672
rect 881 660 885 689
rect 926 688 969 754
rect 976 704 991 738
rect 950 675 969 688
rect 935 660 969 675
rect 840 647 886 660
rect 950 647 971 660
rect 840 634 971 647
rect 840 629 874 634
rect 880 629 971 634
rect 840 626 971 629
rect 840 619 886 626
rect 840 598 925 619
rect 840 579 912 598
rect 840 548 886 579
rect 950 563 971 626
rect 1037 573 1380 836
rect 840 522 874 548
rect 721 510 886 511
rect 721 482 740 510
rect 798 488 828 510
rect 939 500 991 511
rect 950 488 980 500
rect 787 482 839 488
rect 721 477 839 482
rect 939 477 991 488
rect 1051 477 1380 573
rect 1054 388 1380 477
rect 1423 883 1494 898
rect 2343 889 2401 895
rect 1423 424 1493 883
rect 2343 855 2355 889
rect 2343 849 2401 855
rect 1605 815 1663 821
rect 1605 781 1617 815
rect 1775 792 1809 810
rect 2197 792 2231 810
rect 1605 775 1663 781
rect 1775 756 1845 792
rect 1792 722 1863 756
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1423 388 1476 424
rect 1423 354 1634 388
rect 1792 371 1862 722
rect 1974 654 2032 660
rect 1974 620 1986 654
rect 1974 614 2032 620
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1423 335 1600 354
rect 1792 335 1845 371
rect 2161 318 2231 792
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2161 282 2214 318
rect 2532 265 2547 938
rect 2566 904 2601 938
rect 2566 265 2600 904
rect 2712 836 2770 842
rect 2712 802 2724 836
rect 2712 796 2770 802
rect 2882 633 2916 651
rect 4726 639 4761 673
rect 2882 597 2952 633
rect 4727 620 4761 639
rect 2899 563 2970 597
rect 3250 563 3285 597
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2566 231 2581 265
rect -28 204 228 228
rect 2899 212 2969 563
rect 3251 544 3285 563
rect 3081 495 3139 501
rect 3081 461 3093 495
rect 3081 455 3139 461
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 0 176 200 200
rect 2899 176 2952 212
rect 176 54 200 176
rect 204 82 228 172
rect 3270 159 3285 544
rect 3304 510 3339 544
rect 3619 510 3654 544
rect 4042 527 4077 545
rect 3304 159 3338 510
rect 3620 491 3654 510
rect 4006 512 4077 527
rect 3450 442 3508 448
rect 3450 408 3462 442
rect 3450 402 3508 408
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 491
rect 3673 457 3708 491
rect 3673 106 3707 457
rect 3819 389 3877 395
rect 3819 355 3831 389
rect 3819 349 3877 355
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 182 16 200 54
rect 210 16 228 82
rect 3673 72 3688 106
rect 4006 53 4076 512
rect 4188 444 4246 450
rect 4188 410 4200 444
rect 4188 404 4246 410
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4006 17 4059 53
rect 4377 0 4392 546
rect 4411 0 4445 600
rect 4557 571 4615 577
rect 4557 537 4569 571
rect 4557 531 4615 537
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 620
rect 4780 586 4815 620
rect 4780 -53 4814 586
rect 4926 518 4984 524
rect 4926 484 4938 518
rect 4926 478 4984 484
rect 5096 315 5130 333
rect 5096 279 5166 315
rect 5113 245 5184 279
rect 5464 245 5499 279
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5113 -106 5183 245
rect 5465 226 5499 245
rect 5295 177 5353 183
rect 5295 143 5307 177
rect 5295 137 5353 143
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5113 -142 5166 -106
rect 5484 -159 5499 226
rect 5518 192 5553 226
rect 5833 192 5868 226
rect 6256 209 6291 227
rect 5518 -159 5552 192
rect 5834 173 5868 192
rect 6220 194 6291 209
rect 5664 124 5722 130
rect 5664 90 5676 124
rect 5664 84 5722 90
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5518 -193 5533 -159
rect 5853 -212 5868 173
rect 5887 139 5922 173
rect 5887 -212 5921 139
rect 6033 71 6091 77
rect 6033 37 6045 71
rect 6033 31 6091 37
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5887 -246 5902 -212
rect 6220 -265 6290 194
rect 6402 126 6460 132
rect 6402 92 6414 126
rect 6572 103 6606 121
rect 6994 103 7029 121
rect 6402 86 6460 92
rect 6572 67 6642 103
rect 6958 88 7029 103
rect 6589 33 6660 67
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6220 -301 6273 -265
rect 6589 -318 6659 33
rect 6771 -35 6829 -29
rect 6771 -69 6783 -35
rect 6771 -75 6829 -69
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6589 -354 6642 -318
rect 6958 -371 7028 88
rect 7140 20 7198 26
rect 7140 -14 7152 20
rect 7310 -3 7344 15
rect 7732 -3 7767 15
rect 7140 -20 7198 -14
rect 7310 -39 7380 -3
rect 7696 -18 7767 -3
rect 7327 -73 7398 -39
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6958 -407 7011 -371
rect 7327 -424 7397 -73
rect 7509 -141 7567 -135
rect 7509 -175 7521 -141
rect 7509 -181 7567 -175
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7327 -460 7380 -424
rect 7696 -477 7766 -18
rect 7878 -86 7936 -80
rect 7878 -120 7890 -86
rect 7878 -126 7936 -120
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7696 -513 7749 -477
<< nwell >>
rect -676 816 1380 906
rect -676 486 1328 816
rect 1344 486 1380 816
rect -676 366 1380 486
rect -168 354 1380 366
rect -168 328 1346 354
rect -168 262 140 328
rect 150 314 1346 328
rect 150 262 338 314
rect -168 242 338 262
rect -142 228 66 242
<< psubdiff >>
rect -632 -66 -608 -32
rect 1266 -66 1290 -32
<< nsubdiff >>
rect -612 836 -492 870
rect 1062 836 1264 870
<< psubdiffcont >>
rect -608 -66 1266 -32
<< nsubdiffcont >>
rect -492 836 1062 870
<< poly >>
rect -450 788 740 818
rect -554 556 -524 584
rect -574 526 -524 556
rect -574 376 -544 526
rect -450 484 -420 788
rect -486 468 -420 484
rect -486 434 -470 468
rect -436 434 -420 468
rect -486 418 -420 434
rect -346 420 -316 788
rect -258 716 164 746
rect -258 690 -228 716
rect -258 464 -164 494
rect -346 390 -236 420
rect -574 346 -460 376
rect -676 288 -532 304
rect -676 274 -582 288
rect -598 254 -582 274
rect -548 254 -532 288
rect -598 238 -532 254
rect -594 10 -564 116
rect -490 10 -460 346
rect -266 220 -236 390
rect -298 190 -236 220
rect -386 10 -356 112
rect -194 10 -164 464
rect -686 -20 -164 10
rect -58 10 -28 670
rect 30 220 60 648
rect 134 400 164 716
rect 346 508 376 558
rect 206 492 376 508
rect 206 458 222 492
rect 256 478 376 492
rect 256 458 272 478
rect 206 442 272 458
rect 134 370 302 400
rect 150 312 216 328
rect 150 278 166 312
rect 200 278 216 312
rect 150 262 216 278
rect 272 292 302 370
rect 346 364 376 478
rect 450 436 480 788
rect 622 526 652 690
rect 622 462 652 506
rect 710 482 740 788
rect 926 738 992 754
rect 926 704 942 738
rect 976 704 992 738
rect 450 406 578 436
rect 622 420 670 462
rect 798 438 828 690
rect 926 688 992 704
rect 346 334 494 364
rect 272 262 390 292
rect 150 220 180 262
rect 30 190 286 220
rect 360 82 390 262
rect 464 124 494 334
rect 548 288 578 406
rect 548 258 582 288
rect 552 124 582 258
rect 640 240 670 420
rect 728 408 828 438
rect 728 322 758 408
rect 950 378 980 688
rect 950 344 1164 378
rect 800 322 866 336
rect 728 320 866 322
rect 728 292 816 320
rect 728 218 758 292
rect 800 286 816 292
rect 850 286 866 320
rect 800 270 866 286
rect 640 82 670 160
rect 950 82 980 344
rect 1222 302 1252 406
rect 1038 270 1252 302
rect 360 52 670 82
rect 1038 10 1068 270
rect 1158 210 1224 226
rect 1158 176 1174 210
rect 1208 176 1224 210
rect 1158 160 1224 176
rect 1194 90 1224 160
rect 1194 60 1378 90
rect -58 -20 1336 10
<< polycont >>
rect -470 434 -436 468
rect -582 254 -548 288
rect 222 458 256 492
rect 166 278 200 312
rect 942 704 976 738
rect 816 286 850 320
rect 1174 176 1208 210
<< locali >>
rect 926 704 942 738
rect 976 704 992 738
rect -486 434 -470 468
rect -436 434 -420 468
rect 206 458 222 492
rect 256 458 272 492
rect -598 254 -582 288
rect -548 254 -532 288
rect 150 278 166 312
rect 200 278 216 312
rect 800 286 816 320
rect 850 286 866 320
rect 1158 176 1174 210
rect 1208 176 1224 210
rect -624 -66 -608 -32
rect 1266 -66 1282 -32
<< viali >>
rect -638 836 -492 870
rect -492 836 1062 870
rect 1062 836 1286 870
rect 942 704 976 738
rect -470 434 -436 468
rect 222 458 256 492
rect -582 254 -548 288
rect 166 278 200 312
rect 816 286 850 320
rect 1174 176 1208 210
rect -608 -66 1266 -32
<< metal1 >>
rect -676 870 1388 878
rect -676 836 -638 870
rect 1286 836 1388 870
rect -676 782 1388 836
rect -512 742 -478 782
rect -598 626 -566 732
rect -600 484 -566 626
rect -510 586 -476 742
rect -304 718 240 754
rect -600 468 -420 484
rect -600 448 -470 468
rect -600 366 -566 448
rect -486 434 -470 448
rect -436 434 -420 468
rect -486 418 -420 434
rect -654 332 -566 366
rect -654 210 -626 332
rect -598 292 -532 304
rect -392 292 -358 598
rect -304 482 -270 718
rect -216 604 -70 638
rect -304 448 -138 482
rect -598 288 -358 292
rect -598 254 -582 288
rect -548 258 -358 288
rect -548 254 -532 258
rect -598 238 -532 254
rect -654 174 -606 210
rect -640 58 -606 174
rect -432 156 -398 258
rect -172 230 -138 448
rect -344 202 -138 230
rect -104 234 -70 604
rect 206 508 240 718
rect 206 492 272 508
rect 206 458 222 492
rect 256 458 272 492
rect 206 442 272 458
rect 300 390 334 782
rect 664 738 992 754
rect 664 720 942 738
rect 388 644 610 678
rect 100 356 334 390
rect 150 312 216 328
rect 150 278 166 312
rect 200 302 216 312
rect 388 302 422 640
rect 664 482 698 720
rect 926 704 942 720
rect 976 704 992 738
rect 926 688 992 704
rect 1020 660 1054 782
rect 868 626 1054 660
rect 594 448 698 482
rect 200 278 540 302
rect 150 268 540 278
rect 150 262 216 268
rect -104 204 332 234
rect -344 156 -310 202
rect -104 130 -70 204
rect -552 16 -518 122
rect -256 96 -70 130
rect 0 124 200 200
rect -104 56 -70 96
rect -16 16 200 124
rect 210 16 244 124
rect 298 96 332 204
rect 418 16 452 210
rect 506 162 540 268
rect 594 164 628 448
rect 752 420 786 580
rect 682 386 786 420
rect 904 402 1120 436
rect 1264 406 1298 782
rect 682 162 716 386
rect 800 320 866 336
rect 904 320 940 402
rect 800 286 816 320
rect 850 286 940 320
rect 800 270 866 286
rect 904 230 940 286
rect 770 16 804 228
rect 904 210 1224 230
rect 904 196 1174 210
rect 904 88 940 196
rect 992 16 1026 156
rect 1080 90 1114 196
rect 1158 176 1174 196
rect 1208 176 1224 210
rect 1158 160 1224 176
rect -676 10 1378 16
rect -686 -20 1378 10
rect -676 -32 1378 -20
rect -676 -66 -608 -32
rect 1266 -66 1378 -32
rect -676 -72 1378 -66
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_0
timestamp 1615150785
transform 1 0 -283 0 1 129
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_4
timestamp 1615150785
transform 1 0 -579 0 1 89
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_3
timestamp 1615150785
transform 1 0 -371 0 1 129
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_0
timestamp 1615302329
transform 1 0 45 0 1 466
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_3
timestamp 1615302329
transform 1 0 -43 0 1 466
box -109 -242 109 242
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_6
timestamp 1615150785
transform 1 0 567 0 1 195
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_7
timestamp 1615150785
transform 1 0 655 0 1 195
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_5
timestamp 1615150785
transform 1 0 479 0 1 195
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_2
timestamp 1615150785
transform 1 0 271 0 1 127
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_1
timestamp 1615150785
transform 1 0 -43 0 1 89
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_10
timestamp 1615150785
transform 1 0 1053 0 1 123
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_9
timestamp 1615150785
transform 1 0 965 0 1 123
box -73 -71 73 71
use sky130_fd_pr__nfet_01v8_J836M4  sky130_fd_pr__nfet_01v8_J836M4_8
timestamp 1615150785
transform 1 0 743 0 1 195
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_XYCVAL  XM6
timestamp 1624053917
transform 1 0 2372 0 1 628
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM8
timestamp 1624053917
transform 1 0 3110 0 1 378
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM7
timestamp 1624053917
transform 1 0 2741 0 1 575
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XSLFBL  XM11
timestamp 1624053917
transform 1 0 4217 0 1 273
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM10
timestamp 1624053917
transform 1 0 3848 0 1 272
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM9
timestamp 1624053917
transform 1 0 3479 0 1 325
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XYCVAL  XM13
timestamp 1624053917
transform 1 0 4955 0 1 257
box -211 -399 211 399
use sky130_fd_pr__pfet_01v8_XYCVAL  XM12
timestamp 1624053917
transform 1 0 4586 0 1 310
box -211 -399 211 399
use sky130_fd_pr__nfet_01v8_HVW3BE  XM14
timestamp 1624053917
transform 1 0 5324 0 1 60
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_2
timestamp 1615568138
transform 1 0 -243 0 1 600
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_0
timestamp 1615568138
transform 1 0 -539 0 1 662
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_1
timestamp 1615568138
transform 1 0 -331 0 1 600
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_4
timestamp 1615568138
transform 1 0 637 0 1 600
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_5
timestamp 1615568138
transform 1 0 725 0 1 600
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_3
timestamp 1615568138
transform 1 0 361 0 1 628
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_XSLFBL  XM2
timestamp 1624053917
transform 1 0 527 0 1 803
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM3
timestamp 1624053917
transform 1 0 158 0 1 802
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_2
timestamp 1615302329
transform 1 0 1237 0 1 574
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5CNMEE  sky130_fd_pr__pfet_01v8_5CNMEE_1
timestamp 1615302329
transform 1 0 1149 0 1 574
box -109 -242 109 242
use sky130_fd_pr__pfet_01v8_5UWV5B  sky130_fd_pr__pfet_01v8_5UWV5B_6
timestamp 1615568138
transform 1 0 813 0 1 600
box -109 -152 109 152
use sky130_fd_pr__pfet_01v8_XSLFBL  XM5
timestamp 1624053917
transform 1 0 1634 0 1 644
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM0
timestamp 1624053917
transform 1 0 1265 0 1 643
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM1
timestamp 1624053917
transform 1 0 896 0 1 750
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1624053917
transform 1 0 2003 0 1 537
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM21
timestamp 1624053917
transform 1 0 7907 0 1 -257
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM20
timestamp 1624053917
transform 1 0 7538 0 1 -258
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM19
timestamp 1624053917
transform 1 0 7169 0 1 -151
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM18
timestamp 1624053917
transform 1 0 6800 0 1 -152
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_XSLFBL  XM17
timestamp 1624053917
transform 1 0 6431 0 1 -45
box -211 -309 211 309
use sky130_fd_pr__nfet_01v8_HVW3BE  XM16
timestamp 1624053917
transform 1 0 6062 0 1 -46
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM15
timestamp 1624053917
transform 1 0 5693 0 1 7
box -211 -255 211 255
<< labels >>
rlabel poly -676 274 -582 304 1 D
rlabel poly -58 -20 1336 10 1 clr
rlabel poly -686 -20 -164 10 1 clk
rlabel metal1 1174 176 1208 210 1 Q
rlabel metal1 -608 -66 1266 -32 1 vss
rlabel nwell -492 836 1062 870 1 vdd
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 D
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 clr
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 clk
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 vss
port 6 nsew
<< end >>
