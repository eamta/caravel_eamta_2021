magic
tech sky130A
magscale 1 2
timestamp 1616013451
<< error_p >>
rect -29 135 29 141
rect -29 101 -17 135
rect -29 95 29 101
<< nwell >>
rect -109 -188 109 154
<< pmos >>
rect -15 -126 15 54
<< pdiff >>
rect -73 42 -15 54
rect -73 -114 -61 42
rect -27 -114 -15 42
rect -73 -126 -15 -114
rect 15 42 73 54
rect 15 -114 27 42
rect 61 -114 73 42
rect 15 -126 73 -114
<< pdiffc >>
rect -61 -114 -27 42
rect 27 -114 61 42
<< poly >>
rect -33 135 33 151
rect -33 101 -17 135
rect 17 101 33 135
rect -33 85 33 101
rect -15 54 15 85
rect -15 -152 15 -126
<< polycont >>
rect -17 101 17 135
<< locali >>
rect -33 101 -17 135
rect 17 101 33 135
rect -61 42 -27 58
rect -61 -130 -27 -114
rect 27 42 61 58
rect 27 -130 61 -114
<< viali >>
rect -17 101 17 135
rect -61 -114 -27 42
rect 27 -114 61 42
<< metal1 >>
rect -29 135 29 141
rect -29 101 -17 135
rect 17 101 29 135
rect -29 95 29 101
rect -67 42 -21 54
rect -67 -114 -61 42
rect -27 -114 -21 42
rect -67 -126 -21 -114
rect 21 42 67 54
rect 21 -114 27 42
rect 61 -114 67 42
rect 21 -126 67 -114
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.9 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
