magic
tech sky130A
magscale 1 2
timestamp 1615600491
<< error_s >>
rect 1468 2608 1871 2609
rect 1449 2452 1871 2608
rect 1617 2441 1890 2452
rect 2569 2451 2801 2452
rect 1617 2440 1636 2441
rect 1703 2373 1890 2441
rect 1310 1963 1409 2131
rect 1478 1963 1516 2183
rect 1629 1963 1663 2183
rect 1478 1929 1883 1963
rect 2234 1858 2274 2090
rect 2519 1922 2523 1923
rect 2547 1922 2551 1923
rect 2249 1841 2488 1858
rect 2274 1836 2488 1841
<< nwell >>
rect 1409 2451 2287 2452
rect 2290 2451 2547 2452
rect 2569 2451 2869 2452
rect 1409 2450 2869 2451
rect 1409 2444 2482 2450
rect 1409 2441 2485 2444
rect 1409 2440 1636 2441
rect 1703 2440 2485 2441
rect 2489 2440 2869 2450
rect 1409 2374 1617 2440
rect 1409 2373 1636 2374
rect 1703 2373 2869 2440
rect 1409 2152 2869 2373
rect 1409 2056 1467 2152
rect 1468 2056 2869 2152
rect 1409 1963 2869 2056
rect 1409 1929 1478 1963
rect 1516 1929 1629 1963
rect 1663 1929 2712 1963
rect 2773 1929 2869 1963
rect 1409 1858 2869 1929
rect 1409 1836 2234 1858
rect 2274 1836 2869 1858
rect 1409 1440 2869 1836
<< pwell >>
rect 1403 2692 2869 2781
rect 1403 2660 1645 2692
rect 1651 2660 2869 2692
rect 1403 2608 2869 2660
rect 1403 2602 1645 2608
rect 1651 2602 2869 2608
rect 1403 2527 2869 2602
rect 1403 2525 2427 2527
rect 2458 2525 2869 2527
rect 1403 2452 2869 2525
rect 1409 1118 1733 1440
rect 1874 1242 1946 1321
rect 2479 1240 2532 1321
rect 2548 1118 2869 1440
<< poly >>
rect 1651 2661 1851 2691
rect 1651 2652 1711 2661
rect 1651 2618 1667 2652
rect 1701 2618 1711 2652
rect 1651 2602 1711 2618
rect 1437 1409 1467 2459
rect 1468 2406 1483 2436
rect 1541 2245 1853 2279
rect 1666 2068 1732 2084
rect 1666 2034 1682 2068
rect 1716 2034 1732 2068
rect 1666 2018 1732 2034
rect 1509 1866 1539 1867
rect 1672 1866 1702 2018
rect 1509 1836 1702 1866
rect 1509 1501 1539 1836
rect 1587 1663 1653 1679
rect 1587 1629 1603 1663
rect 1637 1647 1653 1663
rect 1637 1629 1853 1647
rect 1587 1613 1853 1629
rect 2235 1615 2437 1645
rect 1509 1467 2046 1501
rect 2235 1423 2265 1615
rect 1437 1378 1853 1409
rect 2215 1407 2281 1423
rect 2215 1373 2231 1407
rect 2265 1373 2281 1407
rect 2215 1357 2281 1373
<< polycont >>
rect 1667 2618 1701 2652
rect 1682 2034 1716 2068
rect 1603 1629 1637 1663
rect 2231 1373 2265 1407
<< locali >>
rect 1651 2652 1711 2668
rect 1651 2618 1667 2652
rect 1701 2618 1711 2652
rect 1651 2602 1711 2618
rect 1666 2068 1732 2084
rect 1666 2034 1682 2068
rect 1716 2034 1732 2068
rect 1666 2018 1732 2034
rect 1587 1663 1653 1679
rect 1587 1629 1603 1663
rect 1637 1629 1653 1663
rect 1587 1613 1653 1629
rect 2215 1407 2281 1423
rect 2215 1373 2231 1407
rect 2265 1373 2281 1407
rect 2215 1357 2281 1373
<< viali >>
rect 1667 2618 1701 2652
rect 1682 2034 1716 2068
rect 1603 1629 1637 1663
rect 2231 1373 2265 1407
<< metal1 >>
rect 1503 2763 2555 2769
rect 1503 2729 1515 2763
rect 1954 2729 2325 2763
rect 2521 2729 2555 2763
rect 1503 2723 2555 2729
rect 2848 2723 2980 2770
rect 2525 2722 2555 2723
rect 2928 2718 2980 2723
rect 1651 2652 1717 2668
rect 1583 2618 1667 2652
rect 1701 2618 1717 2652
rect 1651 2602 1717 2618
rect 1800 2471 1810 2523
rect 1862 2471 1872 2523
rect 1927 2515 2027 2549
rect 2386 2524 2389 2525
rect 2427 2524 2458 2525
rect 1426 2389 1502 2460
rect 1609 2402 1617 2440
rect 2054 2425 2064 2477
rect 2116 2425 2126 2477
rect 2162 2425 2172 2477
rect 2224 2425 2234 2477
rect 2386 2472 2396 2524
rect 2448 2472 2458 2524
rect 2649 2504 2869 2538
rect 1596 2374 1617 2402
rect 2317 2361 2327 2413
rect 2379 2361 2389 2413
rect 2482 2399 2678 2440
rect 2774 2398 2784 2450
rect 2836 2398 2846 2450
rect 1800 2236 1810 2289
rect 1862 2236 1872 2289
rect 2386 2286 2389 2288
rect 2427 2286 2458 2288
rect 2386 2234 2396 2286
rect 2448 2234 2458 2286
rect 1666 2068 1762 2084
rect 1666 2034 1682 2068
rect 1716 2034 1762 2068
rect 1666 2018 1762 2034
rect 1466 1963 1675 1969
rect 1466 1929 1478 1963
rect 1516 1929 1662 1963
rect 1663 1929 1675 1963
rect 1466 1925 1675 1929
rect 1704 1963 2832 1969
rect 1704 1929 1749 1963
rect 1924 1929 2677 1963
rect 2707 1929 2719 1963
rect 2773 1929 2785 1963
rect 2820 1929 2832 1963
rect 1704 1925 2832 1929
rect 1466 1923 2832 1925
rect 1663 1922 1709 1923
rect 2140 1806 2220 1858
rect 2272 1806 2346 1858
rect 2140 1802 2346 1806
rect 1587 1672 1653 1679
rect 1577 1620 1587 1672
rect 1639 1620 1653 1672
rect 1587 1613 1653 1620
rect 1800 1604 1810 1656
rect 1862 1604 1872 1656
rect 2382 1604 2392 1656
rect 2444 1604 2454 1656
rect 1440 1502 1775 1536
rect 2451 1499 2461 1551
rect 2513 1499 2523 1551
rect 1897 1442 2053 1494
rect 2215 1417 2281 1423
rect 1800 1365 1810 1417
rect 1862 1365 1872 1417
rect 2212 1365 2222 1417
rect 2274 1365 2284 1417
rect 2382 1365 2392 1417
rect 2444 1365 2454 1417
rect 2623 1415 2633 1467
rect 2685 1415 2695 1467
rect 2730 1413 2740 1465
rect 2792 1413 2802 1465
rect 2828 1377 2838 1395
rect 2215 1357 2281 1365
rect 2663 1343 2838 1377
rect 2890 1343 2900 1395
rect 2928 1169 2980 1175
rect 1408 1123 1718 1169
rect 2284 1123 2305 1169
rect 2535 1123 2556 1169
rect 2860 1123 2980 1169
<< via1 >>
rect 1810 2471 1862 2523
rect 2064 2425 2116 2477
rect 2172 2425 2224 2477
rect 2396 2472 2448 2524
rect 2327 2361 2379 2413
rect 2784 2398 2836 2450
rect 1810 2237 1862 2289
rect 2396 2234 2448 2286
rect 2220 1806 2272 1858
rect 1587 1663 1639 1672
rect 1587 1629 1603 1663
rect 1603 1629 1637 1663
rect 1637 1629 1639 1663
rect 1587 1620 1639 1629
rect 1810 1604 1862 1656
rect 2461 1499 2513 1551
rect 1810 1365 1862 1417
rect 2222 1407 2274 1417
rect 2222 1373 2231 1407
rect 2231 1373 2265 1407
rect 2265 1373 2274 1407
rect 2222 1365 2274 1373
rect 2392 1365 2444 1417
rect 2633 1415 2685 1467
rect 2740 1413 2792 1465
rect 2838 1343 2890 1395
<< metal2 >>
rect 1819 2577 2544 2611
rect 1819 2533 1853 2577
rect 1810 2523 1862 2533
rect 1587 2481 1810 2517
rect 1587 1682 1621 2481
rect 1810 2461 1862 2471
rect 1988 2524 2448 2549
rect 1988 2515 2396 2524
rect 1988 2445 2022 2515
rect 2064 2477 2116 2487
rect 1988 2314 2023 2445
rect 1810 2289 1862 2299
rect 1989 2279 2023 2314
rect 1862 2245 2023 2279
rect 2064 2398 2116 2425
rect 2172 2477 2224 2487
rect 2396 2462 2448 2472
rect 2172 2415 2224 2425
rect 1810 2227 1862 2237
rect 2064 2146 2098 2398
rect 1670 2112 2098 2146
rect 1587 1672 1639 1682
rect 1587 1610 1639 1620
rect 1670 1327 1704 2112
rect 2179 1868 2213 2415
rect 2327 2413 2379 2423
rect 2310 2361 2327 2413
rect 2310 2351 2379 2361
rect 2310 2064 2344 2351
rect 2396 2286 2448 2296
rect 2510 2282 2544 2577
rect 2776 2450 2890 2460
rect 2776 2398 2784 2450
rect 2836 2398 2890 2450
rect 2776 2388 2890 2398
rect 2448 2236 2544 2282
rect 2396 2224 2448 2234
rect 2310 2030 2572 2064
rect 2179 1858 2272 1868
rect 2179 1806 2220 1858
rect 2220 1796 2272 1806
rect 1810 1657 1862 1666
rect 1809 1656 1869 1657
rect 1809 1604 1810 1656
rect 1862 1604 1869 1656
rect 1809 1600 1869 1604
rect 1809 1566 2433 1600
rect 2399 1427 2433 1566
rect 2538 1561 2572 2030
rect 2461 1551 2572 1561
rect 2513 1499 2685 1551
rect 2461 1489 2513 1499
rect 2633 1467 2685 1499
rect 1810 1417 1862 1427
rect 2222 1417 2274 1427
rect 1862 1375 2222 1409
rect 1810 1355 1862 1365
rect 2222 1355 2274 1365
rect 2392 1417 2444 1427
rect 2444 1374 2448 1408
rect 2633 1405 2685 1415
rect 2740 1465 2792 1475
rect 2740 1403 2792 1413
rect 2392 1355 2444 1365
rect 2750 1327 2784 1403
rect 2838 1395 2890 2388
rect 2838 1333 2890 1343
rect 1435 1293 2785 1327
use tg  tg_3
timestamp 1615600491
transform 1 0 1747 0 1 1429
box -35 -326 258 621
use tg  tg_1
timestamp 1615600491
transform -1 0 2507 0 -1 2462
box -35 -326 258 621
use tg  tg_2
timestamp 1615600491
transform 1 0 2328 0 1 1429
box -35 -326 258 621
use tg  tg_0
timestamp 1615600491
transform -1 0 1926 0 -1 2462
box -35 -326 258 621
use nor  nor_1
timestamp 1615600491
transform -1 0 2844 0 1 1134
box -17 -20 296 869
use nor  nor_0
timestamp 1615600491
transform -1 0 2273 0 -1 2758
box -17 -20 296 869
use inverter  inverter_1
timestamp 1615600491
transform -1 0 2503 0 -1 2611
box -369 -159 -44 689
use inverter  inverter_2
timestamp 1615600491
transform 1 0 2332 0 1 1281
box -369 -159 -44 689
use inverter  inverter_0
timestamp 1615600491
transform 1 0 1769 0 -1 2611
box -369 -159 -44 689
<< labels >>
rlabel metal2 1435 1293 2785 1327 1 CLR
rlabel metal1 1426 2389 1502 2460 1 CLK
rlabel metal1 2649 2504 2869 2538 1 Qb
rlabel metal1 1440 1502 1775 1536 1 D
rlabel metal2 2776 2388 2890 2460 1 Q
<< end >>
