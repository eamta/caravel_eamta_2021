magic
tech sky130A
magscale 1 2
timestamp 1615910487
<< nwell >>
rect -1550 -764 1550 798
<< pmos >>
rect -1456 -664 -1316 736
rect -1258 -664 -1118 736
rect -1060 -664 -920 736
rect -862 -664 -722 736
rect -664 -664 -524 736
rect -466 -664 -326 736
rect -268 -664 -128 736
rect -70 -664 70 736
rect 128 -664 268 736
rect 326 -664 466 736
rect 524 -664 664 736
rect 722 -664 862 736
rect 920 -664 1060 736
rect 1118 -664 1258 736
rect 1316 -664 1456 736
<< pdiff >>
rect -1514 724 -1456 736
rect -1514 -652 -1502 724
rect -1468 -652 -1456 724
rect -1514 -664 -1456 -652
rect -1316 724 -1258 736
rect -1316 -652 -1304 724
rect -1270 -652 -1258 724
rect -1316 -664 -1258 -652
rect -1118 724 -1060 736
rect -1118 -652 -1106 724
rect -1072 -652 -1060 724
rect -1118 -664 -1060 -652
rect -920 724 -862 736
rect -920 -652 -908 724
rect -874 -652 -862 724
rect -920 -664 -862 -652
rect -722 724 -664 736
rect -722 -652 -710 724
rect -676 -652 -664 724
rect -722 -664 -664 -652
rect -524 724 -466 736
rect -524 -652 -512 724
rect -478 -652 -466 724
rect -524 -664 -466 -652
rect -326 724 -268 736
rect -326 -652 -314 724
rect -280 -652 -268 724
rect -326 -664 -268 -652
rect -128 724 -70 736
rect -128 -652 -116 724
rect -82 -652 -70 724
rect -128 -664 -70 -652
rect 70 724 128 736
rect 70 -652 82 724
rect 116 -652 128 724
rect 70 -664 128 -652
rect 268 724 326 736
rect 268 -652 280 724
rect 314 -652 326 724
rect 268 -664 326 -652
rect 466 724 524 736
rect 466 -652 478 724
rect 512 -652 524 724
rect 466 -664 524 -652
rect 664 724 722 736
rect 664 -652 676 724
rect 710 -652 722 724
rect 664 -664 722 -652
rect 862 724 920 736
rect 862 -652 874 724
rect 908 -652 920 724
rect 862 -664 920 -652
rect 1060 724 1118 736
rect 1060 -652 1072 724
rect 1106 -652 1118 724
rect 1060 -664 1118 -652
rect 1258 724 1316 736
rect 1258 -652 1270 724
rect 1304 -652 1316 724
rect 1258 -664 1316 -652
rect 1456 724 1514 736
rect 1456 -652 1468 724
rect 1502 -652 1514 724
rect 1456 -664 1514 -652
<< pdiffc >>
rect -1502 -652 -1468 724
rect -1304 -652 -1270 724
rect -1106 -652 -1072 724
rect -908 -652 -874 724
rect -710 -652 -676 724
rect -512 -652 -478 724
rect -314 -652 -280 724
rect -116 -652 -82 724
rect 82 -652 116 724
rect 280 -652 314 724
rect 478 -652 512 724
rect 676 -652 710 724
rect 874 -652 908 724
rect 1072 -652 1106 724
rect 1270 -652 1304 724
rect 1468 -652 1502 724
<< poly >>
rect -1456 736 -1316 762
rect -1258 736 -1118 762
rect -1060 736 -920 762
rect -862 736 -722 762
rect -664 736 -524 762
rect -466 736 -326 762
rect -268 736 -128 762
rect -70 736 70 762
rect 128 736 268 762
rect 326 736 466 762
rect 524 736 664 762
rect 722 736 862 762
rect 920 736 1060 762
rect 1118 736 1258 762
rect 1316 736 1456 762
rect -1456 -711 -1316 -664
rect -1456 -745 -1440 -711
rect -1332 -745 -1316 -711
rect -1456 -761 -1316 -745
rect -1258 -711 -1118 -664
rect -1258 -745 -1242 -711
rect -1134 -745 -1118 -711
rect -1258 -761 -1118 -745
rect -1060 -711 -920 -664
rect -1060 -745 -1044 -711
rect -936 -745 -920 -711
rect -1060 -761 -920 -745
rect -862 -711 -722 -664
rect -862 -745 -846 -711
rect -738 -745 -722 -711
rect -862 -761 -722 -745
rect -664 -711 -524 -664
rect -664 -745 -648 -711
rect -540 -745 -524 -711
rect -664 -761 -524 -745
rect -466 -711 -326 -664
rect -466 -745 -450 -711
rect -342 -745 -326 -711
rect -466 -761 -326 -745
rect -268 -711 -128 -664
rect -268 -745 -252 -711
rect -144 -745 -128 -711
rect -268 -761 -128 -745
rect -70 -711 70 -664
rect -70 -745 -54 -711
rect 54 -745 70 -711
rect -70 -761 70 -745
rect 128 -711 268 -664
rect 128 -745 144 -711
rect 252 -745 268 -711
rect 128 -761 268 -745
rect 326 -711 466 -664
rect 326 -745 342 -711
rect 450 -745 466 -711
rect 326 -761 466 -745
rect 524 -711 664 -664
rect 524 -745 540 -711
rect 648 -745 664 -711
rect 524 -761 664 -745
rect 722 -711 862 -664
rect 722 -745 738 -711
rect 846 -745 862 -711
rect 722 -761 862 -745
rect 920 -711 1060 -664
rect 920 -745 936 -711
rect 1044 -745 1060 -711
rect 920 -761 1060 -745
rect 1118 -711 1258 -664
rect 1118 -745 1134 -711
rect 1242 -745 1258 -711
rect 1118 -761 1258 -745
rect 1316 -711 1456 -664
rect 1316 -745 1332 -711
rect 1440 -745 1456 -711
rect 1316 -761 1456 -745
<< polycont >>
rect -1440 -745 -1332 -711
rect -1242 -745 -1134 -711
rect -1044 -745 -936 -711
rect -846 -745 -738 -711
rect -648 -745 -540 -711
rect -450 -745 -342 -711
rect -252 -745 -144 -711
rect -54 -745 54 -711
rect 144 -745 252 -711
rect 342 -745 450 -711
rect 540 -745 648 -711
rect 738 -745 846 -711
rect 936 -745 1044 -711
rect 1134 -745 1242 -711
rect 1332 -745 1440 -711
<< locali >>
rect -1502 724 -1468 740
rect -1502 -668 -1468 -652
rect -1304 724 -1270 740
rect -1304 -668 -1270 -652
rect -1106 724 -1072 740
rect -1106 -668 -1072 -652
rect -908 724 -874 740
rect -908 -668 -874 -652
rect -710 724 -676 740
rect -710 -668 -676 -652
rect -512 724 -478 740
rect -512 -668 -478 -652
rect -314 724 -280 740
rect -314 -668 -280 -652
rect -116 724 -82 740
rect -116 -668 -82 -652
rect 82 724 116 740
rect 82 -668 116 -652
rect 280 724 314 740
rect 280 -668 314 -652
rect 478 724 512 740
rect 478 -668 512 -652
rect 676 724 710 740
rect 676 -668 710 -652
rect 874 724 908 740
rect 874 -668 908 -652
rect 1072 724 1106 740
rect 1072 -668 1106 -652
rect 1270 724 1304 740
rect 1270 -668 1304 -652
rect 1468 724 1502 740
rect 1468 -668 1502 -652
rect -1456 -745 -1440 -711
rect -1332 -745 -1316 -711
rect -1258 -745 -1242 -711
rect -1134 -745 -1118 -711
rect -1060 -745 -1044 -711
rect -936 -745 -920 -711
rect -862 -745 -846 -711
rect -738 -745 -722 -711
rect -664 -745 -648 -711
rect -540 -745 -524 -711
rect -466 -745 -450 -711
rect -342 -745 -326 -711
rect -268 -745 -252 -711
rect -144 -745 -128 -711
rect -70 -745 -54 -711
rect 54 -745 70 -711
rect 128 -745 144 -711
rect 252 -745 268 -711
rect 326 -745 342 -711
rect 450 -745 466 -711
rect 524 -745 540 -711
rect 648 -745 664 -711
rect 722 -745 738 -711
rect 846 -745 862 -711
rect 920 -745 936 -711
rect 1044 -745 1060 -711
rect 1118 -745 1134 -711
rect 1242 -745 1258 -711
rect 1316 -745 1332 -711
rect 1440 -745 1456 -711
<< viali >>
rect -1502 -652 -1468 724
rect -1304 -652 -1270 724
rect -1106 -652 -1072 724
rect -908 -652 -874 724
rect -710 -652 -676 724
rect -512 -652 -478 724
rect -314 -652 -280 724
rect -116 -652 -82 724
rect 82 -652 116 724
rect 280 -652 314 724
rect 478 -652 512 724
rect 676 -652 710 724
rect 874 -652 908 724
rect 1072 -652 1106 724
rect 1270 -652 1304 724
rect 1468 -652 1502 724
rect -1440 -745 -1332 -711
rect -1242 -745 -1134 -711
rect -1044 -745 -936 -711
rect -846 -745 -738 -711
rect -648 -745 -540 -711
rect -450 -745 -342 -711
rect -252 -745 -144 -711
rect -54 -745 54 -711
rect 144 -745 252 -711
rect 342 -745 450 -711
rect 540 -745 648 -711
rect 738 -745 846 -711
rect 936 -745 1044 -711
rect 1134 -745 1242 -711
rect 1332 -745 1440 -711
<< metal1 >>
rect -1508 724 -1462 736
rect -1508 -652 -1502 724
rect -1468 -652 -1462 724
rect -1508 -664 -1462 -652
rect -1310 724 -1264 736
rect -1310 -652 -1304 724
rect -1270 -652 -1264 724
rect -1310 -664 -1264 -652
rect -1112 724 -1066 736
rect -1112 -652 -1106 724
rect -1072 -652 -1066 724
rect -1112 -664 -1066 -652
rect -914 724 -868 736
rect -914 -652 -908 724
rect -874 -652 -868 724
rect -914 -664 -868 -652
rect -716 724 -670 736
rect -716 -652 -710 724
rect -676 -652 -670 724
rect -716 -664 -670 -652
rect -518 724 -472 736
rect -518 -652 -512 724
rect -478 -652 -472 724
rect -518 -664 -472 -652
rect -320 724 -274 736
rect -320 -652 -314 724
rect -280 -652 -274 724
rect -320 -664 -274 -652
rect -122 724 -76 736
rect -122 -652 -116 724
rect -82 -652 -76 724
rect -122 -664 -76 -652
rect 76 724 122 736
rect 76 -652 82 724
rect 116 -652 122 724
rect 76 -664 122 -652
rect 274 724 320 736
rect 274 -652 280 724
rect 314 -652 320 724
rect 274 -664 320 -652
rect 472 724 518 736
rect 472 -652 478 724
rect 512 -652 518 724
rect 472 -664 518 -652
rect 670 724 716 736
rect 670 -652 676 724
rect 710 -652 716 724
rect 670 -664 716 -652
rect 868 724 914 736
rect 868 -652 874 724
rect 908 -652 914 724
rect 868 -664 914 -652
rect 1066 724 1112 736
rect 1066 -652 1072 724
rect 1106 -652 1112 724
rect 1066 -664 1112 -652
rect 1264 724 1310 736
rect 1264 -652 1270 724
rect 1304 -652 1310 724
rect 1264 -664 1310 -652
rect 1462 724 1508 736
rect 1462 -652 1468 724
rect 1502 -652 1508 724
rect 1462 -664 1508 -652
rect -1452 -711 -1320 -705
rect -1452 -745 -1440 -711
rect -1332 -745 -1320 -711
rect -1452 -751 -1320 -745
rect -1254 -711 -1122 -705
rect -1254 -745 -1242 -711
rect -1134 -745 -1122 -711
rect -1254 -751 -1122 -745
rect -1056 -711 -924 -705
rect -1056 -745 -1044 -711
rect -936 -745 -924 -711
rect -1056 -751 -924 -745
rect -858 -711 -726 -705
rect -858 -745 -846 -711
rect -738 -745 -726 -711
rect -858 -751 -726 -745
rect -660 -711 -528 -705
rect -660 -745 -648 -711
rect -540 -745 -528 -711
rect -660 -751 -528 -745
rect -462 -711 -330 -705
rect -462 -745 -450 -711
rect -342 -745 -330 -711
rect -462 -751 -330 -745
rect -264 -711 -132 -705
rect -264 -745 -252 -711
rect -144 -745 -132 -711
rect -264 -751 -132 -745
rect -66 -711 66 -705
rect -66 -745 -54 -711
rect 54 -745 66 -711
rect -66 -751 66 -745
rect 132 -711 264 -705
rect 132 -745 144 -711
rect 252 -745 264 -711
rect 132 -751 264 -745
rect 330 -711 462 -705
rect 330 -745 342 -711
rect 450 -745 462 -711
rect 330 -751 462 -745
rect 528 -711 660 -705
rect 528 -745 540 -711
rect 648 -745 660 -711
rect 528 -751 660 -745
rect 726 -711 858 -705
rect 726 -745 738 -711
rect 846 -745 858 -711
rect 726 -751 858 -745
rect 924 -711 1056 -705
rect 924 -745 936 -711
rect 1044 -745 1056 -711
rect 924 -751 1056 -745
rect 1122 -711 1254 -705
rect 1122 -745 1134 -711
rect 1242 -745 1254 -711
rect 1122 -751 1254 -745
rect 1320 -711 1452 -705
rect 1320 -745 1332 -711
rect 1440 -745 1452 -711
rect 1320 -751 1452 -745
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 1 nf 15 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
