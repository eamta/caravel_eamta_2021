magic
tech sky130A
magscale 1 2
timestamp 1624138001
<< error_s >>
rect 1837 756 1850 784
rect 1077 720 1088 748
rect 1124 686 1135 720
rect 1196 686 1205 748
rect 1884 722 1897 756
rect 1944 722 1965 784
rect 2069 756 2090 784
rect 2333 756 2354 784
rect 2116 722 2137 756
rect 2380 722 2401 756
rect 2404 722 2424 756
rect 2440 722 2461 784
rect 2857 756 2878 784
rect 2922 766 2938 772
rect 2894 756 2948 766
rect 3123 756 3144 784
rect 3188 766 3204 772
rect 3160 756 3214 766
rect 2888 746 2954 756
rect 2888 740 2925 746
rect 2904 722 2925 740
rect 2928 740 2954 746
rect 3154 746 3220 756
rect 3154 740 3191 746
rect 2928 722 2948 740
rect 3170 722 3191 740
rect 3194 740 3220 746
rect 3194 722 3214 740
rect 3230 722 3251 784
rect 3353 756 3376 784
rect 3418 766 3434 772
rect 3390 756 3444 766
rect 3384 746 3450 756
rect 3384 740 3423 746
rect 3400 722 3423 740
rect 3424 740 3450 746
rect 3424 722 3444 740
rect 3462 722 3481 784
rect 3589 756 3608 784
rect 3654 766 3670 772
rect 3626 756 3680 766
rect 3620 746 3686 756
rect 3620 740 3655 746
rect 3636 722 3655 740
rect 3660 740 3686 746
rect 3660 722 3680 740
rect 3694 722 3717 784
rect 1953 604 2081 625
rect 2147 594 2148 636
rect 2208 604 2266 625
rect 2998 604 3056 625
rect 3239 604 3367 625
rect 2000 578 2002 588
rect 2032 578 2034 588
rect 2000 568 2012 578
rect 2022 568 2034 578
rect 2189 578 2190 594
rect 2998 588 3014 594
rect 3318 588 3320 594
rect 2970 578 3024 588
rect 3276 578 3288 588
rect 3318 578 3330 588
rect 2189 554 2199 578
rect 2000 544 2034 552
rect 2189 544 2201 554
rect 2213 544 2233 578
rect 2964 568 3030 578
rect 2964 562 2990 568
rect 2980 544 2990 562
rect 3004 562 3030 568
rect 3270 568 3298 578
rect 3308 568 3336 578
rect 3270 562 3296 568
rect 3004 544 3024 562
rect 3286 554 3296 562
rect 3310 562 3336 568
rect 3310 554 3330 562
rect 3286 544 3330 554
rect 2296 510 2298 516
rect 2254 500 2266 510
rect 2296 500 2308 510
rect 3012 500 3014 542
rect 3304 534 3330 544
rect 3304 528 3320 534
rect 3086 510 3088 516
rect 3304 510 3320 516
rect 3044 500 3056 510
rect 3086 500 3098 510
rect 3276 500 3288 510
rect 3304 502 3330 510
rect 3318 500 3330 502
rect 2248 490 2276 500
rect 2286 490 2314 500
rect 2248 484 2274 490
rect 2264 466 2274 484
rect 2288 484 2314 490
rect 3038 490 3066 500
rect 3076 490 3104 500
rect 3038 484 3064 490
rect 2288 466 2308 484
rect 3054 476 3064 484
rect 3078 484 3104 490
rect 3270 492 3336 500
rect 3270 490 3298 492
rect 3308 490 3336 492
rect 3270 484 3296 490
rect 3078 476 3098 484
rect 3054 466 3098 476
rect 3286 476 3296 484
rect 3310 484 3336 490
rect 3310 476 3330 484
rect 3286 466 3298 476
rect 3308 466 3330 476
rect 2264 450 2298 460
rect 3072 456 3098 466
rect 3318 456 3330 466
rect 2449 424 2577 455
rect 3072 450 3088 456
rect 3318 450 3320 456
rect 3791 424 3919 455
rect 2528 418 2530 424
rect 3870 418 3872 424
rect 2486 408 2498 418
rect 2528 408 2540 418
rect 3828 408 3840 418
rect 3870 408 3882 418
rect 2480 398 2508 408
rect 2518 398 2546 408
rect 2480 392 2506 398
rect 2496 384 2506 392
rect 2520 392 2546 398
rect 3822 398 3850 408
rect 3860 398 3888 408
rect 3822 392 3848 398
rect 2520 384 2540 392
rect 2496 374 2508 384
rect 2518 374 2540 384
rect 3838 384 3848 392
rect 3862 392 3888 398
rect 3862 384 3882 392
rect 3838 374 3850 384
rect 3860 374 3882 384
rect 2528 364 2540 374
rect 3870 364 3882 374
rect 2528 358 2530 364
rect 3870 358 3872 364
rect 2820 350 2822 356
rect 3782 350 3786 356
rect 1340 340 1374 346
rect 2778 340 2790 350
rect 2820 340 2832 350
rect 3782 340 3796 350
rect 2114 306 2124 340
rect 2138 306 2158 340
rect 2772 330 2800 340
rect 2810 330 2838 340
rect 2772 324 2798 330
rect 2788 316 2798 324
rect 2812 324 2838 330
rect 2812 316 2832 324
rect 2788 306 2800 316
rect 2810 306 2832 316
rect 3170 306 3180 340
rect 3194 306 3214 340
rect 3752 306 3762 340
rect 3772 330 3802 340
rect 3776 324 3802 330
rect 3776 316 3796 324
rect 3772 306 3796 316
rect 2820 296 2832 306
rect 3782 296 3796 306
rect 2820 290 2822 296
rect 3782 290 3786 296
rect 2732 282 2748 288
rect 2714 272 2758 282
rect 2714 262 2764 272
rect 2738 256 2764 262
rect 2738 254 2758 256
rect 2714 238 2758 254
rect 2904 254 2914 272
rect 2904 238 2916 254
rect 2928 238 2948 272
rect 2732 228 2758 238
rect 2732 222 2748 228
rect 1846 188 1850 216
rect 1884 164 1894 188
rect 1908 164 1928 188
rect 1884 154 1928 164
rect 1944 154 1956 216
rect 2076 188 2090 216
rect 2342 188 2354 216
rect 2114 164 2128 188
rect 2138 164 2158 188
rect 2114 154 2158 164
rect 2380 164 2392 188
rect 2404 164 2424 188
rect 2380 154 2424 164
rect 2440 154 2452 216
rect 2866 188 2878 216
rect 3132 188 3144 216
rect 2904 164 2916 188
rect 2928 164 2948 188
rect 2904 154 2948 164
rect 3170 164 3182 188
rect 3194 164 3214 188
rect 3170 154 3214 164
rect 3230 154 3242 216
rect 3362 188 3376 216
rect 3400 164 3414 188
rect 3424 164 3444 188
rect 3400 154 3444 164
rect 3462 154 3472 216
rect 3598 188 3608 216
rect 3636 164 3646 188
rect 3660 164 3680 188
rect 3636 154 3680 164
rect 3694 154 3708 216
rect 1902 144 1928 154
rect 2132 144 2158 154
rect 2398 144 2424 154
rect 2922 144 2948 154
rect 3188 144 3214 154
rect 3418 144 3444 154
rect 3654 144 3680 154
rect 1902 138 1918 144
rect 2132 138 2148 144
rect 2398 138 2414 144
rect 2922 138 2938 144
rect 3188 138 3204 144
rect 3418 138 3434 144
rect 3654 138 3670 144
rect 1846 -154 1850 -126
rect 1902 -144 1918 -138
rect 1874 -154 1928 -144
rect 1868 -164 1934 -154
rect 1868 -170 1894 -164
rect 1884 -188 1894 -170
rect 1908 -170 1934 -164
rect 1908 -188 1928 -170
rect 1944 -188 1956 -126
rect 2076 -154 2090 -126
rect 2132 -144 2148 -138
rect 2104 -154 2158 -144
rect 2342 -154 2354 -126
rect 2398 -144 2414 -138
rect 2370 -154 2424 -144
rect 2098 -164 2164 -154
rect 2098 -170 2128 -164
rect 2114 -188 2128 -170
rect 2138 -170 2164 -164
rect 2364 -164 2430 -154
rect 2364 -170 2392 -164
rect 2138 -188 2158 -170
rect 2380 -188 2392 -170
rect 2404 -170 2430 -164
rect 2404 -188 2424 -170
rect 2440 -188 2452 -126
rect 2866 -154 2878 -126
rect 2922 -144 2938 -138
rect 2894 -154 2948 -144
rect 3132 -154 3144 -126
rect 3188 -144 3204 -138
rect 3160 -154 3214 -144
rect 2888 -164 2954 -154
rect 2888 -170 2916 -164
rect 2904 -188 2916 -170
rect 2928 -170 2954 -164
rect 3154 -164 3220 -154
rect 3154 -170 3182 -164
rect 2928 -188 2948 -170
rect 3170 -188 3182 -170
rect 3194 -170 3220 -164
rect 3194 -188 3214 -170
rect 3230 -188 3242 -126
rect 3362 -154 3376 -126
rect 3418 -144 3434 -138
rect 3390 -154 3444 -144
rect 3384 -164 3450 -154
rect 3384 -170 3414 -164
rect 3400 -188 3414 -170
rect 3424 -170 3450 -164
rect 3424 -188 3444 -170
rect 3462 -188 3472 -126
rect 3598 -154 3608 -126
rect 3654 -144 3670 -138
rect 3626 -154 3680 -144
rect 3620 -164 3686 -154
rect 3620 -170 3646 -164
rect 3636 -188 3646 -170
rect 3660 -170 3686 -164
rect 3660 -188 3680 -170
rect 3694 -188 3708 -126
rect 2732 -216 2786 -200
rect 2866 -216 2878 -200
rect 2732 -228 2748 -222
rect 2714 -238 2758 -228
rect 2714 -248 2764 -238
rect 2738 -254 2764 -248
rect 2738 -262 2758 -254
rect 2714 -272 2758 -262
rect 2904 -272 2914 -238
rect 2928 -272 2948 -238
rect 2732 -282 2758 -272
rect 2732 -288 2748 -282
rect 2820 -296 2822 -290
rect 3782 -296 3786 -290
rect 1302 -308 1412 -302
rect 2778 -306 2790 -296
rect 2820 -306 2832 -296
rect 3782 -306 3796 -296
rect 2114 -340 2124 -306
rect 2138 -340 2158 -306
rect 2772 -316 2800 -306
rect 2810 -316 2838 -306
rect 2772 -322 2798 -316
rect 2788 -330 2798 -322
rect 2812 -322 2838 -316
rect 2812 -330 2832 -322
rect 2788 -340 2800 -330
rect 2810 -340 2832 -330
rect 3170 -340 3180 -306
rect 3194 -340 3214 -306
rect 3752 -340 3762 -306
rect 3772 -316 3802 -306
rect 3776 -322 3802 -316
rect 3776 -330 3796 -322
rect 3772 -340 3796 -330
rect 2820 -350 2832 -340
rect 3782 -350 3796 -340
rect 2820 -356 2822 -350
rect 3782 -356 3786 -350
rect 2528 -364 2530 -358
rect 3870 -364 3872 -358
rect 2486 -374 2498 -364
rect 2528 -374 2540 -364
rect 3828 -374 3840 -364
rect 3870 -374 3882 -364
rect 2480 -377 2508 -374
rect 2518 -377 2546 -374
rect 2480 -390 2546 -377
rect 3822 -377 3850 -374
rect 3860 -377 3888 -374
rect 3822 -390 3888 -377
rect 2496 -408 2540 -390
rect 3838 -408 3882 -390
rect 2222 -418 2296 -408
rect 2528 -418 2540 -408
rect 3870 -418 3882 -408
rect 2528 -424 2530 -418
rect 3870 -424 3872 -418
rect 3012 -466 3014 -424
rect 3072 -456 3088 -450
rect 3318 -456 3320 -450
rect 3044 -466 3098 -456
rect 3276 -466 3288 -456
rect 3318 -466 3330 -456
rect 2264 -490 2274 -466
rect 2288 -490 2308 -466
rect 3038 -476 3104 -466
rect 3038 -482 3064 -476
rect 2264 -500 2276 -490
rect 2286 -500 2308 -490
rect 3054 -490 3064 -482
rect 3078 -482 3104 -476
rect 3270 -476 3298 -466
rect 3308 -476 3336 -466
rect 3270 -482 3296 -476
rect 3078 -490 3098 -482
rect 3286 -484 3296 -482
rect 3054 -500 3066 -490
rect 3076 -500 3098 -490
rect 3272 -490 3296 -484
rect 3310 -482 3336 -476
rect 3310 -484 3330 -482
rect 3310 -490 3334 -484
rect 3272 -492 3298 -490
rect 3308 -492 3334 -490
rect 3272 -500 3334 -492
rect 2147 -544 2148 -502
rect 2296 -510 2308 -500
rect 3086 -510 3098 -500
rect 3318 -502 3330 -500
rect 3304 -510 3330 -502
rect 2296 -516 2298 -510
rect 3086 -516 3088 -510
rect 3304 -516 3320 -510
rect 3304 -534 3320 -528
rect 2179 -544 2191 -534
rect 3276 -544 3330 -534
rect 2000 -552 2034 -544
rect 2173 -554 2201 -544
rect 2173 -557 2199 -554
rect 2213 -557 2233 -544
rect 2000 -578 2034 -557
rect 2173 -560 2233 -557
rect 2189 -578 2233 -560
rect 2980 -557 2990 -544
rect 3004 -557 3024 -544
rect 2980 -578 3024 -557
rect 3270 -554 3336 -544
rect 3270 -557 3296 -554
rect 3310 -557 3336 -554
rect 3270 -560 3336 -557
rect 3286 -578 3330 -560
rect 2189 -594 2190 -578
rect 2998 -588 3024 -578
rect 3318 -588 3330 -578
rect 2998 -594 3014 -588
rect 3318 -594 3320 -588
rect 2208 -609 2238 -604
rect 1077 -686 1088 -639
rect 1124 -720 1135 -686
rect 1196 -720 1205 -639
rect 1837 -722 1850 -675
rect 1884 -756 1897 -722
rect 1944 -756 1965 -675
rect 2069 -722 2090 -675
rect 2333 -722 2354 -675
rect 2116 -756 2137 -722
rect 2380 -756 2401 -722
rect 2404 -756 2424 -722
rect 2440 -756 2461 -675
rect 2857 -722 2878 -675
rect 3123 -722 3144 -675
rect 2904 -746 2925 -722
rect 2928 -746 2948 -722
rect 2904 -756 2948 -746
rect 3170 -746 3191 -722
rect 3194 -746 3214 -722
rect 3170 -756 3214 -746
rect 3230 -756 3251 -675
rect 3353 -722 3376 -675
rect 3400 -746 3423 -722
rect 3424 -746 3444 -722
rect 3400 -756 3444 -746
rect 3462 -756 3481 -675
rect 3589 -722 3608 -675
rect 3636 -746 3655 -722
rect 3660 -746 3680 -722
rect 3636 -756 3680 -746
rect 3694 -756 3717 -675
rect 2922 -766 2948 -756
rect 3188 -766 3214 -756
rect 3418 -766 3444 -756
rect 3654 -766 3680 -756
rect 2922 -772 2938 -766
rect 3188 -772 3204 -766
rect 3418 -772 3434 -766
rect 3654 -772 3670 -766
rect 1837 -1064 1850 -1036
rect 1077 -1100 1088 -1072
rect 1124 -1134 1135 -1100
rect 1196 -1134 1205 -1072
rect 1884 -1098 1897 -1064
rect 1944 -1098 1965 -1036
rect 2069 -1064 2090 -1036
rect 2333 -1064 2354 -1036
rect 2116 -1098 2137 -1064
rect 2380 -1098 2401 -1064
rect 2404 -1098 2424 -1064
rect 2440 -1098 2461 -1036
rect 2857 -1064 2878 -1036
rect 2922 -1054 2938 -1048
rect 2894 -1064 2948 -1054
rect 3123 -1064 3144 -1036
rect 3188 -1054 3204 -1048
rect 3160 -1064 3214 -1054
rect 2888 -1074 2954 -1064
rect 2888 -1080 2925 -1074
rect 2904 -1098 2925 -1080
rect 2928 -1080 2954 -1074
rect 3154 -1074 3220 -1064
rect 3154 -1080 3191 -1074
rect 2928 -1098 2948 -1080
rect 3170 -1098 3191 -1080
rect 3194 -1080 3220 -1074
rect 3194 -1098 3214 -1080
rect 3230 -1098 3251 -1036
rect 3353 -1064 3376 -1036
rect 3418 -1054 3434 -1048
rect 3390 -1064 3444 -1054
rect 3384 -1074 3450 -1064
rect 3384 -1080 3423 -1074
rect 3400 -1098 3423 -1080
rect 3424 -1080 3450 -1074
rect 3424 -1098 3444 -1080
rect 3462 -1098 3481 -1036
rect 3589 -1064 3608 -1036
rect 3654 -1054 3670 -1048
rect 3626 -1064 3680 -1054
rect 3620 -1074 3686 -1064
rect 3620 -1080 3655 -1074
rect 3636 -1098 3655 -1080
rect 3660 -1080 3686 -1074
rect 3660 -1098 3680 -1080
rect 3694 -1098 3717 -1036
rect 1953 -1216 2081 -1195
rect 2147 -1226 2148 -1184
rect 2208 -1216 2266 -1195
rect 2998 -1216 3056 -1195
rect 3239 -1216 3367 -1195
rect 2000 -1242 2002 -1232
rect 2032 -1242 2034 -1232
rect 2000 -1252 2012 -1242
rect 2022 -1252 2034 -1242
rect 2189 -1242 2190 -1226
rect 2998 -1232 3014 -1226
rect 3318 -1232 3320 -1226
rect 2970 -1242 3024 -1232
rect 3276 -1242 3288 -1232
rect 3318 -1242 3330 -1232
rect 2189 -1266 2199 -1242
rect 2000 -1276 2034 -1268
rect 2189 -1276 2201 -1266
rect 2213 -1276 2233 -1242
rect 2964 -1252 3030 -1242
rect 2964 -1258 2990 -1252
rect 2980 -1276 2990 -1258
rect 3004 -1258 3030 -1252
rect 3270 -1252 3298 -1242
rect 3308 -1252 3336 -1242
rect 3270 -1258 3296 -1252
rect 3004 -1276 3024 -1258
rect 3286 -1266 3296 -1258
rect 3310 -1258 3336 -1252
rect 3310 -1266 3330 -1258
rect 3286 -1276 3330 -1266
rect 2296 -1310 2298 -1304
rect 2254 -1320 2266 -1310
rect 2296 -1320 2308 -1310
rect 3012 -1320 3014 -1278
rect 3304 -1286 3330 -1276
rect 3304 -1292 3320 -1286
rect 3086 -1310 3088 -1304
rect 3304 -1310 3320 -1304
rect 3044 -1320 3056 -1310
rect 3086 -1320 3098 -1310
rect 3276 -1320 3288 -1310
rect 3304 -1318 3330 -1310
rect 3318 -1320 3330 -1318
rect 2248 -1330 2276 -1320
rect 2286 -1330 2314 -1320
rect 2248 -1336 2274 -1330
rect 2264 -1354 2274 -1336
rect 2288 -1336 2314 -1330
rect 3038 -1330 3066 -1320
rect 3076 -1330 3104 -1320
rect 3038 -1336 3064 -1330
rect 2288 -1354 2308 -1336
rect 3054 -1344 3064 -1336
rect 3078 -1336 3104 -1330
rect 3270 -1328 3336 -1320
rect 3270 -1330 3298 -1328
rect 3308 -1330 3336 -1328
rect 3270 -1336 3296 -1330
rect 3078 -1344 3098 -1336
rect 3054 -1354 3098 -1344
rect 3286 -1344 3296 -1336
rect 3310 -1336 3336 -1330
rect 3310 -1344 3330 -1336
rect 3286 -1354 3298 -1344
rect 3308 -1354 3330 -1344
rect 2264 -1370 2298 -1360
rect 3072 -1364 3098 -1354
rect 3318 -1364 3330 -1354
rect 2449 -1396 2577 -1365
rect 3072 -1370 3088 -1364
rect 3318 -1370 3320 -1364
rect 3791 -1396 3919 -1365
rect 2528 -1402 2530 -1396
rect 3870 -1402 3872 -1396
rect 2486 -1412 2498 -1402
rect 2528 -1412 2540 -1402
rect 3828 -1412 3840 -1402
rect 3870 -1412 3882 -1402
rect 2480 -1422 2508 -1412
rect 2518 -1422 2546 -1412
rect 2480 -1428 2506 -1422
rect 2496 -1436 2506 -1428
rect 2520 -1428 2546 -1422
rect 3822 -1422 3850 -1412
rect 3860 -1422 3888 -1412
rect 3822 -1428 3848 -1422
rect 2520 -1436 2540 -1428
rect 2496 -1446 2508 -1436
rect 2518 -1446 2540 -1436
rect 3838 -1436 3848 -1428
rect 3862 -1428 3888 -1422
rect 3862 -1436 3882 -1428
rect 3838 -1446 3850 -1436
rect 3860 -1446 3882 -1436
rect 2528 -1456 2540 -1446
rect 3870 -1456 3882 -1446
rect 2528 -1462 2530 -1456
rect 3870 -1462 3872 -1456
rect 2820 -1470 2822 -1464
rect 3782 -1470 3786 -1464
rect 1340 -1480 1374 -1474
rect 2778 -1480 2790 -1470
rect 2820 -1480 2832 -1470
rect 3782 -1480 3796 -1470
rect 2114 -1514 2124 -1480
rect 2138 -1514 2158 -1480
rect 2772 -1490 2800 -1480
rect 2810 -1490 2838 -1480
rect 2772 -1496 2798 -1490
rect 2788 -1504 2798 -1496
rect 2812 -1496 2838 -1490
rect 2812 -1504 2832 -1496
rect 2788 -1514 2800 -1504
rect 2810 -1514 2832 -1504
rect 3170 -1514 3180 -1480
rect 3194 -1514 3214 -1480
rect 3752 -1514 3762 -1480
rect 3772 -1490 3802 -1480
rect 3776 -1496 3802 -1490
rect 3776 -1504 3796 -1496
rect 3772 -1514 3796 -1504
rect 2820 -1524 2832 -1514
rect 3782 -1524 3796 -1514
rect 2820 -1530 2822 -1524
rect 3782 -1530 3786 -1524
rect 2732 -1538 2748 -1532
rect 2714 -1548 2758 -1538
rect 2714 -1558 2764 -1548
rect 2738 -1564 2764 -1558
rect 2738 -1566 2758 -1564
rect 2714 -1582 2758 -1566
rect 2904 -1566 2914 -1548
rect 2904 -1582 2916 -1566
rect 2928 -1582 2948 -1548
rect 2732 -1592 2758 -1582
rect 2732 -1598 2748 -1592
rect 1846 -1632 1850 -1604
rect 1884 -1656 1894 -1632
rect 1908 -1656 1928 -1632
rect 1884 -1666 1928 -1656
rect 1944 -1666 1956 -1604
rect 2076 -1632 2090 -1604
rect 2342 -1632 2354 -1604
rect 2114 -1656 2128 -1632
rect 2138 -1656 2158 -1632
rect 2114 -1666 2158 -1656
rect 2380 -1656 2392 -1632
rect 2404 -1656 2424 -1632
rect 2380 -1666 2424 -1656
rect 2440 -1666 2452 -1604
rect 2866 -1632 2878 -1604
rect 3132 -1632 3144 -1604
rect 2904 -1656 2916 -1632
rect 2928 -1656 2948 -1632
rect 2904 -1666 2948 -1656
rect 3170 -1656 3182 -1632
rect 3194 -1656 3214 -1632
rect 3170 -1666 3214 -1656
rect 3230 -1666 3242 -1604
rect 3362 -1632 3376 -1604
rect 3400 -1656 3414 -1632
rect 3424 -1656 3444 -1632
rect 3400 -1666 3444 -1656
rect 3462 -1666 3472 -1604
rect 3598 -1632 3608 -1604
rect 3636 -1656 3646 -1632
rect 3660 -1656 3680 -1632
rect 3636 -1666 3680 -1656
rect 3694 -1666 3708 -1604
rect 1902 -1676 1928 -1666
rect 2132 -1676 2158 -1666
rect 2398 -1676 2424 -1666
rect 2922 -1676 2948 -1666
rect 3188 -1676 3214 -1666
rect 3418 -1676 3444 -1666
rect 3654 -1676 3680 -1666
rect 1902 -1682 1918 -1676
rect 2132 -1682 2148 -1676
rect 2398 -1682 2414 -1676
rect 2922 -1682 2938 -1676
rect 3188 -1682 3204 -1676
rect 3418 -1682 3434 -1676
rect 3654 -1682 3670 -1676
rect 1846 -1974 1850 -1946
rect 1902 -1964 1918 -1958
rect 1874 -1974 1928 -1964
rect 1868 -1984 1934 -1974
rect 1868 -1990 1894 -1984
rect 1884 -2008 1894 -1990
rect 1908 -1990 1934 -1984
rect 1908 -2008 1928 -1990
rect 1944 -2008 1956 -1946
rect 2076 -1974 2090 -1946
rect 2132 -1964 2148 -1958
rect 2104 -1974 2158 -1964
rect 2342 -1974 2354 -1946
rect 2398 -1964 2414 -1958
rect 2370 -1974 2424 -1964
rect 2098 -1984 2164 -1974
rect 2098 -1990 2128 -1984
rect 2114 -2008 2128 -1990
rect 2138 -1990 2164 -1984
rect 2364 -1984 2430 -1974
rect 2364 -1990 2392 -1984
rect 2138 -2008 2158 -1990
rect 2380 -2008 2392 -1990
rect 2404 -1990 2430 -1984
rect 2404 -2008 2424 -1990
rect 2440 -2008 2452 -1946
rect 2866 -1974 2878 -1946
rect 2922 -1964 2938 -1958
rect 2894 -1974 2948 -1964
rect 3132 -1974 3144 -1946
rect 3188 -1964 3204 -1958
rect 3160 -1974 3214 -1964
rect 2888 -1984 2954 -1974
rect 2888 -1990 2916 -1984
rect 2904 -2008 2916 -1990
rect 2928 -1990 2954 -1984
rect 3154 -1984 3220 -1974
rect 3154 -1990 3182 -1984
rect 2928 -2008 2948 -1990
rect 3170 -2008 3182 -1990
rect 3194 -1990 3220 -1984
rect 3194 -2008 3214 -1990
rect 3230 -2008 3242 -1946
rect 3362 -1974 3376 -1946
rect 3418 -1964 3434 -1958
rect 3390 -1974 3444 -1964
rect 3384 -1984 3450 -1974
rect 3384 -1990 3414 -1984
rect 3400 -2008 3414 -1990
rect 3424 -1990 3450 -1984
rect 3424 -2008 3444 -1990
rect 3462 -2008 3472 -1946
rect 3598 -1974 3608 -1946
rect 3654 -1964 3670 -1958
rect 3626 -1974 3680 -1964
rect 3620 -1984 3686 -1974
rect 3620 -1990 3646 -1984
rect 3636 -2008 3646 -1990
rect 3660 -1990 3686 -1984
rect 3660 -2008 3680 -1990
rect 3694 -2008 3708 -1946
rect 2732 -2036 2786 -2020
rect 2866 -2036 2878 -2020
rect 2732 -2048 2748 -2042
rect 2714 -2058 2758 -2048
rect 2714 -2068 2764 -2058
rect 2738 -2074 2764 -2068
rect 2738 -2082 2758 -2074
rect 2714 -2092 2758 -2082
rect 2904 -2092 2914 -2058
rect 2928 -2092 2948 -2058
rect 2732 -2102 2758 -2092
rect 2732 -2108 2748 -2102
rect 2820 -2116 2822 -2110
rect 3782 -2116 3786 -2110
rect 1302 -2128 1412 -2122
rect 2778 -2126 2790 -2116
rect 2820 -2126 2832 -2116
rect 3782 -2126 3796 -2116
rect 2114 -2160 2124 -2126
rect 2138 -2160 2158 -2126
rect 2772 -2136 2800 -2126
rect 2810 -2136 2838 -2126
rect 2772 -2142 2798 -2136
rect 2788 -2150 2798 -2142
rect 2812 -2142 2838 -2136
rect 2812 -2150 2832 -2142
rect 2788 -2160 2800 -2150
rect 2810 -2160 2832 -2150
rect 3170 -2160 3180 -2126
rect 3194 -2160 3214 -2126
rect 3752 -2160 3762 -2126
rect 3772 -2136 3802 -2126
rect 3776 -2142 3802 -2136
rect 3776 -2150 3796 -2142
rect 3772 -2160 3796 -2150
rect 2820 -2170 2832 -2160
rect 3782 -2170 3796 -2160
rect 2820 -2176 2822 -2170
rect 3782 -2176 3786 -2170
rect 2528 -2184 2530 -2178
rect 3870 -2184 3872 -2178
rect 2486 -2194 2498 -2184
rect 2528 -2194 2540 -2184
rect 3828 -2194 3840 -2184
rect 3870 -2194 3882 -2184
rect 2480 -2197 2508 -2194
rect 2518 -2197 2546 -2194
rect 2480 -2210 2546 -2197
rect 3822 -2197 3850 -2194
rect 3860 -2197 3888 -2194
rect 3822 -2210 3888 -2197
rect 2496 -2228 2540 -2210
rect 3838 -2228 3882 -2210
rect 2222 -2238 2296 -2228
rect 2528 -2238 2540 -2228
rect 3870 -2238 3882 -2228
rect 2528 -2244 2530 -2238
rect 3870 -2244 3872 -2238
rect 3012 -2286 3014 -2244
rect 3072 -2276 3088 -2270
rect 3318 -2276 3320 -2270
rect 3044 -2286 3098 -2276
rect 3276 -2286 3288 -2276
rect 3318 -2286 3330 -2276
rect 2264 -2310 2274 -2286
rect 2288 -2310 2308 -2286
rect 3038 -2296 3104 -2286
rect 3038 -2302 3064 -2296
rect 2264 -2320 2276 -2310
rect 2286 -2320 2308 -2310
rect 3054 -2310 3064 -2302
rect 3078 -2302 3104 -2296
rect 3270 -2296 3298 -2286
rect 3308 -2296 3336 -2286
rect 3270 -2302 3296 -2296
rect 3078 -2310 3098 -2302
rect 3286 -2304 3296 -2302
rect 3054 -2320 3066 -2310
rect 3076 -2320 3098 -2310
rect 3272 -2310 3296 -2304
rect 3310 -2302 3336 -2296
rect 3310 -2304 3330 -2302
rect 3310 -2310 3334 -2304
rect 3272 -2312 3298 -2310
rect 3308 -2312 3334 -2310
rect 3272 -2320 3334 -2312
rect 2147 -2364 2148 -2322
rect 2296 -2330 2308 -2320
rect 3086 -2330 3098 -2320
rect 3318 -2322 3330 -2320
rect 3304 -2330 3330 -2322
rect 2296 -2336 2298 -2330
rect 3086 -2336 3088 -2330
rect 3304 -2336 3320 -2330
rect 3304 -2354 3320 -2348
rect 2179 -2364 2191 -2354
rect 3276 -2364 3330 -2354
rect 2000 -2372 2034 -2364
rect 2173 -2374 2201 -2364
rect 2173 -2377 2199 -2374
rect 2213 -2377 2233 -2364
rect 2000 -2398 2034 -2377
rect 2173 -2380 2233 -2377
rect 2189 -2398 2233 -2380
rect 2980 -2377 2990 -2364
rect 3004 -2377 3024 -2364
rect 2980 -2398 3024 -2377
rect 3270 -2374 3336 -2364
rect 3270 -2377 3296 -2374
rect 3310 -2377 3336 -2374
rect 3270 -2380 3336 -2377
rect 3286 -2398 3330 -2380
rect 2189 -2414 2190 -2398
rect 2998 -2408 3024 -2398
rect 3318 -2408 3330 -2398
rect 2998 -2414 3014 -2408
rect 3318 -2414 3320 -2408
rect 2208 -2429 2238 -2424
rect 1077 -2506 1088 -2459
rect 1124 -2540 1135 -2506
rect 1196 -2540 1205 -2459
rect 1837 -2542 1850 -2495
rect 1884 -2576 1897 -2542
rect 1944 -2576 1965 -2495
rect 2069 -2542 2090 -2495
rect 2333 -2542 2354 -2495
rect 2116 -2576 2137 -2542
rect 2380 -2576 2401 -2542
rect 2404 -2576 2424 -2542
rect 2440 -2576 2461 -2495
rect 2857 -2542 2878 -2495
rect 3123 -2542 3144 -2495
rect 2904 -2566 2925 -2542
rect 2928 -2566 2948 -2542
rect 2904 -2576 2948 -2566
rect 3170 -2566 3191 -2542
rect 3194 -2566 3214 -2542
rect 3170 -2576 3214 -2566
rect 3230 -2576 3251 -2495
rect 3353 -2542 3376 -2495
rect 3400 -2566 3423 -2542
rect 3424 -2566 3444 -2542
rect 3400 -2576 3444 -2566
rect 3462 -2576 3481 -2495
rect 3589 -2542 3608 -2495
rect 3636 -2566 3655 -2542
rect 3660 -2566 3680 -2542
rect 3636 -2576 3680 -2566
rect 3694 -2576 3717 -2495
rect 2922 -2586 2948 -2576
rect 3188 -2586 3214 -2576
rect 3418 -2586 3444 -2576
rect 3654 -2586 3680 -2576
rect 2922 -2592 2938 -2586
rect 3188 -2592 3204 -2586
rect 3418 -2592 3434 -2586
rect 3654 -2592 3670 -2586
<< metal1 >>
rect 0 872 3964 910
rect 0 -18 3964 20
rect 0 -929 3964 -891
rect 0 -1839 3964 -1801
rect 0 -2730 3964 -2692
<< metal2 >>
rect 386 429 456 499
rect 1788 448 1858 518
rect 552 -206 622 383
rect 2478 303 2548 373
rect 3894 254 3964 324
rect 386 -276 622 -206
rect 386 -466 456 -276
rect 3894 -324 3964 -254
rect 552 -1251 622 -383
rect 386 -1321 622 -1251
rect 386 -1364 456 -1321
rect 552 -2018 622 -1458
rect 3894 -1566 3964 -1496
rect 386 -2088 622 -2018
rect 386 -2251 456 -2088
rect 3894 -2144 3964 -2074
use counter1b  counter1b_3
timestamp 1624138001
transform 1 0 1668 0 -1 -1820
box -1668 0 2296 910
use counter1b  counter1b_2
timestamp 1624138001
transform 1 0 1668 0 1 -1820
box -1668 0 2296 910
use counter1b  counter1b_1
timestamp 1624138001
transform 1 0 1668 0 -1 0
box -1668 0 2296 910
use counter1b  counter1b_0
timestamp 1624138001
transform 1 0 1668 0 1 0
box -1668 0 2296 910
<< labels >>
rlabel metal2 420 429 420 429 5 CE
rlabel metal1 0 -2710 0 -2710 7 VDD
rlabel metal1 0 -1819 0 -1819 7 VSS
rlabel metal1 0 -907 0 -907 7 VDD
rlabel metal1 0 0 0 0 7 VSS
rlabel metal1 0 891 0 891 7 VDD
rlabel metal2 1823 448 1823 448 5 CLK
rlabel metal2 2513 303 2513 303 5 CLR
rlabel metal2 3929 254 3929 254 5 Q0
rlabel metal2 3930 -1566 3930 -1566 5 Q2
rlabel metal2 3929 -324 3929 -324 5 Q1
rlabel metal2 3929 -2144 3929 -2144 5 Q3
rlabel metal1 0 -2730 0 -2730 7 VDD
rlabel metal1 0 -929 0 -929 7 VDD
rlabel metal1 0 872 0 872 7 VDD
rlabel metal1 0 -18 0 -18 7 VSS
rlabel metal1 0 -1839 0 -1839 7 VSS
<< end >>
