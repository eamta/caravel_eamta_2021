magic
tech sky130A
magscale 1 2
timestamp 1623094427
<< pwell >>
rect -1127 -1710 1127 1710
<< nmos >>
rect -927 -1500 -897 1500
rect -831 -1500 -801 1500
rect -735 -1500 -705 1500
rect -639 -1500 -609 1500
rect -543 -1500 -513 1500
rect -447 -1500 -417 1500
rect -351 -1500 -321 1500
rect -255 -1500 -225 1500
rect -159 -1500 -129 1500
rect -63 -1500 -33 1500
rect 33 -1500 63 1500
rect 129 -1500 159 1500
rect 225 -1500 255 1500
rect 321 -1500 351 1500
rect 417 -1500 447 1500
rect 513 -1500 543 1500
rect 609 -1500 639 1500
rect 705 -1500 735 1500
rect 801 -1500 831 1500
rect 897 -1500 927 1500
<< ndiff >>
rect -989 1488 -927 1500
rect -989 -1488 -977 1488
rect -943 -1488 -927 1488
rect -989 -1500 -927 -1488
rect -897 1488 -831 1500
rect -897 -1488 -881 1488
rect -847 -1488 -831 1488
rect -897 -1500 -831 -1488
rect -801 1488 -735 1500
rect -801 -1488 -785 1488
rect -751 -1488 -735 1488
rect -801 -1500 -735 -1488
rect -705 1488 -639 1500
rect -705 -1488 -689 1488
rect -655 -1488 -639 1488
rect -705 -1500 -639 -1488
rect -609 1488 -543 1500
rect -609 -1488 -593 1488
rect -559 -1488 -543 1488
rect -609 -1500 -543 -1488
rect -513 1488 -447 1500
rect -513 -1488 -497 1488
rect -463 -1488 -447 1488
rect -513 -1500 -447 -1488
rect -417 1488 -351 1500
rect -417 -1488 -401 1488
rect -367 -1488 -351 1488
rect -417 -1500 -351 -1488
rect -321 1488 -255 1500
rect -321 -1488 -305 1488
rect -271 -1488 -255 1488
rect -321 -1500 -255 -1488
rect -225 1488 -159 1500
rect -225 -1488 -209 1488
rect -175 -1488 -159 1488
rect -225 -1500 -159 -1488
rect -129 1488 -63 1500
rect -129 -1488 -113 1488
rect -79 -1488 -63 1488
rect -129 -1500 -63 -1488
rect -33 1488 33 1500
rect -33 -1488 -17 1488
rect 17 -1488 33 1488
rect -33 -1500 33 -1488
rect 63 1488 129 1500
rect 63 -1488 79 1488
rect 113 -1488 129 1488
rect 63 -1500 129 -1488
rect 159 1488 225 1500
rect 159 -1488 175 1488
rect 209 -1488 225 1488
rect 159 -1500 225 -1488
rect 255 1488 321 1500
rect 255 -1488 271 1488
rect 305 -1488 321 1488
rect 255 -1500 321 -1488
rect 351 1488 417 1500
rect 351 -1488 367 1488
rect 401 -1488 417 1488
rect 351 -1500 417 -1488
rect 447 1488 513 1500
rect 447 -1488 463 1488
rect 497 -1488 513 1488
rect 447 -1500 513 -1488
rect 543 1488 609 1500
rect 543 -1488 559 1488
rect 593 -1488 609 1488
rect 543 -1500 609 -1488
rect 639 1488 705 1500
rect 639 -1488 655 1488
rect 689 -1488 705 1488
rect 639 -1500 705 -1488
rect 735 1488 801 1500
rect 735 -1488 751 1488
rect 785 -1488 801 1488
rect 735 -1500 801 -1488
rect 831 1488 897 1500
rect 831 -1488 847 1488
rect 881 -1488 897 1488
rect 831 -1500 897 -1488
rect 927 1488 989 1500
rect 927 -1488 943 1488
rect 977 -1488 989 1488
rect 927 -1500 989 -1488
<< ndiffc >>
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
<< psubdiff >>
rect -1091 -1640 -1057 1640
rect 1057 1578 1091 1640
rect 1057 -1640 1091 -1578
rect -1091 -1674 1091 -1640
<< psubdiffcont >>
rect 1057 -1578 1091 1578
<< poly >>
rect -927 1589 945 1614
rect -927 1554 -908 1589
rect 927 1554 945 1589
rect -927 1522 945 1554
rect -927 1500 -897 1522
rect -831 1500 -801 1522
rect -735 1500 -705 1522
rect -639 1500 -609 1522
rect -543 1500 -513 1522
rect -447 1500 -417 1522
rect -351 1500 -321 1522
rect -255 1500 -225 1522
rect -159 1500 -129 1522
rect -63 1500 -33 1522
rect 33 1500 63 1522
rect 129 1500 159 1522
rect 225 1500 255 1522
rect 321 1500 351 1522
rect 417 1500 447 1522
rect 513 1500 543 1522
rect 609 1500 639 1522
rect 705 1500 735 1522
rect 801 1500 831 1522
rect 897 1500 927 1522
rect -927 -1526 -897 -1500
rect -831 -1526 -801 -1500
rect -735 -1526 -705 -1500
rect -639 -1526 -609 -1500
rect -543 -1526 -513 -1500
rect -447 -1526 -417 -1500
rect -351 -1526 -321 -1500
rect -255 -1526 -225 -1500
rect -159 -1526 -129 -1500
rect -63 -1526 -33 -1500
rect 33 -1526 63 -1500
rect 129 -1526 159 -1500
rect 225 -1526 255 -1500
rect 321 -1526 351 -1500
rect 417 -1526 447 -1500
rect 513 -1526 543 -1500
rect 609 -1526 639 -1500
rect 705 -1526 735 -1500
rect 801 -1526 831 -1500
rect 897 -1526 927 -1500
<< polycont >>
rect -908 1554 927 1589
<< locali >>
rect -1091 -1640 -1057 1640
rect -924 1589 943 1605
rect -924 1554 -908 1589
rect 927 1554 943 1589
rect -924 1538 943 1554
rect 1057 1578 1091 1640
rect -977 1488 -943 1504
rect -977 -1504 -943 -1488
rect -881 1488 -847 1504
rect -881 -1504 -847 -1488
rect -785 1488 -751 1504
rect -785 -1504 -751 -1488
rect -689 1488 -655 1504
rect -689 -1504 -655 -1488
rect -593 1488 -559 1504
rect -593 -1504 -559 -1488
rect -497 1488 -463 1504
rect -497 -1504 -463 -1488
rect -401 1488 -367 1504
rect -401 -1504 -367 -1488
rect -305 1488 -271 1504
rect -305 -1504 -271 -1488
rect -209 1488 -175 1504
rect -209 -1504 -175 -1488
rect -113 1488 -79 1504
rect -113 -1504 -79 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 79 1488 113 1504
rect 79 -1504 113 -1488
rect 175 1488 209 1504
rect 175 -1504 209 -1488
rect 271 1488 305 1504
rect 271 -1504 305 -1488
rect 367 1488 401 1504
rect 367 -1504 401 -1488
rect 463 1488 497 1504
rect 463 -1504 497 -1488
rect 559 1488 593 1504
rect 559 -1504 593 -1488
rect 655 1488 689 1504
rect 655 -1504 689 -1488
rect 751 1488 785 1504
rect 751 -1504 785 -1488
rect 847 1488 881 1504
rect 847 -1504 881 -1488
rect 943 1488 977 1504
rect 943 -1504 977 -1488
rect 1057 -1640 1091 -1578
rect -1091 -1674 1091 -1640
<< viali >>
rect -908 1554 927 1589
rect -977 -1488 -943 1488
rect -881 -1488 -847 1488
rect -785 -1488 -751 1488
rect -689 -1488 -655 1488
rect -593 -1488 -559 1488
rect -497 -1488 -463 1488
rect -401 -1488 -367 1488
rect -305 -1488 -271 1488
rect -209 -1488 -175 1488
rect -113 -1488 -79 1488
rect -17 -1488 17 1488
rect 79 -1488 113 1488
rect 175 -1488 209 1488
rect 271 -1488 305 1488
rect 367 -1488 401 1488
rect 463 -1488 497 1488
rect 559 -1488 593 1488
rect 655 -1488 689 1488
rect 751 -1488 785 1488
rect 847 -1488 881 1488
rect 943 -1488 977 1488
<< metal1 >>
rect -926 1589 946 1614
rect -926 1554 -908 1589
rect 927 1554 946 1589
rect -926 1536 946 1554
rect -1002 -1504 -992 1504
rect -928 -1504 -918 1504
rect -887 1488 -841 1500
rect -887 -1488 -881 1488
rect -847 -1488 -841 1488
rect -887 -1568 -841 -1488
rect -810 -1504 -800 1504
rect -736 -1504 -726 1504
rect -695 1488 -649 1500
rect -695 -1488 -689 1488
rect -655 -1488 -649 1488
rect -695 -1568 -649 -1488
rect -618 -1504 -608 1504
rect -544 -1504 -534 1504
rect -503 1488 -457 1500
rect -503 -1488 -497 1488
rect -463 -1488 -457 1488
rect -503 -1568 -457 -1488
rect -426 -1504 -416 1504
rect -352 -1504 -342 1504
rect -311 1488 -265 1500
rect -311 -1488 -305 1488
rect -271 -1488 -265 1488
rect -311 -1568 -265 -1488
rect -234 -1504 -224 1504
rect -160 -1504 -150 1504
rect -119 1488 -73 1500
rect -119 -1488 -113 1488
rect -79 -1488 -73 1488
rect -119 -1568 -73 -1488
rect -42 -1504 -32 1504
rect 32 -1504 42 1504
rect 73 1488 119 1500
rect 73 -1488 79 1488
rect 113 -1488 119 1488
rect 73 -1568 119 -1488
rect 150 -1504 160 1504
rect 224 -1504 234 1504
rect 265 1488 311 1500
rect 265 -1488 271 1488
rect 305 -1488 311 1488
rect 265 -1568 311 -1488
rect 342 -1504 352 1504
rect 416 -1504 426 1504
rect 457 1488 503 1500
rect 457 -1488 463 1488
rect 497 -1488 503 1488
rect 457 -1568 503 -1488
rect 534 -1504 544 1504
rect 608 -1504 618 1504
rect 649 1488 695 1500
rect 649 -1488 655 1488
rect 689 -1488 695 1488
rect 649 -1568 695 -1488
rect 726 -1504 736 1504
rect 800 -1504 810 1504
rect 841 1488 887 1500
rect 841 -1488 847 1488
rect 881 -1488 887 1488
rect 841 -1568 887 -1488
rect 918 -1504 928 1504
rect 992 -1504 1002 1504
rect -887 -1573 887 -1568
rect -893 -1668 -883 -1573
rect 882 -1668 892 -1573
rect -887 -1674 887 -1668
<< via1 >>
rect -992 1488 -928 1504
rect -992 -1488 -977 1488
rect -977 -1488 -943 1488
rect -943 -1488 -928 1488
rect -992 -1504 -928 -1488
rect -800 1488 -736 1504
rect -800 -1488 -785 1488
rect -785 -1488 -751 1488
rect -751 -1488 -736 1488
rect -800 -1504 -736 -1488
rect -608 1488 -544 1504
rect -608 -1488 -593 1488
rect -593 -1488 -559 1488
rect -559 -1488 -544 1488
rect -608 -1504 -544 -1488
rect -416 1488 -352 1504
rect -416 -1488 -401 1488
rect -401 -1488 -367 1488
rect -367 -1488 -352 1488
rect -416 -1504 -352 -1488
rect -224 1488 -160 1504
rect -224 -1488 -209 1488
rect -209 -1488 -175 1488
rect -175 -1488 -160 1488
rect -224 -1504 -160 -1488
rect -32 1488 32 1504
rect -32 -1488 -17 1488
rect -17 -1488 17 1488
rect 17 -1488 32 1488
rect -32 -1504 32 -1488
rect 160 1488 224 1504
rect 160 -1488 175 1488
rect 175 -1488 209 1488
rect 209 -1488 224 1488
rect 160 -1504 224 -1488
rect 352 1488 416 1504
rect 352 -1488 367 1488
rect 367 -1488 401 1488
rect 401 -1488 416 1488
rect 352 -1504 416 -1488
rect 544 1488 608 1504
rect 544 -1488 559 1488
rect 559 -1488 593 1488
rect 593 -1488 608 1488
rect 544 -1504 608 -1488
rect 736 1488 800 1504
rect 736 -1488 751 1488
rect 751 -1488 785 1488
rect 785 -1488 800 1488
rect 736 -1504 800 -1488
rect 928 1488 992 1504
rect 928 -1488 943 1488
rect 943 -1488 977 1488
rect 977 -1488 992 1488
rect 928 -1504 992 -1488
rect -883 -1668 882 -1573
<< metal2 >>
rect -992 1514 992 1675
rect -992 1504 -928 1514
rect -992 -1514 -928 -1504
rect -800 1504 -736 1514
rect -800 -1514 -736 -1504
rect -608 1504 -544 1514
rect -608 -1514 -544 -1504
rect -416 1504 -352 1514
rect -416 -1514 -352 -1504
rect -224 1504 -160 1514
rect -224 -1514 -160 -1504
rect -32 1504 32 1514
rect -32 -1514 32 -1504
rect 160 1504 224 1514
rect 160 -1514 224 -1504
rect 352 1504 416 1514
rect 352 -1514 416 -1504
rect 544 1504 608 1514
rect 544 -1514 608 -1504
rect 736 1504 800 1514
rect 736 -1514 800 -1504
rect 928 1504 992 1514
rect 928 -1514 992 -1504
rect -883 -1573 882 -1563
rect -883 -1678 882 -1668
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -1074 -1657 1074 1657
string parameters w 15 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 0 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
