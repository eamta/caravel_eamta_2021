magic
tech sky130A
timestamp 1624052787
<< end >>
