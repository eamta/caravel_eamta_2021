magic
tech sky130A
magscale 1 2
timestamp 1616605166
<< error_p >>
rect -4685 222 -4627 228
rect -4493 222 -4435 228
rect -4301 222 -4243 228
rect -4109 222 -4051 228
rect -3917 222 -3859 228
rect -3725 222 -3667 228
rect -3533 222 -3475 228
rect -3341 222 -3283 228
rect -3149 222 -3091 228
rect -2957 222 -2899 228
rect -2765 222 -2707 228
rect -2573 222 -2515 228
rect -2381 222 -2323 228
rect -2189 222 -2131 228
rect -1997 222 -1939 228
rect -1805 222 -1747 228
rect -1613 222 -1555 228
rect -1421 222 -1363 228
rect -1229 222 -1171 228
rect -1037 222 -979 228
rect -845 222 -787 228
rect -653 222 -595 228
rect -461 222 -403 228
rect -269 222 -211 228
rect -77 222 -19 228
rect 115 222 173 228
rect 307 222 365 228
rect 499 222 557 228
rect 691 222 749 228
rect 883 222 941 228
rect 1075 222 1133 228
rect 1267 222 1325 228
rect 1459 222 1517 228
rect 1651 222 1709 228
rect 1843 222 1901 228
rect 2035 222 2093 228
rect 2227 222 2285 228
rect 2419 222 2477 228
rect 2611 222 2669 228
rect 2803 222 2861 228
rect 2995 222 3053 228
rect 3187 222 3245 228
rect 3379 222 3437 228
rect 3571 222 3629 228
rect 3763 222 3821 228
rect 3955 222 4013 228
rect 4147 222 4205 228
rect 4339 222 4397 228
rect 4531 222 4589 228
rect 4723 222 4781 228
rect -4685 188 -4673 222
rect -4493 188 -4481 222
rect -4301 188 -4289 222
rect -4109 188 -4097 222
rect -3917 188 -3905 222
rect -3725 188 -3713 222
rect -3533 188 -3521 222
rect -3341 188 -3329 222
rect -3149 188 -3137 222
rect -2957 188 -2945 222
rect -2765 188 -2753 222
rect -2573 188 -2561 222
rect -2381 188 -2369 222
rect -2189 188 -2177 222
rect -1997 188 -1985 222
rect -1805 188 -1793 222
rect -1613 188 -1601 222
rect -1421 188 -1409 222
rect -1229 188 -1217 222
rect -1037 188 -1025 222
rect -845 188 -833 222
rect -653 188 -641 222
rect -461 188 -449 222
rect -269 188 -257 222
rect -77 188 -65 222
rect 115 188 127 222
rect 307 188 319 222
rect 499 188 511 222
rect 691 188 703 222
rect 883 188 895 222
rect 1075 188 1087 222
rect 1267 188 1279 222
rect 1459 188 1471 222
rect 1651 188 1663 222
rect 1843 188 1855 222
rect 2035 188 2047 222
rect 2227 188 2239 222
rect 2419 188 2431 222
rect 2611 188 2623 222
rect 2803 188 2815 222
rect 2995 188 3007 222
rect 3187 188 3199 222
rect 3379 188 3391 222
rect 3571 188 3583 222
rect 3763 188 3775 222
rect 3955 188 3967 222
rect 4147 188 4159 222
rect 4339 188 4351 222
rect 4531 188 4543 222
rect 4723 188 4735 222
rect -4685 182 -4627 188
rect -4493 182 -4435 188
rect -4301 182 -4243 188
rect -4109 182 -4051 188
rect -3917 182 -3859 188
rect -3725 182 -3667 188
rect -3533 182 -3475 188
rect -3341 182 -3283 188
rect -3149 182 -3091 188
rect -2957 182 -2899 188
rect -2765 182 -2707 188
rect -2573 182 -2515 188
rect -2381 182 -2323 188
rect -2189 182 -2131 188
rect -1997 182 -1939 188
rect -1805 182 -1747 188
rect -1613 182 -1555 188
rect -1421 182 -1363 188
rect -1229 182 -1171 188
rect -1037 182 -979 188
rect -845 182 -787 188
rect -653 182 -595 188
rect -461 182 -403 188
rect -269 182 -211 188
rect -77 182 -19 188
rect 115 182 173 188
rect 307 182 365 188
rect 499 182 557 188
rect 691 182 749 188
rect 883 182 941 188
rect 1075 182 1133 188
rect 1267 182 1325 188
rect 1459 182 1517 188
rect 1651 182 1709 188
rect 1843 182 1901 188
rect 2035 182 2093 188
rect 2227 182 2285 188
rect 2419 182 2477 188
rect 2611 182 2669 188
rect 2803 182 2861 188
rect 2995 182 3053 188
rect 3187 182 3245 188
rect 3379 182 3437 188
rect 3571 182 3629 188
rect 3763 182 3821 188
rect 3955 182 4013 188
rect 4147 182 4205 188
rect 4339 182 4397 188
rect 4531 182 4589 188
rect 4723 182 4781 188
rect -4781 -188 -4723 -182
rect -4589 -188 -4531 -182
rect -4397 -188 -4339 -182
rect -4205 -188 -4147 -182
rect -4013 -188 -3955 -182
rect -3821 -188 -3763 -182
rect -3629 -188 -3571 -182
rect -3437 -188 -3379 -182
rect -3245 -188 -3187 -182
rect -3053 -188 -2995 -182
rect -2861 -188 -2803 -182
rect -2669 -188 -2611 -182
rect -2477 -188 -2419 -182
rect -2285 -188 -2227 -182
rect -2093 -188 -2035 -182
rect -1901 -188 -1843 -182
rect -1709 -188 -1651 -182
rect -1517 -188 -1459 -182
rect -1325 -188 -1267 -182
rect -1133 -188 -1075 -182
rect -941 -188 -883 -182
rect -749 -188 -691 -182
rect -557 -188 -499 -182
rect -365 -188 -307 -182
rect -173 -188 -115 -182
rect 19 -188 77 -182
rect 211 -188 269 -182
rect 403 -188 461 -182
rect 595 -188 653 -182
rect 787 -188 845 -182
rect 979 -188 1037 -182
rect 1171 -188 1229 -182
rect 1363 -188 1421 -182
rect 1555 -188 1613 -182
rect 1747 -188 1805 -182
rect 1939 -188 1997 -182
rect 2131 -188 2189 -182
rect 2323 -188 2381 -182
rect 2515 -188 2573 -182
rect 2707 -188 2765 -182
rect 2899 -188 2957 -182
rect 3091 -188 3149 -182
rect 3283 -188 3341 -182
rect 3475 -188 3533 -182
rect 3667 -188 3725 -182
rect 3859 -188 3917 -182
rect 4051 -188 4109 -182
rect 4243 -188 4301 -182
rect 4435 -188 4493 -182
rect 4627 -188 4685 -182
rect -4781 -222 -4769 -188
rect -4589 -222 -4577 -188
rect -4397 -222 -4385 -188
rect -4205 -222 -4193 -188
rect -4013 -222 -4001 -188
rect -3821 -222 -3809 -188
rect -3629 -222 -3617 -188
rect -3437 -222 -3425 -188
rect -3245 -222 -3233 -188
rect -3053 -222 -3041 -188
rect -2861 -222 -2849 -188
rect -2669 -222 -2657 -188
rect -2477 -222 -2465 -188
rect -2285 -222 -2273 -188
rect -2093 -222 -2081 -188
rect -1901 -222 -1889 -188
rect -1709 -222 -1697 -188
rect -1517 -222 -1505 -188
rect -1325 -222 -1313 -188
rect -1133 -222 -1121 -188
rect -941 -222 -929 -188
rect -749 -222 -737 -188
rect -557 -222 -545 -188
rect -365 -222 -353 -188
rect -173 -222 -161 -188
rect 19 -222 31 -188
rect 211 -222 223 -188
rect 403 -222 415 -188
rect 595 -222 607 -188
rect 787 -222 799 -188
rect 979 -222 991 -188
rect 1171 -222 1183 -188
rect 1363 -222 1375 -188
rect 1555 -222 1567 -188
rect 1747 -222 1759 -188
rect 1939 -222 1951 -188
rect 2131 -222 2143 -188
rect 2323 -222 2335 -188
rect 2515 -222 2527 -188
rect 2707 -222 2719 -188
rect 2899 -222 2911 -188
rect 3091 -222 3103 -188
rect 3283 -222 3295 -188
rect 3475 -222 3487 -188
rect 3667 -222 3679 -188
rect 3859 -222 3871 -188
rect 4051 -222 4063 -188
rect 4243 -222 4255 -188
rect 4435 -222 4447 -188
rect 4627 -222 4639 -188
rect -4781 -228 -4723 -222
rect -4589 -228 -4531 -222
rect -4397 -228 -4339 -222
rect -4205 -228 -4147 -222
rect -4013 -228 -3955 -222
rect -3821 -228 -3763 -222
rect -3629 -228 -3571 -222
rect -3437 -228 -3379 -222
rect -3245 -228 -3187 -222
rect -3053 -228 -2995 -222
rect -2861 -228 -2803 -222
rect -2669 -228 -2611 -222
rect -2477 -228 -2419 -222
rect -2285 -228 -2227 -222
rect -2093 -228 -2035 -222
rect -1901 -228 -1843 -222
rect -1709 -228 -1651 -222
rect -1517 -228 -1459 -222
rect -1325 -228 -1267 -222
rect -1133 -228 -1075 -222
rect -941 -228 -883 -222
rect -749 -228 -691 -222
rect -557 -228 -499 -222
rect -365 -228 -307 -222
rect -173 -228 -115 -222
rect 19 -228 77 -222
rect 211 -228 269 -222
rect 403 -228 461 -222
rect 595 -228 653 -222
rect 787 -228 845 -222
rect 979 -228 1037 -222
rect 1171 -228 1229 -222
rect 1363 -228 1421 -222
rect 1555 -228 1613 -222
rect 1747 -228 1805 -222
rect 1939 -228 1997 -222
rect 2131 -228 2189 -222
rect 2323 -228 2381 -222
rect 2515 -228 2573 -222
rect 2707 -228 2765 -222
rect 2899 -228 2957 -222
rect 3091 -228 3149 -222
rect 3283 -228 3341 -222
rect 3475 -228 3533 -222
rect 3667 -228 3725 -222
rect 3859 -228 3917 -222
rect 4051 -228 4109 -222
rect 4243 -228 4301 -222
rect 4435 -228 4493 -222
rect 4627 -228 4685 -222
<< pwell >>
rect -4967 -360 4967 360
<< nmos >>
rect -4767 -150 -4737 150
rect -4671 -150 -4641 150
rect -4575 -150 -4545 150
rect -4479 -150 -4449 150
rect -4383 -150 -4353 150
rect -4287 -150 -4257 150
rect -4191 -150 -4161 150
rect -4095 -150 -4065 150
rect -3999 -150 -3969 150
rect -3903 -150 -3873 150
rect -3807 -150 -3777 150
rect -3711 -150 -3681 150
rect -3615 -150 -3585 150
rect -3519 -150 -3489 150
rect -3423 -150 -3393 150
rect -3327 -150 -3297 150
rect -3231 -150 -3201 150
rect -3135 -150 -3105 150
rect -3039 -150 -3009 150
rect -2943 -150 -2913 150
rect -2847 -150 -2817 150
rect -2751 -150 -2721 150
rect -2655 -150 -2625 150
rect -2559 -150 -2529 150
rect -2463 -150 -2433 150
rect -2367 -150 -2337 150
rect -2271 -150 -2241 150
rect -2175 -150 -2145 150
rect -2079 -150 -2049 150
rect -1983 -150 -1953 150
rect -1887 -150 -1857 150
rect -1791 -150 -1761 150
rect -1695 -150 -1665 150
rect -1599 -150 -1569 150
rect -1503 -150 -1473 150
rect -1407 -150 -1377 150
rect -1311 -150 -1281 150
rect -1215 -150 -1185 150
rect -1119 -150 -1089 150
rect -1023 -150 -993 150
rect -927 -150 -897 150
rect -831 -150 -801 150
rect -735 -150 -705 150
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
rect 705 -150 735 150
rect 801 -150 831 150
rect 897 -150 927 150
rect 993 -150 1023 150
rect 1089 -150 1119 150
rect 1185 -150 1215 150
rect 1281 -150 1311 150
rect 1377 -150 1407 150
rect 1473 -150 1503 150
rect 1569 -150 1599 150
rect 1665 -150 1695 150
rect 1761 -150 1791 150
rect 1857 -150 1887 150
rect 1953 -150 1983 150
rect 2049 -150 2079 150
rect 2145 -150 2175 150
rect 2241 -150 2271 150
rect 2337 -150 2367 150
rect 2433 -150 2463 150
rect 2529 -150 2559 150
rect 2625 -150 2655 150
rect 2721 -150 2751 150
rect 2817 -150 2847 150
rect 2913 -150 2943 150
rect 3009 -150 3039 150
rect 3105 -150 3135 150
rect 3201 -150 3231 150
rect 3297 -150 3327 150
rect 3393 -150 3423 150
rect 3489 -150 3519 150
rect 3585 -150 3615 150
rect 3681 -150 3711 150
rect 3777 -150 3807 150
rect 3873 -150 3903 150
rect 3969 -150 3999 150
rect 4065 -150 4095 150
rect 4161 -150 4191 150
rect 4257 -150 4287 150
rect 4353 -150 4383 150
rect 4449 -150 4479 150
rect 4545 -150 4575 150
rect 4641 -150 4671 150
rect 4737 -150 4767 150
<< ndiff >>
rect -4829 138 -4767 150
rect -4829 -138 -4817 138
rect -4783 -138 -4767 138
rect -4829 -150 -4767 -138
rect -4737 138 -4671 150
rect -4737 -138 -4721 138
rect -4687 -138 -4671 138
rect -4737 -150 -4671 -138
rect -4641 138 -4575 150
rect -4641 -138 -4625 138
rect -4591 -138 -4575 138
rect -4641 -150 -4575 -138
rect -4545 138 -4479 150
rect -4545 -138 -4529 138
rect -4495 -138 -4479 138
rect -4545 -150 -4479 -138
rect -4449 138 -4383 150
rect -4449 -138 -4433 138
rect -4399 -138 -4383 138
rect -4449 -150 -4383 -138
rect -4353 138 -4287 150
rect -4353 -138 -4337 138
rect -4303 -138 -4287 138
rect -4353 -150 -4287 -138
rect -4257 138 -4191 150
rect -4257 -138 -4241 138
rect -4207 -138 -4191 138
rect -4257 -150 -4191 -138
rect -4161 138 -4095 150
rect -4161 -138 -4145 138
rect -4111 -138 -4095 138
rect -4161 -150 -4095 -138
rect -4065 138 -3999 150
rect -4065 -138 -4049 138
rect -4015 -138 -3999 138
rect -4065 -150 -3999 -138
rect -3969 138 -3903 150
rect -3969 -138 -3953 138
rect -3919 -138 -3903 138
rect -3969 -150 -3903 -138
rect -3873 138 -3807 150
rect -3873 -138 -3857 138
rect -3823 -138 -3807 138
rect -3873 -150 -3807 -138
rect -3777 138 -3711 150
rect -3777 -138 -3761 138
rect -3727 -138 -3711 138
rect -3777 -150 -3711 -138
rect -3681 138 -3615 150
rect -3681 -138 -3665 138
rect -3631 -138 -3615 138
rect -3681 -150 -3615 -138
rect -3585 138 -3519 150
rect -3585 -138 -3569 138
rect -3535 -138 -3519 138
rect -3585 -150 -3519 -138
rect -3489 138 -3423 150
rect -3489 -138 -3473 138
rect -3439 -138 -3423 138
rect -3489 -150 -3423 -138
rect -3393 138 -3327 150
rect -3393 -138 -3377 138
rect -3343 -138 -3327 138
rect -3393 -150 -3327 -138
rect -3297 138 -3231 150
rect -3297 -138 -3281 138
rect -3247 -138 -3231 138
rect -3297 -150 -3231 -138
rect -3201 138 -3135 150
rect -3201 -138 -3185 138
rect -3151 -138 -3135 138
rect -3201 -150 -3135 -138
rect -3105 138 -3039 150
rect -3105 -138 -3089 138
rect -3055 -138 -3039 138
rect -3105 -150 -3039 -138
rect -3009 138 -2943 150
rect -3009 -138 -2993 138
rect -2959 -138 -2943 138
rect -3009 -150 -2943 -138
rect -2913 138 -2847 150
rect -2913 -138 -2897 138
rect -2863 -138 -2847 138
rect -2913 -150 -2847 -138
rect -2817 138 -2751 150
rect -2817 -138 -2801 138
rect -2767 -138 -2751 138
rect -2817 -150 -2751 -138
rect -2721 138 -2655 150
rect -2721 -138 -2705 138
rect -2671 -138 -2655 138
rect -2721 -150 -2655 -138
rect -2625 138 -2559 150
rect -2625 -138 -2609 138
rect -2575 -138 -2559 138
rect -2625 -150 -2559 -138
rect -2529 138 -2463 150
rect -2529 -138 -2513 138
rect -2479 -138 -2463 138
rect -2529 -150 -2463 -138
rect -2433 138 -2367 150
rect -2433 -138 -2417 138
rect -2383 -138 -2367 138
rect -2433 -150 -2367 -138
rect -2337 138 -2271 150
rect -2337 -138 -2321 138
rect -2287 -138 -2271 138
rect -2337 -150 -2271 -138
rect -2241 138 -2175 150
rect -2241 -138 -2225 138
rect -2191 -138 -2175 138
rect -2241 -150 -2175 -138
rect -2145 138 -2079 150
rect -2145 -138 -2129 138
rect -2095 -138 -2079 138
rect -2145 -150 -2079 -138
rect -2049 138 -1983 150
rect -2049 -138 -2033 138
rect -1999 -138 -1983 138
rect -2049 -150 -1983 -138
rect -1953 138 -1887 150
rect -1953 -138 -1937 138
rect -1903 -138 -1887 138
rect -1953 -150 -1887 -138
rect -1857 138 -1791 150
rect -1857 -138 -1841 138
rect -1807 -138 -1791 138
rect -1857 -150 -1791 -138
rect -1761 138 -1695 150
rect -1761 -138 -1745 138
rect -1711 -138 -1695 138
rect -1761 -150 -1695 -138
rect -1665 138 -1599 150
rect -1665 -138 -1649 138
rect -1615 -138 -1599 138
rect -1665 -150 -1599 -138
rect -1569 138 -1503 150
rect -1569 -138 -1553 138
rect -1519 -138 -1503 138
rect -1569 -150 -1503 -138
rect -1473 138 -1407 150
rect -1473 -138 -1457 138
rect -1423 -138 -1407 138
rect -1473 -150 -1407 -138
rect -1377 138 -1311 150
rect -1377 -138 -1361 138
rect -1327 -138 -1311 138
rect -1377 -150 -1311 -138
rect -1281 138 -1215 150
rect -1281 -138 -1265 138
rect -1231 -138 -1215 138
rect -1281 -150 -1215 -138
rect -1185 138 -1119 150
rect -1185 -138 -1169 138
rect -1135 -138 -1119 138
rect -1185 -150 -1119 -138
rect -1089 138 -1023 150
rect -1089 -138 -1073 138
rect -1039 -138 -1023 138
rect -1089 -150 -1023 -138
rect -993 138 -927 150
rect -993 -138 -977 138
rect -943 -138 -927 138
rect -993 -150 -927 -138
rect -897 138 -831 150
rect -897 -138 -881 138
rect -847 -138 -831 138
rect -897 -150 -831 -138
rect -801 138 -735 150
rect -801 -138 -785 138
rect -751 -138 -735 138
rect -801 -150 -735 -138
rect -705 138 -639 150
rect -705 -138 -689 138
rect -655 -138 -639 138
rect -705 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 705 150
rect 639 -138 655 138
rect 689 -138 705 138
rect 639 -150 705 -138
rect 735 138 801 150
rect 735 -138 751 138
rect 785 -138 801 138
rect 735 -150 801 -138
rect 831 138 897 150
rect 831 -138 847 138
rect 881 -138 897 138
rect 831 -150 897 -138
rect 927 138 993 150
rect 927 -138 943 138
rect 977 -138 993 138
rect 927 -150 993 -138
rect 1023 138 1089 150
rect 1023 -138 1039 138
rect 1073 -138 1089 138
rect 1023 -150 1089 -138
rect 1119 138 1185 150
rect 1119 -138 1135 138
rect 1169 -138 1185 138
rect 1119 -150 1185 -138
rect 1215 138 1281 150
rect 1215 -138 1231 138
rect 1265 -138 1281 138
rect 1215 -150 1281 -138
rect 1311 138 1377 150
rect 1311 -138 1327 138
rect 1361 -138 1377 138
rect 1311 -150 1377 -138
rect 1407 138 1473 150
rect 1407 -138 1423 138
rect 1457 -138 1473 138
rect 1407 -150 1473 -138
rect 1503 138 1569 150
rect 1503 -138 1519 138
rect 1553 -138 1569 138
rect 1503 -150 1569 -138
rect 1599 138 1665 150
rect 1599 -138 1615 138
rect 1649 -138 1665 138
rect 1599 -150 1665 -138
rect 1695 138 1761 150
rect 1695 -138 1711 138
rect 1745 -138 1761 138
rect 1695 -150 1761 -138
rect 1791 138 1857 150
rect 1791 -138 1807 138
rect 1841 -138 1857 138
rect 1791 -150 1857 -138
rect 1887 138 1953 150
rect 1887 -138 1903 138
rect 1937 -138 1953 138
rect 1887 -150 1953 -138
rect 1983 138 2049 150
rect 1983 -138 1999 138
rect 2033 -138 2049 138
rect 1983 -150 2049 -138
rect 2079 138 2145 150
rect 2079 -138 2095 138
rect 2129 -138 2145 138
rect 2079 -150 2145 -138
rect 2175 138 2241 150
rect 2175 -138 2191 138
rect 2225 -138 2241 138
rect 2175 -150 2241 -138
rect 2271 138 2337 150
rect 2271 -138 2287 138
rect 2321 -138 2337 138
rect 2271 -150 2337 -138
rect 2367 138 2433 150
rect 2367 -138 2383 138
rect 2417 -138 2433 138
rect 2367 -150 2433 -138
rect 2463 138 2529 150
rect 2463 -138 2479 138
rect 2513 -138 2529 138
rect 2463 -150 2529 -138
rect 2559 138 2625 150
rect 2559 -138 2575 138
rect 2609 -138 2625 138
rect 2559 -150 2625 -138
rect 2655 138 2721 150
rect 2655 -138 2671 138
rect 2705 -138 2721 138
rect 2655 -150 2721 -138
rect 2751 138 2817 150
rect 2751 -138 2767 138
rect 2801 -138 2817 138
rect 2751 -150 2817 -138
rect 2847 138 2913 150
rect 2847 -138 2863 138
rect 2897 -138 2913 138
rect 2847 -150 2913 -138
rect 2943 138 3009 150
rect 2943 -138 2959 138
rect 2993 -138 3009 138
rect 2943 -150 3009 -138
rect 3039 138 3105 150
rect 3039 -138 3055 138
rect 3089 -138 3105 138
rect 3039 -150 3105 -138
rect 3135 138 3201 150
rect 3135 -138 3151 138
rect 3185 -138 3201 138
rect 3135 -150 3201 -138
rect 3231 138 3297 150
rect 3231 -138 3247 138
rect 3281 -138 3297 138
rect 3231 -150 3297 -138
rect 3327 138 3393 150
rect 3327 -138 3343 138
rect 3377 -138 3393 138
rect 3327 -150 3393 -138
rect 3423 138 3489 150
rect 3423 -138 3439 138
rect 3473 -138 3489 138
rect 3423 -150 3489 -138
rect 3519 138 3585 150
rect 3519 -138 3535 138
rect 3569 -138 3585 138
rect 3519 -150 3585 -138
rect 3615 138 3681 150
rect 3615 -138 3631 138
rect 3665 -138 3681 138
rect 3615 -150 3681 -138
rect 3711 138 3777 150
rect 3711 -138 3727 138
rect 3761 -138 3777 138
rect 3711 -150 3777 -138
rect 3807 138 3873 150
rect 3807 -138 3823 138
rect 3857 -138 3873 138
rect 3807 -150 3873 -138
rect 3903 138 3969 150
rect 3903 -138 3919 138
rect 3953 -138 3969 138
rect 3903 -150 3969 -138
rect 3999 138 4065 150
rect 3999 -138 4015 138
rect 4049 -138 4065 138
rect 3999 -150 4065 -138
rect 4095 138 4161 150
rect 4095 -138 4111 138
rect 4145 -138 4161 138
rect 4095 -150 4161 -138
rect 4191 138 4257 150
rect 4191 -138 4207 138
rect 4241 -138 4257 138
rect 4191 -150 4257 -138
rect 4287 138 4353 150
rect 4287 -138 4303 138
rect 4337 -138 4353 138
rect 4287 -150 4353 -138
rect 4383 138 4449 150
rect 4383 -138 4399 138
rect 4433 -138 4449 138
rect 4383 -150 4449 -138
rect 4479 138 4545 150
rect 4479 -138 4495 138
rect 4529 -138 4545 138
rect 4479 -150 4545 -138
rect 4575 138 4641 150
rect 4575 -138 4591 138
rect 4625 -138 4641 138
rect 4575 -150 4641 -138
rect 4671 138 4737 150
rect 4671 -138 4687 138
rect 4721 -138 4737 138
rect 4671 -150 4737 -138
rect 4767 138 4829 150
rect 4767 -138 4783 138
rect 4817 -138 4829 138
rect 4767 -150 4829 -138
<< ndiffc >>
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
<< psubdiff >>
rect -4931 290 -4835 324
rect 4835 290 4931 324
rect -4931 228 -4897 290
rect 4897 228 4931 290
rect -4931 -290 -4897 -228
rect 4897 -290 4931 -228
rect -4931 -324 -4835 -290
rect 4835 -324 4931 -290
<< psubdiffcont >>
rect -4835 290 4835 324
rect -4931 -228 -4897 228
rect 4897 -228 4931 228
rect -4835 -324 4835 -290
<< poly >>
rect -4689 222 -4623 238
rect -4689 188 -4673 222
rect -4639 188 -4623 222
rect -4767 150 -4737 176
rect -4689 172 -4623 188
rect -4497 222 -4431 238
rect -4497 188 -4481 222
rect -4447 188 -4431 222
rect -4671 150 -4641 172
rect -4575 150 -4545 176
rect -4497 172 -4431 188
rect -4305 222 -4239 238
rect -4305 188 -4289 222
rect -4255 188 -4239 222
rect -4479 150 -4449 172
rect -4383 150 -4353 176
rect -4305 172 -4239 188
rect -4113 222 -4047 238
rect -4113 188 -4097 222
rect -4063 188 -4047 222
rect -4287 150 -4257 172
rect -4191 150 -4161 176
rect -4113 172 -4047 188
rect -3921 222 -3855 238
rect -3921 188 -3905 222
rect -3871 188 -3855 222
rect -4095 150 -4065 172
rect -3999 150 -3969 176
rect -3921 172 -3855 188
rect -3729 222 -3663 238
rect -3729 188 -3713 222
rect -3679 188 -3663 222
rect -3903 150 -3873 172
rect -3807 150 -3777 176
rect -3729 172 -3663 188
rect -3537 222 -3471 238
rect -3537 188 -3521 222
rect -3487 188 -3471 222
rect -3711 150 -3681 172
rect -3615 150 -3585 176
rect -3537 172 -3471 188
rect -3345 222 -3279 238
rect -3345 188 -3329 222
rect -3295 188 -3279 222
rect -3519 150 -3489 172
rect -3423 150 -3393 176
rect -3345 172 -3279 188
rect -3153 222 -3087 238
rect -3153 188 -3137 222
rect -3103 188 -3087 222
rect -3327 150 -3297 172
rect -3231 150 -3201 176
rect -3153 172 -3087 188
rect -2961 222 -2895 238
rect -2961 188 -2945 222
rect -2911 188 -2895 222
rect -3135 150 -3105 172
rect -3039 150 -3009 176
rect -2961 172 -2895 188
rect -2769 222 -2703 238
rect -2769 188 -2753 222
rect -2719 188 -2703 222
rect -2943 150 -2913 172
rect -2847 150 -2817 176
rect -2769 172 -2703 188
rect -2577 222 -2511 238
rect -2577 188 -2561 222
rect -2527 188 -2511 222
rect -2751 150 -2721 172
rect -2655 150 -2625 176
rect -2577 172 -2511 188
rect -2385 222 -2319 238
rect -2385 188 -2369 222
rect -2335 188 -2319 222
rect -2559 150 -2529 172
rect -2463 150 -2433 176
rect -2385 172 -2319 188
rect -2193 222 -2127 238
rect -2193 188 -2177 222
rect -2143 188 -2127 222
rect -2367 150 -2337 172
rect -2271 150 -2241 176
rect -2193 172 -2127 188
rect -2001 222 -1935 238
rect -2001 188 -1985 222
rect -1951 188 -1935 222
rect -2175 150 -2145 172
rect -2079 150 -2049 176
rect -2001 172 -1935 188
rect -1809 222 -1743 238
rect -1809 188 -1793 222
rect -1759 188 -1743 222
rect -1983 150 -1953 172
rect -1887 150 -1857 176
rect -1809 172 -1743 188
rect -1617 222 -1551 238
rect -1617 188 -1601 222
rect -1567 188 -1551 222
rect -1791 150 -1761 172
rect -1695 150 -1665 176
rect -1617 172 -1551 188
rect -1425 222 -1359 238
rect -1425 188 -1409 222
rect -1375 188 -1359 222
rect -1599 150 -1569 172
rect -1503 150 -1473 176
rect -1425 172 -1359 188
rect -1233 222 -1167 238
rect -1233 188 -1217 222
rect -1183 188 -1167 222
rect -1407 150 -1377 172
rect -1311 150 -1281 176
rect -1233 172 -1167 188
rect -1041 222 -975 238
rect -1041 188 -1025 222
rect -991 188 -975 222
rect -1215 150 -1185 172
rect -1119 150 -1089 176
rect -1041 172 -975 188
rect -849 222 -783 238
rect -849 188 -833 222
rect -799 188 -783 222
rect -1023 150 -993 172
rect -927 150 -897 176
rect -849 172 -783 188
rect -657 222 -591 238
rect -657 188 -641 222
rect -607 188 -591 222
rect -831 150 -801 172
rect -735 150 -705 176
rect -657 172 -591 188
rect -465 222 -399 238
rect -465 188 -449 222
rect -415 188 -399 222
rect -639 150 -609 172
rect -543 150 -513 176
rect -465 172 -399 188
rect -273 222 -207 238
rect -273 188 -257 222
rect -223 188 -207 222
rect -447 150 -417 172
rect -351 150 -321 176
rect -273 172 -207 188
rect -81 222 -15 238
rect -81 188 -65 222
rect -31 188 -15 222
rect -255 150 -225 172
rect -159 150 -129 176
rect -81 172 -15 188
rect 111 222 177 238
rect 111 188 127 222
rect 161 188 177 222
rect -63 150 -33 172
rect 33 150 63 176
rect 111 172 177 188
rect 303 222 369 238
rect 303 188 319 222
rect 353 188 369 222
rect 129 150 159 172
rect 225 150 255 176
rect 303 172 369 188
rect 495 222 561 238
rect 495 188 511 222
rect 545 188 561 222
rect 321 150 351 172
rect 417 150 447 176
rect 495 172 561 188
rect 687 222 753 238
rect 687 188 703 222
rect 737 188 753 222
rect 513 150 543 172
rect 609 150 639 176
rect 687 172 753 188
rect 879 222 945 238
rect 879 188 895 222
rect 929 188 945 222
rect 705 150 735 172
rect 801 150 831 176
rect 879 172 945 188
rect 1071 222 1137 238
rect 1071 188 1087 222
rect 1121 188 1137 222
rect 897 150 927 172
rect 993 150 1023 176
rect 1071 172 1137 188
rect 1263 222 1329 238
rect 1263 188 1279 222
rect 1313 188 1329 222
rect 1089 150 1119 172
rect 1185 150 1215 176
rect 1263 172 1329 188
rect 1455 222 1521 238
rect 1455 188 1471 222
rect 1505 188 1521 222
rect 1281 150 1311 172
rect 1377 150 1407 176
rect 1455 172 1521 188
rect 1647 222 1713 238
rect 1647 188 1663 222
rect 1697 188 1713 222
rect 1473 150 1503 172
rect 1569 150 1599 176
rect 1647 172 1713 188
rect 1839 222 1905 238
rect 1839 188 1855 222
rect 1889 188 1905 222
rect 1665 150 1695 172
rect 1761 150 1791 176
rect 1839 172 1905 188
rect 2031 222 2097 238
rect 2031 188 2047 222
rect 2081 188 2097 222
rect 1857 150 1887 172
rect 1953 150 1983 176
rect 2031 172 2097 188
rect 2223 222 2289 238
rect 2223 188 2239 222
rect 2273 188 2289 222
rect 2049 150 2079 172
rect 2145 150 2175 176
rect 2223 172 2289 188
rect 2415 222 2481 238
rect 2415 188 2431 222
rect 2465 188 2481 222
rect 2241 150 2271 172
rect 2337 150 2367 176
rect 2415 172 2481 188
rect 2607 222 2673 238
rect 2607 188 2623 222
rect 2657 188 2673 222
rect 2433 150 2463 172
rect 2529 150 2559 176
rect 2607 172 2673 188
rect 2799 222 2865 238
rect 2799 188 2815 222
rect 2849 188 2865 222
rect 2625 150 2655 172
rect 2721 150 2751 176
rect 2799 172 2865 188
rect 2991 222 3057 238
rect 2991 188 3007 222
rect 3041 188 3057 222
rect 2817 150 2847 172
rect 2913 150 2943 176
rect 2991 172 3057 188
rect 3183 222 3249 238
rect 3183 188 3199 222
rect 3233 188 3249 222
rect 3009 150 3039 172
rect 3105 150 3135 176
rect 3183 172 3249 188
rect 3375 222 3441 238
rect 3375 188 3391 222
rect 3425 188 3441 222
rect 3201 150 3231 172
rect 3297 150 3327 176
rect 3375 172 3441 188
rect 3567 222 3633 238
rect 3567 188 3583 222
rect 3617 188 3633 222
rect 3393 150 3423 172
rect 3489 150 3519 176
rect 3567 172 3633 188
rect 3759 222 3825 238
rect 3759 188 3775 222
rect 3809 188 3825 222
rect 3585 150 3615 172
rect 3681 150 3711 176
rect 3759 172 3825 188
rect 3951 222 4017 238
rect 3951 188 3967 222
rect 4001 188 4017 222
rect 3777 150 3807 172
rect 3873 150 3903 176
rect 3951 172 4017 188
rect 4143 222 4209 238
rect 4143 188 4159 222
rect 4193 188 4209 222
rect 3969 150 3999 172
rect 4065 150 4095 176
rect 4143 172 4209 188
rect 4335 222 4401 238
rect 4335 188 4351 222
rect 4385 188 4401 222
rect 4161 150 4191 172
rect 4257 150 4287 176
rect 4335 172 4401 188
rect 4527 222 4593 238
rect 4527 188 4543 222
rect 4577 188 4593 222
rect 4353 150 4383 172
rect 4449 150 4479 176
rect 4527 172 4593 188
rect 4719 222 4785 238
rect 4719 188 4735 222
rect 4769 188 4785 222
rect 4545 150 4575 172
rect 4641 150 4671 176
rect 4719 172 4785 188
rect 4737 150 4767 172
rect -4767 -172 -4737 -150
rect -4785 -188 -4719 -172
rect -4671 -176 -4641 -150
rect -4575 -172 -4545 -150
rect -4785 -222 -4769 -188
rect -4735 -222 -4719 -188
rect -4785 -238 -4719 -222
rect -4593 -188 -4527 -172
rect -4479 -176 -4449 -150
rect -4383 -172 -4353 -150
rect -4593 -222 -4577 -188
rect -4543 -222 -4527 -188
rect -4593 -238 -4527 -222
rect -4401 -188 -4335 -172
rect -4287 -176 -4257 -150
rect -4191 -172 -4161 -150
rect -4401 -222 -4385 -188
rect -4351 -222 -4335 -188
rect -4401 -238 -4335 -222
rect -4209 -188 -4143 -172
rect -4095 -176 -4065 -150
rect -3999 -172 -3969 -150
rect -4209 -222 -4193 -188
rect -4159 -222 -4143 -188
rect -4209 -238 -4143 -222
rect -4017 -188 -3951 -172
rect -3903 -176 -3873 -150
rect -3807 -172 -3777 -150
rect -4017 -222 -4001 -188
rect -3967 -222 -3951 -188
rect -4017 -238 -3951 -222
rect -3825 -188 -3759 -172
rect -3711 -176 -3681 -150
rect -3615 -172 -3585 -150
rect -3825 -222 -3809 -188
rect -3775 -222 -3759 -188
rect -3825 -238 -3759 -222
rect -3633 -188 -3567 -172
rect -3519 -176 -3489 -150
rect -3423 -172 -3393 -150
rect -3633 -222 -3617 -188
rect -3583 -222 -3567 -188
rect -3633 -238 -3567 -222
rect -3441 -188 -3375 -172
rect -3327 -176 -3297 -150
rect -3231 -172 -3201 -150
rect -3441 -222 -3425 -188
rect -3391 -222 -3375 -188
rect -3441 -238 -3375 -222
rect -3249 -188 -3183 -172
rect -3135 -176 -3105 -150
rect -3039 -172 -3009 -150
rect -3249 -222 -3233 -188
rect -3199 -222 -3183 -188
rect -3249 -238 -3183 -222
rect -3057 -188 -2991 -172
rect -2943 -176 -2913 -150
rect -2847 -172 -2817 -150
rect -3057 -222 -3041 -188
rect -3007 -222 -2991 -188
rect -3057 -238 -2991 -222
rect -2865 -188 -2799 -172
rect -2751 -176 -2721 -150
rect -2655 -172 -2625 -150
rect -2865 -222 -2849 -188
rect -2815 -222 -2799 -188
rect -2865 -238 -2799 -222
rect -2673 -188 -2607 -172
rect -2559 -176 -2529 -150
rect -2463 -172 -2433 -150
rect -2673 -222 -2657 -188
rect -2623 -222 -2607 -188
rect -2673 -238 -2607 -222
rect -2481 -188 -2415 -172
rect -2367 -176 -2337 -150
rect -2271 -172 -2241 -150
rect -2481 -222 -2465 -188
rect -2431 -222 -2415 -188
rect -2481 -238 -2415 -222
rect -2289 -188 -2223 -172
rect -2175 -176 -2145 -150
rect -2079 -172 -2049 -150
rect -2289 -222 -2273 -188
rect -2239 -222 -2223 -188
rect -2289 -238 -2223 -222
rect -2097 -188 -2031 -172
rect -1983 -176 -1953 -150
rect -1887 -172 -1857 -150
rect -2097 -222 -2081 -188
rect -2047 -222 -2031 -188
rect -2097 -238 -2031 -222
rect -1905 -188 -1839 -172
rect -1791 -176 -1761 -150
rect -1695 -172 -1665 -150
rect -1905 -222 -1889 -188
rect -1855 -222 -1839 -188
rect -1905 -238 -1839 -222
rect -1713 -188 -1647 -172
rect -1599 -176 -1569 -150
rect -1503 -172 -1473 -150
rect -1713 -222 -1697 -188
rect -1663 -222 -1647 -188
rect -1713 -238 -1647 -222
rect -1521 -188 -1455 -172
rect -1407 -176 -1377 -150
rect -1311 -172 -1281 -150
rect -1521 -222 -1505 -188
rect -1471 -222 -1455 -188
rect -1521 -238 -1455 -222
rect -1329 -188 -1263 -172
rect -1215 -176 -1185 -150
rect -1119 -172 -1089 -150
rect -1329 -222 -1313 -188
rect -1279 -222 -1263 -188
rect -1329 -238 -1263 -222
rect -1137 -188 -1071 -172
rect -1023 -176 -993 -150
rect -927 -172 -897 -150
rect -1137 -222 -1121 -188
rect -1087 -222 -1071 -188
rect -1137 -238 -1071 -222
rect -945 -188 -879 -172
rect -831 -176 -801 -150
rect -735 -172 -705 -150
rect -945 -222 -929 -188
rect -895 -222 -879 -188
rect -945 -238 -879 -222
rect -753 -188 -687 -172
rect -639 -176 -609 -150
rect -543 -172 -513 -150
rect -753 -222 -737 -188
rect -703 -222 -687 -188
rect -753 -238 -687 -222
rect -561 -188 -495 -172
rect -447 -176 -417 -150
rect -351 -172 -321 -150
rect -561 -222 -545 -188
rect -511 -222 -495 -188
rect -561 -238 -495 -222
rect -369 -188 -303 -172
rect -255 -176 -225 -150
rect -159 -172 -129 -150
rect -369 -222 -353 -188
rect -319 -222 -303 -188
rect -369 -238 -303 -222
rect -177 -188 -111 -172
rect -63 -176 -33 -150
rect 33 -172 63 -150
rect -177 -222 -161 -188
rect -127 -222 -111 -188
rect -177 -238 -111 -222
rect 15 -188 81 -172
rect 129 -176 159 -150
rect 225 -172 255 -150
rect 15 -222 31 -188
rect 65 -222 81 -188
rect 15 -238 81 -222
rect 207 -188 273 -172
rect 321 -176 351 -150
rect 417 -172 447 -150
rect 207 -222 223 -188
rect 257 -222 273 -188
rect 207 -238 273 -222
rect 399 -188 465 -172
rect 513 -176 543 -150
rect 609 -172 639 -150
rect 399 -222 415 -188
rect 449 -222 465 -188
rect 399 -238 465 -222
rect 591 -188 657 -172
rect 705 -176 735 -150
rect 801 -172 831 -150
rect 591 -222 607 -188
rect 641 -222 657 -188
rect 591 -238 657 -222
rect 783 -188 849 -172
rect 897 -176 927 -150
rect 993 -172 1023 -150
rect 783 -222 799 -188
rect 833 -222 849 -188
rect 783 -238 849 -222
rect 975 -188 1041 -172
rect 1089 -176 1119 -150
rect 1185 -172 1215 -150
rect 975 -222 991 -188
rect 1025 -222 1041 -188
rect 975 -238 1041 -222
rect 1167 -188 1233 -172
rect 1281 -176 1311 -150
rect 1377 -172 1407 -150
rect 1167 -222 1183 -188
rect 1217 -222 1233 -188
rect 1167 -238 1233 -222
rect 1359 -188 1425 -172
rect 1473 -176 1503 -150
rect 1569 -172 1599 -150
rect 1359 -222 1375 -188
rect 1409 -222 1425 -188
rect 1359 -238 1425 -222
rect 1551 -188 1617 -172
rect 1665 -176 1695 -150
rect 1761 -172 1791 -150
rect 1551 -222 1567 -188
rect 1601 -222 1617 -188
rect 1551 -238 1617 -222
rect 1743 -188 1809 -172
rect 1857 -176 1887 -150
rect 1953 -172 1983 -150
rect 1743 -222 1759 -188
rect 1793 -222 1809 -188
rect 1743 -238 1809 -222
rect 1935 -188 2001 -172
rect 2049 -176 2079 -150
rect 2145 -172 2175 -150
rect 1935 -222 1951 -188
rect 1985 -222 2001 -188
rect 1935 -238 2001 -222
rect 2127 -188 2193 -172
rect 2241 -176 2271 -150
rect 2337 -172 2367 -150
rect 2127 -222 2143 -188
rect 2177 -222 2193 -188
rect 2127 -238 2193 -222
rect 2319 -188 2385 -172
rect 2433 -176 2463 -150
rect 2529 -172 2559 -150
rect 2319 -222 2335 -188
rect 2369 -222 2385 -188
rect 2319 -238 2385 -222
rect 2511 -188 2577 -172
rect 2625 -176 2655 -150
rect 2721 -172 2751 -150
rect 2511 -222 2527 -188
rect 2561 -222 2577 -188
rect 2511 -238 2577 -222
rect 2703 -188 2769 -172
rect 2817 -176 2847 -150
rect 2913 -172 2943 -150
rect 2703 -222 2719 -188
rect 2753 -222 2769 -188
rect 2703 -238 2769 -222
rect 2895 -188 2961 -172
rect 3009 -176 3039 -150
rect 3105 -172 3135 -150
rect 2895 -222 2911 -188
rect 2945 -222 2961 -188
rect 2895 -238 2961 -222
rect 3087 -188 3153 -172
rect 3201 -176 3231 -150
rect 3297 -172 3327 -150
rect 3087 -222 3103 -188
rect 3137 -222 3153 -188
rect 3087 -238 3153 -222
rect 3279 -188 3345 -172
rect 3393 -176 3423 -150
rect 3489 -172 3519 -150
rect 3279 -222 3295 -188
rect 3329 -222 3345 -188
rect 3279 -238 3345 -222
rect 3471 -188 3537 -172
rect 3585 -176 3615 -150
rect 3681 -172 3711 -150
rect 3471 -222 3487 -188
rect 3521 -222 3537 -188
rect 3471 -238 3537 -222
rect 3663 -188 3729 -172
rect 3777 -176 3807 -150
rect 3873 -172 3903 -150
rect 3663 -222 3679 -188
rect 3713 -222 3729 -188
rect 3663 -238 3729 -222
rect 3855 -188 3921 -172
rect 3969 -176 3999 -150
rect 4065 -172 4095 -150
rect 3855 -222 3871 -188
rect 3905 -222 3921 -188
rect 3855 -238 3921 -222
rect 4047 -188 4113 -172
rect 4161 -176 4191 -150
rect 4257 -172 4287 -150
rect 4047 -222 4063 -188
rect 4097 -222 4113 -188
rect 4047 -238 4113 -222
rect 4239 -188 4305 -172
rect 4353 -176 4383 -150
rect 4449 -172 4479 -150
rect 4239 -222 4255 -188
rect 4289 -222 4305 -188
rect 4239 -238 4305 -222
rect 4431 -188 4497 -172
rect 4545 -176 4575 -150
rect 4641 -172 4671 -150
rect 4431 -222 4447 -188
rect 4481 -222 4497 -188
rect 4431 -238 4497 -222
rect 4623 -188 4689 -172
rect 4737 -176 4767 -150
rect 4623 -222 4639 -188
rect 4673 -222 4689 -188
rect 4623 -238 4689 -222
<< polycont >>
rect -4673 188 -4639 222
rect -4481 188 -4447 222
rect -4289 188 -4255 222
rect -4097 188 -4063 222
rect -3905 188 -3871 222
rect -3713 188 -3679 222
rect -3521 188 -3487 222
rect -3329 188 -3295 222
rect -3137 188 -3103 222
rect -2945 188 -2911 222
rect -2753 188 -2719 222
rect -2561 188 -2527 222
rect -2369 188 -2335 222
rect -2177 188 -2143 222
rect -1985 188 -1951 222
rect -1793 188 -1759 222
rect -1601 188 -1567 222
rect -1409 188 -1375 222
rect -1217 188 -1183 222
rect -1025 188 -991 222
rect -833 188 -799 222
rect -641 188 -607 222
rect -449 188 -415 222
rect -257 188 -223 222
rect -65 188 -31 222
rect 127 188 161 222
rect 319 188 353 222
rect 511 188 545 222
rect 703 188 737 222
rect 895 188 929 222
rect 1087 188 1121 222
rect 1279 188 1313 222
rect 1471 188 1505 222
rect 1663 188 1697 222
rect 1855 188 1889 222
rect 2047 188 2081 222
rect 2239 188 2273 222
rect 2431 188 2465 222
rect 2623 188 2657 222
rect 2815 188 2849 222
rect 3007 188 3041 222
rect 3199 188 3233 222
rect 3391 188 3425 222
rect 3583 188 3617 222
rect 3775 188 3809 222
rect 3967 188 4001 222
rect 4159 188 4193 222
rect 4351 188 4385 222
rect 4543 188 4577 222
rect 4735 188 4769 222
rect -4769 -222 -4735 -188
rect -4577 -222 -4543 -188
rect -4385 -222 -4351 -188
rect -4193 -222 -4159 -188
rect -4001 -222 -3967 -188
rect -3809 -222 -3775 -188
rect -3617 -222 -3583 -188
rect -3425 -222 -3391 -188
rect -3233 -222 -3199 -188
rect -3041 -222 -3007 -188
rect -2849 -222 -2815 -188
rect -2657 -222 -2623 -188
rect -2465 -222 -2431 -188
rect -2273 -222 -2239 -188
rect -2081 -222 -2047 -188
rect -1889 -222 -1855 -188
rect -1697 -222 -1663 -188
rect -1505 -222 -1471 -188
rect -1313 -222 -1279 -188
rect -1121 -222 -1087 -188
rect -929 -222 -895 -188
rect -737 -222 -703 -188
rect -545 -222 -511 -188
rect -353 -222 -319 -188
rect -161 -222 -127 -188
rect 31 -222 65 -188
rect 223 -222 257 -188
rect 415 -222 449 -188
rect 607 -222 641 -188
rect 799 -222 833 -188
rect 991 -222 1025 -188
rect 1183 -222 1217 -188
rect 1375 -222 1409 -188
rect 1567 -222 1601 -188
rect 1759 -222 1793 -188
rect 1951 -222 1985 -188
rect 2143 -222 2177 -188
rect 2335 -222 2369 -188
rect 2527 -222 2561 -188
rect 2719 -222 2753 -188
rect 2911 -222 2945 -188
rect 3103 -222 3137 -188
rect 3295 -222 3329 -188
rect 3487 -222 3521 -188
rect 3679 -222 3713 -188
rect 3871 -222 3905 -188
rect 4063 -222 4097 -188
rect 4255 -222 4289 -188
rect 4447 -222 4481 -188
rect 4639 -222 4673 -188
<< locali >>
rect -4931 290 -4835 324
rect 4835 290 4931 324
rect -4931 228 -4897 290
rect 4897 228 4931 290
rect -4689 188 -4673 222
rect -4639 188 -4623 222
rect -4497 188 -4481 222
rect -4447 188 -4431 222
rect -4305 188 -4289 222
rect -4255 188 -4239 222
rect -4113 188 -4097 222
rect -4063 188 -4047 222
rect -3921 188 -3905 222
rect -3871 188 -3855 222
rect -3729 188 -3713 222
rect -3679 188 -3663 222
rect -3537 188 -3521 222
rect -3487 188 -3471 222
rect -3345 188 -3329 222
rect -3295 188 -3279 222
rect -3153 188 -3137 222
rect -3103 188 -3087 222
rect -2961 188 -2945 222
rect -2911 188 -2895 222
rect -2769 188 -2753 222
rect -2719 188 -2703 222
rect -2577 188 -2561 222
rect -2527 188 -2511 222
rect -2385 188 -2369 222
rect -2335 188 -2319 222
rect -2193 188 -2177 222
rect -2143 188 -2127 222
rect -2001 188 -1985 222
rect -1951 188 -1935 222
rect -1809 188 -1793 222
rect -1759 188 -1743 222
rect -1617 188 -1601 222
rect -1567 188 -1551 222
rect -1425 188 -1409 222
rect -1375 188 -1359 222
rect -1233 188 -1217 222
rect -1183 188 -1167 222
rect -1041 188 -1025 222
rect -991 188 -975 222
rect -849 188 -833 222
rect -799 188 -783 222
rect -657 188 -641 222
rect -607 188 -591 222
rect -465 188 -449 222
rect -415 188 -399 222
rect -273 188 -257 222
rect -223 188 -207 222
rect -81 188 -65 222
rect -31 188 -15 222
rect 111 188 127 222
rect 161 188 177 222
rect 303 188 319 222
rect 353 188 369 222
rect 495 188 511 222
rect 545 188 561 222
rect 687 188 703 222
rect 737 188 753 222
rect 879 188 895 222
rect 929 188 945 222
rect 1071 188 1087 222
rect 1121 188 1137 222
rect 1263 188 1279 222
rect 1313 188 1329 222
rect 1455 188 1471 222
rect 1505 188 1521 222
rect 1647 188 1663 222
rect 1697 188 1713 222
rect 1839 188 1855 222
rect 1889 188 1905 222
rect 2031 188 2047 222
rect 2081 188 2097 222
rect 2223 188 2239 222
rect 2273 188 2289 222
rect 2415 188 2431 222
rect 2465 188 2481 222
rect 2607 188 2623 222
rect 2657 188 2673 222
rect 2799 188 2815 222
rect 2849 188 2865 222
rect 2991 188 3007 222
rect 3041 188 3057 222
rect 3183 188 3199 222
rect 3233 188 3249 222
rect 3375 188 3391 222
rect 3425 188 3441 222
rect 3567 188 3583 222
rect 3617 188 3633 222
rect 3759 188 3775 222
rect 3809 188 3825 222
rect 3951 188 3967 222
rect 4001 188 4017 222
rect 4143 188 4159 222
rect 4193 188 4209 222
rect 4335 188 4351 222
rect 4385 188 4401 222
rect 4527 188 4543 222
rect 4577 188 4593 222
rect 4719 188 4735 222
rect 4769 188 4785 222
rect -4817 138 -4783 154
rect -4817 -154 -4783 -138
rect -4721 138 -4687 154
rect -4721 -154 -4687 -138
rect -4625 138 -4591 154
rect -4625 -154 -4591 -138
rect -4529 138 -4495 154
rect -4529 -154 -4495 -138
rect -4433 138 -4399 154
rect -4433 -154 -4399 -138
rect -4337 138 -4303 154
rect -4337 -154 -4303 -138
rect -4241 138 -4207 154
rect -4241 -154 -4207 -138
rect -4145 138 -4111 154
rect -4145 -154 -4111 -138
rect -4049 138 -4015 154
rect -4049 -154 -4015 -138
rect -3953 138 -3919 154
rect -3953 -154 -3919 -138
rect -3857 138 -3823 154
rect -3857 -154 -3823 -138
rect -3761 138 -3727 154
rect -3761 -154 -3727 -138
rect -3665 138 -3631 154
rect -3665 -154 -3631 -138
rect -3569 138 -3535 154
rect -3569 -154 -3535 -138
rect -3473 138 -3439 154
rect -3473 -154 -3439 -138
rect -3377 138 -3343 154
rect -3377 -154 -3343 -138
rect -3281 138 -3247 154
rect -3281 -154 -3247 -138
rect -3185 138 -3151 154
rect -3185 -154 -3151 -138
rect -3089 138 -3055 154
rect -3089 -154 -3055 -138
rect -2993 138 -2959 154
rect -2993 -154 -2959 -138
rect -2897 138 -2863 154
rect -2897 -154 -2863 -138
rect -2801 138 -2767 154
rect -2801 -154 -2767 -138
rect -2705 138 -2671 154
rect -2705 -154 -2671 -138
rect -2609 138 -2575 154
rect -2609 -154 -2575 -138
rect -2513 138 -2479 154
rect -2513 -154 -2479 -138
rect -2417 138 -2383 154
rect -2417 -154 -2383 -138
rect -2321 138 -2287 154
rect -2321 -154 -2287 -138
rect -2225 138 -2191 154
rect -2225 -154 -2191 -138
rect -2129 138 -2095 154
rect -2129 -154 -2095 -138
rect -2033 138 -1999 154
rect -2033 -154 -1999 -138
rect -1937 138 -1903 154
rect -1937 -154 -1903 -138
rect -1841 138 -1807 154
rect -1841 -154 -1807 -138
rect -1745 138 -1711 154
rect -1745 -154 -1711 -138
rect -1649 138 -1615 154
rect -1649 -154 -1615 -138
rect -1553 138 -1519 154
rect -1553 -154 -1519 -138
rect -1457 138 -1423 154
rect -1457 -154 -1423 -138
rect -1361 138 -1327 154
rect -1361 -154 -1327 -138
rect -1265 138 -1231 154
rect -1265 -154 -1231 -138
rect -1169 138 -1135 154
rect -1169 -154 -1135 -138
rect -1073 138 -1039 154
rect -1073 -154 -1039 -138
rect -977 138 -943 154
rect -977 -154 -943 -138
rect -881 138 -847 154
rect -881 -154 -847 -138
rect -785 138 -751 154
rect -785 -154 -751 -138
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect 751 138 785 154
rect 751 -154 785 -138
rect 847 138 881 154
rect 847 -154 881 -138
rect 943 138 977 154
rect 943 -154 977 -138
rect 1039 138 1073 154
rect 1039 -154 1073 -138
rect 1135 138 1169 154
rect 1135 -154 1169 -138
rect 1231 138 1265 154
rect 1231 -154 1265 -138
rect 1327 138 1361 154
rect 1327 -154 1361 -138
rect 1423 138 1457 154
rect 1423 -154 1457 -138
rect 1519 138 1553 154
rect 1519 -154 1553 -138
rect 1615 138 1649 154
rect 1615 -154 1649 -138
rect 1711 138 1745 154
rect 1711 -154 1745 -138
rect 1807 138 1841 154
rect 1807 -154 1841 -138
rect 1903 138 1937 154
rect 1903 -154 1937 -138
rect 1999 138 2033 154
rect 1999 -154 2033 -138
rect 2095 138 2129 154
rect 2095 -154 2129 -138
rect 2191 138 2225 154
rect 2191 -154 2225 -138
rect 2287 138 2321 154
rect 2287 -154 2321 -138
rect 2383 138 2417 154
rect 2383 -154 2417 -138
rect 2479 138 2513 154
rect 2479 -154 2513 -138
rect 2575 138 2609 154
rect 2575 -154 2609 -138
rect 2671 138 2705 154
rect 2671 -154 2705 -138
rect 2767 138 2801 154
rect 2767 -154 2801 -138
rect 2863 138 2897 154
rect 2863 -154 2897 -138
rect 2959 138 2993 154
rect 2959 -154 2993 -138
rect 3055 138 3089 154
rect 3055 -154 3089 -138
rect 3151 138 3185 154
rect 3151 -154 3185 -138
rect 3247 138 3281 154
rect 3247 -154 3281 -138
rect 3343 138 3377 154
rect 3343 -154 3377 -138
rect 3439 138 3473 154
rect 3439 -154 3473 -138
rect 3535 138 3569 154
rect 3535 -154 3569 -138
rect 3631 138 3665 154
rect 3631 -154 3665 -138
rect 3727 138 3761 154
rect 3727 -154 3761 -138
rect 3823 138 3857 154
rect 3823 -154 3857 -138
rect 3919 138 3953 154
rect 3919 -154 3953 -138
rect 4015 138 4049 154
rect 4015 -154 4049 -138
rect 4111 138 4145 154
rect 4111 -154 4145 -138
rect 4207 138 4241 154
rect 4207 -154 4241 -138
rect 4303 138 4337 154
rect 4303 -154 4337 -138
rect 4399 138 4433 154
rect 4399 -154 4433 -138
rect 4495 138 4529 154
rect 4495 -154 4529 -138
rect 4591 138 4625 154
rect 4591 -154 4625 -138
rect 4687 138 4721 154
rect 4687 -154 4721 -138
rect 4783 138 4817 154
rect 4783 -154 4817 -138
rect -4785 -222 -4769 -188
rect -4735 -222 -4719 -188
rect -4593 -222 -4577 -188
rect -4543 -222 -4527 -188
rect -4401 -222 -4385 -188
rect -4351 -222 -4335 -188
rect -4209 -222 -4193 -188
rect -4159 -222 -4143 -188
rect -4017 -222 -4001 -188
rect -3967 -222 -3951 -188
rect -3825 -222 -3809 -188
rect -3775 -222 -3759 -188
rect -3633 -222 -3617 -188
rect -3583 -222 -3567 -188
rect -3441 -222 -3425 -188
rect -3391 -222 -3375 -188
rect -3249 -222 -3233 -188
rect -3199 -222 -3183 -188
rect -3057 -222 -3041 -188
rect -3007 -222 -2991 -188
rect -2865 -222 -2849 -188
rect -2815 -222 -2799 -188
rect -2673 -222 -2657 -188
rect -2623 -222 -2607 -188
rect -2481 -222 -2465 -188
rect -2431 -222 -2415 -188
rect -2289 -222 -2273 -188
rect -2239 -222 -2223 -188
rect -2097 -222 -2081 -188
rect -2047 -222 -2031 -188
rect -1905 -222 -1889 -188
rect -1855 -222 -1839 -188
rect -1713 -222 -1697 -188
rect -1663 -222 -1647 -188
rect -1521 -222 -1505 -188
rect -1471 -222 -1455 -188
rect -1329 -222 -1313 -188
rect -1279 -222 -1263 -188
rect -1137 -222 -1121 -188
rect -1087 -222 -1071 -188
rect -945 -222 -929 -188
rect -895 -222 -879 -188
rect -753 -222 -737 -188
rect -703 -222 -687 -188
rect -561 -222 -545 -188
rect -511 -222 -495 -188
rect -369 -222 -353 -188
rect -319 -222 -303 -188
rect -177 -222 -161 -188
rect -127 -222 -111 -188
rect 15 -222 31 -188
rect 65 -222 81 -188
rect 207 -222 223 -188
rect 257 -222 273 -188
rect 399 -222 415 -188
rect 449 -222 465 -188
rect 591 -222 607 -188
rect 641 -222 657 -188
rect 783 -222 799 -188
rect 833 -222 849 -188
rect 975 -222 991 -188
rect 1025 -222 1041 -188
rect 1167 -222 1183 -188
rect 1217 -222 1233 -188
rect 1359 -222 1375 -188
rect 1409 -222 1425 -188
rect 1551 -222 1567 -188
rect 1601 -222 1617 -188
rect 1743 -222 1759 -188
rect 1793 -222 1809 -188
rect 1935 -222 1951 -188
rect 1985 -222 2001 -188
rect 2127 -222 2143 -188
rect 2177 -222 2193 -188
rect 2319 -222 2335 -188
rect 2369 -222 2385 -188
rect 2511 -222 2527 -188
rect 2561 -222 2577 -188
rect 2703 -222 2719 -188
rect 2753 -222 2769 -188
rect 2895 -222 2911 -188
rect 2945 -222 2961 -188
rect 3087 -222 3103 -188
rect 3137 -222 3153 -188
rect 3279 -222 3295 -188
rect 3329 -222 3345 -188
rect 3471 -222 3487 -188
rect 3521 -222 3537 -188
rect 3663 -222 3679 -188
rect 3713 -222 3729 -188
rect 3855 -222 3871 -188
rect 3905 -222 3921 -188
rect 4047 -222 4063 -188
rect 4097 -222 4113 -188
rect 4239 -222 4255 -188
rect 4289 -222 4305 -188
rect 4431 -222 4447 -188
rect 4481 -222 4497 -188
rect 4623 -222 4639 -188
rect 4673 -222 4689 -188
rect -4931 -290 -4897 -228
rect 4897 -290 4931 -228
rect -4931 -324 -4835 -290
rect 4835 -324 4931 -290
<< viali >>
rect -4673 188 -4639 222
rect -4481 188 -4447 222
rect -4289 188 -4255 222
rect -4097 188 -4063 222
rect -3905 188 -3871 222
rect -3713 188 -3679 222
rect -3521 188 -3487 222
rect -3329 188 -3295 222
rect -3137 188 -3103 222
rect -2945 188 -2911 222
rect -2753 188 -2719 222
rect -2561 188 -2527 222
rect -2369 188 -2335 222
rect -2177 188 -2143 222
rect -1985 188 -1951 222
rect -1793 188 -1759 222
rect -1601 188 -1567 222
rect -1409 188 -1375 222
rect -1217 188 -1183 222
rect -1025 188 -991 222
rect -833 188 -799 222
rect -641 188 -607 222
rect -449 188 -415 222
rect -257 188 -223 222
rect -65 188 -31 222
rect 127 188 161 222
rect 319 188 353 222
rect 511 188 545 222
rect 703 188 737 222
rect 895 188 929 222
rect 1087 188 1121 222
rect 1279 188 1313 222
rect 1471 188 1505 222
rect 1663 188 1697 222
rect 1855 188 1889 222
rect 2047 188 2081 222
rect 2239 188 2273 222
rect 2431 188 2465 222
rect 2623 188 2657 222
rect 2815 188 2849 222
rect 3007 188 3041 222
rect 3199 188 3233 222
rect 3391 188 3425 222
rect 3583 188 3617 222
rect 3775 188 3809 222
rect 3967 188 4001 222
rect 4159 188 4193 222
rect 4351 188 4385 222
rect 4543 188 4577 222
rect 4735 188 4769 222
rect -4817 -138 -4783 138
rect -4721 -138 -4687 138
rect -4625 -138 -4591 138
rect -4529 -138 -4495 138
rect -4433 -138 -4399 138
rect -4337 -138 -4303 138
rect -4241 -138 -4207 138
rect -4145 -138 -4111 138
rect -4049 -138 -4015 138
rect -3953 -138 -3919 138
rect -3857 -138 -3823 138
rect -3761 -138 -3727 138
rect -3665 -138 -3631 138
rect -3569 -138 -3535 138
rect -3473 -138 -3439 138
rect -3377 -138 -3343 138
rect -3281 -138 -3247 138
rect -3185 -138 -3151 138
rect -3089 -138 -3055 138
rect -2993 -138 -2959 138
rect -2897 -138 -2863 138
rect -2801 -138 -2767 138
rect -2705 -138 -2671 138
rect -2609 -138 -2575 138
rect -2513 -138 -2479 138
rect -2417 -138 -2383 138
rect -2321 -138 -2287 138
rect -2225 -138 -2191 138
rect -2129 -138 -2095 138
rect -2033 -138 -1999 138
rect -1937 -138 -1903 138
rect -1841 -138 -1807 138
rect -1745 -138 -1711 138
rect -1649 -138 -1615 138
rect -1553 -138 -1519 138
rect -1457 -138 -1423 138
rect -1361 -138 -1327 138
rect -1265 -138 -1231 138
rect -1169 -138 -1135 138
rect -1073 -138 -1039 138
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect 1039 -138 1073 138
rect 1135 -138 1169 138
rect 1231 -138 1265 138
rect 1327 -138 1361 138
rect 1423 -138 1457 138
rect 1519 -138 1553 138
rect 1615 -138 1649 138
rect 1711 -138 1745 138
rect 1807 -138 1841 138
rect 1903 -138 1937 138
rect 1999 -138 2033 138
rect 2095 -138 2129 138
rect 2191 -138 2225 138
rect 2287 -138 2321 138
rect 2383 -138 2417 138
rect 2479 -138 2513 138
rect 2575 -138 2609 138
rect 2671 -138 2705 138
rect 2767 -138 2801 138
rect 2863 -138 2897 138
rect 2959 -138 2993 138
rect 3055 -138 3089 138
rect 3151 -138 3185 138
rect 3247 -138 3281 138
rect 3343 -138 3377 138
rect 3439 -138 3473 138
rect 3535 -138 3569 138
rect 3631 -138 3665 138
rect 3727 -138 3761 138
rect 3823 -138 3857 138
rect 3919 -138 3953 138
rect 4015 -138 4049 138
rect 4111 -138 4145 138
rect 4207 -138 4241 138
rect 4303 -138 4337 138
rect 4399 -138 4433 138
rect 4495 -138 4529 138
rect 4591 -138 4625 138
rect 4687 -138 4721 138
rect 4783 -138 4817 138
rect -4769 -222 -4735 -188
rect -4577 -222 -4543 -188
rect -4385 -222 -4351 -188
rect -4193 -222 -4159 -188
rect -4001 -222 -3967 -188
rect -3809 -222 -3775 -188
rect -3617 -222 -3583 -188
rect -3425 -222 -3391 -188
rect -3233 -222 -3199 -188
rect -3041 -222 -3007 -188
rect -2849 -222 -2815 -188
rect -2657 -222 -2623 -188
rect -2465 -222 -2431 -188
rect -2273 -222 -2239 -188
rect -2081 -222 -2047 -188
rect -1889 -222 -1855 -188
rect -1697 -222 -1663 -188
rect -1505 -222 -1471 -188
rect -1313 -222 -1279 -188
rect -1121 -222 -1087 -188
rect -929 -222 -895 -188
rect -737 -222 -703 -188
rect -545 -222 -511 -188
rect -353 -222 -319 -188
rect -161 -222 -127 -188
rect 31 -222 65 -188
rect 223 -222 257 -188
rect 415 -222 449 -188
rect 607 -222 641 -188
rect 799 -222 833 -188
rect 991 -222 1025 -188
rect 1183 -222 1217 -188
rect 1375 -222 1409 -188
rect 1567 -222 1601 -188
rect 1759 -222 1793 -188
rect 1951 -222 1985 -188
rect 2143 -222 2177 -188
rect 2335 -222 2369 -188
rect 2527 -222 2561 -188
rect 2719 -222 2753 -188
rect 2911 -222 2945 -188
rect 3103 -222 3137 -188
rect 3295 -222 3329 -188
rect 3487 -222 3521 -188
rect 3679 -222 3713 -188
rect 3871 -222 3905 -188
rect 4063 -222 4097 -188
rect 4255 -222 4289 -188
rect 4447 -222 4481 -188
rect 4639 -222 4673 -188
<< metal1 >>
rect -4685 222 -4627 228
rect -4685 188 -4673 222
rect -4639 188 -4627 222
rect -4685 182 -4627 188
rect -4493 222 -4435 228
rect -4493 188 -4481 222
rect -4447 188 -4435 222
rect -4493 182 -4435 188
rect -4301 222 -4243 228
rect -4301 188 -4289 222
rect -4255 188 -4243 222
rect -4301 182 -4243 188
rect -4109 222 -4051 228
rect -4109 188 -4097 222
rect -4063 188 -4051 222
rect -4109 182 -4051 188
rect -3917 222 -3859 228
rect -3917 188 -3905 222
rect -3871 188 -3859 222
rect -3917 182 -3859 188
rect -3725 222 -3667 228
rect -3725 188 -3713 222
rect -3679 188 -3667 222
rect -3725 182 -3667 188
rect -3533 222 -3475 228
rect -3533 188 -3521 222
rect -3487 188 -3475 222
rect -3533 182 -3475 188
rect -3341 222 -3283 228
rect -3341 188 -3329 222
rect -3295 188 -3283 222
rect -3341 182 -3283 188
rect -3149 222 -3091 228
rect -3149 188 -3137 222
rect -3103 188 -3091 222
rect -3149 182 -3091 188
rect -2957 222 -2899 228
rect -2957 188 -2945 222
rect -2911 188 -2899 222
rect -2957 182 -2899 188
rect -2765 222 -2707 228
rect -2765 188 -2753 222
rect -2719 188 -2707 222
rect -2765 182 -2707 188
rect -2573 222 -2515 228
rect -2573 188 -2561 222
rect -2527 188 -2515 222
rect -2573 182 -2515 188
rect -2381 222 -2323 228
rect -2381 188 -2369 222
rect -2335 188 -2323 222
rect -2381 182 -2323 188
rect -2189 222 -2131 228
rect -2189 188 -2177 222
rect -2143 188 -2131 222
rect -2189 182 -2131 188
rect -1997 222 -1939 228
rect -1997 188 -1985 222
rect -1951 188 -1939 222
rect -1997 182 -1939 188
rect -1805 222 -1747 228
rect -1805 188 -1793 222
rect -1759 188 -1747 222
rect -1805 182 -1747 188
rect -1613 222 -1555 228
rect -1613 188 -1601 222
rect -1567 188 -1555 222
rect -1613 182 -1555 188
rect -1421 222 -1363 228
rect -1421 188 -1409 222
rect -1375 188 -1363 222
rect -1421 182 -1363 188
rect -1229 222 -1171 228
rect -1229 188 -1217 222
rect -1183 188 -1171 222
rect -1229 182 -1171 188
rect -1037 222 -979 228
rect -1037 188 -1025 222
rect -991 188 -979 222
rect -1037 182 -979 188
rect -845 222 -787 228
rect -845 188 -833 222
rect -799 188 -787 222
rect -845 182 -787 188
rect -653 222 -595 228
rect -653 188 -641 222
rect -607 188 -595 222
rect -653 182 -595 188
rect -461 222 -403 228
rect -461 188 -449 222
rect -415 188 -403 222
rect -461 182 -403 188
rect -269 222 -211 228
rect -269 188 -257 222
rect -223 188 -211 222
rect -269 182 -211 188
rect -77 222 -19 228
rect -77 188 -65 222
rect -31 188 -19 222
rect -77 182 -19 188
rect 115 222 173 228
rect 115 188 127 222
rect 161 188 173 222
rect 115 182 173 188
rect 307 222 365 228
rect 307 188 319 222
rect 353 188 365 222
rect 307 182 365 188
rect 499 222 557 228
rect 499 188 511 222
rect 545 188 557 222
rect 499 182 557 188
rect 691 222 749 228
rect 691 188 703 222
rect 737 188 749 222
rect 691 182 749 188
rect 883 222 941 228
rect 883 188 895 222
rect 929 188 941 222
rect 883 182 941 188
rect 1075 222 1133 228
rect 1075 188 1087 222
rect 1121 188 1133 222
rect 1075 182 1133 188
rect 1267 222 1325 228
rect 1267 188 1279 222
rect 1313 188 1325 222
rect 1267 182 1325 188
rect 1459 222 1517 228
rect 1459 188 1471 222
rect 1505 188 1517 222
rect 1459 182 1517 188
rect 1651 222 1709 228
rect 1651 188 1663 222
rect 1697 188 1709 222
rect 1651 182 1709 188
rect 1843 222 1901 228
rect 1843 188 1855 222
rect 1889 188 1901 222
rect 1843 182 1901 188
rect 2035 222 2093 228
rect 2035 188 2047 222
rect 2081 188 2093 222
rect 2035 182 2093 188
rect 2227 222 2285 228
rect 2227 188 2239 222
rect 2273 188 2285 222
rect 2227 182 2285 188
rect 2419 222 2477 228
rect 2419 188 2431 222
rect 2465 188 2477 222
rect 2419 182 2477 188
rect 2611 222 2669 228
rect 2611 188 2623 222
rect 2657 188 2669 222
rect 2611 182 2669 188
rect 2803 222 2861 228
rect 2803 188 2815 222
rect 2849 188 2861 222
rect 2803 182 2861 188
rect 2995 222 3053 228
rect 2995 188 3007 222
rect 3041 188 3053 222
rect 2995 182 3053 188
rect 3187 222 3245 228
rect 3187 188 3199 222
rect 3233 188 3245 222
rect 3187 182 3245 188
rect 3379 222 3437 228
rect 3379 188 3391 222
rect 3425 188 3437 222
rect 3379 182 3437 188
rect 3571 222 3629 228
rect 3571 188 3583 222
rect 3617 188 3629 222
rect 3571 182 3629 188
rect 3763 222 3821 228
rect 3763 188 3775 222
rect 3809 188 3821 222
rect 3763 182 3821 188
rect 3955 222 4013 228
rect 3955 188 3967 222
rect 4001 188 4013 222
rect 3955 182 4013 188
rect 4147 222 4205 228
rect 4147 188 4159 222
rect 4193 188 4205 222
rect 4147 182 4205 188
rect 4339 222 4397 228
rect 4339 188 4351 222
rect 4385 188 4397 222
rect 4339 182 4397 188
rect 4531 222 4589 228
rect 4531 188 4543 222
rect 4577 188 4589 222
rect 4531 182 4589 188
rect 4723 222 4781 228
rect 4723 188 4735 222
rect 4769 188 4781 222
rect 4723 182 4781 188
rect -4823 138 -4777 150
rect -4823 -138 -4817 138
rect -4783 -138 -4777 138
rect -4823 -150 -4777 -138
rect -4727 138 -4681 150
rect -4727 -138 -4721 138
rect -4687 -138 -4681 138
rect -4727 -150 -4681 -138
rect -4631 138 -4585 150
rect -4631 -138 -4625 138
rect -4591 -138 -4585 138
rect -4631 -150 -4585 -138
rect -4535 138 -4489 150
rect -4535 -138 -4529 138
rect -4495 -138 -4489 138
rect -4535 -150 -4489 -138
rect -4439 138 -4393 150
rect -4439 -138 -4433 138
rect -4399 -138 -4393 138
rect -4439 -150 -4393 -138
rect -4343 138 -4297 150
rect -4343 -138 -4337 138
rect -4303 -138 -4297 138
rect -4343 -150 -4297 -138
rect -4247 138 -4201 150
rect -4247 -138 -4241 138
rect -4207 -138 -4201 138
rect -4247 -150 -4201 -138
rect -4151 138 -4105 150
rect -4151 -138 -4145 138
rect -4111 -138 -4105 138
rect -4151 -150 -4105 -138
rect -4055 138 -4009 150
rect -4055 -138 -4049 138
rect -4015 -138 -4009 138
rect -4055 -150 -4009 -138
rect -3959 138 -3913 150
rect -3959 -138 -3953 138
rect -3919 -138 -3913 138
rect -3959 -150 -3913 -138
rect -3863 138 -3817 150
rect -3863 -138 -3857 138
rect -3823 -138 -3817 138
rect -3863 -150 -3817 -138
rect -3767 138 -3721 150
rect -3767 -138 -3761 138
rect -3727 -138 -3721 138
rect -3767 -150 -3721 -138
rect -3671 138 -3625 150
rect -3671 -138 -3665 138
rect -3631 -138 -3625 138
rect -3671 -150 -3625 -138
rect -3575 138 -3529 150
rect -3575 -138 -3569 138
rect -3535 -138 -3529 138
rect -3575 -150 -3529 -138
rect -3479 138 -3433 150
rect -3479 -138 -3473 138
rect -3439 -138 -3433 138
rect -3479 -150 -3433 -138
rect -3383 138 -3337 150
rect -3383 -138 -3377 138
rect -3343 -138 -3337 138
rect -3383 -150 -3337 -138
rect -3287 138 -3241 150
rect -3287 -138 -3281 138
rect -3247 -138 -3241 138
rect -3287 -150 -3241 -138
rect -3191 138 -3145 150
rect -3191 -138 -3185 138
rect -3151 -138 -3145 138
rect -3191 -150 -3145 -138
rect -3095 138 -3049 150
rect -3095 -138 -3089 138
rect -3055 -138 -3049 138
rect -3095 -150 -3049 -138
rect -2999 138 -2953 150
rect -2999 -138 -2993 138
rect -2959 -138 -2953 138
rect -2999 -150 -2953 -138
rect -2903 138 -2857 150
rect -2903 -138 -2897 138
rect -2863 -138 -2857 138
rect -2903 -150 -2857 -138
rect -2807 138 -2761 150
rect -2807 -138 -2801 138
rect -2767 -138 -2761 138
rect -2807 -150 -2761 -138
rect -2711 138 -2665 150
rect -2711 -138 -2705 138
rect -2671 -138 -2665 138
rect -2711 -150 -2665 -138
rect -2615 138 -2569 150
rect -2615 -138 -2609 138
rect -2575 -138 -2569 138
rect -2615 -150 -2569 -138
rect -2519 138 -2473 150
rect -2519 -138 -2513 138
rect -2479 -138 -2473 138
rect -2519 -150 -2473 -138
rect -2423 138 -2377 150
rect -2423 -138 -2417 138
rect -2383 -138 -2377 138
rect -2423 -150 -2377 -138
rect -2327 138 -2281 150
rect -2327 -138 -2321 138
rect -2287 -138 -2281 138
rect -2327 -150 -2281 -138
rect -2231 138 -2185 150
rect -2231 -138 -2225 138
rect -2191 -138 -2185 138
rect -2231 -150 -2185 -138
rect -2135 138 -2089 150
rect -2135 -138 -2129 138
rect -2095 -138 -2089 138
rect -2135 -150 -2089 -138
rect -2039 138 -1993 150
rect -2039 -138 -2033 138
rect -1999 -138 -1993 138
rect -2039 -150 -1993 -138
rect -1943 138 -1897 150
rect -1943 -138 -1937 138
rect -1903 -138 -1897 138
rect -1943 -150 -1897 -138
rect -1847 138 -1801 150
rect -1847 -138 -1841 138
rect -1807 -138 -1801 138
rect -1847 -150 -1801 -138
rect -1751 138 -1705 150
rect -1751 -138 -1745 138
rect -1711 -138 -1705 138
rect -1751 -150 -1705 -138
rect -1655 138 -1609 150
rect -1655 -138 -1649 138
rect -1615 -138 -1609 138
rect -1655 -150 -1609 -138
rect -1559 138 -1513 150
rect -1559 -138 -1553 138
rect -1519 -138 -1513 138
rect -1559 -150 -1513 -138
rect -1463 138 -1417 150
rect -1463 -138 -1457 138
rect -1423 -138 -1417 138
rect -1463 -150 -1417 -138
rect -1367 138 -1321 150
rect -1367 -138 -1361 138
rect -1327 -138 -1321 138
rect -1367 -150 -1321 -138
rect -1271 138 -1225 150
rect -1271 -138 -1265 138
rect -1231 -138 -1225 138
rect -1271 -150 -1225 -138
rect -1175 138 -1129 150
rect -1175 -138 -1169 138
rect -1135 -138 -1129 138
rect -1175 -150 -1129 -138
rect -1079 138 -1033 150
rect -1079 -138 -1073 138
rect -1039 -138 -1033 138
rect -1079 -150 -1033 -138
rect -983 138 -937 150
rect -983 -138 -977 138
rect -943 -138 -937 138
rect -983 -150 -937 -138
rect -887 138 -841 150
rect -887 -138 -881 138
rect -847 -138 -841 138
rect -887 -150 -841 -138
rect -791 138 -745 150
rect -791 -138 -785 138
rect -751 -138 -745 138
rect -791 -150 -745 -138
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
rect 745 138 791 150
rect 745 -138 751 138
rect 785 -138 791 138
rect 745 -150 791 -138
rect 841 138 887 150
rect 841 -138 847 138
rect 881 -138 887 138
rect 841 -150 887 -138
rect 937 138 983 150
rect 937 -138 943 138
rect 977 -138 983 138
rect 937 -150 983 -138
rect 1033 138 1079 150
rect 1033 -138 1039 138
rect 1073 -138 1079 138
rect 1033 -150 1079 -138
rect 1129 138 1175 150
rect 1129 -138 1135 138
rect 1169 -138 1175 138
rect 1129 -150 1175 -138
rect 1225 138 1271 150
rect 1225 -138 1231 138
rect 1265 -138 1271 138
rect 1225 -150 1271 -138
rect 1321 138 1367 150
rect 1321 -138 1327 138
rect 1361 -138 1367 138
rect 1321 -150 1367 -138
rect 1417 138 1463 150
rect 1417 -138 1423 138
rect 1457 -138 1463 138
rect 1417 -150 1463 -138
rect 1513 138 1559 150
rect 1513 -138 1519 138
rect 1553 -138 1559 138
rect 1513 -150 1559 -138
rect 1609 138 1655 150
rect 1609 -138 1615 138
rect 1649 -138 1655 138
rect 1609 -150 1655 -138
rect 1705 138 1751 150
rect 1705 -138 1711 138
rect 1745 -138 1751 138
rect 1705 -150 1751 -138
rect 1801 138 1847 150
rect 1801 -138 1807 138
rect 1841 -138 1847 138
rect 1801 -150 1847 -138
rect 1897 138 1943 150
rect 1897 -138 1903 138
rect 1937 -138 1943 138
rect 1897 -150 1943 -138
rect 1993 138 2039 150
rect 1993 -138 1999 138
rect 2033 -138 2039 138
rect 1993 -150 2039 -138
rect 2089 138 2135 150
rect 2089 -138 2095 138
rect 2129 -138 2135 138
rect 2089 -150 2135 -138
rect 2185 138 2231 150
rect 2185 -138 2191 138
rect 2225 -138 2231 138
rect 2185 -150 2231 -138
rect 2281 138 2327 150
rect 2281 -138 2287 138
rect 2321 -138 2327 138
rect 2281 -150 2327 -138
rect 2377 138 2423 150
rect 2377 -138 2383 138
rect 2417 -138 2423 138
rect 2377 -150 2423 -138
rect 2473 138 2519 150
rect 2473 -138 2479 138
rect 2513 -138 2519 138
rect 2473 -150 2519 -138
rect 2569 138 2615 150
rect 2569 -138 2575 138
rect 2609 -138 2615 138
rect 2569 -150 2615 -138
rect 2665 138 2711 150
rect 2665 -138 2671 138
rect 2705 -138 2711 138
rect 2665 -150 2711 -138
rect 2761 138 2807 150
rect 2761 -138 2767 138
rect 2801 -138 2807 138
rect 2761 -150 2807 -138
rect 2857 138 2903 150
rect 2857 -138 2863 138
rect 2897 -138 2903 138
rect 2857 -150 2903 -138
rect 2953 138 2999 150
rect 2953 -138 2959 138
rect 2993 -138 2999 138
rect 2953 -150 2999 -138
rect 3049 138 3095 150
rect 3049 -138 3055 138
rect 3089 -138 3095 138
rect 3049 -150 3095 -138
rect 3145 138 3191 150
rect 3145 -138 3151 138
rect 3185 -138 3191 138
rect 3145 -150 3191 -138
rect 3241 138 3287 150
rect 3241 -138 3247 138
rect 3281 -138 3287 138
rect 3241 -150 3287 -138
rect 3337 138 3383 150
rect 3337 -138 3343 138
rect 3377 -138 3383 138
rect 3337 -150 3383 -138
rect 3433 138 3479 150
rect 3433 -138 3439 138
rect 3473 -138 3479 138
rect 3433 -150 3479 -138
rect 3529 138 3575 150
rect 3529 -138 3535 138
rect 3569 -138 3575 138
rect 3529 -150 3575 -138
rect 3625 138 3671 150
rect 3625 -138 3631 138
rect 3665 -138 3671 138
rect 3625 -150 3671 -138
rect 3721 138 3767 150
rect 3721 -138 3727 138
rect 3761 -138 3767 138
rect 3721 -150 3767 -138
rect 3817 138 3863 150
rect 3817 -138 3823 138
rect 3857 -138 3863 138
rect 3817 -150 3863 -138
rect 3913 138 3959 150
rect 3913 -138 3919 138
rect 3953 -138 3959 138
rect 3913 -150 3959 -138
rect 4009 138 4055 150
rect 4009 -138 4015 138
rect 4049 -138 4055 138
rect 4009 -150 4055 -138
rect 4105 138 4151 150
rect 4105 -138 4111 138
rect 4145 -138 4151 138
rect 4105 -150 4151 -138
rect 4201 138 4247 150
rect 4201 -138 4207 138
rect 4241 -138 4247 138
rect 4201 -150 4247 -138
rect 4297 138 4343 150
rect 4297 -138 4303 138
rect 4337 -138 4343 138
rect 4297 -150 4343 -138
rect 4393 138 4439 150
rect 4393 -138 4399 138
rect 4433 -138 4439 138
rect 4393 -150 4439 -138
rect 4489 138 4535 150
rect 4489 -138 4495 138
rect 4529 -138 4535 138
rect 4489 -150 4535 -138
rect 4585 138 4631 150
rect 4585 -138 4591 138
rect 4625 -138 4631 138
rect 4585 -150 4631 -138
rect 4681 138 4727 150
rect 4681 -138 4687 138
rect 4721 -138 4727 138
rect 4681 -150 4727 -138
rect 4777 138 4823 150
rect 4777 -138 4783 138
rect 4817 -138 4823 138
rect 4777 -150 4823 -138
rect -4781 -188 -4723 -182
rect -4781 -222 -4769 -188
rect -4735 -222 -4723 -188
rect -4781 -228 -4723 -222
rect -4589 -188 -4531 -182
rect -4589 -222 -4577 -188
rect -4543 -222 -4531 -188
rect -4589 -228 -4531 -222
rect -4397 -188 -4339 -182
rect -4397 -222 -4385 -188
rect -4351 -222 -4339 -188
rect -4397 -228 -4339 -222
rect -4205 -188 -4147 -182
rect -4205 -222 -4193 -188
rect -4159 -222 -4147 -188
rect -4205 -228 -4147 -222
rect -4013 -188 -3955 -182
rect -4013 -222 -4001 -188
rect -3967 -222 -3955 -188
rect -4013 -228 -3955 -222
rect -3821 -188 -3763 -182
rect -3821 -222 -3809 -188
rect -3775 -222 -3763 -188
rect -3821 -228 -3763 -222
rect -3629 -188 -3571 -182
rect -3629 -222 -3617 -188
rect -3583 -222 -3571 -188
rect -3629 -228 -3571 -222
rect -3437 -188 -3379 -182
rect -3437 -222 -3425 -188
rect -3391 -222 -3379 -188
rect -3437 -228 -3379 -222
rect -3245 -188 -3187 -182
rect -3245 -222 -3233 -188
rect -3199 -222 -3187 -188
rect -3245 -228 -3187 -222
rect -3053 -188 -2995 -182
rect -3053 -222 -3041 -188
rect -3007 -222 -2995 -188
rect -3053 -228 -2995 -222
rect -2861 -188 -2803 -182
rect -2861 -222 -2849 -188
rect -2815 -222 -2803 -188
rect -2861 -228 -2803 -222
rect -2669 -188 -2611 -182
rect -2669 -222 -2657 -188
rect -2623 -222 -2611 -188
rect -2669 -228 -2611 -222
rect -2477 -188 -2419 -182
rect -2477 -222 -2465 -188
rect -2431 -222 -2419 -188
rect -2477 -228 -2419 -222
rect -2285 -188 -2227 -182
rect -2285 -222 -2273 -188
rect -2239 -222 -2227 -188
rect -2285 -228 -2227 -222
rect -2093 -188 -2035 -182
rect -2093 -222 -2081 -188
rect -2047 -222 -2035 -188
rect -2093 -228 -2035 -222
rect -1901 -188 -1843 -182
rect -1901 -222 -1889 -188
rect -1855 -222 -1843 -188
rect -1901 -228 -1843 -222
rect -1709 -188 -1651 -182
rect -1709 -222 -1697 -188
rect -1663 -222 -1651 -188
rect -1709 -228 -1651 -222
rect -1517 -188 -1459 -182
rect -1517 -222 -1505 -188
rect -1471 -222 -1459 -188
rect -1517 -228 -1459 -222
rect -1325 -188 -1267 -182
rect -1325 -222 -1313 -188
rect -1279 -222 -1267 -188
rect -1325 -228 -1267 -222
rect -1133 -188 -1075 -182
rect -1133 -222 -1121 -188
rect -1087 -222 -1075 -188
rect -1133 -228 -1075 -222
rect -941 -188 -883 -182
rect -941 -222 -929 -188
rect -895 -222 -883 -188
rect -941 -228 -883 -222
rect -749 -188 -691 -182
rect -749 -222 -737 -188
rect -703 -222 -691 -188
rect -749 -228 -691 -222
rect -557 -188 -499 -182
rect -557 -222 -545 -188
rect -511 -222 -499 -188
rect -557 -228 -499 -222
rect -365 -188 -307 -182
rect -365 -222 -353 -188
rect -319 -222 -307 -188
rect -365 -228 -307 -222
rect -173 -188 -115 -182
rect -173 -222 -161 -188
rect -127 -222 -115 -188
rect -173 -228 -115 -222
rect 19 -188 77 -182
rect 19 -222 31 -188
rect 65 -222 77 -188
rect 19 -228 77 -222
rect 211 -188 269 -182
rect 211 -222 223 -188
rect 257 -222 269 -188
rect 211 -228 269 -222
rect 403 -188 461 -182
rect 403 -222 415 -188
rect 449 -222 461 -188
rect 403 -228 461 -222
rect 595 -188 653 -182
rect 595 -222 607 -188
rect 641 -222 653 -188
rect 595 -228 653 -222
rect 787 -188 845 -182
rect 787 -222 799 -188
rect 833 -222 845 -188
rect 787 -228 845 -222
rect 979 -188 1037 -182
rect 979 -222 991 -188
rect 1025 -222 1037 -188
rect 979 -228 1037 -222
rect 1171 -188 1229 -182
rect 1171 -222 1183 -188
rect 1217 -222 1229 -188
rect 1171 -228 1229 -222
rect 1363 -188 1421 -182
rect 1363 -222 1375 -188
rect 1409 -222 1421 -188
rect 1363 -228 1421 -222
rect 1555 -188 1613 -182
rect 1555 -222 1567 -188
rect 1601 -222 1613 -188
rect 1555 -228 1613 -222
rect 1747 -188 1805 -182
rect 1747 -222 1759 -188
rect 1793 -222 1805 -188
rect 1747 -228 1805 -222
rect 1939 -188 1997 -182
rect 1939 -222 1951 -188
rect 1985 -222 1997 -188
rect 1939 -228 1997 -222
rect 2131 -188 2189 -182
rect 2131 -222 2143 -188
rect 2177 -222 2189 -188
rect 2131 -228 2189 -222
rect 2323 -188 2381 -182
rect 2323 -222 2335 -188
rect 2369 -222 2381 -188
rect 2323 -228 2381 -222
rect 2515 -188 2573 -182
rect 2515 -222 2527 -188
rect 2561 -222 2573 -188
rect 2515 -228 2573 -222
rect 2707 -188 2765 -182
rect 2707 -222 2719 -188
rect 2753 -222 2765 -188
rect 2707 -228 2765 -222
rect 2899 -188 2957 -182
rect 2899 -222 2911 -188
rect 2945 -222 2957 -188
rect 2899 -228 2957 -222
rect 3091 -188 3149 -182
rect 3091 -222 3103 -188
rect 3137 -222 3149 -188
rect 3091 -228 3149 -222
rect 3283 -188 3341 -182
rect 3283 -222 3295 -188
rect 3329 -222 3341 -188
rect 3283 -228 3341 -222
rect 3475 -188 3533 -182
rect 3475 -222 3487 -188
rect 3521 -222 3533 -188
rect 3475 -228 3533 -222
rect 3667 -188 3725 -182
rect 3667 -222 3679 -188
rect 3713 -222 3725 -188
rect 3667 -228 3725 -222
rect 3859 -188 3917 -182
rect 3859 -222 3871 -188
rect 3905 -222 3917 -188
rect 3859 -228 3917 -222
rect 4051 -188 4109 -182
rect 4051 -222 4063 -188
rect 4097 -222 4109 -188
rect 4051 -228 4109 -222
rect 4243 -188 4301 -182
rect 4243 -222 4255 -188
rect 4289 -222 4301 -188
rect 4243 -228 4301 -222
rect 4435 -188 4493 -182
rect 4435 -222 4447 -188
rect 4481 -222 4493 -188
rect 4435 -228 4493 -222
rect 4627 -188 4685 -182
rect 4627 -222 4639 -188
rect 4673 -222 4685 -188
rect 4627 -228 4685 -222
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -4914 -307 4914 307
string parameters w 1.5 l 0.15 m 1 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
