* NGSPICE file created from /home/eamta/caravel_eamta_2021/mag/user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_DDZS4V VSUBS a_1316_n761# a_1456_n664# a_n524_n664#
+ w_n1652_n884# a_70_n664# a_128_n761# a_n920_n664# a_n1060_n761# a_268_n664# a_n1258_n761#
+ a_524_n761# a_664_n664# a_n466_n761# a_n1118_n664# a_920_n761# a_1118_n761# a_1060_n664#
+ a_1258_n664# a_n862_n761# a_n1514_n664# a_n326_n664# a_n722_n664# a_n70_n761# a_326_n761#
+ a_466_n664# a_n1456_n761# a_n268_n761# a_722_n761# a_862_n664# a_n664_n761# a_n1316_n664#
+ a_n128_n664#
X0 a_n722_n664# a_n862_n761# a_n920_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X1 a_466_n664# a_326_n761# a_268_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X2 a_n920_n664# a_n1060_n761# a_n1118_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X3 a_1456_n664# a_1316_n761# a_1258_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X4 a_1060_n664# a_920_n761# a_862_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X5 a_n326_n664# a_n466_n761# a_n524_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X6 a_664_n664# a_524_n761# a_466_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X7 a_n1118_n664# a_n1258_n761# a_n1316_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X8 a_n524_n664# a_n664_n761# a_n722_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X9 a_268_n664# a_128_n761# a_70_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X10 a_70_n664# a_n70_n761# a_n128_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X11 a_1258_n664# a_1118_n761# a_1060_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X12 a_862_n664# a_722_n761# a_664_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X13 a_n128_n664# a_n268_n761# a_n326_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X14 a_n1316_n664# a_n1456_n761# a_n1514_n664# w_n1652_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
.ends

.subckt M5_B VSUBS a_3389_167# a_9069_167# m1_1675_167# m1_1279_167# a_8673_167# m1_91_167#
+ w_n104_n76# a_8277_167# a_7881_167# m1_883_167# a_7485_167# m1_487_167# a_6161_167#
+ a_7089_167# a_5765_167# a_5369_167# a_6693_167# a_4973_167# a_4577_167# m1_2863_167#
+ a_4181_167# m1_2467_167# a_3447_70# a_3587_167# a_3785_167# a_9465_167# m1_2071_167#
Xsky130_fd_pr__pfet_01v8_DDZS4V_0 VSUBS a_3447_70# a_3587_167# a_3587_167# w_n104_n76#
+ m1_1675_167# a_3447_70# a_3587_167# a_3447_70# a_3587_167# a_3447_70# a_3447_70#
+ a_3587_167# a_3447_70# m1_487_167# a_3447_70# a_3447_70# a_3587_167# m1_2863_167#
+ a_3447_70# m1_91_167# m1_1279_167# m1_883_167# a_3447_70# a_3447_70# m1_2071_167#
+ a_3447_70# a_3447_70# a_3447_70# m1_2467_167# a_3447_70# a_3587_167# a_3587_167#
+ sky130_fd_pr__pfet_01v8_DDZS4V
X0 a_3587_167# a_3447_70# a_7485_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=4.79196e+13p pd=3.44115e+08u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X1 a_3587_167# a_3447_70# a_8673_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X2 a_3587_167# a_3447_70# a_7881_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X3 a_6161_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X4 a_3587_167# a_3447_70# a_3785_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X5 a_5369_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X6 a_7485_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X7 a_8673_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X8 a_9069_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X9 a_3785_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X10 a_4973_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X11 a_3587_167# a_3447_70# a_6161_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X12 a_3587_167# a_3447_70# a_7089_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X13 a_3587_167# a_3447_70# a_8277_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X14 a_3587_167# a_3447_70# a_9465_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X15 a_3587_167# a_3447_70# a_3389_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X16 a_3587_167# a_3447_70# a_4577_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X17 a_3587_167# a_3447_70# a_5765_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X18 a_3587_167# a_3447_70# a_6693_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X19 a_8277_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X20 a_9465_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X21 a_4181_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X22 a_5765_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X23 a_4577_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X24 a_7881_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X25 a_3587_167# a_3447_70# a_9069_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X26 a_7089_167# a_3447_70# a_3587_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X27 a_3587_167# a_3447_70# a_4973_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X28 a_3587_167# a_3447_70# a_4181_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X29 a_3587_167# a_3447_70# a_5369_167# w_n104_n76# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MXMZMC a_367_n801# a_n29_n801# a_227_n827# a_n425_n801#
+ a_n169_n827# a_169_n801# a_29_n827# a_n227_n801# w_n563_n949# a_n367_n827#
X0 a_n227_n801# a_n367_n827# a_n425_n801# w_n563_n949# sky130_fd_pr__nfet_01v8 ad=2.233e+12p pd=1.598e+07u as=2.233e+12p ps=1.598e+07u w=7.7e+06u l=700000u
X1 a_n29_n801# a_n169_n827# a_n227_n801# w_n563_n949# sky130_fd_pr__nfet_01v8 ad=2.233e+12p pd=1.598e+07u as=0p ps=0u w=7.7e+06u l=700000u
X2 a_169_n801# a_29_n827# a_n29_n801# w_n563_n949# sky130_fd_pr__nfet_01v8 ad=2.233e+12p pd=1.598e+07u as=0p ps=0u w=7.7e+06u l=700000u
X3 a_367_n801# a_227_n827# a_169_n801# w_n563_n949# sky130_fd_pr__nfet_01v8 ad=2.233e+12p pd=1.598e+07u as=0p ps=0u w=7.7e+06u l=700000u
.ends

.subckt M3 VSUBS m1_1812_2442# m1_2548_645# m1_2152_645# m1_1756_645#
Xsky130_fd_pr__nfet_01v8_MXMZMC_0 m1_2548_645# m1_2152_645# m1_1812_2442# m1_1756_645#
+ m1_1812_2442# m1_1812_2442# m1_1812_2442# m1_1812_2442# VSUBS m1_1812_2442# sky130_fd_pr__nfet_01v8_MXMZMC
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_2674SJ VSUBS c1_n2450_n2400# m3_n2550_n2500#
X0 c1_n2450_n2400# m3_n2550_n2500# sky130_fd_pr__cap_mim_m3_1 l=2.4e+07u w=2.4e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_DDDKZT VSUBS a_227_n761# a_367_n664# a_n169_n761#
+ a_623_n761# a_n29_n664# a_763_n664# a_n565_n761# w_n1157_n884# a_n961_n761# a_n425_n664#
+ a_29_n761# a_n821_n664# a_169_n664# a_425_n761# a_565_n664# a_n367_n761# a_n1019_n664#
+ a_821_n761# a_961_n664# a_n763_n761# a_n227_n664# a_n623_n664#
X0 a_n227_n664# a_n367_n761# a_n425_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X1 a_n821_n664# a_n961_n761# a_n1019_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X2 a_565_n664# a_425_n761# a_367_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X3 a_n425_n664# a_n565_n761# a_n623_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X4 a_169_n664# a_29_n761# a_n29_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X5 a_763_n664# a_623_n761# a_565_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X6 a_n29_n664# a_n169_n761# a_n227_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X7 a_367_n664# a_227_n761# a_169_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X8 a_n623_n664# a_n763_n761# a_n821_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X9 a_961_n664# a_821_n761# a_763_n664# w_n1157_n884# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
.ends

.subckt M8 VSUBS m1_2077_167# m1_1681_167# m1_1285_167# m1_889_167# m1_493_167# m1_97_179#
+ w_n182_n122# m1_143_80#
Xsky130_fd_pr__pfet_01v8_DDDKZT_0 VSUBS m1_143_80# m1_143_80# m1_143_80# m1_143_80#
+ m1_143_80# m1_143_80# m1_143_80# w_n182_n122# m1_143_80# m1_143_80# m1_143_80# m1_143_80#
+ m1_1285_167# m1_143_80# m1_1681_167# m1_143_80# m1_97_179# m1_143_80# m1_2077_167#
+ m1_143_80# m1_889_167# m1_493_167# sky130_fd_pr__pfet_01v8_DDDKZT
.ends

.subckt sky130_fd_pr__nfet_01v8_93MENK a_n1744_n357# a_1088_n357# VSUBS a_2386_n357#
+ a_3684_n357# a_4982_n357# a_2032_n357# a_734_n357# a_3330_n357# a_n3097_n269# a_5218_n357#
+ a_n5693_n269# a_2095_n269# a_n265_n269# a_n4395_n269# a_n1390_n357# a_4691_n269#
+ a_3393_n269# a_797_n269# a_n4041_n269# a_n4576_n357# a_n3278_n357# a_443_n269# a_n5874_n357#
+ a_n446_n357# a_n4222_n357# a_380_n357# a_n5520_n357# a_n92_n357# a_2858_n357# a_1206_n357#
+ a_2504_n357# a_3802_n357# a_n1681_n269# a_1269_n269# a_n3569_n269# a_n4867_n269#
+ a_3865_n269# a_2567_n269# a_n737_n269# a_n1862_n357# a_n3215_n269# a_n5811_n269#
+ a_2213_n269# a_n4513_n269# a_3511_n269# a_915_n269# a_n918_n357# a_2150_n357# a_852_n357#
+ a_4038_n357# a_5336_n357# a_n383_n269# a_n2098_n357# a_5399_n269# a_n4694_n357#
+ a_n3396_n357# a_561_n269# a_n564_n357# a_5045_n269# a_n4340_n357# a_n3042_n357#
+ a_n210_n357# a_1678_n357# a_2976_n357# a_1324_n357# a_2622_n357# a_3920_n357# a_n2389_n269#
+ a_5808_n357# a_1387_n269# a_n3687_n269# a_n4985_n269# a_3983_n269# a_2685_n269#
+ a_n855_n269# a_n2035_n269# a_n1980_n357# a_1033_n269# a_n3333_n269# a_2331_n269#
+ a_n501_n269# a_n4631_n269# a_n3868_n357# a_4219_n269# a_n3514_n357# a_n2216_n357#
+ a_970_n357# a_5517_n269# a_n4812_n357# a_4156_n357# a_5454_n357# a_5100_n357# a_n682_n357#
+ a_5163_n269# a_n3160_n357# a_1859_n269# a_n5048_n357# a_n1209_n269# a_n2507_n269#
+ a_1796_n357# a_1505_n269# a_n3805_n269# a_2803_n269# a_1442_n357# a_2740_n357# a_4628_n357#
+ a_n973_n269# a_n2153_n269# a_n3451_n269# a_26_n357# a_1151_n269# a_n3986_n357# a_n2688_n357#
+ a_n5339_n269# a_n1036_n357# a_4337_n269# a_3039_n269# a_n2334_n357# a_5635_n269#
+ a_89_n269# a_n4930_n357# a_n3632_n357# a_4274_n357# a_n800_n357# a_5572_n357# a_1914_n357#
+ a_5281_n269# a_n2979_n269# a_1977_n269# a_n5166_n357# a_n1327_n269# a_n2625_n269#
+ a_1623_n269# a_n3923_n269# a_2921_n269# a_1560_n357# a_n1508_n357# a_4809_n269#
+ a_n2806_n357# a_3448_n357# a_n29_n269# a_4746_n357# a_n2271_n269# a_n5457_n269#
+ a_n4159_n269# a_n1154_n357# a_4455_n269# a_3157_n269# a_n2452_n357# a_5753_n269#
+ a_n5103_n269# a_n3750_n357# a_498_n357# a_3094_n357# a_4392_n357# a_4101_n269# a_5690_n357#
+ a_207_n269# a_n5638_n357# a_144_n357# a_n1799_n269# a_n5284_n357# a_n1445_n269#
+ a_n2743_n269# a_1741_n269# a_n5929_n269# a_3629_n269# a_n1626_n357# a_4927_n269#
+ a_n2924_n357# a_2268_n357# a_3566_n357# a_4864_n357# a_3212_n357# a_n1091_n269#
+ a_616_n357# a_4510_n357# a_n5575_n269# a_n147_n269# a_n4277_n269# a_n1272_n357#
+ a_4573_n269# a_3275_n269# a_679_n269# a_n2570_n357# a_5871_n269# a_n5221_n269# a_n4458_n357#
+ a_325_n269# a_n1917_n269# a_n5756_n357# a_n328_n357# a_n4104_n357# a_262_n357# a_n5402_n357#
+ a_n1563_n269# a_n2861_n269# a_n4749_n269# a_3747_n269# a_2449_n269# a_n619_n269#
X0 a_n147_n269# a_n210_n357# a_n265_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X1 a_1623_n269# a_1560_n357# a_1505_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X2 a_4101_n269# a_4038_n357# a_3983_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X3 a_561_n269# a_498_n357# a_443_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X4 a_n1091_n269# a_n1154_n357# a_n1209_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X5 a_4691_n269# a_4628_n357# a_4573_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X6 a_n1681_n269# a_n1744_n357# a_n1799_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X7 a_n3333_n269# a_n3396_n357# a_n3451_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X8 a_1505_n269# a_1442_n357# a_1387_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X9 a_n3923_n269# a_n3986_n357# a_n4041_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X10 a_3157_n269# a_3094_n357# a_3039_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X11 a_n973_n269# a_n1036_n357# a_n1091_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X12 a_3747_n269# a_3684_n357# a_3629_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X13 a_4573_n269# a_4510_n357# a_4455_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X14 a_n1563_n269# a_n1626_n357# a_n1681_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X15 a_n3215_n269# a_n3278_n357# a_n3333_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X16 a_1387_n269# a_1324_n357# a_1269_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X17 a_n3805_n269# a_n3868_n357# a_n3923_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X18 a_n4041_n269# a_n4104_n357# a_n4159_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X19 a_1977_n269# a_1914_n357# a_1859_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X20 a_3629_n269# a_3566_n357# a_3511_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X21 a_n1445_n269# a_n1508_n357# a_n1563_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X22 a_n3097_n269# a_n3160_n357# a_n3215_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X23 a_1269_n269# a_1206_n357# a_1151_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X24 a_n3687_n269# a_n3750_n357# a_n3805_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X25 a_n5339_n269# a_n5402_n357# a_n5457_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X26 a_n737_n269# a_n800_n357# a_n855_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X27 a_n2979_n269# a_n3042_n357# a_n3097_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X28 a_n3569_n269# a_n3632_n357# a_n3687_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X29 a_n619_n269# a_n682_n357# a_n737_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X30 a_2331_n269# a_2268_n357# a_2213_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X31 a_2921_n269# a_2858_n357# a_2803_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X32 a_443_n269# a_380_n357# a_325_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X33 a_1033_n269# a_970_n357# a_915_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X34 a_2213_n269# a_2150_n357# a_2095_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X35 a_n4631_n269# a_n4694_n357# a_n4749_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X36 a_2803_n269# a_2740_n357# a_2685_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X37 a_325_n269# a_262_n357# a_207_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X38 a_915_n269# a_852_n357# a_797_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X39 a_4455_n269# a_4392_n357# a_4337_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X40 a_n2271_n269# a_n2334_n357# a_n2389_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X41 a_5281_n269# a_5218_n357# a_5163_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X42 a_5045_n269# a_4982_n357# a_4927_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X43 a_5871_n269# a_5808_n357# a_5753_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X44 a_n2861_n269# a_n2924_n357# a_n2979_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X45 a_2095_n269# a_2032_n357# a_1977_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X46 a_1859_n269# a_1796_n357# a_1741_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X47 a_n4513_n269# a_n4576_n357# a_n4631_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X48 a_207_n269# a_144_n357# a_89_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X49 a_2685_n269# a_2622_n357# a_2567_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X50 a_4337_n269# a_4274_n357# a_4219_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X51 a_797_n269# a_734_n357# a_679_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X52 a_n1327_n269# a_n1390_n357# a_n1445_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X53 a_n1917_n269# a_n1980_n357# a_n2035_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X54 a_n2153_n269# a_n2216_n357# a_n2271_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X55 a_5163_n269# a_5100_n357# a_5045_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X56 a_4927_n269# a_4864_n357# a_4809_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X57 a_n29_n269# a_n92_n357# a_n147_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X58 a_n2743_n269# a_n2806_n357# a_n2861_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X59 a_n4395_n269# a_n4458_n357# a_n4513_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X60 a_2567_n269# a_2504_n357# a_2449_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X61 a_4219_n269# a_4156_n357# a_4101_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X62 a_679_n269# a_616_n357# a_561_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X63 a_n1209_n269# a_n1272_n357# a_n1327_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X64 a_n1799_n269# a_n1862_n357# a_n1917_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X65 a_4809_n269# a_4746_n357# a_4691_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X66 a_n4277_n269# a_n4340_n357# a_n4395_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X67 a_n4867_n269# a_n4930_n357# a_n4985_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X68 a_n4159_n269# a_n4222_n357# a_n4277_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X69 a_n4749_n269# a_n4812_n357# a_n4867_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X70 a_3511_n269# a_3448_n357# a_3393_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X71 a_89_n269# a_26_n357# a_n29_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X72 a_5753_n269# a_5690_n357# a_5635_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X73 a_n5221_n269# a_n5284_n357# a_n5339_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X74 a_3393_n269# a_3330_n357# a_3275_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X75 a_n5811_n269# a_n5874_n357# a_n5929_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X76 a_n2035_n269# a_n2098_n357# a_n2153_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X77 a_3983_n269# a_3920_n357# a_3865_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X78 a_5635_n269# a_5572_n357# a_5517_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X79 a_n2625_n269# a_n2688_n357# a_n2743_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X80 a_n3451_n269# a_n3514_n357# a_n3569_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X81 a_2449_n269# a_2386_n357# a_2331_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X82 a_n5103_n269# a_n5166_n357# a_n5221_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X83 a_3275_n269# a_3212_n357# a_3157_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X84 a_3039_n269# a_2976_n357# a_2921_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X85 a_n5693_n269# a_n5756_n357# a_n5811_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X86 a_n501_n269# a_n564_n357# a_n619_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X87 a_3865_n269# a_3802_n357# a_3747_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X88 a_5517_n269# a_5454_n357# a_5399_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X89 a_n2507_n269# a_n2570_n357# a_n2625_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X90 a_n4985_n269# a_n5048_n357# a_n5103_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X91 a_n5575_n269# a_n5638_n357# a_n5693_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X92 a_n383_n269# a_n446_n357# a_n501_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X93 a_5399_n269# a_5336_n357# a_5281_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X94 a_n2389_n269# a_n2452_n357# a_n2507_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X95 a_n5457_n269# a_n5520_n357# a_n5575_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X96 a_n265_n269# a_n328_n357# a_n383_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X97 a_n855_n269# a_n918_n357# a_n973_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X98 a_1151_n269# a_1088_n357# a_1033_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X99 a_1741_n269# a_1678_n357# a_1623_n269# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F2M6PM a_n2806_n388# a_n1508_n388# VSUBS a_3448_n388#
+ a_4746_n388# a_1269_n300# a_n3569_n300# a_2567_n300# a_n737_n300# a_n4867_n300#
+ a_3865_n300# a_n3215_n300# a_n5811_n300# a_2213_n300# a_n4513_n300# a_3511_n300#
+ a_915_n300# a_n2452_n388# a_n1154_n388# a_n3750_n388# a_3094_n388# a_498_n388# a_4392_n388#
+ a_5690_n388# a_n5638_n388# a_n383_n300# a_144_n388# a_5399_n300# a_561_n300# a_5045_n300#
+ a_n5284_n388# a_n2924_n388# a_n1626_n388# a_2268_n388# a_n2389_n300# a_3566_n388#
+ a_4864_n388# a_n3687_n300# a_2685_n300# a_1387_n300# a_n855_n300# a_n4985_n300#
+ a_3212_n388# a_3983_n300# a_n2035_n300# a_n3333_n300# a_616_n388# a_4510_n388# a_2331_n300#
+ a_1033_n300# a_n4631_n300# a_n501_n300# a_4219_n300# a_n1272_n388# a_5517_n300#
+ a_n2570_n388# a_n5756_n388# a_n4458_n388# a_n328_n388# a_262_n388# a_n5402_n388#
+ a_n4104_n388# a_5163_n300# a_1859_n300# a_n1209_n300# a_n2507_n300# a_1505_n300#
+ a_n3805_n300# a_2803_n300# a_n1744_n388# a_1088_n388# a_2386_n388# a_3684_n388#
+ a_4982_n388# a_2032_n388# a_n973_n300# a_3330_n388# a_n2153_n300# a_n3451_n300#
+ a_734_n388# a_1151_n300# a_5218_n388# a_n5339_n300# a_4337_n300# a_3039_n300# a_n1390_n388#
+ a_5635_n300# a_89_n300# a_n3278_n388# a_n5874_n388# a_n4576_n388# a_n446_n388# a_380_n388#
+ a_n5520_n388# a_n4222_n388# a_n92_n388# a_5281_n300# a_2858_n388# a_n2979_n300#
+ a_1977_n300# a_1206_n388# a_2504_n388# a_n1327_n300# a_n2625_n300# a_3802_n388#
+ a_1623_n300# a_n3923_n300# a_2921_n300# a_4809_n300# a_n1862_n388# a_n29_n300# a_2150_n388#
+ a_n918_n388# a_n2271_n300# a_852_n388# a_4038_n388# a_5336_n388# a_n5457_n300# a_n4159_n300#
+ a_4455_n300# a_3157_n300# a_5753_n300# a_n2098_n388# a_n5103_n300# a_n3396_n388#
+ a_4101_n300# a_207_n300# a_n4694_n388# a_n564_n388# a_n3042_n388# a_n4340_n388#
+ a_n210_n388# a_1678_n388# a_2976_n388# a_n1799_n300# a_1324_n388# a_2622_n388# a_n1445_n300#
+ a_n2743_n300# a_3920_n388# a_1741_n300# a_5808_n388# a_n5929_n300# a_4927_n300#
+ a_3629_n300# a_n1980_n388# a_n3868_n388# a_n1091_n300# a_n2216_n388# a_n3514_n388#
+ a_970_n388# a_n4812_n388# a_4156_n388# a_5454_n388# a_n5575_n300# a_n4277_n300#
+ a_3275_n300# a_n147_n300# a_5100_n388# a_5871_n300# a_4573_n300# a_679_n300# a_n5221_n300#
+ a_325_n300# a_n682_n388# a_n1917_n300# a_n3160_n388# a_n5048_n388# a_1796_n388#
+ a_1442_n388# a_2740_n388# a_n1563_n300# a_n2861_n300# a_4628_n388# a_2449_n300#
+ a_n619_n300# a_n4749_n300# a_3747_n300# a_26_n388# a_n2688_n388# a_n3986_n388# a_n2334_n388#
+ a_n1036_n388# a_n3632_n388# a_n3097_n300# a_n4930_n388# a_n800_n388# a_4274_n388#
+ a_5572_n388# a_n5693_n300# a_2095_n300# a_n4395_n300# a_3393_n300# a_n265_n300#
+ a_4691_n300# a_797_n300# a_n4041_n300# a_1914_n388# a_443_n300# a_n5166_n388# a_1560_n388#
+ a_n1681_n300#
X0 a_n619_n300# a_n682_n388# a_n737_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X1 a_2331_n300# a_2268_n388# a_2213_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X2 a_443_n300# a_380_n388# a_325_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X3 a_2921_n300# a_2858_n388# a_2803_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X4 a_1033_n300# a_970_n388# a_915_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X5 a_2213_n300# a_2150_n388# a_2095_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X6 a_325_n300# a_262_n388# a_207_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X7 a_n4631_n300# a_n4694_n388# a_n4749_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X8 a_2803_n300# a_2740_n388# a_2685_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X9 a_4455_n300# a_4392_n388# a_4337_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X10 a_915_n300# a_852_n388# a_797_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X11 a_5281_n300# a_5218_n388# a_5163_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X12 a_5045_n300# a_4982_n388# a_4927_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X13 a_n2271_n300# a_n2334_n388# a_n2389_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X14 a_n2861_n300# a_n2924_n388# a_n2979_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X15 a_5871_n300# a_5808_n388# a_5753_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X16 a_2095_n300# a_2032_n388# a_1977_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X17 a_1859_n300# a_1796_n388# a_1741_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X18 a_207_n300# a_144_n388# a_89_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X19 a_n4513_n300# a_n4576_n388# a_n4631_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X20 a_2685_n300# a_2622_n388# a_2567_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X21 a_797_n300# a_734_n388# a_679_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X22 a_n1327_n300# a_n1390_n388# a_n1445_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X23 a_4337_n300# a_4274_n388# a_4219_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X24 a_5163_n300# a_5100_n388# a_5045_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X25 a_4927_n300# a_4864_n388# a_4809_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X26 a_n29_n300# a_n92_n388# a_n147_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X27 a_n1917_n300# a_n1980_n388# a_n2035_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X28 a_n2153_n300# a_n2216_n388# a_n2271_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X29 a_n2743_n300# a_n2806_n388# a_n2861_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X30 a_n4395_n300# a_n4458_n388# a_n4513_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X31 a_2567_n300# a_2504_n388# a_2449_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X32 a_679_n300# a_616_n388# a_561_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X33 a_n1209_n300# a_n1272_n388# a_n1327_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X34 a_4219_n300# a_4156_n388# a_4101_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X35 a_4809_n300# a_4746_n388# a_4691_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X36 a_n1799_n300# a_n1862_n388# a_n1917_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X37 a_n4277_n300# a_n4340_n388# a_n4395_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X38 a_n4867_n300# a_n4930_n388# a_n4985_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X39 a_n4159_n300# a_n4222_n388# a_n4277_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X40 a_n4749_n300# a_n4812_n388# a_n4867_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X41 a_3511_n300# a_3448_n388# a_3393_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X42 a_89_n300# a_26_n388# a_n29_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X43 a_5753_n300# a_5690_n388# a_5635_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X44 a_n5221_n300# a_n5284_n388# a_n5339_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X45 a_3393_n300# a_3330_n388# a_3275_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X46 a_n5811_n300# a_n5874_n388# a_n5929_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X47 a_n2035_n300# a_n2098_n388# a_n2153_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X48 a_3983_n300# a_3920_n388# a_3865_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X49 a_n2625_n300# a_n2688_n388# a_n2743_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X50 a_5635_n300# a_5572_n388# a_5517_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X51 a_n3451_n300# a_n3514_n388# a_n3569_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X52 a_2449_n300# a_2386_n388# a_2331_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X53 a_n5103_n300# a_n5166_n388# a_n5221_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X54 a_3275_n300# a_3212_n388# a_3157_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X55 a_3039_n300# a_2976_n388# a_2921_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X56 a_n5693_n300# a_n5756_n388# a_n5811_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X57 a_n501_n300# a_n564_n388# a_n619_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X58 a_3865_n300# a_3802_n388# a_3747_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X59 a_n2507_n300# a_n2570_n388# a_n2625_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X60 a_5517_n300# a_5454_n388# a_5399_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X61 a_n4985_n300# a_n5048_n388# a_n5103_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X62 a_n5575_n300# a_n5638_n388# a_n5693_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X63 a_n383_n300# a_n446_n388# a_n501_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X64 a_n2389_n300# a_n2452_n388# a_n2507_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X65 a_5399_n300# a_5336_n388# a_5281_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X66 a_n5457_n300# a_n5520_n388# a_n5575_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X67 a_n265_n300# a_n328_n388# a_n383_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X68 a_n855_n300# a_n918_n388# a_n973_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X69 a_1151_n300# a_1088_n388# a_1033_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X70 a_1741_n300# a_1678_n388# a_1623_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X71 a_n147_n300# a_n210_n388# a_n265_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X72 a_1623_n300# a_1560_n388# a_1505_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X73 a_561_n300# a_498_n388# a_443_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X74 a_n1091_n300# a_n1154_n388# a_n1209_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X75 a_4101_n300# a_4038_n388# a_3983_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X76 a_n1681_n300# a_n1744_n388# a_n1799_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X77 a_4691_n300# a_4628_n388# a_4573_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X78 a_n3333_n300# a_n3396_n388# a_n3451_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X79 a_1505_n300# a_1442_n388# a_1387_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X80 a_n3923_n300# a_n3986_n388# a_n4041_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X81 a_3157_n300# a_3094_n388# a_3039_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X82 a_n973_n300# a_n1036_n388# a_n1091_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X83 a_3747_n300# a_3684_n388# a_3629_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X84 a_n1563_n300# a_n1626_n388# a_n1681_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X85 a_4573_n300# a_4510_n388# a_4455_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X86 a_n3215_n300# a_n3278_n388# a_n3333_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X87 a_1387_n300# a_1324_n388# a_1269_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X88 a_n3805_n300# a_n3868_n388# a_n3923_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X89 a_n4041_n300# a_n4104_n388# a_n4159_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X90 a_1977_n300# a_1914_n388# a_1859_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X91 a_3629_n300# a_3566_n388# a_3511_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X92 a_n1445_n300# a_n1508_n388# a_n1563_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X93 a_n3097_n300# a_n3160_n388# a_n3215_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X94 a_1269_n300# a_1206_n388# a_1151_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X95 a_n3687_n300# a_n3750_n388# a_n3805_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X96 a_n5339_n300# a_n5402_n388# a_n5457_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X97 a_n737_n300# a_n800_n388# a_n855_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X98 a_n2979_n300# a_n3042_n388# a_n3097_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X99 a_n3569_n300# a_n3632_n388# a_n3687_n300# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt M6 m1_7781_n610# m1_2825_n610# m1_229_n610# m1_8725_n610# m1_1881_n610# m1_465_n610#
+ m1_4949_n610# m1_10377_n610# m1_7073_n610# m1_8961_n610# m1_11557_n610# m1_4241_n610#
+ m1_2353_n610# m1_4477_n610# m1_1409_n610# m1_n7_n610# m1_10849_n610# m1_7545_n610#
+ m1_1645_n610# m1_9197_n610# m1_11793_n610# m1_701_n610# m1_4005_n610# m1_n115_10#
+ m1_3533_n610# m1_937_n610# m1_3061_n610# m1_2589_n610# m1_1173_n610# m1_9669_n610#
+ m1_5893_n610# m1_8017_n610# m1_5657_n610# m1_10613_n610# m1_6129_n610# m1_4713_n610#
+ m1_2117_n610# m1_111_n610# m1_3769_n610# m1_8489_n610# m1_5185_n610# m1_9433_n610#
+ m1_6601_n610# m1_11321_n610# m1_3297_n610# m1_7309_n610# m1_9905_n610# m1_8253_n610#
+ m1_5421_n610# m1_10141_n610# m1_6365_n610# m1_11085_n610# m1_6837_n610# sky130_fd_pr__nfet_01v8_F2M6PM_0/VSUBS
Xsky130_fd_pr__nfet_01v8_93MENK_0 m1_n115_10# m1_n115_10# sky130_fd_pr__nfet_01v8_F2M6PM_0/VSUBS
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_2825_n610#
+ m1_n115_10# m1_229_n610# m1_8017_n610# m1_5657_n610# m1_111_n610# m1_n115_10# m1_10613_n610#
+ m1_111_n610# m1_111_n610# m1_1881_n610# m1_n115_10# m1_n115_10# m1_6365_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_4241_n610# m1_111_n610# m1_2353_n610# m1_111_n610# m1_111_n610#
+ m1_8489_n610# m1_5185_n610# m1_n115_10# m1_111_n610# m1_111_n610# m1_111_n610# m1_1409_n610#
+ m1_9433_n610# m1_6837_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_11321_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_3533_n610# m1_n115_10# m1_7309_n610# m1_111_n610# m1_937_n610#
+ m1_9905_n610# m1_111_n610# m1_111_n610# m1_111_n610# m1_n115_10# m1_111_n610# m1_2589_n610#
+ m1_8253_n610# m1_5421_n610# m1_111_n610# m1_n115_10# m1_10141_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_11085_n610# m1_n115_10# m1_7781_n610# m1_n115_10# m1_4713_n610# m1_111_n610#
+ m1_n115_10# m1_111_n610# m1_2117_n610# m1_8725_n610# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_4949_n610# m1_3769_n610# m1_111_n610# m1_n115_10# m1_7073_n610# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_111_n610# m1_8961_n610# m1_n115_10# m1_11557_n610# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610#
+ m1_111_n610# m1_111_n610# m1_n115_10# m1_111_n610# m1_3297_n610# m1_7545_n610# m1_111_n610#
+ m1_111_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_n115_10# m1_5893_n610#
+ m1_n115_10# m1_111_n610# m1_465_n610# m1_111_n610# m1_n115_10# m1_10377_n610# m1_111_n610#
+ m1_n115_10# m1_111_n610# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_6129_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_4477_n610# m1_111_n610# m1_111_n610# m1_n7_n610# m1_111_n610# m1_n115_10# m1_10849_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_n115_10# m1_111_n610# m1_111_n610# m1_1645_n610# m1_n115_10# m1_111_n610# m1_9197_n610#
+ m1_6601_n610# m1_n115_10# m1_11793_n610# m1_701_n610# m1_n115_10# m1_111_n610# m1_4005_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_3061_n610#
+ m1_1173_n610# m1_9669_n610# m1_111_n610# m1_111_n610# sky130_fd_pr__nfet_01v8_93MENK
Xsky130_fd_pr__nfet_01v8_93MENK_1 m1_n115_10# m1_n115_10# sky130_fd_pr__nfet_01v8_F2M6PM_0/VSUBS
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_2825_n610#
+ m1_n115_10# m1_229_n610# m1_8017_n610# m1_5657_n610# m1_111_n610# m1_n115_10# m1_10613_n610#
+ m1_111_n610# m1_111_n610# m1_1881_n610# m1_n115_10# m1_n115_10# m1_6365_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_4241_n610# m1_111_n610# m1_2353_n610# m1_111_n610# m1_111_n610#
+ m1_8489_n610# m1_5185_n610# m1_n115_10# m1_111_n610# m1_111_n610# m1_111_n610# m1_1409_n610#
+ m1_9433_n610# m1_6837_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_11321_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_3533_n610# m1_n115_10# m1_7309_n610# m1_111_n610# m1_937_n610#
+ m1_9905_n610# m1_111_n610# m1_111_n610# m1_111_n610# m1_n115_10# m1_111_n610# m1_2589_n610#
+ m1_8253_n610# m1_5421_n610# m1_111_n610# m1_n115_10# m1_10141_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_11085_n610# m1_n115_10# m1_7781_n610# m1_n115_10# m1_4713_n610# m1_111_n610#
+ m1_n115_10# m1_111_n610# m1_2117_n610# m1_8725_n610# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_4949_n610# m1_3769_n610# m1_111_n610# m1_n115_10# m1_7073_n610# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_111_n610# m1_8961_n610# m1_n115_10# m1_11557_n610# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610#
+ m1_111_n610# m1_111_n610# m1_n115_10# m1_111_n610# m1_3297_n610# m1_7545_n610# m1_111_n610#
+ m1_111_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_n115_10# m1_5893_n610#
+ m1_n115_10# m1_111_n610# m1_465_n610# m1_111_n610# m1_n115_10# m1_10377_n610# m1_111_n610#
+ m1_n115_10# m1_111_n610# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_n115_10# m1_6129_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_4477_n610# m1_111_n610# m1_111_n610# m1_n7_n610# m1_111_n610# m1_n115_10# m1_10849_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_n115_10# m1_111_n610# m1_111_n610# m1_1645_n610# m1_n115_10# m1_111_n610# m1_9197_n610#
+ m1_6601_n610# m1_n115_10# m1_11793_n610# m1_701_n610# m1_n115_10# m1_111_n610# m1_4005_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_3061_n610#
+ m1_1173_n610# m1_9669_n610# m1_111_n610# m1_111_n610# sky130_fd_pr__nfet_01v8_93MENK
Xsky130_fd_pr__nfet_01v8_F2M6PM_0 m1_n115_10# m1_n115_10# sky130_fd_pr__nfet_01v8_F2M6PM_0/VSUBS
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_2353_n610# m1_8489_n610# m1_5185_n610# m1_111_n610#
+ m1_111_n610# m1_111_n610# m1_111_n610# m1_111_n610# m1_1409_n610# m1_9433_n610#
+ m1_6837_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_11321_n610# m1_111_n610# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_3533_n610# m1_n115_10# m1_n115_10#
+ m1_111_n610# m1_111_n610# m1_7309_n610# m1_111_n610# m1_937_n610# m1_n115_10# m1_9905_n610#
+ m1_111_n610# m1_2589_n610# m1_n115_10# m1_n115_10# m1_8253_n610# m1_111_n610# m1_111_n610#
+ m1_5421_n610# m1_10141_n610# m1_n115_10# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_11085_n610# m1_7781_n610# m1_4713_n610#
+ m1_111_n610# m1_111_n610# m1_2117_n610# m1_8725_n610# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_4949_n610# m1_n115_10# m1_3769_n610# m1_111_n610#
+ m1_n115_10# m1_7073_n610# m1_n115_10# m1_111_n610# m1_111_n610# m1_8961_n610# m1_n115_10#
+ m1_11557_n610# m1_111_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10# m1_111_n610# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_3297_n610# m1_n115_10# m1_7545_n610# m1_111_n610#
+ m1_111_n610# m1_111_n610# m1_n115_10# m1_5893_n610# m1_n115_10# m1_n115_10# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_465_n610# m1_111_n610# m1_10377_n610# m1_111_n610#
+ m1_111_n610# m1_n115_10# m1_111_n610# m1_n115_10# m1_111_n610# m1_6129_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610#
+ m1_n115_10# m1_n115_10# m1_4477_n610# m1_111_n610# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_n7_n610# m1_10849_n610# m1_111_n610# m1_n115_10# m1_n115_10# m1_111_n610# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_111_n610# m1_1645_n610#
+ m1_9197_n610# m1_111_n610# m1_n115_10# m1_11793_n610# m1_111_n610# m1_6601_n610#
+ m1_701_n610# m1_111_n610# m1_n115_10# m1_4005_n610# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_n115_10# m1_111_n610# m1_3061_n610# m1_n115_10# m1_111_n610# m1_111_n610#
+ m1_1173_n610# m1_9669_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10#
+ m1_n115_10# m1_2825_n610# m1_n115_10# m1_n115_10# m1_n115_10# m1_n115_10# m1_229_n610#
+ m1_8017_n610# m1_111_n610# m1_111_n610# m1_5657_n610# m1_10613_n610# m1_111_n610#
+ m1_1881_n610# m1_n115_10# m1_6365_n610# m1_n115_10# m1_n115_10# m1_4241_n610# sky130_fd_pr__nfet_01v8_F2M6PM
.ends

.subckt M4 VSUBS m1_6155_n92# m1_5419_1637# m1_5759_n92# m1_5363_n92# m1_5548_77#
Xsky130_fd_pr__nfet_01v8_MXMZMC_0 m1_6155_n92# m1_5759_n92# m1_5419_1637# m1_5363_n92#
+ m1_5419_1637# m1_5548_77# m1_5419_1637# m1_5548_77# VSUBS m1_5419_1637# sky130_fd_pr__nfet_01v8_MXMZMC
.ends

.subckt sky130_fd_pr__nfet_01v8_QMU5EQ a_n151_291# w_n1642_n479# a_n1504_n331# a_266_n331#
+ a_1029_291# a_n1150_n331# a_n741_291# a_793_291# a_n206_n331# a_738_n331# a_n33_291#
+ a_30_n331# a_85_291# a_384_n331# a_n1331_291# a_n1095_291# a_1383_291# a_321_291#
+ a_n678_n331# a_n324_n331# a_502_n331# a_856_n331# a_n623_291# a_911_291# a_n387_291#
+ a_675_291# a_1328_n331# a_n796_n331# a_n442_n331# a_974_n331# a_n1213_291# a_n977_291#
+ a_620_n331# a_1265_291# a_203_291# a_1446_n331# a_n914_n331# a_1092_n331# a_n505_291#
+ a_n560_n331# a_n269_291# a_557_291# a_n1268_n331# a_n859_291# a_1147_291# a_1210_n331#
+ a_148_n331# a_n1449_291# a_n1386_n331# a_439_291# a_n1032_n331# a_n88_n331#
X0 a_1092_n331# a_1029_291# a_974_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X1 a_n324_n331# a_n387_291# a_n442_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X2 a_n914_n331# a_n977_291# a_n1032_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X3 a_n206_n331# a_n269_291# a_n324_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X4 a_n796_n331# a_n859_291# a_n914_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X5 a_n678_n331# a_n741_291# a_n796_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X6 a_n88_n331# a_n151_291# a_n206_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X7 a_620_n331# a_557_291# a_502_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X8 a_n1032_n331# a_n1095_291# a_n1150_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X9 a_n560_n331# a_n623_291# a_n678_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X10 a_502_n331# a_439_291# a_384_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X11 a_1446_n331# a_1383_291# a_1328_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X12 a_384_n331# a_321_291# a_266_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X13 a_974_n331# a_911_291# a_856_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X14 a_1328_n331# a_1265_291# a_1210_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X15 a_n1386_n331# a_n1449_291# a_n1504_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X16 a_266_n331# a_203_291# a_148_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X17 a_n1268_n331# a_n1331_291# a_n1386_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X18 a_30_n331# a_n33_291# a_n88_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X19 a_n1150_n331# a_n1213_291# a_n1268_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X20 a_856_n331# a_793_291# a_738_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X21 a_738_n331# a_675_291# a_620_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X22 a_n442_n331# a_n505_291# a_n560_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X23 a_148_n331# a_85_291# a_30_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X24 a_1210_n331# a_1147_291# a_1092_n331# w_n1642_n479# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt M9 m1_n114_n283# m1_n180_n903# m1_n50_n1145# w_n546_n1326#
Xsky130_fd_pr__nfet_01v8_QMU5EQ_0 m1_n114_n283# w_n546_n1326# m1_n180_n903# m1_n50_n1145#
+ m1_n114_n283# m1_n50_n1145# m1_n114_n283# m1_n114_n283# m1_n50_n1145# m1_n50_n1145#
+ m1_n114_n283# m1_n50_n1145# m1_n114_n283# m1_n180_n903# m1_n114_n283# m1_n114_n283#
+ m1_n114_n283# m1_n114_n283# m1_n50_n1145# m1_n180_n903# m1_n50_n1145# m1_n180_n903#
+ m1_n114_n283# m1_n114_n283# m1_n114_n283# m1_n114_n283# m1_n180_n903# m1_n180_n903#
+ m1_n50_n1145# m1_n50_n1145# m1_n114_n283# m1_n114_n283# m1_n180_n903# m1_n114_n283#
+ m1_n114_n283# m1_n50_n1145# m1_n50_n1145# m1_n180_n903# m1_n114_n283# m1_n180_n903#
+ m1_n114_n283# m1_n114_n283# m1_n180_n903# m1_n114_n283# m1_n114_n283# m1_n50_n1145#
+ m1_n180_n903# m1_n114_n283# m1_n50_n1145# m1_n114_n283# m1_n180_n903# m1_n180_n903#
+ sky130_fd_pr__nfet_01v8_QMU5EQ
.ends

.subckt sky130_fd_pr__pfet_01v8_ZYZ5C6 VSUBS a_227_n761# a_3791_n761# a_3931_n664#
+ a_n2149_n761# a_3989_n761# a_367_n664# a_n4129_n761# a_n1357_n761# a_n169_n761#
+ a_n3337_n761# a_623_n761# a_n2545_n761# a_n2009_n664# a_n29_n664# a_763_n664# a_n1753_n761#
+ a_n565_n761# a_n1217_n664# a_n3733_n761# a_2009_n761# a_n2941_n761# a_1217_n761#
+ a_2149_n664# a_n3197_n664# a_n2405_n664# a_1357_n664# a_4129_n664# a_n961_n761#
+ a_2405_n761# a_n1613_n664# a_n425_n664# a_3337_n664# a_3197_n761# a_29_n761# a_1613_n761#
+ a_n3593_n664# a_n2801_n664# a_2545_n664# a_1753_n664# a_2801_n761# a_3593_n761#
+ a_n2999_n664# a_n821_n664# a_3733_n664# w_n4223_n764# a_169_n664# a_2941_n664# a_n1159_n761#
+ a_2999_n761# a_n3139_n761# a_425_n761# a_n2347_n761# a_565_n664# a_n1555_n761# a_n367_n761#
+ a_n1019_n664# a_n3535_n761# a_821_n761# a_1019_n761# a_n2743_n761# a_n2207_n664#
+ a_961_n664# a_1159_n664# a_n1951_n761# a_n763_n761# a_n1415_n664# a_n227_n664# a_3139_n664#
+ a_n3931_n761# a_2207_n761# a_n4187_n664# a_1415_n761# a_n3395_n664# a_n2603_n664#
+ a_2347_n664# a_1555_n664# a_2603_n761# a_3395_n761# a_n1811_n664# a_n623_n664# a_3535_n664#
+ a_2743_n664# a_1811_n761# a_n3791_n664# a_n3989_n664# a_1951_n664#
X0 a_n2999_n664# a_n3139_n761# a_n3197_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X1 a_n227_n664# a_n367_n761# a_n425_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X2 a_3931_n664# a_3791_n761# a_3733_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X3 a_n1415_n664# a_n1555_n761# a_n1613_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X4 a_1951_n664# a_1811_n761# a_1753_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X5 a_3139_n664# a_2999_n761# a_2941_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X6 a_n2009_n664# a_n2149_n761# a_n2207_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X7 a_n3593_n664# a_n3733_n761# a_n3791_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X8 a_n821_n664# a_n961_n761# a_n1019_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X9 a_565_n664# a_425_n761# a_367_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X10 a_2545_n664# a_2405_n761# a_2347_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X11 a_3535_n664# a_3395_n761# a_3337_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X12 a_n2603_n664# a_n2743_n761# a_n2801_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X13 a_n1019_n664# a_n1159_n761# a_n1217_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X14 a_1555_n664# a_1415_n761# a_1357_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X15 a_n3197_n664# a_n3337_n761# a_n3395_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X16 a_n425_n664# a_n565_n761# a_n623_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X17 a_2149_n664# a_2009_n761# a_1951_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X18 a_n1613_n664# a_n1753_n761# a_n1811_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X19 a_n2207_n664# a_n2347_n761# a_n2405_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X20 a_1159_n664# a_1019_n761# a_961_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X21 a_n3791_n664# a_n3931_n761# a_n3989_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X22 a_169_n664# a_29_n761# a_n29_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X23 a_763_n664# a_623_n761# a_565_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X24 a_2743_n664# a_2603_n761# a_2545_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X25 a_n29_n664# a_n169_n761# a_n227_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X26 a_3733_n664# a_3593_n761# a_3535_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X27 a_n1217_n664# a_n1357_n761# a_n1415_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X28 a_n2801_n664# a_n2941_n761# a_n2999_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X29 a_1753_n664# a_1613_n761# a_1555_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X30 a_n3395_n664# a_n3535_n761# a_n3593_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X31 a_367_n664# a_227_n761# a_169_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X32 a_2347_n664# a_2207_n761# a_2149_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X33 a_n623_n664# a_n763_n761# a_n821_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X34 a_n3989_n664# a_n4129_n761# a_n4187_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X35 a_3337_n664# a_3197_n761# a_3139_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X36 a_n1811_n664# a_n1951_n761# a_n2009_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X37 a_1357_n664# a_1217_n761# a_1159_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X38 a_n2405_n664# a_n2545_n761# a_n2603_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X39 a_961_n664# a_821_n761# a_763_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X40 a_2941_n664# a_2801_n761# a_2743_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X41 a_4129_n664# a_3989_n761# a_3931_n664# w_n4223_n764# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
.ends

.subckt sky130_fd_pr__pfet_01v8_9JQ4XZ a_n367_n1615# VSUBS a_n1811_118# a_425_n1615#
+ a_n3791_118# a_n1613_118# a_961_118# a_n821_n1518# a_n565_n1615# a_n169_21# a_623_n1615#
+ a_n3593_118# a_n1415_118# a_763_118# a_n3395_118# a_n1217_118# a_565_118# a_821_n1615#
+ a_n763_n1615# a_n3197_118# a_n1019_118# a_367_118# a_n4129_21# a_n565_21# a_2999_21#
+ a_169_118# a_n961_n1615# a_n2149_21# a_n29_118# a_n3197_n1518# a_169_n1518# a_3197_n1615#
+ a_n2999_118# a_n4187_n1518# a_n3337_21# a_n821_118# a_29_n1615# a_n3395_n1518# a_3395_n1615#
+ a_n1357_21# a_3197_21# a_n623_118# a_367_n1518# a_n961_21# a_n2545_21# a_2009_21#
+ a_n425_118# a_425_21# a_n3593_n1518# a_3593_n1615# a_565_n1518# a_n3733_21# a_n227_118#
+ a_n1753_21# a_1217_21# a_3593_21# a_763_n1518# a_n3791_n1518# a_3791_n1615# a_4129_118#
+ a_n2941_21# a_821_21# a_2405_21# a_961_n1518# a_n1019_n1518# a_1019_n1615# a_n2009_n1518#
+ a_n2999_n1518# a_2999_n1615# a_2009_n1615# a_1613_21# a_n3989_n1518# a_3989_n1615#
+ a_n1217_n1518# a_2801_21# a_1217_n1615# a_n2207_n1518# a_2207_n1615# a_3931_118#
+ a_n1415_n1518# a_1415_n1615# a_n1159_n1615# a_3733_118# a_n2405_n1518# a_2405_n1615#
+ a_n2149_n1615# a_n3139_n1615# a_3535_118# a_n1613_n1518# a_1613_n1615# a_n4129_n1615#
+ a_n2603_n1518# a_n1357_n1615# a_2603_n1615# a_3337_118# w_n4223_n1618# a_n2347_n1615#
+ a_n3337_n1615# a_3139_118# a_n1811_n1518# a_1811_n1615# a_n2801_n1518# a_n1555_n1615#
+ a_2801_n1615# a_n2545_n1615# a_n3535_n1615# a_n1753_n1615# a_n367_21# a_n2743_n1615#
+ a_1159_n1518# a_n3733_n1615# a_2149_n1518# a_3989_21# a_n1951_n1615# a_3139_n1518#
+ a_n3139_21# a_4129_n1518# a_n2941_n1615# a_2941_118# a_1357_n1518# a_29_21# a_n3931_n1615#
+ a_n1159_21# a_2347_n1518# a_2743_118# a_n763_21# a_3337_n1518# a_n2347_21# a_227_21#
+ a_1555_n1518# a_2545_118# a_2545_n1518# a_3535_n1518# a_2347_118# a_n3535_21# a_1019_21#
+ a_1753_n1518# a_n1555_21# a_3395_21# a_2743_n1518# a_2149_118# a_3733_n1518# a_2207_21#
+ a_n2743_21# a_623_21# a_n2801_118# a_1951_n1518# a_2941_n1518# a_n2603_118# a_n3931_21#
+ a_3931_n1518# a_1415_21# a_n1951_21# a_3791_21# a_n2405_118# a_2603_21# a_n2207_118#
+ a_1951_118# a_n4187_118# a_n2009_118# a_1753_118# a_n227_n1518# a_1811_21# a_1555_118#
+ w_n4223_18# a_1357_118# a_n29_n1518# a_n425_n1518# a_n3989_118# a_227_n1615# a_n169_n1615#
+ a_1159_118# a_n623_n1518#
X0 a_2545_n1518# a_2405_n1615# a_2347_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X1 a_n2999_118# a_n3139_21# a_n3197_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X2 a_n2801_118# a_n2941_21# a_n2999_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X3 a_n1613_118# a_n1753_21# a_n1811_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X4 a_n623_118# a_n763_21# a_n821_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X5 a_n2999_n1518# a_n3139_n1615# a_n3197_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X6 a_3337_118# a_3197_21# a_3139_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X7 a_n3593_n1518# a_n3733_n1615# a_n3791_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X8 a_1555_n1518# a_1415_n1615# a_1357_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X9 a_565_n1518# a_425_n1615# a_367_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X10 a_1357_118# a_1217_21# a_1159_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X11 a_2545_118# a_2405_21# a_2347_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X12 a_n2009_n1518# a_n2149_n1615# a_n2207_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X13 a_367_118# a_227_21# a_169_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X14 a_n2603_n1518# a_n2743_n1615# a_n2801_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X15 a_n425_n1518# a_n565_n1615# a_n623_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X16 a_n3989_118# a_n4129_21# a_n4187_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X17 a_n3791_118# a_n3931_21# a_n3989_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X18 a_n2603_118# a_n2743_21# a_n2801_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X19 a_n1415_118# a_n1555_21# a_n1613_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X20 a_3733_n1518# a_3593_n1615# a_3535_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X21 a_n425_118# a_n565_21# a_n623_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X22 a_n1019_n1518# a_n1159_n1615# a_n1217_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X23 a_169_118# a_29_21# a_n29_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X24 a_n1613_n1518# a_n1753_n1615# a_n1811_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X25 a_2347_n1518# a_2207_n1615# a_2149_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X26 a_2941_n1518# a_2801_n1615# a_2743_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X27 a_1159_118# a_1019_21# a_961_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X28 a_2347_118# a_2207_21# a_2149_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X29 a_n3593_118# a_n3733_21# a_n3791_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X30 a_n3395_n1518# a_n3535_n1615# a_n3593_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X31 a_1357_n1518# a_1217_n1615# a_1159_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X32 a_n2405_118# a_n2545_21# a_n2603_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X33 a_n1217_118# a_n1357_21# a_n1415_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X34 a_n227_118# a_n367_21# a_n425_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X35 a_1951_n1518# a_1811_n1615# a_1753_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X36 a_3931_118# a_3791_21# a_3733_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X37 a_169_n1518# a_29_n1615# a_n29_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X38 a_367_n1518# a_227_n1615# a_169_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X39 a_n2405_n1518# a_n2545_n1615# a_n2603_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X40 a_n227_n1518# a_n367_n1615# a_n425_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X41 a_961_n1518# a_821_n1615# a_763_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X42 a_3139_118# a_2999_21# a_2941_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X43 a_n821_n1518# a_n961_n1615# a_n1019_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X44 a_961_118# a_821_21# a_763_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X45 a_1951_118# a_1811_21# a_1753_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X46 a_2149_118# a_2009_21# a_1951_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X47 a_3535_n1518# a_3395_n1615# a_3337_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X48 a_n1415_n1518# a_n1555_n1615# a_n1613_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X49 a_n3395_118# a_n3535_21# a_n3593_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X50 a_n2207_118# a_n2347_21# a_n2405_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X51 a_n1019_118# a_n1159_21# a_n1217_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X52 a_2149_n1518# a_2009_n1615# a_1951_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X53 a_n29_118# a_n169_21# a_n227_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X54 a_2743_n1518# a_2603_n1615# a_2545_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X55 a_3733_118# a_3593_21# a_3535_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X56 a_4129_118# a_3989_21# a_3931_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=700000u
X57 a_n3197_n1518# a_n3337_n1615# a_n3395_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X58 a_1753_118# a_1613_21# a_1555_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X59 a_2941_118# a_2801_21# a_2743_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X60 a_n3791_n1518# a_n3931_n1615# a_n3989_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X61 a_1159_n1518# a_1019_n1615# a_961_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X62 a_1753_n1518# a_1613_n1615# a_1555_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X63 a_763_118# a_623_21# a_565_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X64 a_n3197_118# a_n3337_21# a_n3395_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X65 a_n1811_118# a_n1951_21# a_n2009_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X66 a_763_n1518# a_623_n1615# a_565_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X67 a_4129_n1518# a_3989_n1615# a_3931_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X68 a_n2009_118# a_n2149_21# a_n2207_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X69 a_n821_118# a_n961_21# a_n1019_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X70 a_n2801_n1518# a_n2941_n1615# a_n2999_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X71 a_n2207_n1518# a_n2347_n1615# a_n2405_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X72 a_n29_n1518# a_n169_n1615# a_n227_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X73 a_3535_118# a_3395_21# a_3337_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X74 a_n623_n1518# a_n763_n1615# a_n821_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X75 a_3337_n1518# a_3197_n1615# a_3139_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X76 a_3139_n1518# a_2999_n1615# a_2941_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X77 a_3931_n1518# a_3791_n1615# a_3733_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X78 a_n1217_n1518# a_n1357_n1615# a_n1415_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X79 a_565_118# a_425_21# a_367_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X80 a_1555_118# a_1415_21# a_1357_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X81 a_2743_118# a_2603_21# a_2545_118# w_n4223_18# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X82 a_n3989_n1518# a_n4129_n1615# a_n4187_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=700000u
X83 a_n1811_n1518# a_n1951_n1615# a_n2009_n1518# w_n4223_n1618# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
.ends

.subckt M7 VSUBS m1_7907_n4720# a_23485_n4733# a_11495_n4759# a_11635_n4733# m1_n211_n4721#
+ w_n1784_n5513#
Xsky130_fd_pr__pfet_01v8_ZYZ5C6_1 VSUBS a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_7907_n4720# w_n1784_n5513#
+ m1_7907_n4720# m1_7907_n4720# a_11495_n4759# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759# m1_7907_n4720# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_n211_n4721# sky130_fd_pr__pfet_01v8_ZYZ5C6
Xsky130_fd_pr__pfet_01v8_9JQ4XZ_0 a_11495_n4759# VSUBS m1_7907_n4720# a_11495_n4759#
+ m1_7907_n4720# m1_n211_n4721# m1_7907_n4720# m1_n211_n4721# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_n211_n4721# m1_7907_n4720# m1_n211_n4721# m1_7907_n4720# m1_n211_n4721#
+ m1_7907_n4720# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_7907_n4720# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759#
+ m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# a_11495_n4759# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# m1_n211_n4721# a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ m1_n211_n4721# a_11495_n4759# m1_n211_n4721# a_11495_n4759# m1_7907_n4720# a_11495_n4759#
+ m1_7907_n4720# a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_7907_n4720#
+ a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_7907_n4720#
+ m1_7907_n4720# a_11495_n4759# m1_n211_n4721# m1_7907_n4720# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_n211_n4721# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759#
+ m1_7907_n4720# a_11495_n4759# m1_n211_n4721# m1_7907_n4720# a_11495_n4759# a_11495_n4759#
+ m1_7907_n4720# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759#
+ m1_7907_n4720# w_n1784_n5513# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_7907_n4720#
+ a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# m1_7907_n4720# a_11495_n4759#
+ m1_7907_n4720# m1_7907_n4720# a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ m1_7907_n4720# m1_7907_n4720# m1_n211_n4721# m1_n211_n4721# a_11495_n4759# a_11495_n4759#
+ m1_7907_n4720# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720#
+ m1_7907_n4720# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ m1_n211_n4721# a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_7907_n4720# m1_n211_n4721#
+ m1_7907_n4720# m1_7907_n4720# a_11495_n4759# m1_n211_n4721# w_n1784_n5513# m1_7907_n4720#
+ m1_n211_n4721# m1_n211_n4721# m1_n211_n4721# a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ m1_7907_n4720# sky130_fd_pr__pfet_01v8_9JQ4XZ
Xsky130_fd_pr__pfet_01v8_ZYZ5C6_0 VSUBS a_11495_n4759# a_11495_n4759# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# m1_n211_n4721# m1_n211_n4721# m1_7907_n4720# m1_7907_n4720#
+ a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_7907_n4720# w_n1784_n5513#
+ m1_7907_n4720# m1_7907_n4720# a_11495_n4759# a_11495_n4759# a_11495_n4759# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# a_11495_n4759# a_11495_n4759# m1_7907_n4720# a_11495_n4759#
+ a_11495_n4759# a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721# a_11495_n4759#
+ a_11495_n4759# m1_7907_n4720# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# a_11495_n4759# m1_7907_n4720# m1_7907_n4720# m1_n211_n4721#
+ m1_n211_n4721# a_11495_n4759# m1_7907_n4720# m1_n211_n4721# m1_n211_n4721# sky130_fd_pr__pfet_01v8_ZYZ5C6
X0 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=5.3592e+14p pd=3.84912e+09u as=1.7052e+14p ps=1.22472e+09u w=7e+06u l=700000u
X1 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X2 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X3 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X4 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.7052e+14p ps=1.22472e+09u w=7e+06u l=700000u
X5 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X6 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X7 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X8 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X9 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X10 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X11 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X12 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X13 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X14 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X15 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X16 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X17 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X18 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X19 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X20 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X21 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X22 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X23 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X24 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X25 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X26 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X27 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X28 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X29 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X30 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X31 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X32 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X33 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X34 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X35 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X36 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X37 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X38 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X39 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X40 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X41 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X42 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X43 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X44 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X45 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X46 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X47 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X48 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X49 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X50 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X51 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X52 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X53 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X54 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X55 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X56 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X57 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X58 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X59 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X60 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X61 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X62 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X63 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X64 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X65 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X66 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X67 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X68 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X69 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X70 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X71 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X72 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X73 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X74 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X75 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X76 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X77 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X78 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X79 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X80 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X81 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X82 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X83 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X84 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X85 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X86 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X87 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X88 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X89 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X90 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X91 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X92 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X93 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X94 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X95 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X96 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X97 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X98 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X99 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X100 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X101 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X102 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X103 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X104 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X105 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X106 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X107 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X108 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X109 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X110 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X111 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X112 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X113 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X114 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X115 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X116 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X117 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X118 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X119 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X120 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X121 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X122 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X123 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X124 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X125 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X126 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X127 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X128 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X129 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X130 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X131 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X132 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X133 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X134 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X135 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X136 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X137 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X138 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X139 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X140 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X141 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X142 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X143 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X144 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X145 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X146 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X147 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X148 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X149 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X150 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X151 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X152 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X153 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X154 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X155 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X156 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X157 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X158 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X159 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X160 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X161 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X162 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X163 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X164 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X165 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X166 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X167 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X168 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X169 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X170 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X171 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X172 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X173 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X174 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X175 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X176 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X177 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X178 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X179 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X180 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X181 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X182 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X183 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X184 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X185 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X186 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X187 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X188 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X189 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X190 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X191 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X192 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X193 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X194 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X195 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X196 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X197 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X198 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X199 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X200 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X201 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X202 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X203 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X204 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X205 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X206 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X207 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X208 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X209 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X210 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X211 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X212 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X213 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X214 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X215 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X216 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X217 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X218 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X219 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X220 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X221 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X222 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X223 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X224 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X225 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X226 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X227 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X228 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X229 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X230 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X231 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X232 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X233 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X234 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X235 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X236 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X237 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X238 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X239 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X240 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X241 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X242 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X243 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X244 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X245 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X246 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X247 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X248 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X249 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X250 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X251 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X252 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X253 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X254 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X255 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X256 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X257 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X258 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X259 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X260 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X261 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X262 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X263 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X264 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X265 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X266 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X267 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X268 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X269 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X270 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X271 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X272 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X273 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X274 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X275 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X276 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X277 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X278 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X279 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X280 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X281 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X282 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X283 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X284 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X285 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X286 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X287 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X288 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X289 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X290 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X291 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X292 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X293 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X294 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X295 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X296 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X297 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X298 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X299 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X300 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X301 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X302 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X303 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X304 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X305 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X306 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X307 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X308 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X309 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X310 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X311 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X312 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X313 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X314 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X315 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X316 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X317 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X318 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X319 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X320 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X321 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X322 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X323 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X324 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X325 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X326 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X327 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X328 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X329 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X330 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X331 a_11635_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X332 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X333 m1_7907_n4720# a_11495_n4759# a_11635_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X334 m1_7907_n4720# a_11495_n4759# a_23485_n4733# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
X335 a_23485_n4733# a_11495_n4759# m1_7907_n4720# w_n1784_n5513# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=7e+06u l=700000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SNVJWU a_n5353_n461# a_n6929_n364# VSUBS a_1547_n461#
+ a_n5767_n461# a_1823_n461# a_6239_n461# a_6101_n461# a_n6791_n364# a_6181_n364#
+ a_n2317_n461# a_n385_n461# a_6515_n461# a_6595_n364# a_n3065_n364# a_n799_n461#
+ a_n3479_n364# a_n661_n461# a_6871_n364# a_n3341_n364# a_3145_n364# a_n3755_n364#
+ a_3559_n364# a_3421_n364# a_n2593_n461# a_6791_n461# a_3835_n364# a_3065_n461# a_3479_n461#
+ a_3341_n461# a_3755_n461# a_n29_n364# a_n4249_n461# a_n4111_n461# a_n4525_n461#
+ a_n4939_n461# a_n5273_n364# a_n4801_n461# a_5077_n364# a_n305_n364# a_n5687_n364#
+ a_n719_n364# a_5353_n364# a_n5963_n364# a_5767_n364# a_n2237_n364# a_n1075_n461#
+ a_5273_n461# a_n2513_n364# a_2317_n364# a_n581_n364# a_n1489_n461# a_5687_n461#
+ a_n2927_n364# a_n1351_n461# a_n995_n364# a_n1765_n461# a_5963_n461# a_n6043_n461#
+ a_2237_n461# a_n6457_n461# a_2513_n461# a_n6733_n461# a_2593_n364# a_2927_n461#
+ a_n3007_n461# a_n4031_n364# a_n4169_n364# a_29_n461# a_n4445_n364# a_4249_n364#
+ a_4111_n364# a_n4859_n364# a_n3283_n461# a_n4721_n364# a_4525_n364# a_109_n364#
+ a_n3697_n461# a_4169_n461# a_4939_n364# a_4801_n364# a_n1409_n364# a_n3973_n461#
+ a_4031_n461# a_4445_n461# a_305_n461# a_4859_n461# a_4721_n461# a_385_n364# a_719_n461#
+ a_n1271_n364# a_1075_n364# a_799_n364# a_661_n364# a_n5215_n461# a_1409_n461# a_n1685_n364#
+ a_n5629_n461# a_1489_n364# a_1351_n364# a_n6377_n364# a_n1961_n364# a_1765_n364#
+ a_n5905_n461# a_581_n461# a_6043_n364# a_995_n461# a_n6653_n364# a_n247_n461# a_1271_n461#
+ a_6457_n364# a_n5491_n461# a_1685_n461# a_n523_n461# a_6733_n364# a_n3203_n364#
+ a_3007_n364# a_n2179_n461# a_n937_n461# a_1961_n461# a_6377_n461# a_n3617_n364#
+ a_n2041_n461# a_n2455_n461# a_6653_n461# a_n2869_n461# a_n2731_n461# a_3203_n461#
+ a_3283_n364# a_n3893_n364# a_3617_n461# a_3697_n364# a_3973_n364# a_n5135_n364#
+ a_3893_n461# a_n5411_n364# a_n5549_n364# a_5215_n364# a_n4387_n461# a_n5825_n364#
+ w_n6965_n464# a_5629_n364# a_n4663_n461# a_n167_n364# a_5905_n364# a_5135_n461#
+ a_n443_n364# a_5549_n461# a_n1213_n461# a_5411_n461# a_n857_n364# a_n2099_n364#
+ a_5491_n364# a_n1627_n461# a_5825_n461# a_n2375_n364# a_n6319_n461# a_n1903_n461#
+ a_2179_n364# a_2041_n364# a_n2789_n364# a_n2651_n364# a_2455_n364# a_2099_n461#
+ a_2869_n364# a_2731_n364# a_n6181_n461# a_2375_n461# a_n6595_n461# a_2789_n461#
+ a_2651_n461# a_n4307_n364# a_n6871_n461# a_n3145_n461# a_n3559_n461# a_n3421_n461#
+ a_n3835_n461# a_4307_n461# a_4387_n364# a_n4583_n364# a_n4997_n364# a_247_n364#
+ a_4663_n364# a_n1133_n364# a_523_n364# a_n1547_n364# a_937_n364# a_167_n461# a_4583_n461#
+ a_1213_n364# a_n1823_n364# a_1627_n364# a_n6101_n364# a_n6239_n364# a_443_n461#
+ a_4997_n461# a_n5077_n461# a_n6515_n364# a_1903_n364# a_n109_n461# a_857_n461# a_1133_n461#
+ a_6319_n364#
X0 a_2731_n364# a_2651_n461# a_2593_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X1 a_n3755_n364# a_n3835_n461# a_n3893_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X2 a_n6791_n364# a_n6871_n461# a_n6929_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X3 a_n443_n364# a_n523_n461# a_n581_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X4 a_n1409_n364# a_n1489_n461# a_n1547_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X5 a_5629_n364# a_5549_n461# a_5491_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X6 a_3973_n364# a_3893_n461# a_3835_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X7 a_n2927_n364# a_n3007_n461# a_n3065_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X8 a_n5963_n364# a_n6043_n461# a_n6101_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X9 a_937_n364# a_857_n461# a_799_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X10 a_n1271_n364# a_n1351_n461# a_n1409_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X11 a_5491_n364# a_5411_n461# a_5353_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X12 a_n1823_n364# a_n1903_n461# a_n1961_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X13 a_3145_n364# a_3065_n461# a_3007_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X14 a_n4169_n364# a_n4249_n461# a_n4307_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X15 a_3697_n364# a_3617_n461# a_3559_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X16 a_n2513_n364# a_n2593_n461# a_n2651_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X17 a_6733_n364# a_6653_n461# a_6595_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X18 a_2041_n364# a_1961_n461# a_1903_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X19 a_n4031_n364# a_n4111_n461# a_n4169_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X20 a_4939_n364# a_4859_n461# a_4801_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X21 a_1213_n364# a_1133_n461# a_1075_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X22 a_n2237_n364# a_n2317_n461# a_n2375_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X23 a_n5273_n364# a_n5353_n461# a_n5411_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X24 a_4801_n364# a_4721_n461# a_4663_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X25 a_n5825_n364# a_n5905_n461# a_n5963_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X26 a_2455_n364# a_2375_n461# a_2317_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X27 a_n3479_n364# a_n3559_n461# a_n3617_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X28 a_n6515_n364# a_n6595_n461# a_n6653_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X29 a_109_n364# a_29_n461# a_n29_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X30 a_n167_n364# a_n247_n461# a_n305_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X31 a_6043_n364# a_5963_n461# a_5905_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X32 a_3007_n364# a_2927_n461# a_2869_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X33 a_n3341_n364# a_n3421_n461# a_n3479_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X34 a_n995_n364# a_n1075_n461# a_n1133_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X35 a_5215_n364# a_5135_n461# a_5077_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X36 a_n6239_n364# a_n6319_n461# a_n6377_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X37 a_n1547_n364# a_n1627_n461# a_n1685_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X38 a_n4583_n364# a_n4663_n461# a_n4721_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X39 a_523_n364# a_443_n461# a_385_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X40 a_6457_n364# a_6377_n461# a_6319_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X41 a_1765_n364# a_1685_n461# a_1627_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X42 a_n2789_n364# a_n2869_n461# a_n2927_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X43 a_3283_n364# a_3203_n461# a_3145_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X44 a_n2651_n364# a_n2731_n461# a_n2789_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X45 a_n719_n364# a_n799_n461# a_n857_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X46 a_n4997_n364# a_n5077_n461# a_n5135_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X47 a_4525_n364# a_4445_n461# a_4387_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X48 a_1489_n364# a_1409_n461# a_1351_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X49 a_n5549_n364# a_n5629_n461# a_n5687_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X50 a_n3893_n364# a_n3973_n461# a_n4031_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X51 a_2179_n364# a_2099_n461# a_2041_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X52 a_n581_n364# a_n661_n461# a_n719_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X53 a_5767_n364# a_5687_n461# a_5629_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X54 a_n3065_n364# a_n3145_n461# a_n3203_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X55 a_n6101_n364# a_n6181_n461# a_n6239_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X56 a_2593_n364# a_2513_n461# a_2455_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X57 a_1075_n364# a_995_n461# a_937_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X58 a_n6653_n364# a_n6733_n461# a_n6791_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X59 a_n4307_n364# a_n4387_n461# a_n4445_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X60 a_247_n364# a_167_n461# a_109_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X61 a_6871_n364# a_6791_n461# a_6733_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X62 a_3835_n364# a_3755_n461# a_3697_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X63 a_n4859_n364# a_n4939_n461# a_n4997_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X64 a_799_n364# a_719_n461# a_661_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X65 a_n1133_n364# a_n1213_n461# a_n1271_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X66 a_n4721_n364# a_n4801_n461# a_n4859_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X67 a_5077_n364# a_4997_n461# a_4939_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X68 a_1351_n364# a_1271_n461# a_1213_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X69 a_n2375_n364# a_n2455_n461# a_n2513_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X70 a_6595_n364# a_6515_n461# a_6457_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X71 a_n5411_n364# a_n5491_n461# a_n5549_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X72 a_1903_n364# a_1823_n461# a_1765_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X73 a_4249_n364# a_4169_n461# a_4111_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X74 a_n3617_n364# a_n3697_n461# a_n3755_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X75 a_n305_n364# a_n385_n461# a_n443_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X76 a_4111_n364# a_4031_n461# a_3973_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X77 a_n5135_n364# a_n5215_n461# a_n5273_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X78 a_n857_n364# a_n937_n461# a_n995_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X79 a_n6377_n364# a_n6457_n461# a_n6515_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X80 a_5353_n364# a_5273_n461# a_5215_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X81 a_2317_n364# a_2237_n461# a_2179_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X82 a_n29_n364# a_n109_n461# a_n167_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X83 a_n1685_n364# a_n1765_n461# a_n1823_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X84 a_5905_n364# a_5825_n461# a_5767_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X85 a_661_n364# a_581_n461# a_523_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X86 a_3559_n364# a_3479_n461# a_3421_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X87 a_3421_n364# a_3341_n461# a_3283_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X88 a_n4445_n364# a_n4525_n461# a_n4583_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X89 a_385_n364# a_305_n461# a_247_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X90 a_n2099_n364# a_n2179_n461# a_n2237_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X91 a_6319_n364# a_6239_n461# a_6181_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X92 a_1627_n364# a_1547_n461# a_1489_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X93 a_4663_n364# a_4583_n461# a_4525_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X94 a_n5687_n364# a_n5767_n461# a_n5825_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X95 a_n1961_n364# a_n2041_n461# a_n2099_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X96 a_6181_n364# a_6101_n461# a_6043_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X97 a_2869_n364# a_2789_n461# a_2731_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X98 a_n3203_n364# a_n3283_n461# a_n3341_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X99 a_4387_n364# a_4307_n461# a_4249_n364# w_n6965_n464# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_UNVJW6 a_167_n426# a_4583_n426# VSUBS a_443_n426#
+ a_4997_n426# a_n5077_n426# a_n109_n426# a_857_n426# a_1133_n426# a_2593_n400# a_n5353_n426#
+ a_1547_n426# a_n5767_n426# a_1823_n426# a_6239_n426# a_6101_n426# a_n4169_n400#
+ a_n4031_n400# a_n2317_n426# a_n385_n426# a_6515_n426# a_n4445_n400# a_4249_n400#
+ a_n799_n426# a_4111_n400# a_n4859_n400# a_n661_n426# a_109_n400# a_n4721_n400# a_4525_n400#
+ a_4939_n400# a_4801_n400# a_n1409_n400# a_n2593_n426# a_6791_n426# a_3065_n426#
+ a_3479_n426# a_3341_n426# a_385_n400# a_3755_n426# a_1075_n400# a_799_n400# a_n1271_n400#
+ a_661_n400# a_n1685_n400# a_1489_n400# a_n4249_n426# a_1351_n400# a_n4111_n426#
+ a_n6377_n400# a_1765_n400# a_n1961_n400# a_n4525_n426# a_n6653_n400# a_6043_n400#
+ a_n4939_n426# a_6457_n400# a_n4801_n426# a_6733_n400# a_n3203_n400# a_3007_n400#
+ a_n3617_n400# a_n1075_n426# a_5273_n426# a_n1489_n426# a_5687_n426# a_n1351_n426#
+ a_n1765_n426# a_5963_n426# a_3283_n400# a_n6043_n426# a_n3893_n400# a_2237_n426#
+ a_3697_n400# a_n6457_n426# a_2513_n426# a_3973_n400# a_n6733_n426# a_2927_n426#
+ a_n3007_n426# a_n5135_n400# a_n5549_n400# a_n5411_n400# a_5215_n400# a_n5825_n400#
+ a_29_n426# a_5629_n400# a_n3283_n426# a_n167_n400# a_5905_n400# a_n3697_n426# a_n443_n400#
+ a_4169_n426# a_n3973_n426# a_4031_n426# a_5491_n400# a_n857_n400# a_n2099_n400#
+ a_4445_n426# a_n2375_n400# a_305_n426# a_4859_n426# a_2179_n400# a_4721_n426# a_2041_n400#
+ a_n2789_n400# a_719_n426# a_n2651_n400# a_2455_n400# a_n5215_n426# a_1409_n426#
+ a_2869_n400# a_n5629_n426# a_2731_n400# a_n5905_n426# a_581_n426# a_995_n426# a_n247_n426#
+ a_1271_n426# a_n4307_n400# a_n5491_n426# a_1685_n426# a_n523_n426# a_n2179_n426#
+ a_n937_n426# a_1961_n426# a_6377_n426# a_n2041_n426# a_n2455_n426# a_6653_n426#
+ a_n4583_n400# a_n2869_n426# a_4387_n400# a_n2731_n426# a_n4997_n400# a_3203_n426#
+ a_4663_n400# a_247_n400# a_n1133_n400# a_3617_n426# a_523_n400# a_n1547_n400# a_1213_n400#
+ a_937_n400# a_n1823_n400# a_n6239_n400# a_1627_n400# a_n6101_n400# a_n6515_n400#
+ a_1903_n400# a_3893_n426# a_n6929_n400# a_6319_n400# a_n4387_n426# a_n4663_n426#
+ a_6181_n400# w_n6965_n462# a_n6791_n400# a_5135_n426# a_6595_n400# a_n3065_n400#
+ a_5549_n426# a_n1213_n426# a_5411_n426# a_6871_n400# a_n3479_n400# a_n1627_n426#
+ a_n3341_n400# a_5825_n426# a_3145_n400# a_n3755_n400# a_3559_n400# a_n6319_n426#
+ a_n1903_n426# a_3421_n400# a_3835_n400# a_2099_n426# a_n6181_n426# a_2375_n426#
+ a_n29_n400# a_n6595_n426# a_2789_n426# a_2651_n426# a_n6871_n426# a_n3145_n426#
+ a_n5273_n400# a_n3559_n426# a_5077_n400# a_n305_n400# a_n3421_n426# a_n5687_n400#
+ a_n3835_n426# a_5353_n400# a_n719_n400# a_n5963_n400# a_4307_n426# a_5767_n400#
+ a_n2237_n400# a_n2513_n400# a_2317_n400# a_n581_n400# a_n995_n400# a_n2927_n400#
X0 a_3145_n400# a_3065_n426# a_3007_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X1 a_n4169_n400# a_n4249_n426# a_n4307_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X2 a_3697_n400# a_3617_n426# a_3559_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X3 a_n2513_n400# a_n2593_n426# a_n2651_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X4 a_6733_n400# a_6653_n426# a_6595_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X5 a_2041_n400# a_1961_n426# a_1903_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X6 a_n4031_n400# a_n4111_n426# a_n4169_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X7 a_4939_n400# a_4859_n426# a_4801_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X8 a_1213_n400# a_1133_n426# a_1075_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X9 a_n2237_n400# a_n2317_n426# a_n2375_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X10 a_n5273_n400# a_n5353_n426# a_n5411_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X11 a_4801_n400# a_4721_n426# a_4663_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X12 a_n5825_n400# a_n5905_n426# a_n5963_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X13 a_2455_n400# a_2375_n426# a_2317_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X14 a_n3479_n400# a_n3559_n426# a_n3617_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X15 a_n6515_n400# a_n6595_n426# a_n6653_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X16 a_109_n400# a_29_n426# a_n29_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X17 a_n167_n400# a_n247_n426# a_n305_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X18 a_6043_n400# a_5963_n426# a_5905_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X19 a_3007_n400# a_2927_n426# a_2869_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X20 a_n3341_n400# a_n3421_n426# a_n3479_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X21 a_n995_n400# a_n1075_n426# a_n1133_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X22 a_5215_n400# a_5135_n426# a_5077_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X23 a_n6239_n400# a_n6319_n426# a_n6377_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X24 a_n1547_n400# a_n1627_n426# a_n1685_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X25 a_n4583_n400# a_n4663_n426# a_n4721_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X26 a_523_n400# a_443_n426# a_385_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X27 a_6457_n400# a_6377_n426# a_6319_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X28 a_1765_n400# a_1685_n426# a_1627_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X29 a_n2789_n400# a_n2869_n426# a_n2927_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X30 a_3283_n400# a_3203_n426# a_3145_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X31 a_n2651_n400# a_n2731_n426# a_n2789_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X32 a_n719_n400# a_n799_n426# a_n857_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X33 a_n4997_n400# a_n5077_n426# a_n5135_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X34 a_4525_n400# a_4445_n426# a_4387_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X35 a_1489_n400# a_1409_n426# a_1351_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X36 a_n5549_n400# a_n5629_n426# a_n5687_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X37 a_2179_n400# a_2099_n426# a_2041_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X38 a_n3893_n400# a_n3973_n426# a_n4031_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X39 a_n581_n400# a_n661_n426# a_n719_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X40 a_5767_n400# a_5687_n426# a_5629_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X41 a_n3065_n400# a_n3145_n426# a_n3203_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X42 a_n6101_n400# a_n6181_n426# a_n6239_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X43 a_2593_n400# a_2513_n426# a_2455_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X44 a_1075_n400# a_995_n426# a_937_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X45 a_n6653_n400# a_n6733_n426# a_n6791_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X46 a_n4307_n400# a_n4387_n426# a_n4445_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X47 a_247_n400# a_167_n426# a_109_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X48 a_6871_n400# a_6791_n426# a_6733_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X49 a_3835_n400# a_3755_n426# a_3697_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X50 a_n4859_n400# a_n4939_n426# a_n4997_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X51 a_799_n400# a_719_n426# a_661_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X52 a_n1133_n400# a_n1213_n426# a_n1271_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X53 a_n4721_n400# a_n4801_n426# a_n4859_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X54 a_5077_n400# a_4997_n426# a_4939_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X55 a_1351_n400# a_1271_n426# a_1213_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X56 a_6595_n400# a_6515_n426# a_6457_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X57 a_n2375_n400# a_n2455_n426# a_n2513_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X58 a_n5411_n400# a_n5491_n426# a_n5549_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X59 a_1903_n400# a_1823_n426# a_1765_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X60 a_4249_n400# a_4169_n426# a_4111_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X61 a_n3617_n400# a_n3697_n426# a_n3755_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X62 a_n305_n400# a_n385_n426# a_n443_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X63 a_4111_n400# a_4031_n426# a_3973_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X64 a_n5135_n400# a_n5215_n426# a_n5273_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X65 a_n857_n400# a_n937_n426# a_n995_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X66 a_5353_n400# a_5273_n426# a_5215_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X67 a_2317_n400# a_2237_n426# a_2179_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X68 a_n6377_n400# a_n6457_n426# a_n6515_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X69 a_n29_n400# a_n109_n426# a_n167_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X70 a_n1685_n400# a_n1765_n426# a_n1823_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X71 a_5905_n400# a_5825_n426# a_5767_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X72 a_661_n400# a_581_n426# a_523_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X73 a_3559_n400# a_3479_n426# a_3421_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X74 a_3421_n400# a_3341_n426# a_3283_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X75 a_n4445_n400# a_n4525_n426# a_n4583_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X76 a_385_n400# a_305_n426# a_247_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X77 a_n2099_n400# a_n2179_n426# a_n2237_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X78 a_6319_n400# a_6239_n426# a_6181_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X79 a_1627_n400# a_1547_n426# a_1489_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X80 a_4663_n400# a_4583_n426# a_4525_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X81 a_n5687_n400# a_n5767_n426# a_n5825_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X82 a_n1961_n400# a_n2041_n426# a_n2099_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X83 a_6181_n400# a_6101_n426# a_6043_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X84 a_2869_n400# a_2789_n426# a_2731_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X85 a_4387_n400# a_4307_n426# a_4249_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X86 a_n3203_n400# a_n3283_n426# a_n3341_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X87 a_2731_n400# a_2651_n426# a_2593_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X88 a_n3755_n400# a_n3835_n426# a_n3893_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X89 a_n6791_n400# a_n6871_n426# a_n6929_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X90 a_n443_n400# a_n523_n426# a_n581_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X91 a_n1409_n400# a_n1489_n426# a_n1547_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=400000u
X92 a_5629_n400# a_5549_n426# a_5491_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=400000u
X93 a_3973_n400# a_3893_n426# a_3835_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X94 a_n2927_n400# a_n3007_n426# a_n3065_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X95 a_n5963_n400# a_n6043_n426# a_n6101_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X96 a_937_n400# a_857_n426# a_799_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X97 a_n1271_n400# a_n1351_n426# a_n1409_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X98 a_5491_n400# a_5411_n426# a_5353_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X99 a_n1823_n400# a_n1903_n426# a_n1961_n400# w_n6965_n462# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
.ends

.subckt M1_2 VSUBS m1_216_n771# a_143_n3514# w_n944_n1621# a_143_38# a_223_n3417#
Xsky130_fd_pr__pfet_01v8_lvt_SNVJWU_0 a_143_38# w_n944_n1621# VSUBS a_143_38# a_143_38#
+ a_143_38# a_143_38# a_143_38# m1_216_n771# m1_216_n771# a_143_38# a_143_38# a_143_38#
+ w_n944_n1621# w_n944_n1621# a_143_38# m1_216_n771# a_143_38# w_n944_n1621# w_n944_n1621#
+ m1_216_n771# m1_216_n771# w_n944_n1621# m1_216_n771# a_143_38# a_143_38# w_n944_n1621#
+ a_143_38# a_143_38# a_143_38# a_143_38# w_n944_n1621# a_143_38# a_143_38# a_143_38#
+ a_143_38# w_n944_n1621# a_143_38# m1_216_n771# w_n944_n1621# m1_216_n771# m1_216_n771#
+ m1_216_n771# m1_216_n771# w_n944_n1621# w_n944_n1621# a_143_38# a_143_38# w_n944_n1621#
+ m1_216_n771# w_n944_n1621# a_143_38# a_143_38# m1_216_n771# a_143_38# m1_216_n771#
+ a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# m1_216_n771#
+ a_143_38# a_143_38# m1_216_n771# w_n944_n1621# a_143_38# w_n944_n1621# m1_216_n771#
+ w_n944_n1621# m1_216_n771# a_143_38# w_n944_n1621# m1_216_n771# m1_216_n771# a_143_38#
+ a_143_38# w_n944_n1621# m1_216_n771# w_n944_n1621# a_143_38# a_143_38# a_143_38#
+ a_143_38# a_143_38# a_143_38# m1_216_n771# a_143_38# m1_216_n771# w_n944_n1621#
+ w_n944_n1621# m1_216_n771# a_143_38# a_143_38# w_n944_n1621# a_143_38# m1_216_n771#
+ w_n944_n1621# w_n944_n1621# w_n944_n1621# m1_216_n771# a_143_38# a_143_38# w_n944_n1621#
+ a_143_38# w_n944_n1621# a_143_38# a_143_38# m1_216_n771# a_143_38# a_143_38# a_143_38#
+ m1_216_n771# m1_216_n771# w_n944_n1621# a_143_38# a_143_38# a_143_38# a_143_38#
+ w_n944_n1621# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# w_n944_n1621#
+ w_n944_n1621# a_143_38# m1_216_n771# m1_216_n771# m1_216_n771# a_143_38# m1_216_n771#
+ w_n944_n1621# w_n944_n1621# a_143_38# w_n944_n1621# w_n944_n1621# m1_216_n771# a_143_38#
+ m1_216_n771# m1_216_n771# a_143_38# m1_216_n771# a_143_38# a_143_38# a_143_38# w_n944_n1621#
+ m1_216_n771# w_n944_n1621# a_143_38# a_143_38# m1_216_n771# a_143_38# a_143_38#
+ w_n944_n1621# m1_216_n771# w_n944_n1621# m1_216_n771# w_n944_n1621# a_143_38# m1_216_n771#
+ w_n944_n1621# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# m1_216_n771# a_143_38#
+ a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# w_n944_n1621# m1_216_n771# w_n944_n1621#
+ w_n944_n1621# w_n944_n1621# w_n944_n1621# w_n944_n1621# m1_216_n771# m1_216_n771#
+ a_143_38# a_143_38# m1_216_n771# m1_216_n771# w_n944_n1621# w_n944_n1621# m1_216_n771#
+ a_143_38# a_143_38# a_143_38# m1_216_n771# w_n944_n1621# a_143_38# a_143_38# a_143_38#
+ w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt_SNVJWU
Xsky130_fd_pr__pfet_01v8_lvt_UNVJW6_0 a_143_38# a_143_38# VSUBS a_143_38# a_143_38#
+ a_143_38# a_143_38# a_143_38# a_143_38# m1_216_n771# a_143_38# a_143_38# a_143_38#
+ a_143_38# a_143_38# a_143_38# w_n944_n1621# m1_216_n771# a_143_38# a_143_38# a_143_38#
+ w_n944_n1621# m1_216_n771# a_143_38# w_n944_n1621# m1_216_n771# a_143_38# m1_216_n771#
+ w_n944_n1621# m1_216_n771# w_n944_n1621# m1_216_n771# w_n944_n1621# a_143_38# a_143_38#
+ a_143_38# a_143_38# a_143_38# m1_216_n771# a_143_38# w_n944_n1621# w_n944_n1621#
+ m1_216_n771# m1_216_n771# w_n944_n1621# m1_216_n771# a_143_38# w_n944_n1621# a_143_38#
+ w_n944_n1621# m1_216_n771# w_n944_n1621# a_143_38# w_n944_n1621# w_n944_n1621# a_143_38#
+ m1_216_n771# a_143_38# m1_216_n771# m1_216_n771# w_n944_n1621# w_n944_n1621# a_143_38#
+ a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# w_n944_n1621# a_143_38#
+ w_n944_n1621# a_143_38# m1_216_n771# a_143_38# a_143_38# m1_216_n771# a_143_38#
+ a_143_38# a_143_38# m1_216_n771# w_n944_n1621# m1_216_n771# w_n944_n1621# w_n944_n1621#
+ a_143_38# m1_216_n771# a_143_38# m1_216_n771# m1_216_n771# a_143_38# m1_216_n771#
+ a_143_38# a_143_38# a_143_38# w_n944_n1621# w_n944_n1621# m1_216_n771# a_143_38#
+ m1_216_n771# a_143_38# a_143_38# w_n944_n1621# a_143_38# m1_216_n771# w_n944_n1621#
+ a_143_38# m1_216_n771# w_n944_n1621# a_143_38# a_143_38# m1_216_n771# a_143_38#
+ w_n944_n1621# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# m1_216_n771# a_143_38#
+ a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38#
+ a_143_38# m1_216_n771# a_143_38# w_n944_n1621# a_143_38# w_n944_n1621# a_143_38#
+ w_n944_n1621# w_n944_n1621# w_n944_n1621# a_143_38# w_n944_n1621# m1_216_n771# m1_216_n771#
+ m1_216_n771# m1_216_n771# m1_216_n771# w_n944_n1621# w_n944_n1621# m1_216_n771#
+ w_n944_n1621# a_143_38# w_n944_n1621# w_n944_n1621# a_143_38# a_143_38# m1_216_n771#
+ w_n944_n1621# m1_216_n771# a_143_38# w_n944_n1621# w_n944_n1621# a_143_38# a_143_38#
+ a_143_38# w_n944_n1621# m1_216_n771# a_143_38# w_n944_n1621# a_143_38# m1_216_n771#
+ m1_216_n771# w_n944_n1621# a_143_38# a_143_38# m1_216_n771# w_n944_n1621# a_143_38#
+ a_143_38# a_143_38# w_n944_n1621# a_143_38# a_143_38# a_143_38# a_143_38# a_143_38#
+ w_n944_n1621# a_143_38# m1_216_n771# w_n944_n1621# a_143_38# m1_216_n771# a_143_38#
+ m1_216_n771# m1_216_n771# m1_216_n771# a_143_38# w_n944_n1621# w_n944_n1621# w_n944_n1621#
+ m1_216_n771# w_n944_n1621# m1_216_n771# m1_216_n771# sky130_fd_pr__pfet_01v8_lvt_UNVJW6
X0 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=1.16e+14p pd=8.58e+08u as=2.3664e+14p ps=1.75032e+09u w=4e+06u l=400000u
X1 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X2 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X3 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X4 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X5 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X6 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X7 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X8 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X9 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X10 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X11 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X12 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X13 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X14 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X15 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X16 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X17 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X18 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X19 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X20 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X21 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X22 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X23 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X24 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X25 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X26 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X27 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X28 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X29 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X30 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X31 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X32 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X33 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X34 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X35 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X36 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X37 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X38 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X39 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X40 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X41 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X42 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X43 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X44 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X45 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X46 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X47 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X48 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X49 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X50 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X51 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X52 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X53 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X54 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X55 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X56 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X57 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X58 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X59 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X60 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X61 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X62 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X63 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X64 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X65 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X66 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X67 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X68 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X69 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X70 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X71 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X72 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X73 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X74 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X75 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X76 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X77 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X78 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X79 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X80 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X81 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X82 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X83 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X84 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X85 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X86 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X87 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X88 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X89 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X90 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X91 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X92 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X93 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X94 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X95 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X96 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X97 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X98 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X99 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X100 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X101 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X102 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X103 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X104 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X105 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X106 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X107 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X108 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X109 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X110 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X111 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X112 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X113 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X114 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X115 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X116 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X117 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X118 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X119 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X120 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X121 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X122 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X123 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X124 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X125 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X126 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X127 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X128 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X129 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X130 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X131 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X132 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X133 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X134 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X135 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X136 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X137 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X138 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X139 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X140 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X141 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X142 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X143 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X144 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X145 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X146 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X147 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X148 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X149 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X150 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X151 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X152 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X153 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X154 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X155 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X156 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X157 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X158 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X159 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X160 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X161 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X162 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X163 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X164 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X165 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X166 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X167 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X168 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X169 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X170 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X171 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X172 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X173 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X174 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X175 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X176 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X177 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X178 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X179 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X180 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X181 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X182 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X183 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X184 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X185 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X186 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X187 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X188 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X189 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X190 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X191 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X192 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X193 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X194 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X195 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X196 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X197 w_n944_n1621# a_143_n3514# a_223_n3417# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X198 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
X199 a_223_n3417# a_143_n3514# w_n944_n1621# w_n944_n1621# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=400000u
.ends

.subckt opamp_lucas m2_932_n12357# vin_n vin_p iref vout vss vdd
XM5_B_0 vss vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ vdd vdd vdd vdd iref m2_932_n12357# vdd vdd vdd M5_B
XM3_0 vss m1_5767_n19817# vss vss vss M3
Xsky130_fd_pr__cap_mim_m3_1_2674SJ_0 vss vout m2_17170_n15338# sky130_fd_pr__cap_mim_m3_1_2674SJ
Xsky130_fd_pr__cap_mim_m3_1_2674SJ_1 vss vout m2_17170_n15338# sky130_fd_pr__cap_mim_m3_1_2674SJ
Xsky130_fd_pr__cap_mim_m3_1_2674SJ_2 vss vout m2_17170_n15338# sky130_fd_pr__cap_mim_m3_1_2674SJ
Xsky130_fd_pr__cap_mim_m3_1_2674SJ_3 vss vout m2_17170_n15338# sky130_fd_pr__cap_mim_m3_1_2674SJ
XM8_0 vss vdd vdd vdd vdd vdd vdd vdd iref M8
XM6_0 vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss
+ vss vss vss vss m1_18001_n16633# vss vss vss vss vss vss vss vss vss vss vss vss
+ vss vout vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss vss M6
XM4_0 vss vss m1_5767_n19817# vss vss m1_18001_n16633# M4
XM9_0 vdd m2_17170_n15338# m1_18001_n16633# vss M9
XM7_0 vss vdd vout iref vout vout vdd M7
XM1_2_0 vss m1_5767_n19817# vin_p m2_932_n12357# vin_n m1_18001_n16633# M1_2
.ends

.subckt sky130_fd_pr__nfet_01v8_Z2S3N8 w_n4967_n360# a_2079_n150# a_2463_n150# a_3423_n150#
+ a_n801_n150# a_n417_n150# a_351_n150# a_4383_n150# a_n4449_n150# a_n2913_n150# a_n2529_n150#
+ a_n1569_n150# a_n3873_n150# a_n3489_n150# a_n1953_n150# a_3615_n150# a_n609_n150#
+ a_159_n150# a_543_n150# a_1695_n150# a_2655_n150# a_4575_n150# a_n993_n150# a_2847_n150#
+ a_3807_n150# a_n33_n150# a_735_n150# a_1887_n150# a_4767_n150# a_n4767_n176# a_n3105_n150#
+ a_n4065_n150# a_n2145_n150# a_n1185_n150# a_927_n150# a_1311_n150# a_2271_n150#
+ a_3231_n150# a_3999_n150# a_n225_n150# a_4191_n150# a_n4829_n150# a_n2337_n150#
+ a_n4641_n150# a_n4257_n150# a_n3681_n150# a_n3297_n150# a_n2721_n150# a_n1761_n150#
+ a_n1377_n150# a_1119_n150# a_1503_n150# a_3039_n150#
X0 a_n225_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=2.475e+13p ps=1.83e+08u w=1.5e+06u l=150000u
X1 a_2271_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X2 w_n4967_n360# a_n4767_n176# a_3423_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X3 w_n4967_n360# a_n4767_n176# a_3039_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X4 a_351_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X5 a_n4257_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X6 w_n4967_n360# a_n4767_n176# a_n609_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X7 a_n1569_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_3807_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 w_n4967_n360# a_n4767_n176# a_927_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X10 a_n1185_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X11 w_n4967_n360# a_n4767_n176# a_n4641_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X12 a_n801_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X13 w_n4967_n360# a_n4767_n176# a_n1953_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X14 w_n4967_n360# a_n4767_n176# a_n1569_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X15 w_n4967_n360# a_n4767_n176# a_3231_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X16 a_n4065_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X17 w_n4967_n360# a_n4767_n176# a_n417_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X18 w_n4967_n360# a_n4767_n176# a_n33_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X19 a_3615_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X20 a_n993_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X21 a_3231_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X22 w_n4967_n360# a_n4767_n176# a_n4449_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X23 w_n4967_n360# a_n4767_n176# a_4383_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X24 w_n4967_n360# a_n4767_n176# a_n1761_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X25 w_n4967_n360# a_n4767_n176# a_3807_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X26 w_n4967_n360# a_n4767_n176# a_n1377_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X27 a_n2529_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X28 a_n4641_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X29 a_4767_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.65e+11p pd=3.62e+06u as=0p ps=0u w=1.5e+06u l=150000u
X30 a_n1953_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X31 a_3423_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X32 a_n33_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X33 w_n4967_n360# a_n4767_n176# a_n2913_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X34 w_n4967_n360# a_n4767_n176# a_n2145_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X35 w_n4967_n360# a_n4767_n176# a_n4257_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 w_n4967_n360# a_n4767_n176# a_4191_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X37 w_n4967_n360# a_n4767_n176# a_1503_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X38 w_n4967_n360# a_n4767_n176# a_3615_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X39 a_n2337_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X40 a_4575_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X41 a_n1761_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X42 a_1887_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X43 a_1119_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X44 w_n4967_n360# a_n4767_n176# a_n2721_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X45 w_n4967_n360# a_n4767_n176# a_3999_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X46 a_n3489_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X47 w_n4967_n360# a_n4767_n176# a_1311_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X48 a_n2913_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X49 a_n2145_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X50 a_4383_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X51 w_n4967_n360# a_n4767_n176# a_n3873_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X52 w_n4967_n360# a_n4767_n176# a_n3105_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X53 a_1695_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X54 w_n4967_n360# a_n4767_n176# a_n2529_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 w_n4967_n360# a_n4767_n176# a_4575_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X56 w_n4967_n360# a_n4767_n176# a_2463_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X57 a_n3297_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X58 w_n4967_n360# a_n4767_n176# a_1887_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X59 w_n4967_n360# a_n4767_n176# a_543_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X60 w_n4967_n360# a_n4767_n176# a_1119_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X61 a_n2721_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X62 a_2847_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X63 a_2079_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X64 w_n4967_n360# a_n4767_n176# a_n4065_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X65 a_4191_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X66 w_n4967_n360# a_n4767_n176# a_n3681_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X67 a_1503_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X68 a_159_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X69 w_n4967_n360# a_n4767_n176# a_n2337_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X70 w_n4967_n360# a_n4767_n176# a_2271_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X71 a_n3873_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X72 a_n3105_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X73 w_n4967_n360# a_n4767_n176# a_1695_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X74 w_n4967_n360# a_n4767_n176# a_351_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X75 a_n609_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X76 a_2655_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X77 w_n4967_n360# a_n4767_n176# a_n3489_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X78 a_735_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X79 a_1311_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X80 w_n4967_n360# a_n4767_n176# a_n993_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X81 w_n4967_n360# a_n4767_n176# a_2847_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X82 w_n4967_n360# a_n4767_n176# a_n225_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X83 w_n4967_n360# a_n4767_n176# a_2079_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X84 a_n3681_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X85 a_3039_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X86 w_n4967_n360# a_n4767_n176# a_159_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 a_n417_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X88 a_2463_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X89 a_927_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X90 w_n4967_n360# a_n4767_n176# a_n1185_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X91 w_n4967_n360# a_n4767_n176# a_n3297_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X92 a_543_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X93 a_n4449_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X94 w_n4967_n360# a_n4767_n176# a_n801_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X95 w_n4967_n360# a_n4767_n176# a_2655_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X96 a_3999_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X97 a_n1377_n150# a_n4767_n176# w_n4967_n360# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X98 w_n4967_n360# a_n4767_n176# a_735_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X99 w_n4967_n360# a_n4767_n176# a_n4829_n150# w_n4967_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.65e+11p ps=3.62e+06u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_J9MTE9 a_n417_n150# a_351_n150# a_255_n150# a_n609_n150#
+ a_159_n150# a_543_n150# a_n701_n150# a_447_n150# w_n839_n360# a_n639_n178# a_n33_n150#
+ a_639_n150# a_n321_n150# a_n225_n150# a_63_n150# a_n513_n150# a_n129_n150#
X0 a_n225_n150# a_n639_n178# a_n321_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X1 a_351_n150# a_n639_n178# a_255_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X2 a_n513_n150# a_n639_n178# a_n609_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X3 a_n321_n150# a_n639_n178# a_n417_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X4 a_63_n150# a_n639_n178# a_n33_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X5 a_n33_n150# a_n639_n178# a_n129_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X6 a_639_n150# a_n639_n178# a_543_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.65e+11p pd=3.62e+06u as=4.95e+11p ps=3.66e+06u w=1.5e+06u l=150000u
X7 a_159_n150# a_n639_n178# a_63_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X8 a_447_n150# a_n639_n178# a_351_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=4.95e+11p pd=3.66e+06u as=0p ps=0u w=1.5e+06u l=150000u
X9 a_n609_n150# a_n639_n178# a_n701_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.65e+11p ps=3.62e+06u w=1.5e+06u l=150000u
X10 a_n129_n150# a_n639_n178# a_n225_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X11 a_255_n150# a_n639_n178# a_159_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X12 a_n417_n150# a_n639_n178# a_n513_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X13 a_543_n150# a_n639_n178# a_447_n150# w_n839_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_H98ZZM VSUBS a_1859_n189# a_n1209_n189# a_n2507_n189#
+ a_1505_n189# a_2803_n189# a_1088_n286# a_n1744_n286# a_2386_n286# a_n973_n189# a_2032_n286#
+ a_n2153_n189# a_1151_n189# a_734_n286# a_89_n189# a_n1390_n286# a_n446_n286# a_380_n286#
+ a_n92_n286# a_2858_n286# a_n2979_n189# a_1977_n189# a_1206_n286# a_n1327_n189# a_n2625_n189#
+ a_2504_n286# a_1623_n189# a_2921_n189# a_n1862_n286# a_n29_n189# a_2150_n286# a_n918_n286#
+ a_n2271_n189# a_852_n286# a_n2098_n286# a_207_n189# a_n564_n286# a_n210_n286# a_1678_n286#
+ a_n1799_n189# a_1324_n286# a_n1445_n189# a_n2743_n189# a_2622_n286# a_1741_n189#
+ a_n1980_n286# a_n1091_n189# a_n2216_n286# a_970_n286# a_n147_n189# a_679_n189# a_325_n189#
+ a_n1917_n189# a_n682_n286# a_1796_n286# a_1442_n286# a_n1563_n189# a_n2861_n189#
+ a_2740_n286# a_2449_n189# a_n619_n189# a_26_n286# a_n2688_n286# a_n1036_n286# a_n2334_n286#
+ a_2095_n189# a_n265_n189# a_n800_n286# a_797_n189# a_443_n189# a_1914_n286# a_1560_n286#
+ a_n1681_n189# a_n1508_n286# a_n2806_n286# a_1269_n189# a_2567_n189# a_n737_n189#
+ a_2213_n189# a_915_n189# a_n2452_n286# a_n1154_n286# a_n383_n189# a_498_n286# w_n3117_n409#
+ a_144_n286# a_561_n189# a_n1626_n286# a_n2924_n286# a_n2389_n189# a_2268_n286# a_1387_n189#
+ a_2685_n189# a_n855_n189# a_n2035_n189# a_616_n286# a_2331_n189# a_1033_n189# a_n501_n189#
+ a_n2570_n286# a_n1272_n286# a_n328_n286# a_262_n286#
X0 a_89_n189# a_26_n286# a_n29_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X1 a_n2035_n189# a_n2098_n286# a_n2153_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X2 a_n2625_n189# a_n2688_n286# a_n2743_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X3 a_2449_n189# a_2386_n286# a_2331_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X4 a_n2507_n189# a_n2570_n286# a_n2625_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X5 a_n501_n189# a_n564_n286# a_n619_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X6 a_n2389_n189# a_n2452_n286# a_n2507_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X7 a_n383_n189# a_n446_n286# a_n501_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X8 a_n265_n189# a_n328_n286# a_n383_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X9 a_n855_n189# a_n918_n286# a_n973_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X10 a_n147_n189# a_n210_n286# a_n265_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X11 a_1151_n189# a_1088_n286# a_1033_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X12 a_1741_n189# a_1678_n286# a_1623_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X13 a_n1091_n189# a_n1154_n286# a_n1209_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X14 a_561_n189# a_498_n286# a_443_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X15 a_1623_n189# a_1560_n286# a_1505_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X16 a_n1681_n189# a_n1744_n286# a_n1799_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X17 a_n973_n189# a_n1036_n286# a_n1091_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X18 a_1505_n189# a_1442_n286# a_1387_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X19 a_n1563_n189# a_n1626_n286# a_n1681_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X20 a_1387_n189# a_1324_n286# a_1269_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X21 a_n1445_n189# a_n1508_n286# a_n1563_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X22 a_1977_n189# a_1914_n286# a_1859_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X23 a_1269_n189# a_1206_n286# a_1151_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X24 a_n737_n189# a_n800_n286# a_n855_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X25 a_n619_n189# a_n682_n286# a_n737_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X26 a_2331_n189# a_2268_n286# a_2213_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X27 a_443_n189# a_380_n286# a_325_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X28 a_1033_n189# a_970_n286# a_915_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X29 a_2921_n189# a_2858_n286# a_2803_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X30 a_325_n189# a_262_n286# a_207_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X31 a_2213_n189# a_2150_n286# a_2095_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X32 a_n2271_n189# a_n2334_n286# a_n2389_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X33 a_915_n189# a_852_n286# a_797_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X34 a_2803_n189# a_2740_n286# a_2685_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X35 a_n2861_n189# a_n2924_n286# a_n2979_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X36 a_207_n189# a_144_n286# a_89_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X37 a_1859_n189# a_1796_n286# a_1741_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X38 a_2095_n189# a_2032_n286# a_1977_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X39 a_2685_n189# a_2622_n286# a_2567_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X40 a_n2743_n189# a_n2806_n286# a_n2861_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X41 a_n2153_n189# a_n2216_n286# a_n2271_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X42 a_n1917_n189# a_n1980_n286# a_n2035_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X43 a_n1327_n189# a_n1390_n286# a_n1445_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=6.525e+11p pd=5.08e+06u as=0p ps=0u w=2.25e+06u l=300000u
X44 a_n29_n189# a_n92_n286# a_n147_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X45 a_797_n189# a_734_n286# a_679_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.525e+11p ps=5.08e+06u w=2.25e+06u l=300000u
X46 a_n1209_n189# a_n1272_n286# a_n1327_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X47 a_679_n189# a_616_n286# a_561_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X48 a_2567_n189# a_2504_n286# a_2449_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
X49 a_n1799_n189# a_n1862_n286# a_n1917_n189# w_n3117_n409# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.25e+06u l=300000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_7XCYSC VSUBS a_641_n736# a_2843_n762# a_1177_n736#
+ a_163_n762# a_3111_n762# a_n1771_n736# a_n3321_n762# a_n105_n762# a_699_n762# a_n2575_n736#
+ a_1771_n762# a_n1981_n762# a_n3379_n736# a_2575_n762# a_373_n736# a_909_n736# a_3321_n736#
+ a_n2785_n762# a_n1503_n736# a_n3053_n762# a_n2307_n736# a_1503_n762# a_1981_n736#
+ a_n1713_n762# a_2307_n762# a_105_n736# a_2785_n736# a_n2517_n762# a_3053_n736# a_n1235_n736#
+ a_n431_n736# a_n2039_n736# a_n967_n736# a_1713_n736# a_1235_n762# a_2517_n736# a_n1445_n762#
+ a_n641_n762# a_2039_n762# a_n2249_n762# a_n163_n736# a_n699_n736# a_431_n762# a_1445_n736#
+ w_n3517_n884# a_n1177_n762# a_967_n762# a_2249_n736# a_n909_n762# a_n373_n762# a_n2843_n736#
+ a_n3111_n736#
X0 a_n699_n736# a_n909_n762# a_n967_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X1 a_641_n736# a_431_n762# a_373_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X2 a_n2575_n736# a_n2785_n762# a_n2843_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X3 a_105_n736# a_n105_n762# a_n163_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X4 a_1445_n736# a_1235_n762# a_1177_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X5 a_1713_n736# a_1503_n762# a_1445_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X6 a_n163_n736# a_n373_n762# a_n431_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X7 a_n967_n736# a_n1177_n762# a_n1235_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X8 a_3321_n736# a_3111_n762# a_3053_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X9 a_n1235_n736# a_n1445_n762# a_n1503_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X10 a_n431_n736# a_n641_n762# a_n699_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X11 a_n2843_n736# a_n3053_n762# a_n3111_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X12 a_n1503_n736# a_n1713_n762# a_n1771_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X13 a_2249_n736# a_2039_n762# a_1981_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X14 a_1981_n736# a_1771_n762# a_1713_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X15 a_n3111_n736# a_n3321_n762# a_n3379_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X16 a_2517_n736# a_2307_n762# a_2249_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X17 a_n2039_n736# a_n2249_n762# a_n2307_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X18 a_909_n736# a_699_n762# a_641_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X19 a_n1771_n736# a_n1981_n762# a_n2039_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X20 a_n2307_n736# a_n2517_n762# a_n2575_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X21 a_1177_n736# a_967_n762# a_909_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X22 a_2785_n736# a_2575_n762# a_2517_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X23 a_373_n736# a_163_n762# a_105_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X24 a_3053_n736# a_2843_n762# a_2785_n736# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_QVUSYJ a_n1562_n1081# a_n2380_n1107# a_2380_n1081#
+ a_n628_n1107# a_1562_n1107# a_628_n1081# a_n248_n1081# a_n190_n1107# a_248_n1107#
+ w_n2576_n1229# a_n1504_n1107# a_n2000_n1081# a_190_n1081# a_1504_n1081# a_2000_n1107#
+ a_n1124_n1081# a_n686_n1081# a_1124_n1107# a_n1066_n1107# a_1066_n1081# a_n1942_n1107#
+ a_686_n1107# a_n2438_n1081# a_1942_n1081#
X0 a_n1562_n1081# a_n1942_n1107# a_n2000_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X1 a_n248_n1081# a_n628_n1107# a_n686_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X2 a_628_n1081# a_248_n1107# a_190_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X3 a_n686_n1081# a_n1066_n1107# a_n1124_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X4 a_1504_n1081# a_1124_n1107# a_1066_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X5 a_1066_n1081# a_686_n1107# a_628_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=1.9e+06u
X6 a_2380_n1081# a_2000_n1107# a_1942_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
X7 a_190_n1081# a_n190_n1107# a_n248_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=1.9e+06u
X8 a_1942_n1081# a_1562_n1107# a_1504_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=1.9e+06u
X9 a_n1124_n1081# a_n1504_n1107# a_n1562_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=1.9e+06u
X10 a_n2000_n1081# a_n2380_n1107# a_n2438_n1081# w_n2576_n1229# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=1.9e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_K4PBSX a_26_295# VSUBS a_n1563_n336# a_n2861_n336#
+ a_n2924_295# a_n1036_295# a_2449_n336# a_n619_n336# a_1324_295# a_n2688_295# a_1088_295#
+ a_2095_n336# a_n265_n336# a_797_n336# a_443_n336# a_n1626_295# a_n92_295# a_1914_295#
+ a_1678_295# a_n1681_n336# a_616_295# a_1269_n336# a_n328_295# a_n1390_295# a_n2216_295#
+ a_2567_n336# a_n737_n336# a_2504_295# a_2213_n336# a_2268_295# a_915_n336# a_n383_n336#
+ a_380_295# a_561_n336# a_n2806_295# a_n918_295# a_n1980_295# a_1206_295# a_2858_295#
+ a_n2389_n336# a_n2570_295# a_1387_n336# a_970_295# a_n682_295# a_2685_n336# a_n855_n336#
+ a_n2035_n336# a_2331_n336# a_1033_n336# a_n501_n336# a_n1508_295# a_n1272_295# a_1859_n336#
+ a_1560_295# a_n1209_n336# a_n2507_n336# a_1505_n336# a_2803_n336# a_n210_295# a_262_295#
+ a_n973_n336# a_2150_295# a_n2153_n336# a_1151_n336# w_n3117_n484# a_n1862_295# a_89_n336#
+ a_n800_295# a_n2452_295# a_852_295# a_n564_295# a_n2979_n336# a_1977_n336# a_2740_295#
+ a_n1327_n336# a_n2625_n336# a_1623_n336# a_2921_n336# a_n29_n336# a_n2271_n336#
+ a_n1154_295# a_1442_295# a_207_n336# a_n1799_n336# a_144_295# a_2032_295# a_n1445_n336#
+ a_n2743_n336# a_1741_n336# a_n1744_295# a_1796_295# a_n1091_n336# a_n147_n336# a_734_295#
+ a_n2334_295# a_n446_295# a_679_n336# a_2622_295# a_498_295# a_n2098_295# a_325_n336#
+ a_n1917_n336# a_2386_295#
X0 a_n2743_n336# a_n2806_295# a_n2861_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X1 a_n2153_n336# a_n2216_295# a_n2271_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X2 a_n1917_n336# a_n1980_295# a_n2035_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X3 a_n1327_n336# a_n1390_295# a_n1445_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X4 a_n29_n336# a_n92_295# a_n147_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X5 a_797_n336# a_734_295# a_679_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X6 a_n1209_n336# a_n1272_295# a_n1327_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X7 a_679_n336# a_616_295# a_561_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X8 a_2567_n336# a_2504_295# a_2449_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X9 a_n1799_n336# a_n1862_295# a_n1917_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X10 a_89_n336# a_26_295# a_n29_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X11 a_n2035_n336# a_n2098_295# a_n2153_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X12 a_n2625_n336# a_n2688_295# a_n2743_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X13 a_2449_n336# a_2386_295# a_2331_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X14 a_n2507_n336# a_n2570_295# a_n2625_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X15 a_n501_n336# a_n564_295# a_n619_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X16 a_n2389_n336# a_n2452_295# a_n2507_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X17 a_n383_n336# a_n446_295# a_n501_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X18 a_n855_n336# a_n918_295# a_n973_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X19 a_n265_n336# a_n328_295# a_n383_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X20 a_n147_n336# a_n210_295# a_n265_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X21 a_1151_n336# a_1088_295# a_1033_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X22 a_1741_n336# a_1678_295# a_1623_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X23 a_n1091_n336# a_n1154_295# a_n1209_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X24 a_561_n336# a_498_295# a_443_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X25 a_1623_n336# a_1560_295# a_1505_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X26 a_n1681_n336# a_n1744_295# a_n1799_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X27 a_n973_n336# a_n1036_295# a_n1091_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X28 a_1505_n336# a_1442_295# a_1387_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X29 a_n1563_n336# a_n1626_295# a_n1681_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X30 a_1387_n336# a_1324_295# a_1269_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X31 a_n1445_n336# a_n1508_295# a_n1563_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X32 a_1977_n336# a_1914_295# a_1859_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X33 a_1269_n336# a_1206_295# a_1151_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X34 a_n737_n336# a_n800_295# a_n855_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X35 a_n619_n336# a_n682_295# a_n737_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X36 a_2331_n336# a_2268_295# a_2213_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X37 a_443_n336# a_380_295# a_325_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X38 a_1033_n336# a_970_295# a_915_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X39 a_2921_n336# a_2858_295# a_2803_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X40 a_325_n336# a_262_295# a_207_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X41 a_2213_n336# a_2150_295# a_2095_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X42 a_n2271_n336# a_n2334_295# a_n2389_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X43 a_915_n336# a_852_295# a_797_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X44 a_2803_n336# a_2740_295# a_2685_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X45 a_n2861_n336# a_n2924_295# a_n2979_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X46 a_207_n336# a_144_295# a_89_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X47 a_1859_n336# a_1796_295# a_1741_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X48 a_2095_n336# a_2032_295# a_1977_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X49 a_2685_n336# a_2622_295# a_2567_n336# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__pfet_01v8_698KZZ VSUBS a_n387_n211# a_n33_n211# a_n859_n211#
+ a_793_n211# a_n505_n211# a_n151_n211# a_148_n114# a_n88_n114# a_n623_n211# a_266_n114#
+ a_n206_n114# a_30_n114# a_738_n114# a_n741_n211# a_384_n114# a_n678_n114# a_85_n211#
+ a_439_n211# a_n324_n114# a_856_n114# a_502_n114# w_n1052_n334# a_557_n211# a_n796_n114#
+ a_n442_n114# a_203_n211# a_620_n114# a_n269_n211# a_n914_n114# a_321_n211# a_675_n211#
+ a_n560_n114#
X0 a_n324_n114# a_n387_n211# a_n442_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X1 a_n796_n114# a_n859_n211# a_n914_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X2 a_n206_n114# a_n269_n211# a_n324_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=300000u
X3 a_n678_n114# a_n741_n211# a_n796_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=300000u
X4 a_n88_n114# a_n151_n211# a_n206_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=300000u
X5 a_620_n114# a_557_n211# a_502_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X6 a_n560_n114# a_n623_n211# a_n678_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=300000u
X7 a_502_n114# a_439_n211# a_384_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X8 a_384_n114# a_321_n211# a_266_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X9 a_266_n114# a_203_n211# a_148_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X10 a_30_n114# a_n33_n211# a_n88_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=300000u
X11 a_856_n114# a_793_n211# a_738_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=300000u
X12 a_738_n114# a_675_n211# a_620_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=300000u
X13 a_n442_n114# a_n505_n211# a_n560_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=300000u
X14 a_148_n114# a_85_n211# a_30_n114# w_n1052_n334# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=300000u
.ends

.subckt sky130_fd_pr__pfet_01v8_65PBSZ a_970_n361# a_n2216_n361# VSUBS a_n147_n264#
+ a_679_n264# a_325_n264# a_n1917_n264# a_n682_n361# a_1796_n361# a_n1563_n264# a_2740_n361#
+ a_1442_n361# a_n2861_n264# a_2449_n264# a_n619_n264# a_n2688_n361# a_26_n361# a_n1036_n361#
+ a_n2334_n361# a_n800_n361# a_2095_n264# a_n265_n264# a_797_n264# a_1914_n361# a_443_n264#
+ a_n1681_n264# a_1560_n361# a_n2806_n361# a_n1508_n361# a_2567_n264# a_1269_n264#
+ a_n737_n264# a_2213_n264# a_915_n264# a_n1154_n361# a_n2452_n361# a_498_n361# a_n383_n264#
+ a_144_n361# a_561_n264# a_n2924_n361# a_2268_n361# a_n1626_n361# a_n2389_n264# a_2685_n264#
+ a_1387_n264# a_n855_n264# a_n2035_n264# a_1033_n264# a_616_n361# a_2331_n264# a_n501_n264#
+ a_n1272_n361# a_n2570_n361# a_n328_n361# a_262_n361# a_1859_n264# a_n1209_n264#
+ w_n3117_n484# a_n2507_n264# a_2803_n264# a_1505_n264# a_2386_n361# a_1088_n361#
+ a_n1744_n361# a_n973_n264# a_n2153_n264# a_2032_n361# a_1151_n264# a_734_n361# a_n1390_n361#
+ a_89_n264# a_n446_n361# a_380_n361# a_n92_n361# a_2858_n361# a_n2979_n264# a_1977_n264#
+ a_n1327_n264# a_2504_n361# a_1206_n361# a_n2625_n264# a_2921_n264# a_1623_n264#
+ a_n1862_n361# a_n29_n264# a_n2271_n264# a_2150_n361# a_n918_n361# a_852_n361# a_207_n264#
+ a_n2098_n361# a_n564_n361# a_n210_n361# a_1678_n361# a_n1799_n264# a_n1445_n264#
+ a_2622_n361# a_1324_n361# a_n2743_n264# a_1741_n264# a_n1980_n361# a_n1091_n264#
X0 a_n265_n264# a_n328_n361# a_n383_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X1 a_n855_n264# a_n918_n361# a_n973_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X2 a_1151_n264# a_1088_n361# a_1033_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X3 a_n147_n264# a_n210_n361# a_n265_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X4 a_1741_n264# a_1678_n361# a_1623_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X5 a_n1091_n264# a_n1154_n361# a_n1209_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X6 a_561_n264# a_498_n361# a_443_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X7 a_1623_n264# a_1560_n361# a_1505_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X8 a_n1681_n264# a_n1744_n361# a_n1799_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X9 a_1505_n264# a_1442_n361# a_1387_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X10 a_n1563_n264# a_n1626_n361# a_n1681_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X11 a_n973_n264# a_n1036_n361# a_n1091_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X12 a_1387_n264# a_1324_n361# a_1269_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X13 a_1977_n264# a_1914_n361# a_1859_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X14 a_n1445_n264# a_n1508_n361# a_n1563_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X15 a_1269_n264# a_1206_n361# a_1151_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X16 a_n737_n264# a_n800_n361# a_n855_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X17 a_n619_n264# a_n682_n361# a_n737_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X18 a_443_n264# a_380_n361# a_325_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X19 a_2331_n264# a_2268_n361# a_2213_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X20 a_1033_n264# a_970_n361# a_915_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X21 a_2921_n264# a_2858_n361# a_2803_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X22 a_325_n264# a_262_n361# a_207_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X23 a_2213_n264# a_2150_n361# a_2095_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X24 a_2803_n264# a_2740_n361# a_2685_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X25 a_n2861_n264# a_n2924_n361# a_n2979_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X26 a_n2271_n264# a_n2334_n361# a_n2389_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X27 a_915_n264# a_852_n361# a_797_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X28 a_n1327_n264# a_n1390_n361# a_n1445_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X29 a_207_n264# a_144_n361# a_89_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X30 a_797_n264# a_734_n361# a_679_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X31 a_1859_n264# a_1796_n361# a_1741_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X32 a_2095_n264# a_2032_n361# a_1977_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X33 a_2685_n264# a_2622_n361# a_2567_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X34 a_n2743_n264# a_n2806_n361# a_n2861_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X35 a_n2153_n264# a_n2216_n361# a_n2271_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X36 a_n1917_n264# a_n1980_n361# a_n2035_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X37 a_n29_n264# a_n92_n361# a_n147_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X38 a_n1209_n264# a_n1272_n361# a_n1327_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X39 a_679_n264# a_616_n361# a_561_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X40 a_2567_n264# a_2504_n361# a_2449_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=300000u
X41 a_n1799_n264# a_n1862_n361# a_n1917_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X42 a_89_n264# a_26_n361# a_n29_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X43 a_n2625_n264# a_n2688_n361# a_n2743_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X44 a_n2035_n264# a_n2098_n361# a_n2153_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X45 a_2449_n264# a_2386_n361# a_2331_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X46 a_n2507_n264# a_n2570_n361# a_n2625_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X47 a_n501_n264# a_n564_n361# a_n619_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=300000u
X48 a_n383_n264# a_n446_n361# a_n501_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
X49 a_n2389_n264# a_n2452_n361# a_n2507_n264# w_n3117_n484# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=300000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_XFP5BZ VSUBS m3_n3150_n2850# c1_n3050_n2750#
X0 c1_n3050_n2750# m3_n3150_n2850# sky130_fd_pr__cap_mim_m3_1 l=2.75e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_RTJWSN VSUBS a_2249_n664# a_n2843_n664# a_n3111_n664#
+ a_163_n761# a_2843_n761# a_3111_n761# a_641_n664# a_n3321_n761# a_n105_n761# a_699_n761#
+ a_1177_n664# a_n1771_n664# a_1771_n761# a_n2575_n664# a_n1981_n761# a_2575_n761#
+ a_n2785_n761# a_n3379_n664# a_373_n664# a_909_n664# a_3321_n664# a_n3053_n761# a_n1503_n664#
+ a_1503_n761# a_n2307_n664# a_n1713_n761# a_2307_n761# a_1981_n664# a_n2517_n761#
+ a_105_n664# a_2785_n664# a_3053_n664# a_n1235_n664# a_n431_n664# a_n967_n664# a_n1445_n761#
+ a_1235_n761# a_n2039_n664# a_1713_n664# a_n641_n761# a_2039_n761# a_2517_n664# a_n2249_n761#
+ a_431_n761# a_n163_n664# w_n3517_n884# a_967_n761# a_n699_n664# a_1445_n664# a_n1177_n761#
+ a_n909_n761# a_n373_n761#
X0 a_n2307_n664# a_n2517_n761# a_n2575_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X1 a_1177_n664# a_967_n761# a_909_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X2 a_2785_n664# a_2575_n761# a_2517_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X3 a_373_n664# a_163_n761# a_105_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X4 a_3053_n664# a_2843_n761# a_2785_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X5 a_641_n664# a_431_n761# a_373_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X6 a_n699_n664# a_n909_n761# a_n967_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X7 a_n2575_n664# a_n2785_n761# a_n2843_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X8 a_105_n664# a_n105_n761# a_n163_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X9 a_1445_n664# a_1235_n761# a_1177_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X10 a_1713_n664# a_1503_n761# a_1445_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X11 a_n967_n664# a_n1177_n761# a_n1235_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X12 a_n163_n664# a_n373_n761# a_n431_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X13 a_3321_n664# a_3111_n761# a_3053_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X14 a_n1235_n664# a_n1445_n761# a_n1503_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X15 a_n431_n664# a_n641_n761# a_n699_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X16 a_n2843_n664# a_n3053_n761# a_n3111_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X17 a_n1503_n664# a_n1713_n761# a_n1771_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X18 a_2249_n664# a_2039_n761# a_1981_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X19 a_1981_n664# a_1771_n761# a_1713_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X20 a_n3111_n664# a_n3321_n761# a_n3379_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.458e+07u w=7e+06u l=1.05e+06u
X21 a_2517_n664# a_2307_n761# a_2249_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X22 a_n2039_n664# a_n2249_n761# a_n2307_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+12p pd=1.458e+07u as=0p ps=0u w=7e+06u l=1.05e+06u
X23 a_909_n664# a_699_n761# a_641_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
X24 a_n1771_n664# a_n1981_n761# a_n2039_n664# w_n3517_n884# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=7e+06u l=1.05e+06u
.ends

.subckt opamp_manuel vin_n vin_p iref vout vdd vss
Xsky130_fd_pr__nfet_01v8_Z2S3N8_1 vss vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout a_7669_n7225# vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout sky130_fd_pr__nfet_01v8_Z2S3N8
Xsky130_fd_pr__nfet_01v8_J9MTE9_0 m1_11310_n8195# m1_11310_n8195# a_7669_n7225# m1_11310_n8195#
+ m1_11310_n8195# m1_11310_n8195# a_7669_n7225# a_7669_n7225# vss vdd m1_11310_n8195#
+ a_7669_n7225# a_7669_n7225# m1_11310_n8195# a_7669_n7225# a_7669_n7225# a_7669_n7225#
+ sky130_fd_pr__nfet_01v8_J9MTE9
Xsky130_fd_pr__nfet_01v8_Z2S3N8_2 vss vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout a_7669_n7225# vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout sky130_fd_pr__nfet_01v8_Z2S3N8
Xsky130_fd_pr__nfet_01v8_Z2S3N8_3 vss vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout a_7669_n7225# vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout sky130_fd_pr__nfet_01v8_Z2S3N8
Xsky130_fd_pr__pfet_01v8_H98ZZM_0 vss vdd vdd vp vp vdd iref iref iref vdd iref vdd
+ vdd iref vp iref iref iref iref iref vp vp iref vp vdd iref vdd vp iref vdd iref
+ iref vp iref iref vdd iref iref iref vp iref vdd vp iref vp iref vp iref iref vp
+ vdd vp vdd iref iref iref vp vdd iref vp vp iref iref iref iref vdd vdd iref vp
+ vdd iref iref vdd iref iref vp vdd vdd vp vdd iref iref vp iref vdd iref vp iref
+ iref vdd iref vdd vp vp vp iref vdd vp vdd iref iref iref iref sky130_fd_pr__pfet_01v8_H98ZZM
Xsky130_fd_pr__pfet_01v8_lvt_7XCYSC_0 vss m1_944_n7788# vin_p m1_944_n7788# vin_p
+ vin_p vp vin_p vin_p vin_p m1_944_n7788# vin_p vin_p vp vin_p vp vp m1_944_n7788#
+ vin_p m1_944_n7788# vin_p vp vin_p vp vin_p vin_p m1_944_n7788# m1_944_n7788# vin_p
+ vp vp m1_944_n7788# m1_944_n7788# m1_944_n7788# m1_944_n7788# vin_p vp vin_p vin_p
+ vin_p vin_p vp vp vin_p vp vp vin_p vin_p m1_944_n7788# vin_p vin_p vp m1_944_n7788#
+ sky130_fd_pr__pfet_01v8_lvt_7XCYSC
Xsky130_fd_pr__pfet_01v8_lvt_7XCYSC_1 vss a_7669_n7225# vin_n a_7669_n7225# vin_n
+ vin_n vp vin_n vin_n vin_n a_7669_n7225# vin_n vin_n vp vin_n vp vp a_7669_n7225#
+ vin_n a_7669_n7225# vin_n vp vin_n vp vin_n vin_n a_7669_n7225# a_7669_n7225# vin_n
+ vp vp a_7669_n7225# a_7669_n7225# a_7669_n7225# a_7669_n7225# vin_n vp vin_n vin_n
+ vin_n vin_n vp vp vin_n vp vp vin_n vin_n a_7669_n7225# vin_n vin_n vp a_7669_n7225#
+ sky130_fd_pr__pfet_01v8_lvt_7XCYSC
Xsky130_fd_pr__nfet_01v8_QVUSYJ_0 m1_944_n7788# m1_944_n7788# vss m1_944_n7788# m1_944_n7788#
+ vss vss m1_944_n7788# m1_944_n7788# vss m1_944_n7788# vss m1_944_n7788# vss m1_944_n7788#
+ vss m1_944_n7788# m1_944_n7788# m1_944_n7788# m1_944_n7788# m1_944_n7788# m1_944_n7788#
+ m1_944_n7788# m1_944_n7788# sky130_fd_pr__nfet_01v8_QVUSYJ
Xsky130_fd_pr__pfet_01v8_K4PBSX_0 iref vss vdd vout iref iref vdd vdd iref iref iref
+ vout vout vdd vout iref iref iref iref vout iref vdd iref iref iref vout vout iref
+ vdd iref vout vdd iref vdd iref iref iref iref iref vout iref vout iref iref vdd
+ vdd vdd vout vdd vout iref iref vout iref vout vdd vdd vout iref iref vout iref
+ vout vout vdd iref vdd iref iref iref iref vdd vdd iref vdd vout vout vdd vout vdd
+ iref iref vout vdd iref iref vout vdd vdd iref iref vdd vdd iref iref iref vout
+ iref iref iref vdd vout iref sky130_fd_pr__pfet_01v8_K4PBSX
Xsky130_fd_pr__nfet_01v8_QVUSYJ_1 vss m1_944_n7788# a_7669_n7225# m1_944_n7788# m1_944_n7788#
+ a_7669_n7225# a_7669_n7225# m1_944_n7788# m1_944_n7788# vss m1_944_n7788# a_7669_n7225#
+ vss a_7669_n7225# m1_944_n7788# a_7669_n7225# vss m1_944_n7788# m1_944_n7788# vss
+ m1_944_n7788# m1_944_n7788# vss vss sky130_fd_pr__nfet_01v8_QVUSYJ
Xsky130_fd_pr__pfet_01v8_K4PBSX_1 iref vss vdd vout iref iref vdd vdd iref iref iref
+ vout vout vdd vout iref iref iref iref vout iref vdd iref iref iref vout vout iref
+ vdd iref vout vdd iref vdd iref iref iref iref iref vout iref vout iref iref vdd
+ vdd vdd vout vdd vout iref iref vout iref vout vdd vdd vout iref iref vout iref
+ vout vout vdd iref vdd iref iref iref iref vdd vdd iref vdd vout vout vdd vout vdd
+ iref iref vout vdd iref iref vout vdd vdd iref iref vdd vdd iref iref iref vout
+ iref iref iref vdd vout iref sky130_fd_pr__pfet_01v8_K4PBSX
Xsky130_fd_pr__pfet_01v8_698KZZ_0 vss iref iref iref iref iref iref iref iref iref
+ vdd vdd vdd vdd iref iref vdd iref iref iref iref vdd vdd iref iref vdd iref iref
+ iref vdd iref iref iref sky130_fd_pr__pfet_01v8_698KZZ
Xsky130_fd_pr__pfet_01v8_65PBSZ_1 iref iref vss vdd vout vdd vout iref iref vdd iref
+ iref vout vdd vdd iref iref iref iref iref vout vout vdd iref vout vout iref iref
+ iref vout vdd vout vdd vout iref iref iref vdd iref vdd iref iref iref vout vdd
+ vout vdd vdd vdd iref vout vout iref iref iref iref vout vout vdd vdd vout vdd iref
+ iref iref vout vout iref vout iref iref vdd iref iref iref iref vdd vdd vdd iref
+ iref vout vdd vout iref vout vdd iref iref iref vout iref iref iref iref vdd vout
+ iref iref vdd vdd iref vdd sky130_fd_pr__pfet_01v8_65PBSZ
Xsky130_fd_pr__pfet_01v8_65PBSZ_0 iref iref vss vdd vout vdd vout iref iref vdd iref
+ iref vout vdd vdd iref iref iref iref iref vout vout vdd iref vout vout iref iref
+ iref vout vdd vout vdd vout iref iref iref vdd iref vdd iref iref iref vout vdd
+ vout vdd vdd vdd iref vout vout iref iref iref iref vout vout vdd vdd vout vdd iref
+ iref iref vout vout iref vout iref iref vdd iref iref iref iref vdd vdd vdd iref
+ iref vout vdd vout iref vout vdd iref iref iref vout iref iref iref iref vdd vout
+ iref iref vdd vdd iref vdd sky130_fd_pr__pfet_01v8_65PBSZ
Xsky130_fd_pr__cap_mim_m3_1_XFP5BZ_0 vss m1_11310_n8195# vout sky130_fd_pr__cap_mim_m3_1_XFP5BZ
Xsky130_fd_pr__cap_mim_m3_1_XFP5BZ_1 vss m1_11310_n8195# vout sky130_fd_pr__cap_mim_m3_1_XFP5BZ
Xsky130_fd_pr__pfet_01v8_lvt_RTJWSN_0 vss m1_944_n7788# vp m1_944_n7788# vin_p vin_p
+ vin_p m1_944_n7788# vin_p vin_p vin_p m1_944_n7788# vp vin_p m1_944_n7788# vin_p
+ vin_p vin_p vp vp vp m1_944_n7788# vin_p m1_944_n7788# vin_p vp vin_p vin_p vp vin_p
+ m1_944_n7788# m1_944_n7788# vp vp m1_944_n7788# m1_944_n7788# vin_p vin_p m1_944_n7788#
+ m1_944_n7788# vin_p vin_p vp vin_p vin_p vp vp vin_p vp vp vin_p vin_p vin_p sky130_fd_pr__pfet_01v8_lvt_RTJWSN
Xsky130_fd_pr__pfet_01v8_lvt_RTJWSN_1 vss a_7669_n7225# vp a_7669_n7225# vin_n vin_n
+ vin_n a_7669_n7225# vin_n vin_n vin_n a_7669_n7225# vp vin_n a_7669_n7225# vin_n
+ vin_n vin_n vp vp vp a_7669_n7225# vin_n a_7669_n7225# vin_n vp vin_n vin_n vp vin_n
+ a_7669_n7225# a_7669_n7225# vp vp a_7669_n7225# a_7669_n7225# vin_n vin_n a_7669_n7225#
+ a_7669_n7225# vin_n vin_n vp vin_n vin_n vp vp vin_n vp vp vin_n vin_n vin_n sky130_fd_pr__pfet_01v8_lvt_RTJWSN
Xsky130_fd_pr__nfet_01v8_Z2S3N8_0 vss vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout a_7669_n7225# vout vout vout vout vout vout vout vout vout vout vout
+ vout vout vout vout vout vout vout vout vout vout vout vout sky130_fd_pr__nfet_01v8_Z2S3N8
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NRCKZ4 VSUBS a_n861_n1464# a_n477_n1464# a_477_n1561#
+ a_861_n1561# a_n93_n1464# a_163_n1464# a_547_n1464# a_931_n1464# a_n803_n1561# a_n419_n1561#
+ a_93_n1561# a_n35_n1561# a_n733_n1464# a_n291_n1561# a_n349_n1464# a_n675_n1561#
+ a_733_n1561# w_n1127_n1684# a_349_n1561# a_419_n1464# a_803_n1464# a_n989_n1464#
+ a_291_n1464# a_675_n1464# a_35_n1464# a_n221_n1464# a_n605_n1464# a_n931_n1561#
+ a_n163_n1561# a_221_n1561# a_n547_n1561# a_605_n1561#
X0 a_803_n1464# a_733_n1561# a_675_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X1 a_547_n1464# a_477_n1561# a_419_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X2 a_n93_n1464# a_n163_n1561# a_n221_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X3 a_931_n1464# a_861_n1561# a_803_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X4 a_35_n1464# a_n35_n1561# a_n93_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X5 a_n349_n1464# a_n419_n1561# a_n477_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X6 a_n733_n1464# a_n803_n1561# a_n861_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X7 a_291_n1464# a_221_n1561# a_163_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X8 a_n221_n1464# a_n291_n1561# a_n349_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X9 a_n477_n1464# a_n547_n1561# a_n605_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X10 a_n861_n1464# a_n931_n1561# a_n989_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X11 a_n605_n1464# a_n675_n1561# a_n733_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X12 a_675_n1464# a_605_n1561# a_547_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X13 a_163_n1464# a_93_n1561# a_35_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X14 a_419_n1464# a_349_n1561# a_291_n1464# w_n1127_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NRU274 VSUBS a_n861_n1464# a_n477_n1464# a_477_n1561#
+ a_861_n1561# a_n93_n1464# a_1699_n1464# a_163_n1464# a_547_n1464# a_931_n1464# a_n1315_n1561#
+ a_1245_n1561# a_n1245_n1464# a_n1571_n1561# a_1629_n1561# a_n1629_n1464# a_n1187_n1561#
+ a_n803_n1561# a_n419_n1561# a_93_n1561# a_1315_n1464# a_n35_n1561# a_n733_n1464#
+ a_n291_n1561# a_n1885_n1464# a_n349_n1464# a_n675_n1561# a_733_n1561# a_1187_n1464#
+ a_1571_n1464# a_349_n1561# a_419_n1464# a_803_n1464# a_n989_n1464# a_989_n1561#
+ a_1501_n1561# a_n1501_n1464# a_291_n1464# a_1117_n1561# a_n1117_n1464# a_675_n1464#
+ a_n1443_n1561# a_n1059_n1561# a_n1827_n1561# a_35_n1464# a_n221_n1464# w_n2023_n1684#
+ a_1373_n1561# a_n1757_n1464# a_n1373_n1464# a_n605_n1464# a_n931_n1561# a_n163_n1561#
+ a_221_n1561# a_1757_n1561# a_1059_n1464# a_1443_n1464# a_n1699_n1561# a_n547_n1561#
+ a_605_n1561# a_1827_n1464#
X0 a_1827_n1464# a_1757_n1561# a_1699_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X1 a_803_n1464# a_733_n1561# a_675_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X2 a_547_n1464# a_477_n1561# a_419_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X3 a_n1629_n1464# a_n1699_n1561# a_n1757_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X4 a_1187_n1464# a_1117_n1561# a_1059_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X5 a_n93_n1464# a_n163_n1561# a_n221_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X6 a_931_n1464# a_861_n1561# a_803_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X7 a_35_n1464# a_n35_n1561# a_n93_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X8 a_n1245_n1464# a_n1315_n1561# a_n1373_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X9 a_n349_n1464# a_n419_n1561# a_n477_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X10 a_1571_n1464# a_1501_n1561# a_1443_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X11 a_n733_n1464# a_n803_n1561# a_n861_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X12 a_n989_n1464# a_n1059_n1561# a_n1117_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X13 a_291_n1464# a_221_n1561# a_163_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X14 a_1315_n1464# a_1245_n1561# a_1187_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X15 a_n221_n1464# a_n291_n1561# a_n349_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X16 a_n1373_n1464# a_n1443_n1561# a_n1501_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X17 a_n477_n1464# a_n547_n1561# a_n605_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X18 a_n861_n1464# a_n931_n1561# a_n989_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X19 a_n1117_n1464# a_n1187_n1561# a_n1245_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X20 a_1059_n1464# a_989_n1561# a_931_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X21 a_1443_n1464# a_1373_n1561# a_1315_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X22 a_1699_n1464# a_1629_n1561# a_1571_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X23 a_n605_n1464# a_n675_n1561# a_n733_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X24 a_675_n1464# a_605_n1561# a_547_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X25 a_n1501_n1464# a_n1571_n1561# a_n1629_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X26 a_n1757_n1464# a_n1827_n1561# a_n1885_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X27 a_163_n1464# a_93_n1561# a_35_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X28 a_419_n1464# a_349_n1561# a_291_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
.ends

.subckt bias_reference VSUBS vdd vbias_1 ibias
XM7 VSUBS ibias vbias_1 ibias ibias ibias ibias vbias_1 ibias ibias ibias ibias ibias
+ vbias_1 ibias ibias ibias ibias vbias_1 ibias ibias vbias_1 vbias_1 vbias_1 ibias
+ vbias_1 vbias_1 ibias ibias ibias ibias ibias ibias sky130_fd_pr__pfet_01v8_lvt_NRCKZ4
XM8 VSUBS vbias_1 vdd vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vdd vbias_1 vbias_1
+ vbias_1 vdd vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vdd vbias_1
+ vdd vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vdd vbias_1 vbias_1 vdd vdd
+ vbias_1 vbias_1 vdd vdd vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vdd vdd
+ vdd vbias_1 vdd vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vbias_1 vdd vbias_1 vbias_1
+ vbias_1 vbias_1 vdd sky130_fd_pr__pfet_01v8_lvt_NRU274
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_SNTUMW a_n897_n1500# a_255_n1500# a_351_n1500#
+ a_543_n1500# a_159_n1500# a_447_n1500# a_639_n1500# a_735_n1500# a_831_n1500# a_927_n1500#
+ a_n321_n1500# a_n927_n1526# a_n801_n1500# a_n705_n1500# a_n513_n1500# a_n417_n1500#
+ a_n225_n1500# a_n129_n1500# a_n609_n1500# a_n989_n1500# a_n33_n1500# a_63_n1500#
+ w_n1127_n1710#
X0 a_n225_n1500# a_n927_n1526# a_n321_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X1 a_543_n1500# a_n927_n1526# a_447_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X2 a_n33_n1500# a_n927_n1526# a_n129_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X3 a_n417_n1500# a_n927_n1526# a_n513_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X4 a_735_n1500# a_n927_n1526# a_639_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X5 a_n801_n1500# a_n927_n1526# a_n897_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X6 a_n609_n1500# a_n927_n1526# a_n705_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X7 a_63_n1500# a_n927_n1526# a_n33_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=0p ps=0u w=1.5e+07u l=150000u
X8 a_255_n1500# a_n927_n1526# a_159_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X9 a_n321_n1500# a_n927_n1526# a_n417_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X10 a_n129_n1500# a_n927_n1526# a_n225_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X11 a_447_n1500# a_n927_n1526# a_351_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.95e+12p ps=3.066e+07u w=1.5e+07u l=150000u
X12 a_n513_n1500# a_n927_n1526# a_n609_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X13 a_831_n1500# a_n927_n1526# a_735_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.95e+12p pd=3.066e+07u as=0p ps=0u w=1.5e+07u l=150000u
X14 a_639_n1500# a_n927_n1526# a_543_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X15 a_n705_n1500# a_n927_n1526# a_n801_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X16 a_351_n1500# a_n927_n1526# a_255_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X17 a_159_n1500# a_n927_n1526# a_63_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=150000u
X18 a_n897_n1500# a_n927_n1526# a_n989_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.65e+12p ps=3.062e+07u w=1.5e+07u l=150000u
X19 a_927_n1500# a_n927_n1526# a_831_n1500# w_n1127_n1710# sky130_fd_pr__nfet_01v8_lvt ad=4.65e+12p pd=3.062e+07u as=0p ps=0u w=1.5e+07u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_5U6LBF a_n897_n1875# w_n1127_n2085# a_351_n1875#
+ a_159_n1875# a_255_n1875# a_447_n1875# a_543_n1875# a_735_n1875# a_831_n1875# a_639_n1875#
+ a_927_n1875# a_n321_n1875# a_n801_n1875# a_n705_n1875# a_n513_n1875# a_n417_n1875#
+ a_n225_n1875# a_n129_n1875# a_n609_n1875# a_n33_n1875# a_n989_n1875# a_63_n1875#
+ a_n927_n1901#
X0 a_n513_n1875# a_n927_n1901# a_n609_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X1 a_639_n1875# a_n927_n1901# a_543_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X2 a_831_n1875# a_n927_n1901# a_735_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X3 a_n705_n1875# a_n927_n1901# a_n801_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X4 a_351_n1875# a_n927_n1901# a_255_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X5 a_159_n1875# a_n927_n1901# a_63_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X6 a_n897_n1875# a_n927_n1901# a_n989_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=5.8125e+12p ps=3.812e+07u w=1.875e+07u l=150000u
X7 a_927_n1875# a_n927_n1901# a_831_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=5.8125e+12p pd=3.812e+07u as=0p ps=0u w=1.875e+07u l=150000u
X8 a_n225_n1875# a_n927_n1901# a_n321_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X9 a_543_n1875# a_n927_n1901# a_447_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X10 a_n33_n1875# a_n927_n1901# a_n129_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X11 a_n417_n1875# a_n927_n1901# a_n513_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=0p ps=0u w=1.875e+07u l=150000u
X12 a_735_n1875# a_n927_n1901# a_639_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X13 a_n801_n1875# a_n927_n1901# a_n897_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X14 a_n609_n1875# a_n927_n1901# a_n705_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X15 a_63_n1875# a_n927_n1901# a_n33_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X16 a_255_n1875# a_n927_n1901# a_159_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X17 a_n321_n1875# a_n927_n1901# a_n417_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X18 a_n129_n1875# a_n927_n1901# a_n225_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X19 a_447_n1875# a_n927_n1901# a_351_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_EU6LGP a_n897_n1875# w_n1127_n2085# a_351_n1875#
+ a_159_n1875# a_255_n1875# a_447_n1875# a_543_n1875# a_735_n1875# a_831_n1875# a_639_n1875#
+ a_927_n1875# a_n321_n1875# a_n801_n1875# a_n705_n1875# a_n513_n1875# a_n417_n1875#
+ a_n225_n1875# a_n129_n1875# a_n609_n1875# a_n33_n1875# a_n989_n1875# a_63_n1875#
+ a_n927_n1901#
X0 a_n513_n1875# a_n927_n1901# a_n609_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X1 a_639_n1875# a_n927_n1901# a_543_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X2 a_831_n1875# a_n927_n1901# a_735_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X3 a_n705_n1875# a_n927_n1901# a_n801_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X4 a_351_n1875# a_n927_n1901# a_255_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X5 a_159_n1875# a_n927_n1901# a_63_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X6 a_n897_n1875# a_n927_n1901# a_n989_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=5.8125e+12p ps=3.812e+07u w=1.875e+07u l=150000u
X7 a_927_n1875# a_n927_n1901# a_831_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=5.8125e+12p pd=3.812e+07u as=0p ps=0u w=1.875e+07u l=150000u
X8 a_n225_n1875# a_n927_n1901# a_n321_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X9 a_543_n1875# a_n927_n1901# a_447_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X10 a_n33_n1875# a_n927_n1901# a_n129_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=6.1875e+12p ps=3.816e+07u w=1.875e+07u l=150000u
X11 a_n417_n1875# a_n927_n1901# a_n513_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=6.1875e+12p pd=3.816e+07u as=0p ps=0u w=1.875e+07u l=150000u
X12 a_735_n1875# a_n927_n1901# a_639_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X13 a_n801_n1875# a_n927_n1901# a_n897_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X14 a_n609_n1875# a_n927_n1901# a_n705_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X15 a_63_n1875# a_n927_n1901# a_n33_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X16 a_255_n1875# a_n927_n1901# a_159_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X17 a_n321_n1875# a_n927_n1901# a_n417_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X18 a_n129_n1875# a_n927_n1901# a_n225_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
X19 a_447_n1875# a_n927_n1901# a_351_n1875# w_n1127_n2085# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.875e+07u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_L5XAT6 a_639_n900# a_n927_n926# a_n321_n900# a_927_n900#
+ a_n225_n900# a_63_n900# a_n129_n900# a_n989_n900# a_n513_n900# a_n801_n900# a_n417_n900#
+ a_351_n900# a_255_n900# a_n705_n900# a_n609_n900# a_159_n900# a_543_n900# w_n1127_n1110#
+ a_447_n900# a_831_n900# a_n897_n900# a_n33_n900# a_735_n900#
X0 a_159_n900# a_n927_n926# a_63_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.97e+12p ps=1.866e+07u w=9e+06u l=150000u
X1 a_255_n900# a_n927_n926# a_159_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X2 a_351_n900# a_n927_n926# a_255_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X3 a_639_n900# a_n927_n926# a_543_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.97e+12p ps=1.866e+07u w=9e+06u l=150000u
X4 a_735_n900# a_n927_n926# a_639_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X5 a_831_n900# a_n927_n926# a_735_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X6 a_n33_n900# a_n927_n926# a_n129_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.97e+12p ps=1.866e+07u w=9e+06u l=150000u
X7 a_n513_n900# a_n927_n926# a_n609_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.97e+12p ps=1.866e+07u w=9e+06u l=150000u
X8 a_n417_n900# a_n927_n926# a_n513_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X9 a_n897_n900# a_n927_n926# a_n989_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.79e+12p ps=1.862e+07u w=9e+06u l=150000u
X10 a_447_n900# a_n927_n926# a_351_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X11 a_543_n900# a_n927_n926# a_447_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=150000u
X12 a_63_n900# a_n927_n926# a_n33_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=150000u
X13 a_n225_n900# a_n927_n926# a_n321_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=2.97e+12p ps=1.866e+07u w=9e+06u l=150000u
X14 a_n129_n900# a_n927_n926# a_n225_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=150000u
X15 a_n321_n900# a_n927_n926# a_n417_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=150000u
X16 a_n801_n900# a_n927_n926# a_n897_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X17 a_n705_n900# a_n927_n926# a_n801_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.97e+12p pd=1.866e+07u as=0p ps=0u w=9e+06u l=150000u
X18 a_n609_n900# a_n927_n926# a_n705_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=9e+06u l=150000u
X19 a_927_n900# a_n927_n926# a_831_n900# w_n1127_n1110# sky130_fd_pr__nfet_01v8_lvt ad=2.79e+12p pd=1.862e+07u as=0p ps=0u w=9e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QTSHDD VSUBS a_n989_n1014# a_291_n1014# a_675_n1014#
+ a_35_n1014# a_n221_n1014# a_n605_n1014# a_n163_n1111# a_221_n1111# a_n931_n1111#
+ a_n547_n1111# a_605_n1111# a_n861_n1014# a_n477_n1014# a_861_n1111# a_477_n1111#
+ a_n93_n1014# a_163_n1014# a_547_n1014# a_931_n1014# a_n803_n1111# a_93_n1111# a_n419_n1111#
+ a_n35_n1111# a_n733_n1014# a_n349_n1014# a_n291_n1111# w_n1127_n1234# a_n675_n1111#
+ a_349_n1111# a_733_n1111# a_803_n1014# a_419_n1014#
X0 a_547_n1014# a_477_n1111# a_419_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X1 a_n93_n1014# a_n163_n1111# a_n221_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X2 a_931_n1014# a_861_n1111# a_803_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X3 a_n349_n1014# a_n419_n1111# a_n477_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X4 a_35_n1014# a_n35_n1111# a_n93_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=0p ps=0u w=1.05e+07u l=350000u
X5 a_n733_n1014# a_n803_n1111# a_n861_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X6 a_291_n1014# a_221_n1111# a_163_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X7 a_n221_n1014# a_n291_n1111# a_n349_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=350000u
X8 a_n477_n1014# a_n547_n1111# a_n605_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X9 a_n861_n1014# a_n931_n1111# a_n989_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.045e+12p ps=2.158e+07u w=1.05e+07u l=350000u
X10 a_675_n1014# a_605_n1111# a_547_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=3.045e+12p pd=2.158e+07u as=0p ps=0u w=1.05e+07u l=350000u
X11 a_n605_n1014# a_n675_n1111# a_n733_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=350000u
X12 a_163_n1014# a_93_n1111# a_35_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=350000u
X13 a_419_n1014# a_349_n1111# a_291_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=350000u
X14 a_803_n1014# a_733_n1111# a_675_n1014# w_n1127_n1234# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.05e+07u l=350000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_ND8574 VSUBS a_n861_n1464# a_n477_n1464# a_477_n1561#
+ a_861_n1561# a_n93_n1464# a_1699_n1464# a_163_n1464# a_547_n1464# a_931_n1464# a_n1315_n1561#
+ a_1245_n1561# a_n1245_n1464# a_n1571_n1561# a_1629_n1561# a_n1629_n1464# a_n1187_n1561#
+ a_n803_n1561# a_n419_n1561# a_93_n1561# a_1315_n1464# a_n35_n1561# a_n733_n1464#
+ a_n291_n1561# a_n1885_n1464# a_n349_n1464# a_n675_n1561# a_733_n1561# a_1187_n1464#
+ a_1571_n1464# a_349_n1561# a_419_n1464# a_803_n1464# a_n989_n1464# a_989_n1561#
+ a_1501_n1561# a_n1501_n1464# a_291_n1464# a_1117_n1561# a_n1117_n1464# a_675_n1464#
+ a_n1443_n1561# a_n1059_n1561# a_n1827_n1561# a_35_n1464# a_n221_n1464# w_n2023_n1684#
+ a_1373_n1561# a_n1757_n1464# a_n1373_n1464# a_n605_n1464# a_n931_n1561# a_n163_n1561#
+ a_221_n1561# a_1757_n1561# a_1059_n1464# a_1443_n1464# a_n1699_n1561# a_n547_n1561#
+ a_605_n1561# a_1827_n1464#
X0 a_1827_n1464# a_1757_n1561# a_1699_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X1 a_803_n1464# a_733_n1561# a_675_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X2 a_547_n1464# a_477_n1561# a_419_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X3 a_n1629_n1464# a_n1699_n1561# a_n1757_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X4 a_1187_n1464# a_1117_n1561# a_1059_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X5 a_n93_n1464# a_n163_n1561# a_n221_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X6 a_931_n1464# a_861_n1561# a_803_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X7 a_35_n1464# a_n35_n1561# a_n93_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X8 a_n1245_n1464# a_n1315_n1561# a_n1373_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X9 a_n349_n1464# a_n419_n1561# a_n477_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X10 a_1571_n1464# a_1501_n1561# a_1443_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X11 a_n733_n1464# a_n803_n1561# a_n861_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X12 a_n989_n1464# a_n1059_n1561# a_n1117_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X13 a_291_n1464# a_221_n1561# a_163_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X14 a_1315_n1464# a_1245_n1561# a_1187_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.058e+07u as=0p ps=0u w=1.5e+07u l=350000u
X15 a_n221_n1464# a_n291_n1561# a_n349_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X16 a_n1373_n1464# a_n1443_n1561# a_n1501_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X17 a_n477_n1464# a_n547_n1561# a_n605_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X18 a_n861_n1464# a_n931_n1561# a_n989_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X19 a_n1117_n1464# a_n1187_n1561# a_n1245_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X20 a_1059_n1464# a_989_n1561# a_931_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X21 a_1443_n1464# a_1373_n1561# a_1315_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X22 a_1699_n1464# a_1629_n1561# a_1571_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X23 a_n605_n1464# a_n675_n1561# a_n733_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X24 a_675_n1464# a_605_n1561# a_547_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X25 a_n1501_n1464# a_n1571_n1561# a_n1629_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X26 a_n1757_n1464# a_n1827_n1561# a_n1885_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.058e+07u w=1.5e+07u l=350000u
X27 a_163_n1464# a_93_n1561# a_35_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
X28 a_419_n1464# a_349_n1561# a_291_n1464# w_n2023_n1684# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=350000u
.ends

.subckt bias vbias_1 ibias vbias_2 vss vdd
XM1 m1_3008_n382# m1_3008_n382# ibias ibias ibias m1_3008_n382# m1_3008_n382# ibias
+ m1_3008_n382# ibias m1_3008_n382# m1_764_4882# ibias m1_3008_n382# m1_3008_n382#
+ ibias ibias m1_3008_n382# ibias ibias ibias m1_3008_n382# vss sky130_fd_pr__nfet_01v8_lvt_SNTUMW
XM2 m1_3008_n382# vss vss vss m1_3008_n382# m1_3008_n382# vss vss m1_3008_n382# m1_3008_n382#
+ vss m1_3008_n382# vss m1_3008_n382# m1_3008_n382# vss vss m1_3008_n382# vss vss
+ vss m1_3008_n382# m1_879_3464# sky130_fd_pr__nfet_01v8_lvt_5U6LBF
XM4 m1_879_3464# vss vss vss m1_879_3464# m1_879_3464# vss vss m1_879_3464# m1_879_3464#
+ vss m1_879_3464# vss m1_879_3464# m1_879_3464# vss vss m1_879_3464# vss vss vss
+ m1_879_3464# m1_879_3464# sky130_fd_pr__nfet_01v8_lvt_EU6LGP
XM3 m1_879_3464# m1_764_4882# m1_879_3464# m1_764_4882# m1_764_4882# m1_879_3464#
+ m1_879_3464# m1_764_4882# m1_879_3464# m1_764_4882# m1_764_4882# m1_764_4882# m1_879_3464#
+ m1_879_3464# m1_764_4882# m1_764_4882# m1_764_4882# vss m1_879_3464# m1_879_3464#
+ m1_879_3464# m1_764_4882# m1_764_4882# sky130_fd_pr__nfet_01v8_lvt_L5XAT6
XM5 vss w_605_9716# w_605_9716# m1_764_4882# w_605_9716# w_605_9716# m1_764_4882#
+ vbias_2 vbias_2 vbias_2 vbias_2 vbias_2 m1_764_4882# w_605_9716# vbias_2 vbias_2
+ m1_764_4882# m1_764_4882# w_605_9716# m1_764_4882# vbias_2 vbias_2 vbias_2 vbias_2
+ w_605_9716# m1_764_4882# vbias_2 w_605_9716# vbias_2 vbias_2 vbias_2 w_605_9716#
+ m1_764_4882# sky130_fd_pr__pfet_01v8_lvt_QTSHDD
XM6 vss w_605_9716# vdd vbias_1 vbias_1 w_605_9716# w_605_9716# w_605_9716# vdd w_605_9716#
+ vbias_1 vbias_1 vdd vbias_1 vbias_1 w_605_9716# vbias_1 vbias_1 vbias_1 vbias_1
+ vdd vbias_1 vdd vbias_1 w_605_9716# w_605_9716# vbias_1 vbias_1 w_605_9716# vdd
+ vbias_1 w_605_9716# vdd vdd vbias_1 vbias_1 vdd vdd vbias_1 w_605_9716# w_605_9716#
+ vbias_1 vbias_1 vbias_1 vdd vdd vdd vbias_1 vdd w_605_9716# w_605_9716# vbias_1
+ vbias_1 vbias_1 vbias_1 vdd w_605_9716# vbias_1 vbias_1 vbias_1 vdd sky130_fd_pr__pfet_01v8_lvt_ND8574
.ends

.subckt bias_circuit vss vref vdd ibias_1 ibias_2 ibias_3
Xbias_reference_0 vss vdd bias_2/vbias_1 vref bias_reference
Xbias_1 bias_2/vbias_1 ibias_2 vref vss vdd bias
Xbias_0 bias_2/vbias_1 ibias_1 vref vss vdd bias
Xbias_2 bias_2/vbias_1 ibias_3 vref vss vdd bias
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_CWLY9J VSUBS a_n29_n735# a_269_n735# a_29_n832#
+ a_n327_n735# w_n465_n954# a_n269_n832#
X0 a_n29_n735# a_n269_n832# a_n327_n735# w_n465_n954# sky130_fd_pr__pfet_01v8_lvt ad=2.1315e+12p pd=1.528e+07u as=2.1315e+12p ps=1.528e+07u w=7.35e+06u l=1.2e+06u
X1 a_269_n735# a_29_n832# a_n29_n735# w_n465_n954# sky130_fd_pr__pfet_01v8_lvt ad=2.1315e+12p pd=1.528e+07u as=0p ps=0u w=7.35e+06u l=1.2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZWZ6GW a_n325_n420# a_119_n420# a_325_n508# a_n267_n508#
+ a_563_n420# a_n177_n420# a_177_n508# a_n119_n508# a_n621_n420# a_415_n420# a_n563_n508#
+ w_n759_n630# a_n29_n420# a_29_n508# a_n473_n420# a_473_n508# a_267_n420# a_n415_n508#
X0 a_563_n420# a_473_n508# a_415_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=1.218e+12p pd=8.98e+06u as=1.218e+12p ps=8.98e+06u w=4.2e+06u l=450000u
X1 a_267_n420# a_177_n508# a_119_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=1.218e+12p pd=8.98e+06u as=1.218e+12p ps=8.98e+06u w=4.2e+06u l=450000u
X2 a_n473_n420# a_n563_n508# a_n621_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=1.218e+12p pd=8.98e+06u as=1.218e+12p ps=8.98e+06u w=4.2e+06u l=450000u
X3 a_n177_n420# a_n267_n508# a_n325_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=1.218e+12p pd=8.98e+06u as=1.218e+12p ps=8.98e+06u w=4.2e+06u l=450000u
X4 a_415_n420# a_325_n508# a_267_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.2e+06u l=450000u
X5 a_n325_n420# a_n415_n508# a_n473_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.2e+06u l=450000u
X6 a_n29_n420# a_n119_n508# a_n177_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=1.218e+12p pd=8.98e+06u as=0p ps=0u w=4.2e+06u l=450000u
X7 a_119_n420# a_29_n508# a_n29_n420# w_n759_n630# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.2e+06u l=450000u
.ends

.subckt input vss vin_n vin_p iref vout
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|0] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|0] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|0] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|0] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|0] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|1] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|1] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|1] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|1] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|1] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|2] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|2] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|2] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|2] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|2] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|3] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|3] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|3] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|3] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|3] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|4] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|4] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|4] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|4] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|4] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|5] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|5] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|5] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|5] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|5] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|6] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|6] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|6] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|6] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|6] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[0|7] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[1|7] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[2|7] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[3|7] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__pfet_01v8_lvt_CWLY9J_0[4|7] vss iref vout_n vin_n vout iref vin_p sky130_fd_pr__pfet_01v8_lvt_CWLY9J
Xsky130_fd_pr__nfet_01v8_ZWZ6GW_0 vss vout_n vout_n vout_n vss vout vout_n vout_n
+ vss vout vout_n vss vss vout_n vout_n vout_n vss vout_n sky130_fd_pr__nfet_01v8_ZWZ6GW
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_6BP6N2 VSUBS c1_2209_n5080# c1_n4869_n5080# m3_n1430_n5180#
+ c1_n1330_n5080# m3_2109_n5180# m3_n4969_n5180#
X0 c1_n4869_n5080# m3_n4969_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X1 c1_2209_n5080# m3_2109_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X2 c1_n4869_n5080# m3_n4969_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X3 c1_n4869_n5080# m3_n4969_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X4 c1_n1330_n5080# m3_n1430_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X5 c1_n1330_n5080# m3_n1430_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X6 c1_n1330_n5080# m3_n1430_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X7 c1_2209_n5080# m3_2109_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X8 c1_2209_n5080# m3_2109_n5180# sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_RE4H9G a_399_n587# a_n1905_521# a_783_521# a_n945_1737#
+ a_1455_n1303# a_1311_717# a_783_n587# a_1455_1237# a_15_n1803# a_1647_n1303# a_n993_109#
+ a_303_1237# a_n897_n499# a_1695_717# a_111_n1303# a_831_717# a_n465_n87# a_1839_n1303#
+ a_255_1325# a_n177_629# a_1791_1325# a_303_n1303# a_n705_1325# a_1215_109# a_n33_717#
+ a_1743_629# a_1599_109# a_n993_n1715# a_351_717# a_735_109# a_n945_521# a_n897_n1715#
+ a_n1617_1237# a_n1857_717# a_495_21# a_n465_1129# a_n1569_1325# a_1887_n499# a_n1233_21#
+ a_975_n695# a_735_n499# a_n33_n499# a_255_109# a_n1949_n1107# a_399_1737# a_n1905_629#
+ a_n1377_717# a_783_629# a_1071_n87# a_783_1737# a_n1949_109# a_1791_n1715# a_n513_717#
+ a_1695_n1715# a_n1137_n695# a_159_1325# a_1695_1325# a_1599_n1715# a_n609_1325#
+ a_1887_n1715# a_n897_717# a_n1521_n695# a_207_521# a_543_1325# a_n1041_n1303# a_351_n1715#
+ a_495_n1195# a_1551_521# a_1455_1129# a_n1761_109# a_303_1129# a_n465_21# a_n1233_n1303#
+ a_255_n1715# a_543_n1715# a_n417_109# a_n657_1237# a_831_n1715# a_687_n1195# a_n1233_n87#
+ a_1119_717# a_n945_629# a_159_n1715# a_447_n1715# a_n1425_n1303# a_735_n1715# a_879_n1195#
+ a_639_n1715# a_n1281_109# a_639_717# a_n993_1325# a_n1617_n1303# a_927_n1715# a_n1281_n499#
+ a_1023_n499# a_639_n499# a_n1857_1325# a_n1809_n1303# a_n1713_521# a_1839_n87# a_591_521#
+ a_63_109# a_1647_21# a_n1617_1129# a_1503_109# a_159_717# a_975_n587# a_n177_n695#
+ a_1887_109# a_1647_1237# a_n273_n87# a_n561_n695# a_1599_1325# a_n321_n499# a_1023_109#
+ a_15_n695# a_207_629# a_447_1325# a_15_521# a_n273_n1195# a_1551_629# a_879_n87#
+ a_831_1325# a_543_109# a_n321_n1715# a_n465_n1195# a_n1137_n587# a_n753_521# a_495_1237#
+ a_n1281_n1715# a_n1665_717# a_n225_n1715# a_n513_n1715# a_n657_n1195# a_n1521_n587#
+ a_n801_n1715# a_n1473_n1715# a_n1185_n1715# a_n1761_n1715# a_n1809_1237# a_n897_1325#
+ a_n417_n1715# a_n129_n1715# a_1167_n695# a_n1185_n499# a_n705_n1715# a_n849_n1195#
+ a_n1089_n1715# a_n1377_n1715# a_n801_717# a_n657_1129# a_n1665_n1715# a_1551_n695#
+ a_879_21# a_n609_n1715# w_n2087_n1925# a_n1713_629# a_1359_521# a_1311_n499# a_n1569_n1715#
+ a_n1617_21# a_n1185_717# a_591_629# a_n1857_n1715# a_1071_n1195# a_927_n499# a_n1569_109#
+ a_n81_n87# a_n81_n1195# a_1071_21# a_1263_n1195# a_n1041_1237# a_975_1737# a_n321_717#
+ a_n705_109# a_1407_717# a_1023_n1715# a_1311_n1715# a_1455_n1195# a_n1089_109# a_n33_n1715#
+ a_n225_n499# a_1215_n1715# a_n1329_n695# a_1503_n1715# a_1647_n1195# a_927_717#
+ a_1887_1325# a_111_n1195# a_n1713_n695# a_n177_n587# a_15_629# a_1119_n1715# a_399_521#
+ a_1407_n1715# a_1839_n1195# a_n33_1325# a_735_1325# a_n225_109# a_1647_1129# a_n1041_n87#
+ a_n561_n587# a_303_n1195# a_n1137_1737# a_n753_629# a_n849_1237# a_n1949_n499# a_n849_21#
+ a_n1521_1737# a_n81_1237# a_15_n587# a_447_717# a_n1089_n499# a_1791_717# a_63_n1715#
+ a_n1473_n499# a_n1521_521# a_63_n499# a_1647_n87# a_495_1129# a_1215_n499# a_1311_109#
+ a_1359_629# a_n1809_1129# a_1167_n587# a_n1041_21# a_1695_109# a_1551_n587# a_591_n1803#
+ a_831_109# a_n369_n695# a_1839_1237# a_n129_n499# a_303_n87# a_783_n1803# a_n753_n695#
+ a_n33_109# a_n609_717# a_n1281_1325# a_n513_n499# a_n1809_n87# a_399_n1803# a_975_n1803#
+ a_687_n87# a_1023_1325# a_303_21# a_n177_1737# a_n1041_1129# a_639_1325# a_n993_n1107#
+ a_351_109# a_399_629# a_n561_521# a_n561_1737# a_n897_n1107# a_n1473_717# a_n1041_n1195#
+ a_n1857_109# a_n1329_n587# a_1071_1237# a_n129_717# a_687_1237# a_15_1737# a_n1233_n1195#
+ a_n1713_n587# a_n273_21# a_n81_21# a_1359_n695# a_n1377_n499# a_n1425_n1195# a_n1521_629#
+ a_1167_521# a_n321_1325# a_1119_n499# a_n849_1129# a_207_n695# a_n1377_109# a_n993_717#
+ a_1743_n695# a_n1761_n499# a_n1617_n1195# a_n81_1129# a_1503_n499# a_1791_n1107#
+ a_n849_n87# a_1167_1737# a_n1809_n1195# a_n513_109# a_1695_n1107# a_1215_717# a_1551_1737#
+ a_n1233_1237# a_1455_21# a_1599_n1107# a_1887_n1107# a_n897_109# a_1599_717# a_n561_n1803#
+ a_351_n1107# a_n1185_1325# a_735_717# a_591_n695# a_n417_n499# a_n1329_521# a_n177_n1803#
+ a_n753_n1803# a_351_n499# a_255_n1107# a_543_n1107# a_831_n1107# a_n801_n499# a_1119_109#
+ a_n369_n587# a_n369_n1803# a_n1905_n695# a_1311_1325# a_n561_629# a_n945_n1803#
+ a_159_n1107# a_1839_1129# a_927_1325# a_447_n1107# a_735_n1107# a_n753_n587# a_n1329_1737#
+ a_255_717# a_639_109# a_639_n1107# a_927_n1107# a_n1949_n1715# a_n1713_1737# a_1455_n87#
+ a_n1949_717# a_n225_1325# a_1167_629# a_n1665_n499# a_1071_1129# a_1551_n1803# a_687_1129#
+ a_1407_n499# a_159_109# a_n369_521# a_1167_n1803# a_n273_1237# a_1743_n1803# a_1359_n587#
+ a_687_21# a_n1949_1325# a_1359_n1803# a_207_n587# a_n1761_717# a_111_n87# a_n1425_21#
+ a_1743_n587# a_n417_717# a_n1617_n87# a_n1089_1325# a_495_n87# a_n945_n695# a_n1329_629#
+ a_255_n499# a_n1473_1325# a_1791_n499# a_n705_n499# a_n321_n1107# a_63_1325# a_n369_1737#
+ a_1215_1325# a_n1233_1129# a_207_n1803# a_n1281_n1107# a_n1281_717# a_n1665_109#
+ a_n225_n1107# a_n513_n1107# a_n801_n1107# a_n753_1737# a_n1185_n1107# a_n1473_n1107#
+ a_n1761_n1107# a_591_n587# a_n129_n1107# a_n417_n1107# a_n705_n1107# a_1263_1237#
+ a_975_521# a_63_717# a_n1089_n1107# a_879_1237# a_n1377_n1107# a_n801_109# a_n1665_n1107#
+ a_1503_717# a_111_1237# a_n1905_n587# a_n609_n1107# a_n129_1325# a_n1569_n1107#
+ a_n1185_109# a_n1857_n1107# a_495_n1303# a_n1569_n499# a_1887_717# a_n657_21# a_n513_1325#
+ a_n657_n87# a_687_n1303# a_n369_629# a_n321_109# a_1023_717# a_1407_109# a_1023_n1107#
+ a_1359_1737# a_1311_n1107# a_879_n1303# a_n33_n1107# a_207_1737# a_1215_n1107# a_1743_1737#
+ a_1503_n1107# a_n1425_1237# a_543_717# a_927_109# a_n1137_521# a_399_n695# a_1119_n1107#
+ a_1839_21# a_n273_1129# a_1407_n1107# a_159_n499# a_n1377_1325# a_783_n695# a_1695_n499#
+ a_n609_n499# a_1119_1325# a_543_n499# a_n1761_1325# a_1503_1325# a_n1521_n1803#
+ a_447_109# a_n945_n587# a_591_1737# a_1791_109# a_n1137_n1803# a_63_n1107# a_111_21#
+ a_n1569_717# a_n1713_n1803# a_975_629# a_1263_n87# a_n1905_1737# a_n1329_n1803#
+ a_n1905_n1803# a_n993_n499# a_n273_n1303# a_n705_717# a_n417_1325# a_n177_521# a_n1857_n499#
+ a_1263_1129# a_351_1325# a_n465_n1303# a_n1089_717# a_879_1129# a_n801_1325# a_111_1129#
+ a_1743_521# a_n465_1237# a_n657_n1303# a_n225_717# a_n609_109# a_n849_n1303# a_n1425_n87#
+ a_n1137_629# a_n1809_21# a_1599_n499# a_1071_n1303# a_1263_21# a_447_n499# a_n1473_109#
+ a_n1665_1325# a_n81_n1303# a_1407_1325# a_n1425_1129# a_1263_n1303# a_n129_109#
+ a_831_n499#
X0 a_1695_717# a_1647_1129# a_1599_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X1 a_63_1325# a_15_1737# a_n33_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X2 a_n33_717# a_n81_1129# a_n129_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X3 a_1695_109# a_1647_21# a_1599_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X4 a_1695_n1715# a_1647_n1303# a_1599_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X5 a_1503_n499# a_1455_n87# a_1407_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X6 a_n993_1325# a_n1041_1237# a_n1089_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X7 a_n33_109# a_n81_21# a_n129_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X8 a_159_n499# a_111_n87# a_63_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X9 a_735_n1715# a_687_n1303# a_639_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X10 a_1695_n1107# a_1647_n1195# a_1599_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X11 a_735_n1107# a_687_n1195# a_639_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X12 a_1599_717# a_1551_629# a_1503_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X13 a_1599_109# a_1551_521# a_1503_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X14 a_n1665_1325# a_n1713_1737# a_n1761_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X15 a_1791_n499# a_1743_n587# a_1695_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X16 a_n1281_1325# a_n1329_1737# a_n1377_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X17 a_447_n499# a_399_n587# a_351_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X18 a_n609_n499# a_n657_n87# a_n705_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X19 a_n1377_n1715# a_n1425_n1303# a_n1473_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X20 a_n1377_n1107# a_n1425_n1195# a_n1473_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X21 a_n1281_717# a_n1329_629# a_n1377_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X22 a_n1281_109# a_n1329_521# a_n1377_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X23 a_n33_n1715# a_n81_n1303# a_n129_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X24 a_735_n499# a_687_n87# a_639_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X25 a_n33_n1107# a_n81_n1195# a_n129_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X26 a_1311_n499# a_1263_n87# a_1215_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X27 a_n33_1325# a_n81_1237# a_n129_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X28 a_543_717# a_495_1129# a_447_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X29 a_n897_n499# a_n945_n587# a_n993_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X30 a_n321_717# a_n369_629# a_n417_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X31 a_543_109# a_495_21# a_447_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X32 a_n129_n499# a_n177_n587# a_n225_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X33 a_n705_n1715# a_n753_n1803# a_n801_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X34 a_n1185_717# a_n1233_1129# a_n1281_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X35 a_n321_109# a_n369_521# a_n417_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X36 a_1407_n1715# a_1359_n1803# a_1311_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X37 a_n705_n1107# a_n753_n695# a_n801_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X38 a_n1185_109# a_n1233_21# a_n1281_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X39 a_447_n1715# a_399_n1803# a_351_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X40 a_1407_n1107# a_1359_n695# a_1311_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X41 a_447_n1107# a_399_n695# a_351_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X42 a_447_717# a_399_629# a_351_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X43 a_1599_1325# a_1551_1737# a_1503_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X44 a_n225_717# a_n273_1129# a_n321_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X45 a_447_109# a_399_521# a_351_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X46 a_n1089_717# a_n1137_629# a_n1185_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X47 a_n225_109# a_n273_21# a_n321_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X48 a_255_n499# a_207_n587# a_159_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X49 a_n1089_109# a_n1137_521# a_n1185_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X50 a_n417_n499# a_n465_n87# a_n513_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X51 a_1791_n1715# a_1743_n1803# a_1695_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X52 a_831_n1715# a_783_n1803# a_735_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X53 a_n129_717# a_n177_629# a_n225_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X54 a_1791_n1107# a_1743_n695# a_1695_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X55 a_831_n1107# a_783_n695# a_735_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X56 a_n1761_1325# a_n1809_1237# a_n1857_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X57 a_n129_109# a_n177_521# a_n225_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X58 a_n1089_n499# a_n1137_n587# a_n1185_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X59 a_927_n499# a_879_n87# a_831_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X60 a_1887_1325# a_1839_1237# a_1791_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X61 a_n1089_n1715# a_n1137_n1803# a_n1185_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X62 a_n1089_n1107# a_n1137_n695# a_n1185_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X63 a_543_n499# a_495_n87# a_447_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X64 a_1119_1325# a_1071_1237# a_1023_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X65 a_1311_717# a_1263_1129# a_1215_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X66 a_n705_n499# a_n753_n587# a_n801_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X67 a_n1857_n1715# a_n1905_n1803# a_n1949_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X68 a_n897_717# a_n945_629# a_n993_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X69 a_1311_109# a_1263_21# a_1215_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X70 a_n1857_n1107# a_n1905_n695# a_n1949_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X71 a_n897_109# a_n945_521# a_n993_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X72 a_1215_717# a_1167_629# a_1119_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X73 a_n1377_n499# a_n1425_n87# a_n1473_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X74 a_1215_109# a_1167_521# a_1119_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X75 a_n417_n1715# a_n465_n1303# a_n513_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X76 a_1119_n1715# a_1071_n1303# a_1023_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X77 a_159_n1715# a_111_n1303# a_63_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X78 a_n1473_n1715# a_n1521_n1803# a_n1569_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X79 a_n417_n1107# a_n465_n1195# a_n513_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X80 a_831_n499# a_783_n587# a_735_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X81 a_1407_1325# a_1359_1737# a_1311_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X82 a_1119_n1107# a_1071_n1195# a_1023_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X83 a_159_n1107# a_111_n1195# a_63_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X84 a_n1473_n1107# a_n1521_n695# a_n1569_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X85 a_927_n1715# a_879_n1303# a_831_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X86 a_1119_717# a_1071_1129# a_1023_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X87 a_n225_n499# a_n273_n87# a_n321_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X88 a_927_n1107# a_879_n1195# a_831_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X89 a_1119_109# a_1071_21# a_1023_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X90 a_n1761_717# a_n1809_1129# a_n1857_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X91 a_63_717# a_15_629# a_n33_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X92 a_n1761_109# a_n1809_21# a_n1857_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X93 a_63_109# a_15_521# a_n33_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X94 a_1503_n1715# a_1455_n1303# a_1407_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X95 a_n801_n1715# a_n849_n1303# a_n897_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X96 a_n801_n1107# a_n849_n1195# a_n897_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X97 a_1695_1325# a_1647_1237# a_1599_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X98 a_1023_717# a_975_629# a_927_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X99 a_1887_717# a_1839_1129# a_1791_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X100 a_543_n1715# a_495_n1303# a_447_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X101 a_1503_n1107# a_1455_n1195# a_1407_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X102 a_1023_109# a_975_521# a_927_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X103 a_1887_109# a_1839_21# a_1791_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X104 a_351_n499# a_303_n87# a_255_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X105 a_543_n1107# a_495_n1195# a_447_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X106 a_n1665_717# a_n1713_629# a_n1761_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X107 a_n513_n499# a_n561_n587# a_n609_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X108 a_n1665_109# a_n1713_521# a_n1761_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X109 a_n1569_n499# a_n1617_n87# a_n1665_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X110 a_n1569_n1715# a_n1617_n1303# a_n1665_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X111 a_927_717# a_879_1129# a_831_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X112 a_n1569_n1107# a_n1617_n1195# a_n1665_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X113 a_927_109# a_879_21# a_831_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X114 a_n1185_n499# a_n1233_n87# a_n1281_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X115 a_1023_n499# a_975_n587# a_927_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X116 a_n1569_717# a_n1617_1129# a_n1665_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X117 a_639_1325# a_591_1737# a_543_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X118 a_n1569_109# a_n1617_21# a_n1665_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X119 a_1215_1325# a_1167_1737# a_1119_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X120 a_n801_n499# a_n849_n87# a_n897_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X121 a_n129_n1715# a_n177_n1803# a_n225_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X122 a_n129_n1107# a_n177_n695# a_n225_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X123 a_n1857_n499# a_n1905_n587# a_n1949_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X124 a_n1185_n1715# a_n1233_n1303# a_n1281_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X125 a_n1185_n1107# a_n1233_n1195# a_n1281_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X126 a_n1473_n499# a_n1521_n587# a_n1569_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X127 a_831_717# a_783_629# a_735_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X128 a_831_109# a_783_521# a_735_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X129 a_159_1325# a_111_1237# a_63_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X130 a_1503_1325# a_1455_1237# a_1407_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X131 a_n1473_717# a_n1521_629# a_n1569_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X132 a_n1473_109# a_n1521_521# a_n1569_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X133 a_n513_n1715# a_n561_n1803# a_n609_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X134 a_735_717# a_687_1129# a_639_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X135 a_n321_n499# a_n369_n587# a_n417_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X136 a_1215_n1715# a_1167_n1803# a_1119_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X137 a_n513_n1107# a_n561_n695# a_n609_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X138 a_735_109# a_687_21# a_639_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X139 a_255_n1715# a_207_n1803# a_159_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X140 a_1215_n1107# a_1167_n695# a_1119_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X141 a_n513_717# a_n561_629# a_n609_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X142 a_1023_n1715# a_975_n1803# a_927_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X143 a_255_n1107# a_207_n695# a_159_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X144 a_n1377_717# a_n1425_1129# a_n1473_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X145 a_n1377_109# a_n1425_21# a_n1473_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X146 a_n513_109# a_n561_521# a_n609_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X147 a_63_n499# a_15_n587# a_n33_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X148 a_1023_n1107# a_975_n695# a_927_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X149 a_n993_n499# a_n1041_n87# a_n1089_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X150 a_447_1325# a_399_1737# a_351_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X151 a_1791_1325# a_1743_1737# a_1695_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X152 a_639_717# a_591_629# a_543_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X153 a_63_n1715# a_15_n1803# a_n33_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X154 a_639_109# a_591_521# a_543_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X155 a_63_n1107# a_15_n695# a_n33_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X156 a_n609_1325# a_n657_1237# a_n705_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X157 a_n417_717# a_n465_1129# a_n513_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X158 a_n417_109# a_n465_21# a_n513_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X159 a_n1665_n499# a_n1713_n587# a_n1761_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X160 a_n1281_n499# a_n1329_n587# a_n1377_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X161 a_735_1325# a_687_1237# a_639_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X162 a_1311_1325# a_1263_1237# a_1215_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X163 a_n1665_n1715# a_n1713_n1803# a_n1761_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X164 a_n897_1325# a_n945_1737# a_n993_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X165 a_n1665_n1107# a_n1713_n695# a_n1761_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X166 a_1503_717# a_1455_1129# a_1407_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X167 a_n129_1325# a_n177_1737# a_n225_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X168 a_1503_109# a_1455_21# a_1407_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X169 a_n225_n1715# a_n273_n1303# a_n321_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X170 a_1887_n1715# a_1839_n1303# a_1791_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=0p ps=0u w=1.95e+06u l=150000u
X171 a_n1281_n1715# a_n1329_n1803# a_n1377_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X172 a_n225_n1107# a_n273_n1195# a_n321_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X173 a_1407_717# a_1359_629# a_1311_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X174 a_n33_n499# a_n81_n87# a_n129_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X175 a_1887_n1107# a_1839_n1195# a_1791_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=0p ps=0u w=1.95e+06u l=150000u
X176 a_n1281_n1107# a_n1329_n695# a_n1377_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X177 a_255_1325# a_207_1737# a_159_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X178 a_1407_109# a_1359_521# a_1311_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X179 a_n417_1325# a_n465_1237# a_n513_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X180 a_n1089_1325# a_n1137_1737# a_n1185_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X181 a_927_1325# a_879_1237# a_831_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X182 a_1599_n499# a_1551_n587# a_1503_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X183 a_1311_n1715# a_1263_n1303# a_1215_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X184 a_351_n1715# a_303_n1303# a_255_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X185 a_543_1325# a_495_1237# a_447_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X186 a_1311_n1107# a_1263_n1195# a_1215_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X187 a_351_n1107# a_303_n1195# a_255_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X188 a_n705_1325# a_n753_1737# a_n801_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X189 a_n1857_717# a_n1905_629# a_n1949_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X190 a_n1857_109# a_n1905_521# a_n1949_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X191 a_n1761_n499# a_n1809_n87# a_n1857_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X192 a_351_717# a_303_1129# a_255_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X193 a_1887_n499# a_1839_n87# a_1791_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.045e+11p pd=4.52e+06u as=0p ps=0u w=1.95e+06u l=150000u
X194 a_n1377_1325# a_n1425_1237# a_n1473_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X195 a_351_109# a_303_21# a_255_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X196 a_1119_n499# a_1071_n87# a_1023_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X197 a_831_1325# a_783_1737# a_735_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X198 a_n993_717# a_n1041_1129# a_n1089_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X199 a_n993_109# a_n1041_21# a_n1089_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X200 a_n897_n1715# a_n945_n1803# a_n993_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X201 a_n225_1325# a_n273_1237# a_n321_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X202 a_255_717# a_207_629# a_159_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X203 a_1599_n1715# a_1551_n1803# a_1503_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X204 a_639_n1715# a_591_n1803# a_543_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X205 a_n993_n1715# a_n1041_n1303# a_n1089_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X206 a_n897_n1107# a_n945_n695# a_n993_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X207 a_255_109# a_207_521# a_159_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.435e+11p ps=4.56e+06u w=1.95e+06u l=150000u
X208 a_n1761_n1715# a_n1809_n1303# a_n1857_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X209 a_1599_n1107# a_1551_n695# a_1503_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X210 a_639_n1107# a_591_n695# a_543_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X211 a_n993_n1107# a_n1041_n1195# a_n1089_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X212 a_n1761_n1107# a_n1809_n1195# a_n1857_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X213 a_1407_n499# a_1359_n587# a_1311_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X214 a_159_717# a_111_1129# a_63_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X215 a_351_1325# a_303_1237# a_255_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X216 a_159_109# a_111_21# a_63_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X217 a_n321_n1715# a_n369_n1803# a_n417_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X218 a_n513_1325# a_n561_1737# a_n609_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X219 a_n801_717# a_n849_1129# a_n897_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X220 a_n321_n1107# a_n369_n695# a_n417_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X221 a_n801_109# a_n849_21# a_n897_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X222 a_n1569_1325# a_n1617_1237# a_n1665_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X223 a_n1185_1325# a_n1233_1237# a_n1281_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X224 a_1023_1325# a_975_1737# a_927_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X225 a_1695_n499# a_1647_n87# a_1599_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X226 a_n705_717# a_n753_629# a_n801_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X227 a_n705_109# a_n753_521# a_n801_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=6.435e+11p pd=4.56e+06u as=0p ps=0u w=1.95e+06u l=150000u
X228 a_n801_1325# a_n849_1237# a_n897_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X229 a_n609_717# a_n657_1129# a_n705_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X230 a_n1857_1325# a_n1905_1737# a_n1949_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.045e+11p ps=4.52e+06u w=1.95e+06u l=150000u
X231 a_n609_109# a_n657_21# a_n705_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X232 a_n1473_1325# a_n1521_1737# a_n1569_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X233 a_n609_n1715# a_n657_n1303# a_n705_n1715# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X234 a_n609_n1107# a_n657_n1195# a_n705_n1107# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X235 a_639_n499# a_591_n587# a_543_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X236 a_1215_n499# a_1167_n587# a_1119_n499# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X237 a_1791_717# a_1743_629# a_1695_717# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X238 a_1791_109# a_1743_521# a_1695_109# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
X239 a_n321_1325# a_n369_1737# a_n417_1325# w_n2087_n1925# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.95e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_B8HNLY a_n865_627# a_n807_1057# a_1225_109# a_n1283_n1445#
+ a_n807_n1015# a_447_21# a_1283_1575# a_n1701_1145# a_n2061_21# a_807_n1963# a_n1283_n409#
+ a_389_2181# a_447_n497# a_1643_n2481# a_n1701_627# a_n1225_n497# a_n29_n1445# a_1701_n1015#
+ a_n447_n409# a_n1701_n927# a_389_1663# a_n447_109# a_1643_n1963# a_n865_1145# a_2061_n1445#
+ a_n389_n497# a_1225_n2481# a_n1643_n1015# a_29_1057# a_n2061_n497# a_n865_n927#
+ a_1283_539# a_1225_n1963# a_807_n409# a_2061_627# a_29_n1015# a_n2119_1145# a_1225_1145#
+ a_n1643_539# a_389_n1445# a_n1225_n1015# a_447_2093# a_1643_2181# a_1225_n927# a_n2119_n927#
+ a_1701_n497# a_n1701_n1445# a_n1225_2093# a_n2119_627# a_447_1575# a_1643_1663#
+ a_2061_1145# a_n29_1145# a_29_539# a_n1225_1575# a_n1283_627# a_1701_21# a_2061_n927#
+ a_n389_2093# a_n807_21# a_1643_109# a_n29_n927# a_n2061_2093# a_n1283_2181# a_n447_2181#
+ a_n389_1575# a_865_n2569# a_n2061_1575# a_n1283_1663# a_n865_109# a_n447_1663# a_n29_627#
+ a_n2061_n2569# a_1701_2093# a_1283_21# a_1283_1057# a_n389_21# a_n389_n2569# a_807_n1445#
+ a_447_n2569# a_865_n2051# a_n1701_109# a_n2061_539# a_807_2181# a_1701_1575# a_n1701_n409#
+ a_389_1145# a_807_627# a_1643_n1445# a_865_n1533# a_1283_n2569# a_n2061_n2051# a_807_1663#
+ a_865_n497# a_n389_n2051# a_447_n2051# a_389_n927# a_n1643_n497# a_n2061_n1533#
+ a_n865_n409# a_n865_n2481# a_n807_n497# a_1225_n1445# a_447_n1533# a_n389_n1533#
+ w_n2257_n2691# a_2061_109# a_1283_n2051# a_n865_n1963# a_1283_n1533# a_n447_n2481#
+ a_1225_n409# a_n2119_n409# a_n2119_109# a_n2119_n2481# a_n807_n2569# a_447_1057#
+ a_1643_1145# a_n447_n1963# a_29_n497# a_n1225_1057# a_n1283_109# a_n2119_n1963#
+ a_865_2093# a_1643_n927# a_2061_n409# a_447_539# a_389_627# a_n29_n409# a_n1643_2093#
+ a_1701_n2569# a_n1283_n2481# a_n807_n2051# a_n807_2093# a_865_1575# a_n389_1057#
+ a_n1643_21# a_n1701_2181# a_n1643_1575# a_n2061_1057# a_n807_539# a_n1283_1145#
+ a_29_21# a_n1643_n2569# a_n807_1575# a_1225_627# a_n1283_n1963# a_n807_n1533# a_n29_109#
+ a_n29_n2481# a_1701_n2051# a_n447_1145# a_n1701_1663# a_n1283_n927# a_n865_2181#
+ a_29_n2569# a_n29_n1963# a_1701_n1533# a_n447_n927# a_1701_1057# a_2061_n2481# a_n447_627#
+ a_807_109# a_n1225_n2569# a_n1643_n2051# a_29_2093# a_865_n1015# a_n865_1663# a_2061_n1963#
+ a_807_1145# a_n1643_n1533# a_389_n409# a_29_1575# a_29_n2051# a_n2119_2181# a_1225_2181#
+ a_n1225_21# a_n2061_n1015# a_389_n2481# a_n1225_n2051# a_807_n927# a_447_n1015#
+ a_n389_n1015# a_29_n1533# a_n2119_1663# a_1225_1663# a_1283_n497# a_n1701_n2481#
+ a_389_n1963# a_n865_n1445# a_n1225_n1533# a_2061_2181# a_n389_539# a_1283_n1015#
+ a_865_539# a_865_21# a_n1701_n1963# a_n29_2181# a_2061_1663# a_n29_1663# a_n447_n1445#
+ a_n1225_539# a_n2119_n1445# a_1701_539# a_1643_627# a_1643_n409# a_389_109# a_865_1057#
+ a_1283_2093# a_n1643_1057# a_807_n2481#
X0 a_1643_n2481# a_1283_n2569# a_1225_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X1 a_807_2181# a_447_2093# a_389_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X2 a_n29_n2481# a_n389_n2569# a_n447_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X3 a_807_n409# a_447_n497# a_389_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X4 a_1643_1145# a_1283_1057# a_1225_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X5 a_389_n1445# a_29_n1533# a_n29_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X6 a_807_n927# a_447_n1015# a_389_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X7 a_1643_1663# a_1283_1575# a_1225_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X8 a_389_n1963# a_29_n2051# a_n29_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X9 a_n29_1145# a_n389_1057# a_n447_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X10 a_2061_2181# a_1701_2093# a_1643_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X11 a_2061_n1445# a_1701_n1533# a_1643_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X12 a_n29_1663# a_n389_1575# a_n447_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X13 a_n447_n1445# a_n807_n1533# a_n865_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X14 a_2061_n409# a_1701_n497# a_1643_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X15 a_n447_2181# a_n807_2093# a_n865_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X16 a_1225_n2481# a_865_n2569# a_807_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X17 a_2061_n1963# a_1701_n2051# a_1643_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X18 a_n447_n1963# a_n807_n2051# a_n865_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X19 a_2061_n927# a_1701_n1015# a_1643_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X20 a_n865_n2481# a_n1225_n2569# a_n1283_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X21 a_n447_n409# a_n807_n497# a_n865_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X22 a_n865_1145# a_n1225_1057# a_n1283_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X23 a_n447_n927# a_n807_n1015# a_n865_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X24 a_807_109# a_447_21# a_389_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X25 a_n865_1663# a_n1225_1575# a_n1283_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X26 a_807_627# a_447_539# a_389_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X27 a_1643_n1445# a_1283_n1533# a_1225_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X28 a_807_1145# a_447_1057# a_389_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X29 a_n29_n1445# a_n389_n1533# a_n447_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X30 a_1643_n1963# a_1283_n2051# a_1225_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X31 a_807_1663# a_447_1575# a_389_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X32 a_n29_n1963# a_n389_n2051# a_n447_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X33 a_2061_1145# a_1701_1057# a_1643_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X34 a_n1701_2181# a_n2061_2093# a_n2119_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X35 a_2061_1663# a_1701_1575# a_1643_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X36 a_1225_n1445# a_865_n1533# a_807_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X37 a_n1283_109# a_n1643_21# a_n1701_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X38 a_n447_1145# a_n807_1057# a_n865_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X39 a_n1701_n409# a_n2061_n497# a_n2119_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X40 a_1225_n1963# a_865_n2051# a_807_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X41 a_n1283_627# a_n1643_539# a_n1701_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X42 a_n447_1663# a_n807_1575# a_n865_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X43 a_n865_n1445# a_n1225_n1533# a_n1283_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X44 a_n1701_n927# a_n2061_n1015# a_n2119_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X45 a_n865_n1963# a_n1225_n2051# a_n1283_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X46 a_n1283_2181# a_n1643_2093# a_n1701_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X47 a_n1701_n2481# a_n2061_n2569# a_n2119_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X48 a_n1283_n409# a_n1643_n497# a_n1701_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X49 a_n1283_n927# a_n1643_n1015# a_n1701_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X50 a_389_109# a_29_21# a_n29_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X51 a_1225_2181# a_865_2093# a_807_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X52 a_389_627# a_29_539# a_n29_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X53 a_1225_n409# a_865_n497# a_807_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X54 a_1225_n927# a_865_n1015# a_807_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X55 a_807_n2481# a_447_n2569# a_389_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X56 a_n1701_1145# a_n2061_1057# a_n2119_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X57 a_389_2181# a_29_2093# a_n29_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X58 a_n1701_1663# a_n2061_1575# a_n2119_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X59 a_n29_109# a_n389_21# a_n447_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X60 a_n1283_n2481# a_n1643_n2569# a_n1701_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X61 a_389_n409# a_29_n497# a_n29_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X62 a_n29_627# a_n389_539# a_n447_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X63 a_389_n927# a_29_n1015# a_n29_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X64 a_n447_109# a_n807_21# a_n865_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X65 a_n1701_109# a_n2061_21# a_n2119_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X66 a_n1283_1145# a_n1643_1057# a_n1701_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X67 a_n1701_n1445# a_n2061_n1533# a_n2119_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X68 a_n447_627# a_n807_539# a_n865_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X69 a_1225_109# a_865_21# a_807_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X70 a_n1701_627# a_n2061_539# a_n2119_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X71 a_n1283_1663# a_n1643_1575# a_n1701_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X72 a_1643_2181# a_1283_2093# a_1225_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X73 a_n1701_n1963# a_n2061_n2051# a_n2119_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=1.8e+06u
X74 a_389_n2481# a_29_n2569# a_n29_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X75 a_1225_627# a_865_539# a_807_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X76 a_1643_n409# a_1283_n497# a_1225_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X77 a_1225_1145# a_865_1057# a_807_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X78 a_n29_2181# a_n389_2093# a_n447_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X79 a_1643_n927# a_1283_n1015# a_1225_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X80 a_n865_109# a_n1225_21# a_n1283_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X81 a_2061_n2481# a_1701_n2569# a_1643_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X82 a_1225_1663# a_865_1575# a_807_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X83 a_n29_n409# a_n389_n497# a_n447_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X84 a_n447_n2481# a_n807_n2569# a_n865_n2481# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X85 a_n865_627# a_n1225_539# a_n1283_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X86 a_n29_n927# a_n389_n1015# a_n447_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X87 a_1643_109# a_1283_21# a_1225_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X88 a_807_n1445# a_447_n1533# a_389_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X89 a_n865_2181# a_n1225_2093# a_n1283_2181# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X90 a_1643_627# a_1283_539# a_1225_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X91 a_389_1145# a_29_1057# a_n29_1145# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X92 a_807_n1963# a_447_n2051# a_389_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X93 a_2061_109# a_1701_21# a_1643_109# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X94 a_389_1663# a_29_1575# a_n29_1663# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X95 a_n1283_n1445# a_n1643_n1533# a_n1701_n1445# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X96 a_n865_n409# a_n1225_n497# a_n1283_n409# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X97 a_2061_627# a_1701_539# a_1643_627# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X98 a_n1283_n1963# a_n1643_n2051# a_n1701_n1963# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
X99 a_n865_n927# a_n1225_n1015# a_n1283_n927# w_n2257_n2691# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=1.8e+06u
.ends

.subckt output vss vout vdd vin
Xsky130_fd_pr__cap_mim_m3_1_6BP6N2_0 vss vout vout net1 vout net1 net1 sky130_fd_pr__cap_mim_m3_1_6BP6N2
Xsky130_fd_pr__nfet_01v8_RE4H9G_0 vin vin vin vin vin vss vin vin vin vin vss vin
+ vout vss vin vout vin vin vout vin vout vin vout vout vss vin vout vss vss vss vin
+ vout vin vout vin vin vss vss vin vin vss vss vout vss vin vin vss vin vin vin vss
+ vout vout vss vin vss vss vout vss vss vout vin vin vss vin vss vin vin vin vss
+ vin vin vin vout vss vss vin vout vin vin vss vin vss vout vin vss vin vout vout
+ vout vss vin vss vout vout vout vout vin vin vin vin vout vin vin vss vss vin vin
+ vss vin vin vin vout vout vout vin vin vout vin vin vin vin vout vss vout vin vin
+ vin vin vout vout vss vout vin vin vss vout vss vss vin vout vss vout vin vss vout
+ vin vout vss vss vin vout vin vin vss vss vin vin vss vss vin vss vin vout vin vss
+ vss vin vin vin vin vin vin vout vout vout vout vss vin vout vss vss vout vin vss
+ vin vss vss vin vin vin vin vss vin vout vin vss vss vss vin vin vin vin vin vin
+ vin vss vin vin vin vin vout vout vout vout vout vin vout vin vin vout vss vin vin
+ vin vin vss vin vin vout vin vin vout vin vin vin vss vss vout vout vin vin vin
+ vin vout vin vin vin vout vss vss vin vin vin vout vout vin vout vin vin vout vin
+ vin vin vin vin vin vin vss vin vin vin vout vss vin vin vss vss vin vss vin vin
+ vss vout vin vin vin vout vss vout vin vin vin vout vss vout vout vin vss vss vss
+ vin vss vin vin vin vss vout vss vout vss vss vin vin vin vss vin vin vss vin vss
+ vout vss vin vin vout vout vout vss vss vin vin vss vss vin vout vin vin vin vout
+ vss vin vin vin vin vin vin vss vin vin vss vin vin vin vss vin vout vin vin vin
+ vout vout vout vout vout vout vin vout vin vin vout vout vout vss vout vss vin vss
+ vout vss vin vout vss vout vin vin vout vout vin vss vss vout vss vin vin vss vout
+ vss vss vout vin vss vss vin vout vin vin vin vout vout vout vout vin vss vin vss
+ vin vout vin vss vin vss vss vin vin vss vin vin vout vss vss vin vss vss vss vss
+ vss vss vin vout vin vin vout vin vout vin vss vin vin vin vin vin vin vss vin vout
+ vss vin vout vin vss vin vout vin vss vin vin vin vin vss vss vin vin vin vin vout
+ vin vin vout vout vout vin vout vin vin vout vout sky130_fd_pr__nfet_01v8_RE4H9G
Xsky130_fd_pr__nfet_01v8_B8HNLY_0 net1 vdd vin vin vdd vdd vdd net1 vdd net1 vin vin
+ vdd net1 net1 vdd net1 vdd vin net1 vin vin net1 net1 vin vdd vin vdd vdd vdd net1
+ vdd vin net1 vin vdd vin vin vdd vin vdd vdd net1 vin vin vdd net1 vdd vin vdd net1
+ vin net1 vdd vdd vin vdd vin vdd vdd net1 net1 vdd vin vin vdd vdd vdd vin net1
+ vin net1 vdd vdd vdd vdd vdd vdd net1 vdd vdd net1 vdd net1 vdd net1 vin net1 net1
+ vdd vdd vdd net1 vdd vdd vdd vin vdd vdd net1 net1 vdd vin vdd vdd vss vin vdd net1
+ vdd vin vin vin vin vin vdd vdd net1 vin vdd vdd vin vin vdd net1 vin vdd vin net1
+ vdd vdd vin vdd vdd vdd vdd vdd net1 vdd vdd vdd vin vdd vdd vdd vin vin vdd net1
+ net1 vdd vin net1 vin net1 vdd net1 vdd vin vdd vin vin net1 vdd vdd vdd vdd net1
+ vin net1 vdd vin vdd vdd vin vin vdd vdd vin vdd net1 vdd vdd vdd vin vin vdd net1
+ vin net1 vdd vin vdd vdd vdd vdd net1 net1 vin net1 vin vdd vin vdd net1 net1 vin
+ vdd vdd vdd net1 sky130_fd_pr__nfet_01v8_B8HNLY
.ends

.subckt sky130_fd_pr__pfet_01v8_9CZQJE VSUBS a_n267_n637# a_n29_n540# a_1007_n540#
+ a_n1509_n540# a_n1007_n637# a_n711_n637# a_1451_n540# a_n473_n540# a_n1451_n637#
+ a_917_n637# a_267_n540# a_n1213_n540# a_711_n540# a_n859_n637# a_1361_n637# a_177_n637#
+ a_n119_n637# a_621_n637# a_n563_n637# a_859_n540# a_1303_n540# a_n1303_n637# a_n325_n540#
+ a_119_n540# a_29_n637# a_769_n637# a_1213_n637# a_n1065_n540# a_563_n540# a_n917_n540#
+ a_473_n637# a_n415_n637# a_1155_n540# a_n177_n540# a_n1155_n637# a_n621_n540# a_415_n540#
+ a_1065_n637# a_n1361_n540# w_n1647_n759# a_325_n637# a_n769_n540#
X0 a_n917_n540# a_n1007_n637# a_n1065_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X1 a_n473_n540# a_n563_n637# a_n621_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X2 a_n177_n540# a_n267_n637# a_n325_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X3 a_711_n540# a_621_n637# a_563_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X4 a_1303_n540# a_1213_n637# a_1155_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X5 a_415_n540# a_325_n637# a_267_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X6 a_859_n540# a_769_n637# a_711_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=0p ps=0u w=5.4e+06u l=450000u
X7 a_n621_n540# a_n711_n637# a_n769_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X8 a_n325_n540# a_n415_n637# a_n473_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
X9 a_n769_n540# a_n859_n637# a_n917_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
X10 a_n1361_n540# a_n1451_n637# a_n1509_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X11 a_n29_n540# a_n119_n637# a_n177_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=0p ps=0u w=5.4e+06u l=450000u
X12 a_n1065_n540# a_n1155_n637# a_n1213_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.566e+12p ps=1.138e+07u w=5.4e+06u l=450000u
X13 a_119_n540# a_29_n637# a_n29_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=0p ps=0u w=5.4e+06u l=450000u
X14 a_1007_n540# a_917_n637# a_859_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=0p ps=0u w=5.4e+06u l=450000u
X15 a_1451_n540# a_1361_n637# a_1303_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=1.566e+12p pd=1.138e+07u as=0p ps=0u w=5.4e+06u l=450000u
X16 a_563_n540# a_473_n637# a_415_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
X17 a_1155_n540# a_1065_n637# a_1007_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
X18 a_n1213_n540# a_n1303_n637# a_n1361_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
X19 a_267_n540# a_177_n637# a_119_n540# w_n1647_n759# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.4e+06u l=450000u
.ends

.subckt mirror VSUBS idif iout iref vdd
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[0|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[1|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[2|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[3|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[4|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[5|0] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[0|1] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[1|1] VSUBS iref vdd vdd vdd iref iref vdd vdd iref
+ iref vdd vdd vdd iref iref iref iref iref iref vdd vdd iref vdd vdd iref iref iref
+ vdd vdd vdd iref iref vdd vdd iref vdd vdd iref vdd vdd iref vdd sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[2|1] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[3|1] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[4|1] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[5|1] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[0|2] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[1|2] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[2|2] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[3|2] VSUBS iref vdd iref vdd iref iref vdd iref
+ iref iref vdd vdd iref iref iref iref iref iref iref vdd iref iref vdd iref iref
+ iref iref iref vdd vdd iref iref vdd iref iref vdd iref iref iref vdd iref iref
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[4|2] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[5|2] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[0|3] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[1|3] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[2|3] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[3|3] VSUBS iref vdd idif vdd iref iref vdd idif
+ iref iref vdd vdd idif iref iref iref iref iref iref vdd idif iref vdd idif iref
+ iref iref idif vdd vdd iref iref vdd idif iref vdd idif iref idif vdd iref idif
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[4|3] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[5|3] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[0|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[1|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[2|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[3|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[4|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
Xsky130_fd_pr__pfet_01v8_9CZQJE_0[5|4] VSUBS iref vdd iout vdd iref iref vdd iout
+ iref iref vdd vdd iout iref iref iref iref iref iref vdd iout iref vdd iout iref
+ iref iref iout vdd vdd iref iref vdd iout iref vdd iout iref iout vdd iref iout
+ sky130_fd_pr__pfet_01v8_9CZQJE
.ends

.subckt opamp_ramiro vss vin_n vin_p iref vdd output_0/vout
Xinput_0 vss vin_n vin_p input_0/iref output_0/vin input
Xoutput_0 vss output_0/vout vdd output_0/vin output
Xmirror_0 vss input_0/iref output_0/vout iref vdd mirror
.ends

Xopamp_lucas_0 m2_115869_595817# io_analog[8] io_analog[9] opamp_lucas_0/iref io_analog[10]
+ vssa1 opamp_lucas_0/vdd opamp_lucas
Xopamp_manuel_0 io_analog[3] io_analog[2] opamp_manuel_0/iref io_clamp_low[0] opamp_lucas_0/vdd
+ vssa1 opamp_manuel
Xbias_circuit_0 vssa1 io_analog[1] opamp_lucas_0/vdd opamp_lucas_0/iref opamp_ramiro_0/iref
+ opamp_manuel_0/iref bias_circuit
Xopamp_ramiro_0 vssa1 io_clamp_low[2] io_analog[7] opamp_ramiro_0/iref opamp_lucas_0/vdd
+ io_clamp_low[1] opamp_ramiro
.end

