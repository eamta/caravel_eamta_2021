magic
tech sky130A
timestamp 1620674245
<< nwell >>
rect 353 215 878 404
<< nmos >>
rect 400 14 415 59
rect 500 13 515 103
rect 544 13 559 103
rect 671 13 686 103
rect 715 13 730 103
rect 816 14 831 59
<< pmos >>
rect 400 233 415 323
rect 500 233 515 323
rect 544 233 559 323
rect 671 233 686 323
rect 715 233 730 323
rect 816 233 831 323
<< ndiff >>
rect 371 44 400 59
rect 371 27 377 44
rect 394 27 400 44
rect 371 14 400 27
rect 415 44 444 59
rect 415 27 421 44
rect 438 27 444 44
rect 415 14 444 27
rect 471 44 500 103
rect 471 27 477 44
rect 494 27 500 44
rect 471 13 500 27
rect 515 44 544 103
rect 515 27 521 44
rect 538 27 544 44
rect 515 13 544 27
rect 559 44 588 103
rect 559 27 565 44
rect 582 27 588 44
rect 559 13 588 27
rect 642 44 671 103
rect 642 27 648 44
rect 665 27 671 44
rect 642 13 671 27
rect 686 13 715 103
rect 730 44 759 103
rect 730 27 736 44
rect 753 27 759 44
rect 730 13 759 27
rect 787 44 816 59
rect 787 27 793 44
rect 810 27 816 44
rect 787 14 816 27
rect 831 44 860 59
rect 831 27 837 44
rect 854 27 860 44
rect 831 14 860 27
<< pdiff >>
rect 371 309 400 323
rect 371 292 377 309
rect 394 292 400 309
rect 371 233 400 292
rect 415 309 444 323
rect 415 292 421 309
rect 438 292 444 309
rect 415 233 444 292
rect 471 309 500 323
rect 471 292 477 309
rect 494 292 500 309
rect 471 233 500 292
rect 515 309 544 323
rect 515 292 521 309
rect 538 292 544 309
rect 515 233 544 292
rect 559 309 588 323
rect 559 292 565 309
rect 582 292 588 309
rect 559 233 588 292
rect 642 309 671 323
rect 642 292 648 309
rect 665 292 671 309
rect 642 233 671 292
rect 686 309 715 323
rect 686 292 692 309
rect 709 292 715 309
rect 686 233 715 292
rect 730 309 759 323
rect 730 292 736 309
rect 753 292 759 309
rect 730 233 759 292
rect 787 309 816 323
rect 787 292 793 309
rect 810 292 816 309
rect 787 233 816 292
rect 831 309 860 323
rect 831 292 837 309
rect 854 292 860 309
rect 831 233 860 292
<< ndiffc >>
rect 377 27 394 44
rect 421 27 438 44
rect 477 27 494 44
rect 521 27 538 44
rect 565 27 582 44
rect 648 27 665 44
rect 736 27 753 44
rect 793 27 810 44
rect 837 27 854 44
<< pdiffc >>
rect 377 292 394 309
rect 421 292 438 309
rect 477 292 494 309
rect 521 292 538 309
rect 565 292 582 309
rect 648 292 665 309
rect 692 292 709 309
rect 736 292 753 309
rect 793 292 810 309
rect 837 292 854 309
<< psubdiff >>
rect 381 -32 393 -15
rect 839 -32 851 -15
<< nsubdiff >>
rect 381 368 393 385
rect 838 368 850 385
<< psubdiffcont >>
rect 393 -32 839 -15
<< nsubdiffcont >>
rect 393 368 838 385
<< poly >>
rect 400 323 415 336
rect 500 323 515 336
rect 544 323 559 336
rect 671 323 686 336
rect 715 323 730 336
rect 816 323 831 336
rect 598 309 631 316
rect 598 292 606 309
rect 623 292 631 309
rect 598 283 631 292
rect 400 144 415 233
rect 500 215 515 233
rect 485 207 519 215
rect 485 190 495 207
rect 510 190 519 207
rect 485 182 519 190
rect 400 136 461 144
rect 400 119 437 136
rect 452 119 461 136
rect 400 111 461 119
rect 400 59 415 111
rect 500 103 515 182
rect 544 179 559 233
rect 540 171 573 179
rect 540 154 549 171
rect 565 154 573 171
rect 540 146 573 154
rect 544 103 559 146
rect 400 1 415 14
rect 606 52 623 283
rect 671 215 686 233
rect 661 207 694 215
rect 661 190 669 207
rect 686 190 694 207
rect 661 182 694 190
rect 671 103 686 182
rect 715 144 730 233
rect 816 215 831 233
rect 783 207 831 215
rect 783 190 791 207
rect 808 190 831 207
rect 783 182 831 190
rect 707 136 739 144
rect 707 119 715 136
rect 731 119 739 136
rect 707 111 739 119
rect 715 103 730 111
rect 598 45 631 52
rect 598 27 606 45
rect 623 27 631 45
rect 598 19 631 27
rect 816 59 831 182
rect 500 0 515 13
rect 544 0 559 13
rect 671 0 686 13
rect 715 0 730 13
rect 816 1 831 14
<< polycont >>
rect 606 292 623 309
rect 495 190 510 207
rect 437 119 452 136
rect 549 154 565 171
rect 669 190 686 207
rect 791 190 808 207
rect 715 119 731 136
rect 606 27 623 45
<< locali >>
rect 377 368 393 385
rect 838 368 846 385
rect 377 309 394 317
rect 377 207 394 292
rect 421 309 438 368
rect 421 284 438 292
rect 477 309 494 317
rect 477 267 494 292
rect 521 309 538 368
rect 606 334 753 351
rect 521 284 538 292
rect 565 309 582 317
rect 565 267 582 292
rect 606 309 623 334
rect 606 284 623 292
rect 648 309 665 334
rect 648 284 665 292
rect 692 309 709 317
rect 692 267 709 292
rect 736 309 753 334
rect 736 284 753 292
rect 793 309 810 368
rect 793 284 810 292
rect 837 309 854 317
rect 477 250 709 267
rect 377 190 495 207
rect 510 190 520 207
rect 661 190 669 207
rect 686 190 791 207
rect 808 190 816 207
rect 377 44 394 190
rect 837 171 854 292
rect 540 154 549 171
rect 565 154 854 171
rect 427 119 437 136
rect 452 119 714 136
rect 731 119 739 136
rect 377 19 394 27
rect 421 44 438 52
rect 421 -15 438 27
rect 477 44 494 52
rect 477 -15 494 27
rect 521 44 544 52
rect 538 27 544 44
rect 521 19 544 27
rect 565 45 665 52
rect 565 44 606 45
rect 582 27 606 44
rect 623 44 665 45
rect 623 27 648 44
rect 565 19 665 27
rect 736 44 753 52
rect 736 -15 753 27
rect 793 44 810 52
rect 793 -15 810 27
rect 837 44 854 154
rect 837 19 854 27
rect 377 -32 393 -15
rect 839 -32 847 -15
<< viali >>
rect 393 368 838 385
rect 669 190 686 207
rect 714 119 715 136
rect 715 119 731 136
rect 606 27 623 45
rect 393 -32 838 -15
<< metal1 >>
rect 353 385 878 404
rect 353 368 393 385
rect 838 368 878 385
rect 353 349 878 368
rect 661 207 694 215
rect 661 190 669 207
rect 686 190 694 207
rect 661 182 694 190
rect 707 136 739 144
rect 707 119 714 136
rect 731 119 739 136
rect 707 111 739 119
rect 598 45 631 52
rect 598 27 606 45
rect 623 27 631 45
rect 598 19 631 27
rect 353 -15 878 4
rect 353 -32 393 -15
rect 838 -32 878 -15
rect 353 -51 878 -32
<< labels >>
rlabel metal1 598 19 631 27 5 Z
rlabel metal1 614 404 614 404 1 VDD
rlabel metal1 614 -51 614 -51 5 VSS
rlabel metal1 723 111 723 111 5 B
rlabel metal1 661 182 694 190 5 A
<< end >>
