magic
tech sky130A
magscale 1 2
timestamp 1615920820
<< error_p >>
rect -4223 18 4223 236
<< nwell >>
rect -4223 18 4223 1618
rect -4223 -1618 4223 -18
<< pmos >>
rect -4129 118 -3989 1518
rect -3931 118 -3791 1518
rect -3733 118 -3593 1518
rect -3535 118 -3395 1518
rect -3337 118 -3197 1518
rect -3139 118 -2999 1518
rect -2941 118 -2801 1518
rect -2743 118 -2603 1518
rect -2545 118 -2405 1518
rect -2347 118 -2207 1518
rect -2149 118 -2009 1518
rect -1951 118 -1811 1518
rect -1753 118 -1613 1518
rect -1555 118 -1415 1518
rect -1357 118 -1217 1518
rect -1159 118 -1019 1518
rect -961 118 -821 1518
rect -763 118 -623 1518
rect -565 118 -425 1518
rect -367 118 -227 1518
rect -169 118 -29 1518
rect 29 118 169 1518
rect 227 118 367 1518
rect 425 118 565 1518
rect 623 118 763 1518
rect 821 118 961 1518
rect 1019 118 1159 1518
rect 1217 118 1357 1518
rect 1415 118 1555 1518
rect 1613 118 1753 1518
rect 1811 118 1951 1518
rect 2009 118 2149 1518
rect 2207 118 2347 1518
rect 2405 118 2545 1518
rect 2603 118 2743 1518
rect 2801 118 2941 1518
rect 2999 118 3139 1518
rect 3197 118 3337 1518
rect 3395 118 3535 1518
rect 3593 118 3733 1518
rect 3791 118 3931 1518
rect 3989 118 4129 1518
rect -4129 -1518 -3989 -118
rect -3931 -1518 -3791 -118
rect -3733 -1518 -3593 -118
rect -3535 -1518 -3395 -118
rect -3337 -1518 -3197 -118
rect -3139 -1518 -2999 -118
rect -2941 -1518 -2801 -118
rect -2743 -1518 -2603 -118
rect -2545 -1518 -2405 -118
rect -2347 -1518 -2207 -118
rect -2149 -1518 -2009 -118
rect -1951 -1518 -1811 -118
rect -1753 -1518 -1613 -118
rect -1555 -1518 -1415 -118
rect -1357 -1518 -1217 -118
rect -1159 -1518 -1019 -118
rect -961 -1518 -821 -118
rect -763 -1518 -623 -118
rect -565 -1518 -425 -118
rect -367 -1518 -227 -118
rect -169 -1518 -29 -118
rect 29 -1518 169 -118
rect 227 -1518 367 -118
rect 425 -1518 565 -118
rect 623 -1518 763 -118
rect 821 -1518 961 -118
rect 1019 -1518 1159 -118
rect 1217 -1518 1357 -118
rect 1415 -1518 1555 -118
rect 1613 -1518 1753 -118
rect 1811 -1518 1951 -118
rect 2009 -1518 2149 -118
rect 2207 -1518 2347 -118
rect 2405 -1518 2545 -118
rect 2603 -1518 2743 -118
rect 2801 -1518 2941 -118
rect 2999 -1518 3139 -118
rect 3197 -1518 3337 -118
rect 3395 -1518 3535 -118
rect 3593 -1518 3733 -118
rect 3791 -1518 3931 -118
rect 3989 -1518 4129 -118
<< pdiff >>
rect -4187 1506 -4129 1518
rect -4187 130 -4175 1506
rect -4141 130 -4129 1506
rect -4187 118 -4129 130
rect -3989 1506 -3931 1518
rect -3989 130 -3977 1506
rect -3943 130 -3931 1506
rect -3989 118 -3931 130
rect -3791 1506 -3733 1518
rect -3791 130 -3779 1506
rect -3745 130 -3733 1506
rect -3791 118 -3733 130
rect -3593 1506 -3535 1518
rect -3593 130 -3581 1506
rect -3547 130 -3535 1506
rect -3593 118 -3535 130
rect -3395 1506 -3337 1518
rect -3395 130 -3383 1506
rect -3349 130 -3337 1506
rect -3395 118 -3337 130
rect -3197 1506 -3139 1518
rect -3197 130 -3185 1506
rect -3151 130 -3139 1506
rect -3197 118 -3139 130
rect -2999 1506 -2941 1518
rect -2999 130 -2987 1506
rect -2953 130 -2941 1506
rect -2999 118 -2941 130
rect -2801 1506 -2743 1518
rect -2801 130 -2789 1506
rect -2755 130 -2743 1506
rect -2801 118 -2743 130
rect -2603 1506 -2545 1518
rect -2603 130 -2591 1506
rect -2557 130 -2545 1506
rect -2603 118 -2545 130
rect -2405 1506 -2347 1518
rect -2405 130 -2393 1506
rect -2359 130 -2347 1506
rect -2405 118 -2347 130
rect -2207 1506 -2149 1518
rect -2207 130 -2195 1506
rect -2161 130 -2149 1506
rect -2207 118 -2149 130
rect -2009 1506 -1951 1518
rect -2009 130 -1997 1506
rect -1963 130 -1951 1506
rect -2009 118 -1951 130
rect -1811 1506 -1753 1518
rect -1811 130 -1799 1506
rect -1765 130 -1753 1506
rect -1811 118 -1753 130
rect -1613 1506 -1555 1518
rect -1613 130 -1601 1506
rect -1567 130 -1555 1506
rect -1613 118 -1555 130
rect -1415 1506 -1357 1518
rect -1415 130 -1403 1506
rect -1369 130 -1357 1506
rect -1415 118 -1357 130
rect -1217 1506 -1159 1518
rect -1217 130 -1205 1506
rect -1171 130 -1159 1506
rect -1217 118 -1159 130
rect -1019 1506 -961 1518
rect -1019 130 -1007 1506
rect -973 130 -961 1506
rect -1019 118 -961 130
rect -821 1506 -763 1518
rect -821 130 -809 1506
rect -775 130 -763 1506
rect -821 118 -763 130
rect -623 1506 -565 1518
rect -623 130 -611 1506
rect -577 130 -565 1506
rect -623 118 -565 130
rect -425 1506 -367 1518
rect -425 130 -413 1506
rect -379 130 -367 1506
rect -425 118 -367 130
rect -227 1506 -169 1518
rect -227 130 -215 1506
rect -181 130 -169 1506
rect -227 118 -169 130
rect -29 1506 29 1518
rect -29 130 -17 1506
rect 17 130 29 1506
rect -29 118 29 130
rect 169 1506 227 1518
rect 169 130 181 1506
rect 215 130 227 1506
rect 169 118 227 130
rect 367 1506 425 1518
rect 367 130 379 1506
rect 413 130 425 1506
rect 367 118 425 130
rect 565 1506 623 1518
rect 565 130 577 1506
rect 611 130 623 1506
rect 565 118 623 130
rect 763 1506 821 1518
rect 763 130 775 1506
rect 809 130 821 1506
rect 763 118 821 130
rect 961 1506 1019 1518
rect 961 130 973 1506
rect 1007 130 1019 1506
rect 961 118 1019 130
rect 1159 1506 1217 1518
rect 1159 130 1171 1506
rect 1205 130 1217 1506
rect 1159 118 1217 130
rect 1357 1506 1415 1518
rect 1357 130 1369 1506
rect 1403 130 1415 1506
rect 1357 118 1415 130
rect 1555 1506 1613 1518
rect 1555 130 1567 1506
rect 1601 130 1613 1506
rect 1555 118 1613 130
rect 1753 1506 1811 1518
rect 1753 130 1765 1506
rect 1799 130 1811 1506
rect 1753 118 1811 130
rect 1951 1506 2009 1518
rect 1951 130 1963 1506
rect 1997 130 2009 1506
rect 1951 118 2009 130
rect 2149 1506 2207 1518
rect 2149 130 2161 1506
rect 2195 130 2207 1506
rect 2149 118 2207 130
rect 2347 1506 2405 1518
rect 2347 130 2359 1506
rect 2393 130 2405 1506
rect 2347 118 2405 130
rect 2545 1506 2603 1518
rect 2545 130 2557 1506
rect 2591 130 2603 1506
rect 2545 118 2603 130
rect 2743 1506 2801 1518
rect 2743 130 2755 1506
rect 2789 130 2801 1506
rect 2743 118 2801 130
rect 2941 1506 2999 1518
rect 2941 130 2953 1506
rect 2987 130 2999 1506
rect 2941 118 2999 130
rect 3139 1506 3197 1518
rect 3139 130 3151 1506
rect 3185 130 3197 1506
rect 3139 118 3197 130
rect 3337 1506 3395 1518
rect 3337 130 3349 1506
rect 3383 130 3395 1506
rect 3337 118 3395 130
rect 3535 1506 3593 1518
rect 3535 130 3547 1506
rect 3581 130 3593 1506
rect 3535 118 3593 130
rect 3733 1506 3791 1518
rect 3733 130 3745 1506
rect 3779 130 3791 1506
rect 3733 118 3791 130
rect 3931 1506 3989 1518
rect 3931 130 3943 1506
rect 3977 130 3989 1506
rect 3931 118 3989 130
rect 4129 1506 4187 1518
rect 4129 130 4141 1506
rect 4175 130 4187 1506
rect 4129 118 4187 130
rect -4187 -130 -4129 -118
rect -4187 -1506 -4175 -130
rect -4141 -1506 -4129 -130
rect -4187 -1518 -4129 -1506
rect -3989 -130 -3931 -118
rect -3989 -1506 -3977 -130
rect -3943 -1506 -3931 -130
rect -3989 -1518 -3931 -1506
rect -3791 -130 -3733 -118
rect -3791 -1506 -3779 -130
rect -3745 -1506 -3733 -130
rect -3791 -1518 -3733 -1506
rect -3593 -130 -3535 -118
rect -3593 -1506 -3581 -130
rect -3547 -1506 -3535 -130
rect -3593 -1518 -3535 -1506
rect -3395 -130 -3337 -118
rect -3395 -1506 -3383 -130
rect -3349 -1506 -3337 -130
rect -3395 -1518 -3337 -1506
rect -3197 -130 -3139 -118
rect -3197 -1506 -3185 -130
rect -3151 -1506 -3139 -130
rect -3197 -1518 -3139 -1506
rect -2999 -130 -2941 -118
rect -2999 -1506 -2987 -130
rect -2953 -1506 -2941 -130
rect -2999 -1518 -2941 -1506
rect -2801 -130 -2743 -118
rect -2801 -1506 -2789 -130
rect -2755 -1506 -2743 -130
rect -2801 -1518 -2743 -1506
rect -2603 -130 -2545 -118
rect -2603 -1506 -2591 -130
rect -2557 -1506 -2545 -130
rect -2603 -1518 -2545 -1506
rect -2405 -130 -2347 -118
rect -2405 -1506 -2393 -130
rect -2359 -1506 -2347 -130
rect -2405 -1518 -2347 -1506
rect -2207 -130 -2149 -118
rect -2207 -1506 -2195 -130
rect -2161 -1506 -2149 -130
rect -2207 -1518 -2149 -1506
rect -2009 -130 -1951 -118
rect -2009 -1506 -1997 -130
rect -1963 -1506 -1951 -130
rect -2009 -1518 -1951 -1506
rect -1811 -130 -1753 -118
rect -1811 -1506 -1799 -130
rect -1765 -1506 -1753 -130
rect -1811 -1518 -1753 -1506
rect -1613 -130 -1555 -118
rect -1613 -1506 -1601 -130
rect -1567 -1506 -1555 -130
rect -1613 -1518 -1555 -1506
rect -1415 -130 -1357 -118
rect -1415 -1506 -1403 -130
rect -1369 -1506 -1357 -130
rect -1415 -1518 -1357 -1506
rect -1217 -130 -1159 -118
rect -1217 -1506 -1205 -130
rect -1171 -1506 -1159 -130
rect -1217 -1518 -1159 -1506
rect -1019 -130 -961 -118
rect -1019 -1506 -1007 -130
rect -973 -1506 -961 -130
rect -1019 -1518 -961 -1506
rect -821 -130 -763 -118
rect -821 -1506 -809 -130
rect -775 -1506 -763 -130
rect -821 -1518 -763 -1506
rect -623 -130 -565 -118
rect -623 -1506 -611 -130
rect -577 -1506 -565 -130
rect -623 -1518 -565 -1506
rect -425 -130 -367 -118
rect -425 -1506 -413 -130
rect -379 -1506 -367 -130
rect -425 -1518 -367 -1506
rect -227 -130 -169 -118
rect -227 -1506 -215 -130
rect -181 -1506 -169 -130
rect -227 -1518 -169 -1506
rect -29 -130 29 -118
rect -29 -1506 -17 -130
rect 17 -1506 29 -130
rect -29 -1518 29 -1506
rect 169 -130 227 -118
rect 169 -1506 181 -130
rect 215 -1506 227 -130
rect 169 -1518 227 -1506
rect 367 -130 425 -118
rect 367 -1506 379 -130
rect 413 -1506 425 -130
rect 367 -1518 425 -1506
rect 565 -130 623 -118
rect 565 -1506 577 -130
rect 611 -1506 623 -130
rect 565 -1518 623 -1506
rect 763 -130 821 -118
rect 763 -1506 775 -130
rect 809 -1506 821 -130
rect 763 -1518 821 -1506
rect 961 -130 1019 -118
rect 961 -1506 973 -130
rect 1007 -1506 1019 -130
rect 961 -1518 1019 -1506
rect 1159 -130 1217 -118
rect 1159 -1506 1171 -130
rect 1205 -1506 1217 -130
rect 1159 -1518 1217 -1506
rect 1357 -130 1415 -118
rect 1357 -1506 1369 -130
rect 1403 -1506 1415 -130
rect 1357 -1518 1415 -1506
rect 1555 -130 1613 -118
rect 1555 -1506 1567 -130
rect 1601 -1506 1613 -130
rect 1555 -1518 1613 -1506
rect 1753 -130 1811 -118
rect 1753 -1506 1765 -130
rect 1799 -1506 1811 -130
rect 1753 -1518 1811 -1506
rect 1951 -130 2009 -118
rect 1951 -1506 1963 -130
rect 1997 -1506 2009 -130
rect 1951 -1518 2009 -1506
rect 2149 -130 2207 -118
rect 2149 -1506 2161 -130
rect 2195 -1506 2207 -130
rect 2149 -1518 2207 -1506
rect 2347 -130 2405 -118
rect 2347 -1506 2359 -130
rect 2393 -1506 2405 -130
rect 2347 -1518 2405 -1506
rect 2545 -130 2603 -118
rect 2545 -1506 2557 -130
rect 2591 -1506 2603 -130
rect 2545 -1518 2603 -1506
rect 2743 -130 2801 -118
rect 2743 -1506 2755 -130
rect 2789 -1506 2801 -130
rect 2743 -1518 2801 -1506
rect 2941 -130 2999 -118
rect 2941 -1506 2953 -130
rect 2987 -1506 2999 -130
rect 2941 -1518 2999 -1506
rect 3139 -130 3197 -118
rect 3139 -1506 3151 -130
rect 3185 -1506 3197 -130
rect 3139 -1518 3197 -1506
rect 3337 -130 3395 -118
rect 3337 -1506 3349 -130
rect 3383 -1506 3395 -130
rect 3337 -1518 3395 -1506
rect 3535 -130 3593 -118
rect 3535 -1506 3547 -130
rect 3581 -1506 3593 -130
rect 3535 -1518 3593 -1506
rect 3733 -130 3791 -118
rect 3733 -1506 3745 -130
rect 3779 -1506 3791 -130
rect 3733 -1518 3791 -1506
rect 3931 -130 3989 -118
rect 3931 -1506 3943 -130
rect 3977 -1506 3989 -130
rect 3931 -1518 3989 -1506
rect 4129 -130 4187 -118
rect 4129 -1506 4141 -130
rect 4175 -1506 4187 -130
rect 4129 -1518 4187 -1506
<< pdiffc >>
rect -4175 130 -4141 1506
rect -3977 130 -3943 1506
rect -3779 130 -3745 1506
rect -3581 130 -3547 1506
rect -3383 130 -3349 1506
rect -3185 130 -3151 1506
rect -2987 130 -2953 1506
rect -2789 130 -2755 1506
rect -2591 130 -2557 1506
rect -2393 130 -2359 1506
rect -2195 130 -2161 1506
rect -1997 130 -1963 1506
rect -1799 130 -1765 1506
rect -1601 130 -1567 1506
rect -1403 130 -1369 1506
rect -1205 130 -1171 1506
rect -1007 130 -973 1506
rect -809 130 -775 1506
rect -611 130 -577 1506
rect -413 130 -379 1506
rect -215 130 -181 1506
rect -17 130 17 1506
rect 181 130 215 1506
rect 379 130 413 1506
rect 577 130 611 1506
rect 775 130 809 1506
rect 973 130 1007 1506
rect 1171 130 1205 1506
rect 1369 130 1403 1506
rect 1567 130 1601 1506
rect 1765 130 1799 1506
rect 1963 130 1997 1506
rect 2161 130 2195 1506
rect 2359 130 2393 1506
rect 2557 130 2591 1506
rect 2755 130 2789 1506
rect 2953 130 2987 1506
rect 3151 130 3185 1506
rect 3349 130 3383 1506
rect 3547 130 3581 1506
rect 3745 130 3779 1506
rect 3943 130 3977 1506
rect 4141 130 4175 1506
rect -4175 -1506 -4141 -130
rect -3977 -1506 -3943 -130
rect -3779 -1506 -3745 -130
rect -3581 -1506 -3547 -130
rect -3383 -1506 -3349 -130
rect -3185 -1506 -3151 -130
rect -2987 -1506 -2953 -130
rect -2789 -1506 -2755 -130
rect -2591 -1506 -2557 -130
rect -2393 -1506 -2359 -130
rect -2195 -1506 -2161 -130
rect -1997 -1506 -1963 -130
rect -1799 -1506 -1765 -130
rect -1601 -1506 -1567 -130
rect -1403 -1506 -1369 -130
rect -1205 -1506 -1171 -130
rect -1007 -1506 -973 -130
rect -809 -1506 -775 -130
rect -611 -1506 -577 -130
rect -413 -1506 -379 -130
rect -215 -1506 -181 -130
rect -17 -1506 17 -130
rect 181 -1506 215 -130
rect 379 -1506 413 -130
rect 577 -1506 611 -130
rect 775 -1506 809 -130
rect 973 -1506 1007 -130
rect 1171 -1506 1205 -130
rect 1369 -1506 1403 -130
rect 1567 -1506 1601 -130
rect 1765 -1506 1799 -130
rect 1963 -1506 1997 -130
rect 2161 -1506 2195 -130
rect 2359 -1506 2393 -130
rect 2557 -1506 2591 -130
rect 2755 -1506 2789 -130
rect 2953 -1506 2987 -130
rect 3151 -1506 3185 -130
rect 3349 -1506 3383 -130
rect 3547 -1506 3581 -130
rect 3745 -1506 3779 -130
rect 3943 -1506 3977 -130
rect 4141 -1506 4175 -130
<< poly >>
rect -4129 1599 -3989 1615
rect -4129 1565 -4113 1599
rect -4005 1565 -3989 1599
rect -4129 1518 -3989 1565
rect -3931 1599 -3791 1615
rect -3931 1565 -3915 1599
rect -3807 1565 -3791 1599
rect -3931 1518 -3791 1565
rect -3733 1599 -3593 1615
rect -3733 1565 -3717 1599
rect -3609 1565 -3593 1599
rect -3733 1518 -3593 1565
rect -3535 1599 -3395 1615
rect -3535 1565 -3519 1599
rect -3411 1565 -3395 1599
rect -3535 1518 -3395 1565
rect -3337 1599 -3197 1615
rect -3337 1565 -3321 1599
rect -3213 1565 -3197 1599
rect -3337 1518 -3197 1565
rect -3139 1599 -2999 1615
rect -3139 1565 -3123 1599
rect -3015 1565 -2999 1599
rect -3139 1518 -2999 1565
rect -2941 1599 -2801 1615
rect -2941 1565 -2925 1599
rect -2817 1565 -2801 1599
rect -2941 1518 -2801 1565
rect -2743 1599 -2603 1615
rect -2743 1565 -2727 1599
rect -2619 1565 -2603 1599
rect -2743 1518 -2603 1565
rect -2545 1599 -2405 1615
rect -2545 1565 -2529 1599
rect -2421 1565 -2405 1599
rect -2545 1518 -2405 1565
rect -2347 1599 -2207 1615
rect -2347 1565 -2331 1599
rect -2223 1565 -2207 1599
rect -2347 1518 -2207 1565
rect -2149 1599 -2009 1615
rect -2149 1565 -2133 1599
rect -2025 1565 -2009 1599
rect -2149 1518 -2009 1565
rect -1951 1599 -1811 1615
rect -1951 1565 -1935 1599
rect -1827 1565 -1811 1599
rect -1951 1518 -1811 1565
rect -1753 1599 -1613 1615
rect -1753 1565 -1737 1599
rect -1629 1565 -1613 1599
rect -1753 1518 -1613 1565
rect -1555 1599 -1415 1615
rect -1555 1565 -1539 1599
rect -1431 1565 -1415 1599
rect -1555 1518 -1415 1565
rect -1357 1599 -1217 1615
rect -1357 1565 -1341 1599
rect -1233 1565 -1217 1599
rect -1357 1518 -1217 1565
rect -1159 1599 -1019 1615
rect -1159 1565 -1143 1599
rect -1035 1565 -1019 1599
rect -1159 1518 -1019 1565
rect -961 1599 -821 1615
rect -961 1565 -945 1599
rect -837 1565 -821 1599
rect -961 1518 -821 1565
rect -763 1599 -623 1615
rect -763 1565 -747 1599
rect -639 1565 -623 1599
rect -763 1518 -623 1565
rect -565 1599 -425 1615
rect -565 1565 -549 1599
rect -441 1565 -425 1599
rect -565 1518 -425 1565
rect -367 1599 -227 1615
rect -367 1565 -351 1599
rect -243 1565 -227 1599
rect -367 1518 -227 1565
rect -169 1599 -29 1615
rect -169 1565 -153 1599
rect -45 1565 -29 1599
rect -169 1518 -29 1565
rect 29 1599 169 1615
rect 29 1565 45 1599
rect 153 1565 169 1599
rect 29 1518 169 1565
rect 227 1599 367 1615
rect 227 1565 243 1599
rect 351 1565 367 1599
rect 227 1518 367 1565
rect 425 1599 565 1615
rect 425 1565 441 1599
rect 549 1565 565 1599
rect 425 1518 565 1565
rect 623 1599 763 1615
rect 623 1565 639 1599
rect 747 1565 763 1599
rect 623 1518 763 1565
rect 821 1599 961 1615
rect 821 1565 837 1599
rect 945 1565 961 1599
rect 821 1518 961 1565
rect 1019 1599 1159 1615
rect 1019 1565 1035 1599
rect 1143 1565 1159 1599
rect 1019 1518 1159 1565
rect 1217 1599 1357 1615
rect 1217 1565 1233 1599
rect 1341 1565 1357 1599
rect 1217 1518 1357 1565
rect 1415 1599 1555 1615
rect 1415 1565 1431 1599
rect 1539 1565 1555 1599
rect 1415 1518 1555 1565
rect 1613 1599 1753 1615
rect 1613 1565 1629 1599
rect 1737 1565 1753 1599
rect 1613 1518 1753 1565
rect 1811 1599 1951 1615
rect 1811 1565 1827 1599
rect 1935 1565 1951 1599
rect 1811 1518 1951 1565
rect 2009 1599 2149 1615
rect 2009 1565 2025 1599
rect 2133 1565 2149 1599
rect 2009 1518 2149 1565
rect 2207 1599 2347 1615
rect 2207 1565 2223 1599
rect 2331 1565 2347 1599
rect 2207 1518 2347 1565
rect 2405 1599 2545 1615
rect 2405 1565 2421 1599
rect 2529 1565 2545 1599
rect 2405 1518 2545 1565
rect 2603 1599 2743 1615
rect 2603 1565 2619 1599
rect 2727 1565 2743 1599
rect 2603 1518 2743 1565
rect 2801 1599 2941 1615
rect 2801 1565 2817 1599
rect 2925 1565 2941 1599
rect 2801 1518 2941 1565
rect 2999 1599 3139 1615
rect 2999 1565 3015 1599
rect 3123 1565 3139 1599
rect 2999 1518 3139 1565
rect 3197 1599 3337 1615
rect 3197 1565 3213 1599
rect 3321 1565 3337 1599
rect 3197 1518 3337 1565
rect 3395 1599 3535 1615
rect 3395 1565 3411 1599
rect 3519 1565 3535 1599
rect 3395 1518 3535 1565
rect 3593 1599 3733 1615
rect 3593 1565 3609 1599
rect 3717 1565 3733 1599
rect 3593 1518 3733 1565
rect 3791 1599 3931 1615
rect 3791 1565 3807 1599
rect 3915 1565 3931 1599
rect 3791 1518 3931 1565
rect 3989 1599 4129 1615
rect 3989 1565 4005 1599
rect 4113 1565 4129 1599
rect 3989 1518 4129 1565
rect -4129 71 -3989 118
rect -4129 37 -4113 71
rect -4005 37 -3989 71
rect -4129 21 -3989 37
rect -3931 71 -3791 118
rect -3931 37 -3915 71
rect -3807 37 -3791 71
rect -3931 21 -3791 37
rect -3733 71 -3593 118
rect -3733 37 -3717 71
rect -3609 37 -3593 71
rect -3733 21 -3593 37
rect -3535 71 -3395 118
rect -3535 37 -3519 71
rect -3411 37 -3395 71
rect -3535 21 -3395 37
rect -3337 71 -3197 118
rect -3337 37 -3321 71
rect -3213 37 -3197 71
rect -3337 21 -3197 37
rect -3139 71 -2999 118
rect -3139 37 -3123 71
rect -3015 37 -2999 71
rect -3139 21 -2999 37
rect -2941 71 -2801 118
rect -2941 37 -2925 71
rect -2817 37 -2801 71
rect -2941 21 -2801 37
rect -2743 71 -2603 118
rect -2743 37 -2727 71
rect -2619 37 -2603 71
rect -2743 21 -2603 37
rect -2545 71 -2405 118
rect -2545 37 -2529 71
rect -2421 37 -2405 71
rect -2545 21 -2405 37
rect -2347 71 -2207 118
rect -2347 37 -2331 71
rect -2223 37 -2207 71
rect -2347 21 -2207 37
rect -2149 71 -2009 118
rect -2149 37 -2133 71
rect -2025 37 -2009 71
rect -2149 21 -2009 37
rect -1951 71 -1811 118
rect -1951 37 -1935 71
rect -1827 37 -1811 71
rect -1951 21 -1811 37
rect -1753 71 -1613 118
rect -1753 37 -1737 71
rect -1629 37 -1613 71
rect -1753 21 -1613 37
rect -1555 71 -1415 118
rect -1555 37 -1539 71
rect -1431 37 -1415 71
rect -1555 21 -1415 37
rect -1357 71 -1217 118
rect -1357 37 -1341 71
rect -1233 37 -1217 71
rect -1357 21 -1217 37
rect -1159 71 -1019 118
rect -1159 37 -1143 71
rect -1035 37 -1019 71
rect -1159 21 -1019 37
rect -961 71 -821 118
rect -961 37 -945 71
rect -837 37 -821 71
rect -961 21 -821 37
rect -763 71 -623 118
rect -763 37 -747 71
rect -639 37 -623 71
rect -763 21 -623 37
rect -565 71 -425 118
rect -565 37 -549 71
rect -441 37 -425 71
rect -565 21 -425 37
rect -367 71 -227 118
rect -367 37 -351 71
rect -243 37 -227 71
rect -367 21 -227 37
rect -169 71 -29 118
rect -169 37 -153 71
rect -45 37 -29 71
rect -169 21 -29 37
rect 29 71 169 118
rect 29 37 45 71
rect 153 37 169 71
rect 29 21 169 37
rect 227 71 367 118
rect 227 37 243 71
rect 351 37 367 71
rect 227 21 367 37
rect 425 71 565 118
rect 425 37 441 71
rect 549 37 565 71
rect 425 21 565 37
rect 623 71 763 118
rect 623 37 639 71
rect 747 37 763 71
rect 623 21 763 37
rect 821 71 961 118
rect 821 37 837 71
rect 945 37 961 71
rect 821 21 961 37
rect 1019 71 1159 118
rect 1019 37 1035 71
rect 1143 37 1159 71
rect 1019 21 1159 37
rect 1217 71 1357 118
rect 1217 37 1233 71
rect 1341 37 1357 71
rect 1217 21 1357 37
rect 1415 71 1555 118
rect 1415 37 1431 71
rect 1539 37 1555 71
rect 1415 21 1555 37
rect 1613 71 1753 118
rect 1613 37 1629 71
rect 1737 37 1753 71
rect 1613 21 1753 37
rect 1811 71 1951 118
rect 1811 37 1827 71
rect 1935 37 1951 71
rect 1811 21 1951 37
rect 2009 71 2149 118
rect 2009 37 2025 71
rect 2133 37 2149 71
rect 2009 21 2149 37
rect 2207 71 2347 118
rect 2207 37 2223 71
rect 2331 37 2347 71
rect 2207 21 2347 37
rect 2405 71 2545 118
rect 2405 37 2421 71
rect 2529 37 2545 71
rect 2405 21 2545 37
rect 2603 71 2743 118
rect 2603 37 2619 71
rect 2727 37 2743 71
rect 2603 21 2743 37
rect 2801 71 2941 118
rect 2801 37 2817 71
rect 2925 37 2941 71
rect 2801 21 2941 37
rect 2999 71 3139 118
rect 2999 37 3015 71
rect 3123 37 3139 71
rect 2999 21 3139 37
rect 3197 71 3337 118
rect 3197 37 3213 71
rect 3321 37 3337 71
rect 3197 21 3337 37
rect 3395 71 3535 118
rect 3395 37 3411 71
rect 3519 37 3535 71
rect 3395 21 3535 37
rect 3593 71 3733 118
rect 3593 37 3609 71
rect 3717 37 3733 71
rect 3593 21 3733 37
rect 3791 71 3931 118
rect 3791 37 3807 71
rect 3915 37 3931 71
rect 3791 21 3931 37
rect 3989 71 4129 118
rect 3989 37 4005 71
rect 4113 37 4129 71
rect 3989 21 4129 37
rect -4129 -37 -3989 -21
rect -4129 -71 -4113 -37
rect -4005 -71 -3989 -37
rect -4129 -118 -3989 -71
rect -3931 -37 -3791 -21
rect -3931 -71 -3915 -37
rect -3807 -71 -3791 -37
rect -3931 -118 -3791 -71
rect -3733 -37 -3593 -21
rect -3733 -71 -3717 -37
rect -3609 -71 -3593 -37
rect -3733 -118 -3593 -71
rect -3535 -37 -3395 -21
rect -3535 -71 -3519 -37
rect -3411 -71 -3395 -37
rect -3535 -118 -3395 -71
rect -3337 -37 -3197 -21
rect -3337 -71 -3321 -37
rect -3213 -71 -3197 -37
rect -3337 -118 -3197 -71
rect -3139 -37 -2999 -21
rect -3139 -71 -3123 -37
rect -3015 -71 -2999 -37
rect -3139 -118 -2999 -71
rect -2941 -37 -2801 -21
rect -2941 -71 -2925 -37
rect -2817 -71 -2801 -37
rect -2941 -118 -2801 -71
rect -2743 -37 -2603 -21
rect -2743 -71 -2727 -37
rect -2619 -71 -2603 -37
rect -2743 -118 -2603 -71
rect -2545 -37 -2405 -21
rect -2545 -71 -2529 -37
rect -2421 -71 -2405 -37
rect -2545 -118 -2405 -71
rect -2347 -37 -2207 -21
rect -2347 -71 -2331 -37
rect -2223 -71 -2207 -37
rect -2347 -118 -2207 -71
rect -2149 -37 -2009 -21
rect -2149 -71 -2133 -37
rect -2025 -71 -2009 -37
rect -2149 -118 -2009 -71
rect -1951 -37 -1811 -21
rect -1951 -71 -1935 -37
rect -1827 -71 -1811 -37
rect -1951 -118 -1811 -71
rect -1753 -37 -1613 -21
rect -1753 -71 -1737 -37
rect -1629 -71 -1613 -37
rect -1753 -118 -1613 -71
rect -1555 -37 -1415 -21
rect -1555 -71 -1539 -37
rect -1431 -71 -1415 -37
rect -1555 -118 -1415 -71
rect -1357 -37 -1217 -21
rect -1357 -71 -1341 -37
rect -1233 -71 -1217 -37
rect -1357 -118 -1217 -71
rect -1159 -37 -1019 -21
rect -1159 -71 -1143 -37
rect -1035 -71 -1019 -37
rect -1159 -118 -1019 -71
rect -961 -37 -821 -21
rect -961 -71 -945 -37
rect -837 -71 -821 -37
rect -961 -118 -821 -71
rect -763 -37 -623 -21
rect -763 -71 -747 -37
rect -639 -71 -623 -37
rect -763 -118 -623 -71
rect -565 -37 -425 -21
rect -565 -71 -549 -37
rect -441 -71 -425 -37
rect -565 -118 -425 -71
rect -367 -37 -227 -21
rect -367 -71 -351 -37
rect -243 -71 -227 -37
rect -367 -118 -227 -71
rect -169 -37 -29 -21
rect -169 -71 -153 -37
rect -45 -71 -29 -37
rect -169 -118 -29 -71
rect 29 -37 169 -21
rect 29 -71 45 -37
rect 153 -71 169 -37
rect 29 -118 169 -71
rect 227 -37 367 -21
rect 227 -71 243 -37
rect 351 -71 367 -37
rect 227 -118 367 -71
rect 425 -37 565 -21
rect 425 -71 441 -37
rect 549 -71 565 -37
rect 425 -118 565 -71
rect 623 -37 763 -21
rect 623 -71 639 -37
rect 747 -71 763 -37
rect 623 -118 763 -71
rect 821 -37 961 -21
rect 821 -71 837 -37
rect 945 -71 961 -37
rect 821 -118 961 -71
rect 1019 -37 1159 -21
rect 1019 -71 1035 -37
rect 1143 -71 1159 -37
rect 1019 -118 1159 -71
rect 1217 -37 1357 -21
rect 1217 -71 1233 -37
rect 1341 -71 1357 -37
rect 1217 -118 1357 -71
rect 1415 -37 1555 -21
rect 1415 -71 1431 -37
rect 1539 -71 1555 -37
rect 1415 -118 1555 -71
rect 1613 -37 1753 -21
rect 1613 -71 1629 -37
rect 1737 -71 1753 -37
rect 1613 -118 1753 -71
rect 1811 -37 1951 -21
rect 1811 -71 1827 -37
rect 1935 -71 1951 -37
rect 1811 -118 1951 -71
rect 2009 -37 2149 -21
rect 2009 -71 2025 -37
rect 2133 -71 2149 -37
rect 2009 -118 2149 -71
rect 2207 -37 2347 -21
rect 2207 -71 2223 -37
rect 2331 -71 2347 -37
rect 2207 -118 2347 -71
rect 2405 -37 2545 -21
rect 2405 -71 2421 -37
rect 2529 -71 2545 -37
rect 2405 -118 2545 -71
rect 2603 -37 2743 -21
rect 2603 -71 2619 -37
rect 2727 -71 2743 -37
rect 2603 -118 2743 -71
rect 2801 -37 2941 -21
rect 2801 -71 2817 -37
rect 2925 -71 2941 -37
rect 2801 -118 2941 -71
rect 2999 -37 3139 -21
rect 2999 -71 3015 -37
rect 3123 -71 3139 -37
rect 2999 -118 3139 -71
rect 3197 -37 3337 -21
rect 3197 -71 3213 -37
rect 3321 -71 3337 -37
rect 3197 -118 3337 -71
rect 3395 -37 3535 -21
rect 3395 -71 3411 -37
rect 3519 -71 3535 -37
rect 3395 -118 3535 -71
rect 3593 -37 3733 -21
rect 3593 -71 3609 -37
rect 3717 -71 3733 -37
rect 3593 -118 3733 -71
rect 3791 -37 3931 -21
rect 3791 -71 3807 -37
rect 3915 -71 3931 -37
rect 3791 -118 3931 -71
rect 3989 -37 4129 -21
rect 3989 -71 4005 -37
rect 4113 -71 4129 -37
rect 3989 -118 4129 -71
rect -4129 -1565 -3989 -1518
rect -4129 -1599 -4113 -1565
rect -4005 -1599 -3989 -1565
rect -4129 -1615 -3989 -1599
rect -3931 -1565 -3791 -1518
rect -3931 -1599 -3915 -1565
rect -3807 -1599 -3791 -1565
rect -3931 -1615 -3791 -1599
rect -3733 -1565 -3593 -1518
rect -3733 -1599 -3717 -1565
rect -3609 -1599 -3593 -1565
rect -3733 -1615 -3593 -1599
rect -3535 -1565 -3395 -1518
rect -3535 -1599 -3519 -1565
rect -3411 -1599 -3395 -1565
rect -3535 -1615 -3395 -1599
rect -3337 -1565 -3197 -1518
rect -3337 -1599 -3321 -1565
rect -3213 -1599 -3197 -1565
rect -3337 -1615 -3197 -1599
rect -3139 -1565 -2999 -1518
rect -3139 -1599 -3123 -1565
rect -3015 -1599 -2999 -1565
rect -3139 -1615 -2999 -1599
rect -2941 -1565 -2801 -1518
rect -2941 -1599 -2925 -1565
rect -2817 -1599 -2801 -1565
rect -2941 -1615 -2801 -1599
rect -2743 -1565 -2603 -1518
rect -2743 -1599 -2727 -1565
rect -2619 -1599 -2603 -1565
rect -2743 -1615 -2603 -1599
rect -2545 -1565 -2405 -1518
rect -2545 -1599 -2529 -1565
rect -2421 -1599 -2405 -1565
rect -2545 -1615 -2405 -1599
rect -2347 -1565 -2207 -1518
rect -2347 -1599 -2331 -1565
rect -2223 -1599 -2207 -1565
rect -2347 -1615 -2207 -1599
rect -2149 -1565 -2009 -1518
rect -2149 -1599 -2133 -1565
rect -2025 -1599 -2009 -1565
rect -2149 -1615 -2009 -1599
rect -1951 -1565 -1811 -1518
rect -1951 -1599 -1935 -1565
rect -1827 -1599 -1811 -1565
rect -1951 -1615 -1811 -1599
rect -1753 -1565 -1613 -1518
rect -1753 -1599 -1737 -1565
rect -1629 -1599 -1613 -1565
rect -1753 -1615 -1613 -1599
rect -1555 -1565 -1415 -1518
rect -1555 -1599 -1539 -1565
rect -1431 -1599 -1415 -1565
rect -1555 -1615 -1415 -1599
rect -1357 -1565 -1217 -1518
rect -1357 -1599 -1341 -1565
rect -1233 -1599 -1217 -1565
rect -1357 -1615 -1217 -1599
rect -1159 -1565 -1019 -1518
rect -1159 -1599 -1143 -1565
rect -1035 -1599 -1019 -1565
rect -1159 -1615 -1019 -1599
rect -961 -1565 -821 -1518
rect -961 -1599 -945 -1565
rect -837 -1599 -821 -1565
rect -961 -1615 -821 -1599
rect -763 -1565 -623 -1518
rect -763 -1599 -747 -1565
rect -639 -1599 -623 -1565
rect -763 -1615 -623 -1599
rect -565 -1565 -425 -1518
rect -565 -1599 -549 -1565
rect -441 -1599 -425 -1565
rect -565 -1615 -425 -1599
rect -367 -1565 -227 -1518
rect -367 -1599 -351 -1565
rect -243 -1599 -227 -1565
rect -367 -1615 -227 -1599
rect -169 -1565 -29 -1518
rect -169 -1599 -153 -1565
rect -45 -1599 -29 -1565
rect -169 -1615 -29 -1599
rect 29 -1565 169 -1518
rect 29 -1599 45 -1565
rect 153 -1599 169 -1565
rect 29 -1615 169 -1599
rect 227 -1565 367 -1518
rect 227 -1599 243 -1565
rect 351 -1599 367 -1565
rect 227 -1615 367 -1599
rect 425 -1565 565 -1518
rect 425 -1599 441 -1565
rect 549 -1599 565 -1565
rect 425 -1615 565 -1599
rect 623 -1565 763 -1518
rect 623 -1599 639 -1565
rect 747 -1599 763 -1565
rect 623 -1615 763 -1599
rect 821 -1565 961 -1518
rect 821 -1599 837 -1565
rect 945 -1599 961 -1565
rect 821 -1615 961 -1599
rect 1019 -1565 1159 -1518
rect 1019 -1599 1035 -1565
rect 1143 -1599 1159 -1565
rect 1019 -1615 1159 -1599
rect 1217 -1565 1357 -1518
rect 1217 -1599 1233 -1565
rect 1341 -1599 1357 -1565
rect 1217 -1615 1357 -1599
rect 1415 -1565 1555 -1518
rect 1415 -1599 1431 -1565
rect 1539 -1599 1555 -1565
rect 1415 -1615 1555 -1599
rect 1613 -1565 1753 -1518
rect 1613 -1599 1629 -1565
rect 1737 -1599 1753 -1565
rect 1613 -1615 1753 -1599
rect 1811 -1565 1951 -1518
rect 1811 -1599 1827 -1565
rect 1935 -1599 1951 -1565
rect 1811 -1615 1951 -1599
rect 2009 -1565 2149 -1518
rect 2009 -1599 2025 -1565
rect 2133 -1599 2149 -1565
rect 2009 -1615 2149 -1599
rect 2207 -1565 2347 -1518
rect 2207 -1599 2223 -1565
rect 2331 -1599 2347 -1565
rect 2207 -1615 2347 -1599
rect 2405 -1565 2545 -1518
rect 2405 -1599 2421 -1565
rect 2529 -1599 2545 -1565
rect 2405 -1615 2545 -1599
rect 2603 -1565 2743 -1518
rect 2603 -1599 2619 -1565
rect 2727 -1599 2743 -1565
rect 2603 -1615 2743 -1599
rect 2801 -1565 2941 -1518
rect 2801 -1599 2817 -1565
rect 2925 -1599 2941 -1565
rect 2801 -1615 2941 -1599
rect 2999 -1565 3139 -1518
rect 2999 -1599 3015 -1565
rect 3123 -1599 3139 -1565
rect 2999 -1615 3139 -1599
rect 3197 -1565 3337 -1518
rect 3197 -1599 3213 -1565
rect 3321 -1599 3337 -1565
rect 3197 -1615 3337 -1599
rect 3395 -1565 3535 -1518
rect 3395 -1599 3411 -1565
rect 3519 -1599 3535 -1565
rect 3395 -1615 3535 -1599
rect 3593 -1565 3733 -1518
rect 3593 -1599 3609 -1565
rect 3717 -1599 3733 -1565
rect 3593 -1615 3733 -1599
rect 3791 -1565 3931 -1518
rect 3791 -1599 3807 -1565
rect 3915 -1599 3931 -1565
rect 3791 -1615 3931 -1599
rect 3989 -1565 4129 -1518
rect 3989 -1599 4005 -1565
rect 4113 -1599 4129 -1565
rect 3989 -1615 4129 -1599
<< polycont >>
rect -4113 1565 -4005 1599
rect -3915 1565 -3807 1599
rect -3717 1565 -3609 1599
rect -3519 1565 -3411 1599
rect -3321 1565 -3213 1599
rect -3123 1565 -3015 1599
rect -2925 1565 -2817 1599
rect -2727 1565 -2619 1599
rect -2529 1565 -2421 1599
rect -2331 1565 -2223 1599
rect -2133 1565 -2025 1599
rect -1935 1565 -1827 1599
rect -1737 1565 -1629 1599
rect -1539 1565 -1431 1599
rect -1341 1565 -1233 1599
rect -1143 1565 -1035 1599
rect -945 1565 -837 1599
rect -747 1565 -639 1599
rect -549 1565 -441 1599
rect -351 1565 -243 1599
rect -153 1565 -45 1599
rect 45 1565 153 1599
rect 243 1565 351 1599
rect 441 1565 549 1599
rect 639 1565 747 1599
rect 837 1565 945 1599
rect 1035 1565 1143 1599
rect 1233 1565 1341 1599
rect 1431 1565 1539 1599
rect 1629 1565 1737 1599
rect 1827 1565 1935 1599
rect 2025 1565 2133 1599
rect 2223 1565 2331 1599
rect 2421 1565 2529 1599
rect 2619 1565 2727 1599
rect 2817 1565 2925 1599
rect 3015 1565 3123 1599
rect 3213 1565 3321 1599
rect 3411 1565 3519 1599
rect 3609 1565 3717 1599
rect 3807 1565 3915 1599
rect 4005 1565 4113 1599
rect -4113 37 -4005 71
rect -3915 37 -3807 71
rect -3717 37 -3609 71
rect -3519 37 -3411 71
rect -3321 37 -3213 71
rect -3123 37 -3015 71
rect -2925 37 -2817 71
rect -2727 37 -2619 71
rect -2529 37 -2421 71
rect -2331 37 -2223 71
rect -2133 37 -2025 71
rect -1935 37 -1827 71
rect -1737 37 -1629 71
rect -1539 37 -1431 71
rect -1341 37 -1233 71
rect -1143 37 -1035 71
rect -945 37 -837 71
rect -747 37 -639 71
rect -549 37 -441 71
rect -351 37 -243 71
rect -153 37 -45 71
rect 45 37 153 71
rect 243 37 351 71
rect 441 37 549 71
rect 639 37 747 71
rect 837 37 945 71
rect 1035 37 1143 71
rect 1233 37 1341 71
rect 1431 37 1539 71
rect 1629 37 1737 71
rect 1827 37 1935 71
rect 2025 37 2133 71
rect 2223 37 2331 71
rect 2421 37 2529 71
rect 2619 37 2727 71
rect 2817 37 2925 71
rect 3015 37 3123 71
rect 3213 37 3321 71
rect 3411 37 3519 71
rect 3609 37 3717 71
rect 3807 37 3915 71
rect 4005 37 4113 71
rect -4113 -71 -4005 -37
rect -3915 -71 -3807 -37
rect -3717 -71 -3609 -37
rect -3519 -71 -3411 -37
rect -3321 -71 -3213 -37
rect -3123 -71 -3015 -37
rect -2925 -71 -2817 -37
rect -2727 -71 -2619 -37
rect -2529 -71 -2421 -37
rect -2331 -71 -2223 -37
rect -2133 -71 -2025 -37
rect -1935 -71 -1827 -37
rect -1737 -71 -1629 -37
rect -1539 -71 -1431 -37
rect -1341 -71 -1233 -37
rect -1143 -71 -1035 -37
rect -945 -71 -837 -37
rect -747 -71 -639 -37
rect -549 -71 -441 -37
rect -351 -71 -243 -37
rect -153 -71 -45 -37
rect 45 -71 153 -37
rect 243 -71 351 -37
rect 441 -71 549 -37
rect 639 -71 747 -37
rect 837 -71 945 -37
rect 1035 -71 1143 -37
rect 1233 -71 1341 -37
rect 1431 -71 1539 -37
rect 1629 -71 1737 -37
rect 1827 -71 1935 -37
rect 2025 -71 2133 -37
rect 2223 -71 2331 -37
rect 2421 -71 2529 -37
rect 2619 -71 2727 -37
rect 2817 -71 2925 -37
rect 3015 -71 3123 -37
rect 3213 -71 3321 -37
rect 3411 -71 3519 -37
rect 3609 -71 3717 -37
rect 3807 -71 3915 -37
rect 4005 -71 4113 -37
rect -4113 -1599 -4005 -1565
rect -3915 -1599 -3807 -1565
rect -3717 -1599 -3609 -1565
rect -3519 -1599 -3411 -1565
rect -3321 -1599 -3213 -1565
rect -3123 -1599 -3015 -1565
rect -2925 -1599 -2817 -1565
rect -2727 -1599 -2619 -1565
rect -2529 -1599 -2421 -1565
rect -2331 -1599 -2223 -1565
rect -2133 -1599 -2025 -1565
rect -1935 -1599 -1827 -1565
rect -1737 -1599 -1629 -1565
rect -1539 -1599 -1431 -1565
rect -1341 -1599 -1233 -1565
rect -1143 -1599 -1035 -1565
rect -945 -1599 -837 -1565
rect -747 -1599 -639 -1565
rect -549 -1599 -441 -1565
rect -351 -1599 -243 -1565
rect -153 -1599 -45 -1565
rect 45 -1599 153 -1565
rect 243 -1599 351 -1565
rect 441 -1599 549 -1565
rect 639 -1599 747 -1565
rect 837 -1599 945 -1565
rect 1035 -1599 1143 -1565
rect 1233 -1599 1341 -1565
rect 1431 -1599 1539 -1565
rect 1629 -1599 1737 -1565
rect 1827 -1599 1935 -1565
rect 2025 -1599 2133 -1565
rect 2223 -1599 2331 -1565
rect 2421 -1599 2529 -1565
rect 2619 -1599 2727 -1565
rect 2817 -1599 2925 -1565
rect 3015 -1599 3123 -1565
rect 3213 -1599 3321 -1565
rect 3411 -1599 3519 -1565
rect 3609 -1599 3717 -1565
rect 3807 -1599 3915 -1565
rect 4005 -1599 4113 -1565
<< locali >>
rect -4129 1565 -4113 1599
rect -4005 1565 -3989 1599
rect -3931 1565 -3915 1599
rect -3807 1565 -3791 1599
rect -3733 1565 -3717 1599
rect -3609 1565 -3593 1599
rect -3535 1565 -3519 1599
rect -3411 1565 -3395 1599
rect -3337 1565 -3321 1599
rect -3213 1565 -3197 1599
rect -3139 1565 -3123 1599
rect -3015 1565 -2999 1599
rect -2941 1565 -2925 1599
rect -2817 1565 -2801 1599
rect -2743 1565 -2727 1599
rect -2619 1565 -2603 1599
rect -2545 1565 -2529 1599
rect -2421 1565 -2405 1599
rect -2347 1565 -2331 1599
rect -2223 1565 -2207 1599
rect -2149 1565 -2133 1599
rect -2025 1565 -2009 1599
rect -1951 1565 -1935 1599
rect -1827 1565 -1811 1599
rect -1753 1565 -1737 1599
rect -1629 1565 -1613 1599
rect -1555 1565 -1539 1599
rect -1431 1565 -1415 1599
rect -1357 1565 -1341 1599
rect -1233 1565 -1217 1599
rect -1159 1565 -1143 1599
rect -1035 1565 -1019 1599
rect -961 1565 -945 1599
rect -837 1565 -821 1599
rect -763 1565 -747 1599
rect -639 1565 -623 1599
rect -565 1565 -549 1599
rect -441 1565 -425 1599
rect -367 1565 -351 1599
rect -243 1565 -227 1599
rect -169 1565 -153 1599
rect -45 1565 -29 1599
rect 29 1565 45 1599
rect 153 1565 169 1599
rect 227 1565 243 1599
rect 351 1565 367 1599
rect 425 1565 441 1599
rect 549 1565 565 1599
rect 623 1565 639 1599
rect 747 1565 763 1599
rect 821 1565 837 1599
rect 945 1565 961 1599
rect 1019 1565 1035 1599
rect 1143 1565 1159 1599
rect 1217 1565 1233 1599
rect 1341 1565 1357 1599
rect 1415 1565 1431 1599
rect 1539 1565 1555 1599
rect 1613 1565 1629 1599
rect 1737 1565 1753 1599
rect 1811 1565 1827 1599
rect 1935 1565 1951 1599
rect 2009 1565 2025 1599
rect 2133 1565 2149 1599
rect 2207 1565 2223 1599
rect 2331 1565 2347 1599
rect 2405 1565 2421 1599
rect 2529 1565 2545 1599
rect 2603 1565 2619 1599
rect 2727 1565 2743 1599
rect 2801 1565 2817 1599
rect 2925 1565 2941 1599
rect 2999 1565 3015 1599
rect 3123 1565 3139 1599
rect 3197 1565 3213 1599
rect 3321 1565 3337 1599
rect 3395 1565 3411 1599
rect 3519 1565 3535 1599
rect 3593 1565 3609 1599
rect 3717 1565 3733 1599
rect 3791 1565 3807 1599
rect 3915 1565 3931 1599
rect 3989 1565 4005 1599
rect 4113 1565 4129 1599
rect -4175 1506 -4141 1522
rect -4175 114 -4141 130
rect -3977 1506 -3943 1522
rect -3977 114 -3943 130
rect -3779 1506 -3745 1522
rect -3779 114 -3745 130
rect -3581 1506 -3547 1522
rect -3581 114 -3547 130
rect -3383 1506 -3349 1522
rect -3383 114 -3349 130
rect -3185 1506 -3151 1522
rect -3185 114 -3151 130
rect -2987 1506 -2953 1522
rect -2987 114 -2953 130
rect -2789 1506 -2755 1522
rect -2789 114 -2755 130
rect -2591 1506 -2557 1522
rect -2591 114 -2557 130
rect -2393 1506 -2359 1522
rect -2393 114 -2359 130
rect -2195 1506 -2161 1522
rect -2195 114 -2161 130
rect -1997 1506 -1963 1522
rect -1997 114 -1963 130
rect -1799 1506 -1765 1522
rect -1799 114 -1765 130
rect -1601 1506 -1567 1522
rect -1601 114 -1567 130
rect -1403 1506 -1369 1522
rect -1403 114 -1369 130
rect -1205 1506 -1171 1522
rect -1205 114 -1171 130
rect -1007 1506 -973 1522
rect -1007 114 -973 130
rect -809 1506 -775 1522
rect -809 114 -775 130
rect -611 1506 -577 1522
rect -611 114 -577 130
rect -413 1506 -379 1522
rect -413 114 -379 130
rect -215 1506 -181 1522
rect -215 114 -181 130
rect -17 1506 17 1522
rect -17 114 17 130
rect 181 1506 215 1522
rect 181 114 215 130
rect 379 1506 413 1522
rect 379 114 413 130
rect 577 1506 611 1522
rect 577 114 611 130
rect 775 1506 809 1522
rect 775 114 809 130
rect 973 1506 1007 1522
rect 973 114 1007 130
rect 1171 1506 1205 1522
rect 1171 114 1205 130
rect 1369 1506 1403 1522
rect 1369 114 1403 130
rect 1567 1506 1601 1522
rect 1567 114 1601 130
rect 1765 1506 1799 1522
rect 1765 114 1799 130
rect 1963 1506 1997 1522
rect 1963 114 1997 130
rect 2161 1506 2195 1522
rect 2161 114 2195 130
rect 2359 1506 2393 1522
rect 2359 114 2393 130
rect 2557 1506 2591 1522
rect 2557 114 2591 130
rect 2755 1506 2789 1522
rect 2755 114 2789 130
rect 2953 1506 2987 1522
rect 2953 114 2987 130
rect 3151 1506 3185 1522
rect 3151 114 3185 130
rect 3349 1506 3383 1522
rect 3349 114 3383 130
rect 3547 1506 3581 1522
rect 3547 114 3581 130
rect 3745 1506 3779 1522
rect 3745 114 3779 130
rect 3943 1506 3977 1522
rect 3943 114 3977 130
rect 4141 1506 4175 1522
rect 4141 114 4175 130
rect -4129 37 -4113 71
rect -4005 37 -3989 71
rect -3931 37 -3915 71
rect -3807 37 -3791 71
rect -3733 37 -3717 71
rect -3609 37 -3593 71
rect -3535 37 -3519 71
rect -3411 37 -3395 71
rect -3337 37 -3321 71
rect -3213 37 -3197 71
rect -3139 37 -3123 71
rect -3015 37 -2999 71
rect -2941 37 -2925 71
rect -2817 37 -2801 71
rect -2743 37 -2727 71
rect -2619 37 -2603 71
rect -2545 37 -2529 71
rect -2421 37 -2405 71
rect -2347 37 -2331 71
rect -2223 37 -2207 71
rect -2149 37 -2133 71
rect -2025 37 -2009 71
rect -1951 37 -1935 71
rect -1827 37 -1811 71
rect -1753 37 -1737 71
rect -1629 37 -1613 71
rect -1555 37 -1539 71
rect -1431 37 -1415 71
rect -1357 37 -1341 71
rect -1233 37 -1217 71
rect -1159 37 -1143 71
rect -1035 37 -1019 71
rect -961 37 -945 71
rect -837 37 -821 71
rect -763 37 -747 71
rect -639 37 -623 71
rect -565 37 -549 71
rect -441 37 -425 71
rect -367 37 -351 71
rect -243 37 -227 71
rect -169 37 -153 71
rect -45 37 -29 71
rect 29 37 45 71
rect 153 37 169 71
rect 227 37 243 71
rect 351 37 367 71
rect 425 37 441 71
rect 549 37 565 71
rect 623 37 639 71
rect 747 37 763 71
rect 821 37 837 71
rect 945 37 961 71
rect 1019 37 1035 71
rect 1143 37 1159 71
rect 1217 37 1233 71
rect 1341 37 1357 71
rect 1415 37 1431 71
rect 1539 37 1555 71
rect 1613 37 1629 71
rect 1737 37 1753 71
rect 1811 37 1827 71
rect 1935 37 1951 71
rect 2009 37 2025 71
rect 2133 37 2149 71
rect 2207 37 2223 71
rect 2331 37 2347 71
rect 2405 37 2421 71
rect 2529 37 2545 71
rect 2603 37 2619 71
rect 2727 37 2743 71
rect 2801 37 2817 71
rect 2925 37 2941 71
rect 2999 37 3015 71
rect 3123 37 3139 71
rect 3197 37 3213 71
rect 3321 37 3337 71
rect 3395 37 3411 71
rect 3519 37 3535 71
rect 3593 37 3609 71
rect 3717 37 3733 71
rect 3791 37 3807 71
rect 3915 37 3931 71
rect 3989 37 4005 71
rect 4113 37 4129 71
rect -4129 -71 -4113 -37
rect -4005 -71 -3989 -37
rect -3931 -71 -3915 -37
rect -3807 -71 -3791 -37
rect -3733 -71 -3717 -37
rect -3609 -71 -3593 -37
rect -3535 -71 -3519 -37
rect -3411 -71 -3395 -37
rect -3337 -71 -3321 -37
rect -3213 -71 -3197 -37
rect -3139 -71 -3123 -37
rect -3015 -71 -2999 -37
rect -2941 -71 -2925 -37
rect -2817 -71 -2801 -37
rect -2743 -71 -2727 -37
rect -2619 -71 -2603 -37
rect -2545 -71 -2529 -37
rect -2421 -71 -2405 -37
rect -2347 -71 -2331 -37
rect -2223 -71 -2207 -37
rect -2149 -71 -2133 -37
rect -2025 -71 -2009 -37
rect -1951 -71 -1935 -37
rect -1827 -71 -1811 -37
rect -1753 -71 -1737 -37
rect -1629 -71 -1613 -37
rect -1555 -71 -1539 -37
rect -1431 -71 -1415 -37
rect -1357 -71 -1341 -37
rect -1233 -71 -1217 -37
rect -1159 -71 -1143 -37
rect -1035 -71 -1019 -37
rect -961 -71 -945 -37
rect -837 -71 -821 -37
rect -763 -71 -747 -37
rect -639 -71 -623 -37
rect -565 -71 -549 -37
rect -441 -71 -425 -37
rect -367 -71 -351 -37
rect -243 -71 -227 -37
rect -169 -71 -153 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 153 -71 169 -37
rect 227 -71 243 -37
rect 351 -71 367 -37
rect 425 -71 441 -37
rect 549 -71 565 -37
rect 623 -71 639 -37
rect 747 -71 763 -37
rect 821 -71 837 -37
rect 945 -71 961 -37
rect 1019 -71 1035 -37
rect 1143 -71 1159 -37
rect 1217 -71 1233 -37
rect 1341 -71 1357 -37
rect 1415 -71 1431 -37
rect 1539 -71 1555 -37
rect 1613 -71 1629 -37
rect 1737 -71 1753 -37
rect 1811 -71 1827 -37
rect 1935 -71 1951 -37
rect 2009 -71 2025 -37
rect 2133 -71 2149 -37
rect 2207 -71 2223 -37
rect 2331 -71 2347 -37
rect 2405 -71 2421 -37
rect 2529 -71 2545 -37
rect 2603 -71 2619 -37
rect 2727 -71 2743 -37
rect 2801 -71 2817 -37
rect 2925 -71 2941 -37
rect 2999 -71 3015 -37
rect 3123 -71 3139 -37
rect 3197 -71 3213 -37
rect 3321 -71 3337 -37
rect 3395 -71 3411 -37
rect 3519 -71 3535 -37
rect 3593 -71 3609 -37
rect 3717 -71 3733 -37
rect 3791 -71 3807 -37
rect 3915 -71 3931 -37
rect 3989 -71 4005 -37
rect 4113 -71 4129 -37
rect -4175 -130 -4141 -114
rect -4175 -1522 -4141 -1506
rect -3977 -130 -3943 -114
rect -3977 -1522 -3943 -1506
rect -3779 -130 -3745 -114
rect -3779 -1522 -3745 -1506
rect -3581 -130 -3547 -114
rect -3581 -1522 -3547 -1506
rect -3383 -130 -3349 -114
rect -3383 -1522 -3349 -1506
rect -3185 -130 -3151 -114
rect -3185 -1522 -3151 -1506
rect -2987 -130 -2953 -114
rect -2987 -1522 -2953 -1506
rect -2789 -130 -2755 -114
rect -2789 -1522 -2755 -1506
rect -2591 -130 -2557 -114
rect -2591 -1522 -2557 -1506
rect -2393 -130 -2359 -114
rect -2393 -1522 -2359 -1506
rect -2195 -130 -2161 -114
rect -2195 -1522 -2161 -1506
rect -1997 -130 -1963 -114
rect -1997 -1522 -1963 -1506
rect -1799 -130 -1765 -114
rect -1799 -1522 -1765 -1506
rect -1601 -130 -1567 -114
rect -1601 -1522 -1567 -1506
rect -1403 -130 -1369 -114
rect -1403 -1522 -1369 -1506
rect -1205 -130 -1171 -114
rect -1205 -1522 -1171 -1506
rect -1007 -130 -973 -114
rect -1007 -1522 -973 -1506
rect -809 -130 -775 -114
rect -809 -1522 -775 -1506
rect -611 -130 -577 -114
rect -611 -1522 -577 -1506
rect -413 -130 -379 -114
rect -413 -1522 -379 -1506
rect -215 -130 -181 -114
rect -215 -1522 -181 -1506
rect -17 -130 17 -114
rect -17 -1522 17 -1506
rect 181 -130 215 -114
rect 181 -1522 215 -1506
rect 379 -130 413 -114
rect 379 -1522 413 -1506
rect 577 -130 611 -114
rect 577 -1522 611 -1506
rect 775 -130 809 -114
rect 775 -1522 809 -1506
rect 973 -130 1007 -114
rect 973 -1522 1007 -1506
rect 1171 -130 1205 -114
rect 1171 -1522 1205 -1506
rect 1369 -130 1403 -114
rect 1369 -1522 1403 -1506
rect 1567 -130 1601 -114
rect 1567 -1522 1601 -1506
rect 1765 -130 1799 -114
rect 1765 -1522 1799 -1506
rect 1963 -130 1997 -114
rect 1963 -1522 1997 -1506
rect 2161 -130 2195 -114
rect 2161 -1522 2195 -1506
rect 2359 -130 2393 -114
rect 2359 -1522 2393 -1506
rect 2557 -130 2591 -114
rect 2557 -1522 2591 -1506
rect 2755 -130 2789 -114
rect 2755 -1522 2789 -1506
rect 2953 -130 2987 -114
rect 2953 -1522 2987 -1506
rect 3151 -130 3185 -114
rect 3151 -1522 3185 -1506
rect 3349 -130 3383 -114
rect 3349 -1522 3383 -1506
rect 3547 -130 3581 -114
rect 3547 -1522 3581 -1506
rect 3745 -130 3779 -114
rect 3745 -1522 3779 -1506
rect 3943 -130 3977 -114
rect 3943 -1522 3977 -1506
rect 4141 -130 4175 -114
rect 4141 -1522 4175 -1506
rect -4129 -1599 -4113 -1565
rect -4005 -1599 -3989 -1565
rect -3931 -1599 -3915 -1565
rect -3807 -1599 -3791 -1565
rect -3733 -1599 -3717 -1565
rect -3609 -1599 -3593 -1565
rect -3535 -1599 -3519 -1565
rect -3411 -1599 -3395 -1565
rect -3337 -1599 -3321 -1565
rect -3213 -1599 -3197 -1565
rect -3139 -1599 -3123 -1565
rect -3015 -1599 -2999 -1565
rect -2941 -1599 -2925 -1565
rect -2817 -1599 -2801 -1565
rect -2743 -1599 -2727 -1565
rect -2619 -1599 -2603 -1565
rect -2545 -1599 -2529 -1565
rect -2421 -1599 -2405 -1565
rect -2347 -1599 -2331 -1565
rect -2223 -1599 -2207 -1565
rect -2149 -1599 -2133 -1565
rect -2025 -1599 -2009 -1565
rect -1951 -1599 -1935 -1565
rect -1827 -1599 -1811 -1565
rect -1753 -1599 -1737 -1565
rect -1629 -1599 -1613 -1565
rect -1555 -1599 -1539 -1565
rect -1431 -1599 -1415 -1565
rect -1357 -1599 -1341 -1565
rect -1233 -1599 -1217 -1565
rect -1159 -1599 -1143 -1565
rect -1035 -1599 -1019 -1565
rect -961 -1599 -945 -1565
rect -837 -1599 -821 -1565
rect -763 -1599 -747 -1565
rect -639 -1599 -623 -1565
rect -565 -1599 -549 -1565
rect -441 -1599 -425 -1565
rect -367 -1599 -351 -1565
rect -243 -1599 -227 -1565
rect -169 -1599 -153 -1565
rect -45 -1599 -29 -1565
rect 29 -1599 45 -1565
rect 153 -1599 169 -1565
rect 227 -1599 243 -1565
rect 351 -1599 367 -1565
rect 425 -1599 441 -1565
rect 549 -1599 565 -1565
rect 623 -1599 639 -1565
rect 747 -1599 763 -1565
rect 821 -1599 837 -1565
rect 945 -1599 961 -1565
rect 1019 -1599 1035 -1565
rect 1143 -1599 1159 -1565
rect 1217 -1599 1233 -1565
rect 1341 -1599 1357 -1565
rect 1415 -1599 1431 -1565
rect 1539 -1599 1555 -1565
rect 1613 -1599 1629 -1565
rect 1737 -1599 1753 -1565
rect 1811 -1599 1827 -1565
rect 1935 -1599 1951 -1565
rect 2009 -1599 2025 -1565
rect 2133 -1599 2149 -1565
rect 2207 -1599 2223 -1565
rect 2331 -1599 2347 -1565
rect 2405 -1599 2421 -1565
rect 2529 -1599 2545 -1565
rect 2603 -1599 2619 -1565
rect 2727 -1599 2743 -1565
rect 2801 -1599 2817 -1565
rect 2925 -1599 2941 -1565
rect 2999 -1599 3015 -1565
rect 3123 -1599 3139 -1565
rect 3197 -1599 3213 -1565
rect 3321 -1599 3337 -1565
rect 3395 -1599 3411 -1565
rect 3519 -1599 3535 -1565
rect 3593 -1599 3609 -1565
rect 3717 -1599 3733 -1565
rect 3791 -1599 3807 -1565
rect 3915 -1599 3931 -1565
rect 3989 -1599 4005 -1565
rect 4113 -1599 4129 -1565
<< viali >>
rect -4113 1565 -4005 1599
rect -3915 1565 -3807 1599
rect -3717 1565 -3609 1599
rect -3519 1565 -3411 1599
rect -3321 1565 -3213 1599
rect -3123 1565 -3015 1599
rect -2925 1565 -2817 1599
rect -2727 1565 -2619 1599
rect -2529 1565 -2421 1599
rect -2331 1565 -2223 1599
rect -2133 1565 -2025 1599
rect -1935 1565 -1827 1599
rect -1737 1565 -1629 1599
rect -1539 1565 -1431 1599
rect -1341 1565 -1233 1599
rect -1143 1565 -1035 1599
rect -945 1565 -837 1599
rect -747 1565 -639 1599
rect -549 1565 -441 1599
rect -351 1565 -243 1599
rect -153 1565 -45 1599
rect 45 1565 153 1599
rect 243 1565 351 1599
rect 441 1565 549 1599
rect 639 1565 747 1599
rect 837 1565 945 1599
rect 1035 1565 1143 1599
rect 1233 1565 1341 1599
rect 1431 1565 1539 1599
rect 1629 1565 1737 1599
rect 1827 1565 1935 1599
rect 2025 1565 2133 1599
rect 2223 1565 2331 1599
rect 2421 1565 2529 1599
rect 2619 1565 2727 1599
rect 2817 1565 2925 1599
rect 3015 1565 3123 1599
rect 3213 1565 3321 1599
rect 3411 1565 3519 1599
rect 3609 1565 3717 1599
rect 3807 1565 3915 1599
rect 4005 1565 4113 1599
rect -4175 130 -4141 1506
rect -3977 130 -3943 1506
rect -3779 130 -3745 1506
rect -3581 130 -3547 1506
rect -3383 130 -3349 1506
rect -3185 130 -3151 1506
rect -2987 130 -2953 1506
rect -2789 130 -2755 1506
rect -2591 130 -2557 1506
rect -2393 130 -2359 1506
rect -2195 130 -2161 1506
rect -1997 130 -1963 1506
rect -1799 130 -1765 1506
rect -1601 130 -1567 1506
rect -1403 130 -1369 1506
rect -1205 130 -1171 1506
rect -1007 130 -973 1506
rect -809 130 -775 1506
rect -611 130 -577 1506
rect -413 130 -379 1506
rect -215 130 -181 1506
rect -17 130 17 1506
rect 181 130 215 1506
rect 379 130 413 1506
rect 577 130 611 1506
rect 775 130 809 1506
rect 973 130 1007 1506
rect 1171 130 1205 1506
rect 1369 130 1403 1506
rect 1567 130 1601 1506
rect 1765 130 1799 1506
rect 1963 130 1997 1506
rect 2161 130 2195 1506
rect 2359 130 2393 1506
rect 2557 130 2591 1506
rect 2755 130 2789 1506
rect 2953 130 2987 1506
rect 3151 130 3185 1506
rect 3349 130 3383 1506
rect 3547 130 3581 1506
rect 3745 130 3779 1506
rect 3943 130 3977 1506
rect 4141 130 4175 1506
rect -4113 37 -4005 71
rect -3915 37 -3807 71
rect -3717 37 -3609 71
rect -3519 37 -3411 71
rect -3321 37 -3213 71
rect -3123 37 -3015 71
rect -2925 37 -2817 71
rect -2727 37 -2619 71
rect -2529 37 -2421 71
rect -2331 37 -2223 71
rect -2133 37 -2025 71
rect -1935 37 -1827 71
rect -1737 37 -1629 71
rect -1539 37 -1431 71
rect -1341 37 -1233 71
rect -1143 37 -1035 71
rect -945 37 -837 71
rect -747 37 -639 71
rect -549 37 -441 71
rect -351 37 -243 71
rect -153 37 -45 71
rect 45 37 153 71
rect 243 37 351 71
rect 441 37 549 71
rect 639 37 747 71
rect 837 37 945 71
rect 1035 37 1143 71
rect 1233 37 1341 71
rect 1431 37 1539 71
rect 1629 37 1737 71
rect 1827 37 1935 71
rect 2025 37 2133 71
rect 2223 37 2331 71
rect 2421 37 2529 71
rect 2619 37 2727 71
rect 2817 37 2925 71
rect 3015 37 3123 71
rect 3213 37 3321 71
rect 3411 37 3519 71
rect 3609 37 3717 71
rect 3807 37 3915 71
rect 4005 37 4113 71
rect -4113 -71 -4005 -37
rect -3915 -71 -3807 -37
rect -3717 -71 -3609 -37
rect -3519 -71 -3411 -37
rect -3321 -71 -3213 -37
rect -3123 -71 -3015 -37
rect -2925 -71 -2817 -37
rect -2727 -71 -2619 -37
rect -2529 -71 -2421 -37
rect -2331 -71 -2223 -37
rect -2133 -71 -2025 -37
rect -1935 -71 -1827 -37
rect -1737 -71 -1629 -37
rect -1539 -71 -1431 -37
rect -1341 -71 -1233 -37
rect -1143 -71 -1035 -37
rect -945 -71 -837 -37
rect -747 -71 -639 -37
rect -549 -71 -441 -37
rect -351 -71 -243 -37
rect -153 -71 -45 -37
rect 45 -71 153 -37
rect 243 -71 351 -37
rect 441 -71 549 -37
rect 639 -71 747 -37
rect 837 -71 945 -37
rect 1035 -71 1143 -37
rect 1233 -71 1341 -37
rect 1431 -71 1539 -37
rect 1629 -71 1737 -37
rect 1827 -71 1935 -37
rect 2025 -71 2133 -37
rect 2223 -71 2331 -37
rect 2421 -71 2529 -37
rect 2619 -71 2727 -37
rect 2817 -71 2925 -37
rect 3015 -71 3123 -37
rect 3213 -71 3321 -37
rect 3411 -71 3519 -37
rect 3609 -71 3717 -37
rect 3807 -71 3915 -37
rect 4005 -71 4113 -37
rect -4175 -1506 -4141 -130
rect -3977 -1506 -3943 -130
rect -3779 -1506 -3745 -130
rect -3581 -1506 -3547 -130
rect -3383 -1506 -3349 -130
rect -3185 -1506 -3151 -130
rect -2987 -1506 -2953 -130
rect -2789 -1506 -2755 -130
rect -2591 -1506 -2557 -130
rect -2393 -1506 -2359 -130
rect -2195 -1506 -2161 -130
rect -1997 -1506 -1963 -130
rect -1799 -1506 -1765 -130
rect -1601 -1506 -1567 -130
rect -1403 -1506 -1369 -130
rect -1205 -1506 -1171 -130
rect -1007 -1506 -973 -130
rect -809 -1506 -775 -130
rect -611 -1506 -577 -130
rect -413 -1506 -379 -130
rect -215 -1506 -181 -130
rect -17 -1506 17 -130
rect 181 -1506 215 -130
rect 379 -1506 413 -130
rect 577 -1506 611 -130
rect 775 -1506 809 -130
rect 973 -1506 1007 -130
rect 1171 -1506 1205 -130
rect 1369 -1506 1403 -130
rect 1567 -1506 1601 -130
rect 1765 -1506 1799 -130
rect 1963 -1506 1997 -130
rect 2161 -1506 2195 -130
rect 2359 -1506 2393 -130
rect 2557 -1506 2591 -130
rect 2755 -1506 2789 -130
rect 2953 -1506 2987 -130
rect 3151 -1506 3185 -130
rect 3349 -1506 3383 -130
rect 3547 -1506 3581 -130
rect 3745 -1506 3779 -130
rect 3943 -1506 3977 -130
rect 4141 -1506 4175 -130
rect -4113 -1599 -4005 -1565
rect -3915 -1599 -3807 -1565
rect -3717 -1599 -3609 -1565
rect -3519 -1599 -3411 -1565
rect -3321 -1599 -3213 -1565
rect -3123 -1599 -3015 -1565
rect -2925 -1599 -2817 -1565
rect -2727 -1599 -2619 -1565
rect -2529 -1599 -2421 -1565
rect -2331 -1599 -2223 -1565
rect -2133 -1599 -2025 -1565
rect -1935 -1599 -1827 -1565
rect -1737 -1599 -1629 -1565
rect -1539 -1599 -1431 -1565
rect -1341 -1599 -1233 -1565
rect -1143 -1599 -1035 -1565
rect -945 -1599 -837 -1565
rect -747 -1599 -639 -1565
rect -549 -1599 -441 -1565
rect -351 -1599 -243 -1565
rect -153 -1599 -45 -1565
rect 45 -1599 153 -1565
rect 243 -1599 351 -1565
rect 441 -1599 549 -1565
rect 639 -1599 747 -1565
rect 837 -1599 945 -1565
rect 1035 -1599 1143 -1565
rect 1233 -1599 1341 -1565
rect 1431 -1599 1539 -1565
rect 1629 -1599 1737 -1565
rect 1827 -1599 1935 -1565
rect 2025 -1599 2133 -1565
rect 2223 -1599 2331 -1565
rect 2421 -1599 2529 -1565
rect 2619 -1599 2727 -1565
rect 2817 -1599 2925 -1565
rect 3015 -1599 3123 -1565
rect 3213 -1599 3321 -1565
rect 3411 -1599 3519 -1565
rect 3609 -1599 3717 -1565
rect 3807 -1599 3915 -1565
rect 4005 -1599 4113 -1565
<< metal1 >>
rect -4125 1599 -3993 1605
rect -4125 1565 -4113 1599
rect -4005 1565 -3993 1599
rect -4125 1559 -3993 1565
rect -3927 1599 -3795 1605
rect -3927 1565 -3915 1599
rect -3807 1565 -3795 1599
rect -3927 1559 -3795 1565
rect -3729 1599 -3597 1605
rect -3729 1565 -3717 1599
rect -3609 1565 -3597 1599
rect -3729 1559 -3597 1565
rect -3531 1599 -3399 1605
rect -3531 1565 -3519 1599
rect -3411 1565 -3399 1599
rect -3531 1559 -3399 1565
rect -3333 1599 -3201 1605
rect -3333 1565 -3321 1599
rect -3213 1565 -3201 1599
rect -3333 1559 -3201 1565
rect -3135 1599 -3003 1605
rect -3135 1565 -3123 1599
rect -3015 1565 -3003 1599
rect -3135 1559 -3003 1565
rect -2937 1599 -2805 1605
rect -2937 1565 -2925 1599
rect -2817 1565 -2805 1599
rect -2937 1559 -2805 1565
rect -2739 1599 -2607 1605
rect -2739 1565 -2727 1599
rect -2619 1565 -2607 1599
rect -2739 1559 -2607 1565
rect -2541 1599 -2409 1605
rect -2541 1565 -2529 1599
rect -2421 1565 -2409 1599
rect -2541 1559 -2409 1565
rect -2343 1599 -2211 1605
rect -2343 1565 -2331 1599
rect -2223 1565 -2211 1599
rect -2343 1559 -2211 1565
rect -2145 1599 -2013 1605
rect -2145 1565 -2133 1599
rect -2025 1565 -2013 1599
rect -2145 1559 -2013 1565
rect -1947 1599 -1815 1605
rect -1947 1565 -1935 1599
rect -1827 1565 -1815 1599
rect -1947 1559 -1815 1565
rect -1749 1599 -1617 1605
rect -1749 1565 -1737 1599
rect -1629 1565 -1617 1599
rect -1749 1559 -1617 1565
rect -1551 1599 -1419 1605
rect -1551 1565 -1539 1599
rect -1431 1565 -1419 1599
rect -1551 1559 -1419 1565
rect -1353 1599 -1221 1605
rect -1353 1565 -1341 1599
rect -1233 1565 -1221 1599
rect -1353 1559 -1221 1565
rect -1155 1599 -1023 1605
rect -1155 1565 -1143 1599
rect -1035 1565 -1023 1599
rect -1155 1559 -1023 1565
rect -957 1599 -825 1605
rect -957 1565 -945 1599
rect -837 1565 -825 1599
rect -957 1559 -825 1565
rect -759 1599 -627 1605
rect -759 1565 -747 1599
rect -639 1565 -627 1599
rect -759 1559 -627 1565
rect -561 1599 -429 1605
rect -561 1565 -549 1599
rect -441 1565 -429 1599
rect -561 1559 -429 1565
rect -363 1599 -231 1605
rect -363 1565 -351 1599
rect -243 1565 -231 1599
rect -363 1559 -231 1565
rect -165 1599 -33 1605
rect -165 1565 -153 1599
rect -45 1565 -33 1599
rect -165 1559 -33 1565
rect 33 1599 165 1605
rect 33 1565 45 1599
rect 153 1565 165 1599
rect 33 1559 165 1565
rect 231 1599 363 1605
rect 231 1565 243 1599
rect 351 1565 363 1599
rect 231 1559 363 1565
rect 429 1599 561 1605
rect 429 1565 441 1599
rect 549 1565 561 1599
rect 429 1559 561 1565
rect 627 1599 759 1605
rect 627 1565 639 1599
rect 747 1565 759 1599
rect 627 1559 759 1565
rect 825 1599 957 1605
rect 825 1565 837 1599
rect 945 1565 957 1599
rect 825 1559 957 1565
rect 1023 1599 1155 1605
rect 1023 1565 1035 1599
rect 1143 1565 1155 1599
rect 1023 1559 1155 1565
rect 1221 1599 1353 1605
rect 1221 1565 1233 1599
rect 1341 1565 1353 1599
rect 1221 1559 1353 1565
rect 1419 1599 1551 1605
rect 1419 1565 1431 1599
rect 1539 1565 1551 1599
rect 1419 1559 1551 1565
rect 1617 1599 1749 1605
rect 1617 1565 1629 1599
rect 1737 1565 1749 1599
rect 1617 1559 1749 1565
rect 1815 1599 1947 1605
rect 1815 1565 1827 1599
rect 1935 1565 1947 1599
rect 1815 1559 1947 1565
rect 2013 1599 2145 1605
rect 2013 1565 2025 1599
rect 2133 1565 2145 1599
rect 2013 1559 2145 1565
rect 2211 1599 2343 1605
rect 2211 1565 2223 1599
rect 2331 1565 2343 1599
rect 2211 1559 2343 1565
rect 2409 1599 2541 1605
rect 2409 1565 2421 1599
rect 2529 1565 2541 1599
rect 2409 1559 2541 1565
rect 2607 1599 2739 1605
rect 2607 1565 2619 1599
rect 2727 1565 2739 1599
rect 2607 1559 2739 1565
rect 2805 1599 2937 1605
rect 2805 1565 2817 1599
rect 2925 1565 2937 1599
rect 2805 1559 2937 1565
rect 3003 1599 3135 1605
rect 3003 1565 3015 1599
rect 3123 1565 3135 1599
rect 3003 1559 3135 1565
rect 3201 1599 3333 1605
rect 3201 1565 3213 1599
rect 3321 1565 3333 1599
rect 3201 1559 3333 1565
rect 3399 1599 3531 1605
rect 3399 1565 3411 1599
rect 3519 1565 3531 1599
rect 3399 1559 3531 1565
rect 3597 1599 3729 1605
rect 3597 1565 3609 1599
rect 3717 1565 3729 1599
rect 3597 1559 3729 1565
rect 3795 1599 3927 1605
rect 3795 1565 3807 1599
rect 3915 1565 3927 1599
rect 3795 1559 3927 1565
rect 3993 1599 4125 1605
rect 3993 1565 4005 1599
rect 4113 1565 4125 1599
rect 3993 1559 4125 1565
rect -4181 1506 -4135 1518
rect -4181 130 -4175 1506
rect -4141 130 -4135 1506
rect -4181 118 -4135 130
rect -3983 1506 -3937 1518
rect -3983 130 -3977 1506
rect -3943 130 -3937 1506
rect -3983 118 -3937 130
rect -3785 1506 -3739 1518
rect -3785 130 -3779 1506
rect -3745 130 -3739 1506
rect -3785 118 -3739 130
rect -3587 1506 -3541 1518
rect -3587 130 -3581 1506
rect -3547 130 -3541 1506
rect -3587 118 -3541 130
rect -3389 1506 -3343 1518
rect -3389 130 -3383 1506
rect -3349 130 -3343 1506
rect -3389 118 -3343 130
rect -3191 1506 -3145 1518
rect -3191 130 -3185 1506
rect -3151 130 -3145 1506
rect -3191 118 -3145 130
rect -2993 1506 -2947 1518
rect -2993 130 -2987 1506
rect -2953 130 -2947 1506
rect -2993 118 -2947 130
rect -2795 1506 -2749 1518
rect -2795 130 -2789 1506
rect -2755 130 -2749 1506
rect -2795 118 -2749 130
rect -2597 1506 -2551 1518
rect -2597 130 -2591 1506
rect -2557 130 -2551 1506
rect -2597 118 -2551 130
rect -2399 1506 -2353 1518
rect -2399 130 -2393 1506
rect -2359 130 -2353 1506
rect -2399 118 -2353 130
rect -2201 1506 -2155 1518
rect -2201 130 -2195 1506
rect -2161 130 -2155 1506
rect -2201 118 -2155 130
rect -2003 1506 -1957 1518
rect -2003 130 -1997 1506
rect -1963 130 -1957 1506
rect -2003 118 -1957 130
rect -1805 1506 -1759 1518
rect -1805 130 -1799 1506
rect -1765 130 -1759 1506
rect -1805 118 -1759 130
rect -1607 1506 -1561 1518
rect -1607 130 -1601 1506
rect -1567 130 -1561 1506
rect -1607 118 -1561 130
rect -1409 1506 -1363 1518
rect -1409 130 -1403 1506
rect -1369 130 -1363 1506
rect -1409 118 -1363 130
rect -1211 1506 -1165 1518
rect -1211 130 -1205 1506
rect -1171 130 -1165 1506
rect -1211 118 -1165 130
rect -1013 1506 -967 1518
rect -1013 130 -1007 1506
rect -973 130 -967 1506
rect -1013 118 -967 130
rect -815 1506 -769 1518
rect -815 130 -809 1506
rect -775 130 -769 1506
rect -815 118 -769 130
rect -617 1506 -571 1518
rect -617 130 -611 1506
rect -577 130 -571 1506
rect -617 118 -571 130
rect -419 1506 -373 1518
rect -419 130 -413 1506
rect -379 130 -373 1506
rect -419 118 -373 130
rect -221 1506 -175 1518
rect -221 130 -215 1506
rect -181 130 -175 1506
rect -221 118 -175 130
rect -23 1506 23 1518
rect -23 130 -17 1506
rect 17 130 23 1506
rect -23 118 23 130
rect 175 1506 221 1518
rect 175 130 181 1506
rect 215 130 221 1506
rect 175 118 221 130
rect 373 1506 419 1518
rect 373 130 379 1506
rect 413 130 419 1506
rect 373 118 419 130
rect 571 1506 617 1518
rect 571 130 577 1506
rect 611 130 617 1506
rect 571 118 617 130
rect 769 1506 815 1518
rect 769 130 775 1506
rect 809 130 815 1506
rect 769 118 815 130
rect 967 1506 1013 1518
rect 967 130 973 1506
rect 1007 130 1013 1506
rect 967 118 1013 130
rect 1165 1506 1211 1518
rect 1165 130 1171 1506
rect 1205 130 1211 1506
rect 1165 118 1211 130
rect 1363 1506 1409 1518
rect 1363 130 1369 1506
rect 1403 130 1409 1506
rect 1363 118 1409 130
rect 1561 1506 1607 1518
rect 1561 130 1567 1506
rect 1601 130 1607 1506
rect 1561 118 1607 130
rect 1759 1506 1805 1518
rect 1759 130 1765 1506
rect 1799 130 1805 1506
rect 1759 118 1805 130
rect 1957 1506 2003 1518
rect 1957 130 1963 1506
rect 1997 130 2003 1506
rect 1957 118 2003 130
rect 2155 1506 2201 1518
rect 2155 130 2161 1506
rect 2195 130 2201 1506
rect 2155 118 2201 130
rect 2353 1506 2399 1518
rect 2353 130 2359 1506
rect 2393 130 2399 1506
rect 2353 118 2399 130
rect 2551 1506 2597 1518
rect 2551 130 2557 1506
rect 2591 130 2597 1506
rect 2551 118 2597 130
rect 2749 1506 2795 1518
rect 2749 130 2755 1506
rect 2789 130 2795 1506
rect 2749 118 2795 130
rect 2947 1506 2993 1518
rect 2947 130 2953 1506
rect 2987 130 2993 1506
rect 2947 118 2993 130
rect 3145 1506 3191 1518
rect 3145 130 3151 1506
rect 3185 130 3191 1506
rect 3145 118 3191 130
rect 3343 1506 3389 1518
rect 3343 130 3349 1506
rect 3383 130 3389 1506
rect 3343 118 3389 130
rect 3541 1506 3587 1518
rect 3541 130 3547 1506
rect 3581 130 3587 1506
rect 3541 118 3587 130
rect 3739 1506 3785 1518
rect 3739 130 3745 1506
rect 3779 130 3785 1506
rect 3739 118 3785 130
rect 3937 1506 3983 1518
rect 3937 130 3943 1506
rect 3977 130 3983 1506
rect 3937 118 3983 130
rect 4135 1506 4181 1518
rect 4135 130 4141 1506
rect 4175 130 4181 1506
rect 4135 118 4181 130
rect -4125 71 -3993 77
rect -4125 37 -4113 71
rect -4005 37 -3993 71
rect -4125 31 -3993 37
rect -3927 71 -3795 77
rect -3927 37 -3915 71
rect -3807 37 -3795 71
rect -3927 31 -3795 37
rect -3729 71 -3597 77
rect -3729 37 -3717 71
rect -3609 37 -3597 71
rect -3729 31 -3597 37
rect -3531 71 -3399 77
rect -3531 37 -3519 71
rect -3411 37 -3399 71
rect -3531 31 -3399 37
rect -3333 71 -3201 77
rect -3333 37 -3321 71
rect -3213 37 -3201 71
rect -3333 31 -3201 37
rect -3135 71 -3003 77
rect -3135 37 -3123 71
rect -3015 37 -3003 71
rect -3135 31 -3003 37
rect -2937 71 -2805 77
rect -2937 37 -2925 71
rect -2817 37 -2805 71
rect -2937 31 -2805 37
rect -2739 71 -2607 77
rect -2739 37 -2727 71
rect -2619 37 -2607 71
rect -2739 31 -2607 37
rect -2541 71 -2409 77
rect -2541 37 -2529 71
rect -2421 37 -2409 71
rect -2541 31 -2409 37
rect -2343 71 -2211 77
rect -2343 37 -2331 71
rect -2223 37 -2211 71
rect -2343 31 -2211 37
rect -2145 71 -2013 77
rect -2145 37 -2133 71
rect -2025 37 -2013 71
rect -2145 31 -2013 37
rect -1947 71 -1815 77
rect -1947 37 -1935 71
rect -1827 37 -1815 71
rect -1947 31 -1815 37
rect -1749 71 -1617 77
rect -1749 37 -1737 71
rect -1629 37 -1617 71
rect -1749 31 -1617 37
rect -1551 71 -1419 77
rect -1551 37 -1539 71
rect -1431 37 -1419 71
rect -1551 31 -1419 37
rect -1353 71 -1221 77
rect -1353 37 -1341 71
rect -1233 37 -1221 71
rect -1353 31 -1221 37
rect -1155 71 -1023 77
rect -1155 37 -1143 71
rect -1035 37 -1023 71
rect -1155 31 -1023 37
rect -957 71 -825 77
rect -957 37 -945 71
rect -837 37 -825 71
rect -957 31 -825 37
rect -759 71 -627 77
rect -759 37 -747 71
rect -639 37 -627 71
rect -759 31 -627 37
rect -561 71 -429 77
rect -561 37 -549 71
rect -441 37 -429 71
rect -561 31 -429 37
rect -363 71 -231 77
rect -363 37 -351 71
rect -243 37 -231 71
rect -363 31 -231 37
rect -165 71 -33 77
rect -165 37 -153 71
rect -45 37 -33 71
rect -165 31 -33 37
rect 33 71 165 77
rect 33 37 45 71
rect 153 37 165 71
rect 33 31 165 37
rect 231 71 363 77
rect 231 37 243 71
rect 351 37 363 71
rect 231 31 363 37
rect 429 71 561 77
rect 429 37 441 71
rect 549 37 561 71
rect 429 31 561 37
rect 627 71 759 77
rect 627 37 639 71
rect 747 37 759 71
rect 627 31 759 37
rect 825 71 957 77
rect 825 37 837 71
rect 945 37 957 71
rect 825 31 957 37
rect 1023 71 1155 77
rect 1023 37 1035 71
rect 1143 37 1155 71
rect 1023 31 1155 37
rect 1221 71 1353 77
rect 1221 37 1233 71
rect 1341 37 1353 71
rect 1221 31 1353 37
rect 1419 71 1551 77
rect 1419 37 1431 71
rect 1539 37 1551 71
rect 1419 31 1551 37
rect 1617 71 1749 77
rect 1617 37 1629 71
rect 1737 37 1749 71
rect 1617 31 1749 37
rect 1815 71 1947 77
rect 1815 37 1827 71
rect 1935 37 1947 71
rect 1815 31 1947 37
rect 2013 71 2145 77
rect 2013 37 2025 71
rect 2133 37 2145 71
rect 2013 31 2145 37
rect 2211 71 2343 77
rect 2211 37 2223 71
rect 2331 37 2343 71
rect 2211 31 2343 37
rect 2409 71 2541 77
rect 2409 37 2421 71
rect 2529 37 2541 71
rect 2409 31 2541 37
rect 2607 71 2739 77
rect 2607 37 2619 71
rect 2727 37 2739 71
rect 2607 31 2739 37
rect 2805 71 2937 77
rect 2805 37 2817 71
rect 2925 37 2937 71
rect 2805 31 2937 37
rect 3003 71 3135 77
rect 3003 37 3015 71
rect 3123 37 3135 71
rect 3003 31 3135 37
rect 3201 71 3333 77
rect 3201 37 3213 71
rect 3321 37 3333 71
rect 3201 31 3333 37
rect 3399 71 3531 77
rect 3399 37 3411 71
rect 3519 37 3531 71
rect 3399 31 3531 37
rect 3597 71 3729 77
rect 3597 37 3609 71
rect 3717 37 3729 71
rect 3597 31 3729 37
rect 3795 71 3927 77
rect 3795 37 3807 71
rect 3915 37 3927 71
rect 3795 31 3927 37
rect 3993 71 4125 77
rect 3993 37 4005 71
rect 4113 37 4125 71
rect 3993 31 4125 37
rect -4125 -37 -3993 -31
rect -4125 -71 -4113 -37
rect -4005 -71 -3993 -37
rect -4125 -77 -3993 -71
rect -3927 -37 -3795 -31
rect -3927 -71 -3915 -37
rect -3807 -71 -3795 -37
rect -3927 -77 -3795 -71
rect -3729 -37 -3597 -31
rect -3729 -71 -3717 -37
rect -3609 -71 -3597 -37
rect -3729 -77 -3597 -71
rect -3531 -37 -3399 -31
rect -3531 -71 -3519 -37
rect -3411 -71 -3399 -37
rect -3531 -77 -3399 -71
rect -3333 -37 -3201 -31
rect -3333 -71 -3321 -37
rect -3213 -71 -3201 -37
rect -3333 -77 -3201 -71
rect -3135 -37 -3003 -31
rect -3135 -71 -3123 -37
rect -3015 -71 -3003 -37
rect -3135 -77 -3003 -71
rect -2937 -37 -2805 -31
rect -2937 -71 -2925 -37
rect -2817 -71 -2805 -37
rect -2937 -77 -2805 -71
rect -2739 -37 -2607 -31
rect -2739 -71 -2727 -37
rect -2619 -71 -2607 -37
rect -2739 -77 -2607 -71
rect -2541 -37 -2409 -31
rect -2541 -71 -2529 -37
rect -2421 -71 -2409 -37
rect -2541 -77 -2409 -71
rect -2343 -37 -2211 -31
rect -2343 -71 -2331 -37
rect -2223 -71 -2211 -37
rect -2343 -77 -2211 -71
rect -2145 -37 -2013 -31
rect -2145 -71 -2133 -37
rect -2025 -71 -2013 -37
rect -2145 -77 -2013 -71
rect -1947 -37 -1815 -31
rect -1947 -71 -1935 -37
rect -1827 -71 -1815 -37
rect -1947 -77 -1815 -71
rect -1749 -37 -1617 -31
rect -1749 -71 -1737 -37
rect -1629 -71 -1617 -37
rect -1749 -77 -1617 -71
rect -1551 -37 -1419 -31
rect -1551 -71 -1539 -37
rect -1431 -71 -1419 -37
rect -1551 -77 -1419 -71
rect -1353 -37 -1221 -31
rect -1353 -71 -1341 -37
rect -1233 -71 -1221 -37
rect -1353 -77 -1221 -71
rect -1155 -37 -1023 -31
rect -1155 -71 -1143 -37
rect -1035 -71 -1023 -37
rect -1155 -77 -1023 -71
rect -957 -37 -825 -31
rect -957 -71 -945 -37
rect -837 -71 -825 -37
rect -957 -77 -825 -71
rect -759 -37 -627 -31
rect -759 -71 -747 -37
rect -639 -71 -627 -37
rect -759 -77 -627 -71
rect -561 -37 -429 -31
rect -561 -71 -549 -37
rect -441 -71 -429 -37
rect -561 -77 -429 -71
rect -363 -37 -231 -31
rect -363 -71 -351 -37
rect -243 -71 -231 -37
rect -363 -77 -231 -71
rect -165 -37 -33 -31
rect -165 -71 -153 -37
rect -45 -71 -33 -37
rect -165 -77 -33 -71
rect 33 -37 165 -31
rect 33 -71 45 -37
rect 153 -71 165 -37
rect 33 -77 165 -71
rect 231 -37 363 -31
rect 231 -71 243 -37
rect 351 -71 363 -37
rect 231 -77 363 -71
rect 429 -37 561 -31
rect 429 -71 441 -37
rect 549 -71 561 -37
rect 429 -77 561 -71
rect 627 -37 759 -31
rect 627 -71 639 -37
rect 747 -71 759 -37
rect 627 -77 759 -71
rect 825 -37 957 -31
rect 825 -71 837 -37
rect 945 -71 957 -37
rect 825 -77 957 -71
rect 1023 -37 1155 -31
rect 1023 -71 1035 -37
rect 1143 -71 1155 -37
rect 1023 -77 1155 -71
rect 1221 -37 1353 -31
rect 1221 -71 1233 -37
rect 1341 -71 1353 -37
rect 1221 -77 1353 -71
rect 1419 -37 1551 -31
rect 1419 -71 1431 -37
rect 1539 -71 1551 -37
rect 1419 -77 1551 -71
rect 1617 -37 1749 -31
rect 1617 -71 1629 -37
rect 1737 -71 1749 -37
rect 1617 -77 1749 -71
rect 1815 -37 1947 -31
rect 1815 -71 1827 -37
rect 1935 -71 1947 -37
rect 1815 -77 1947 -71
rect 2013 -37 2145 -31
rect 2013 -71 2025 -37
rect 2133 -71 2145 -37
rect 2013 -77 2145 -71
rect 2211 -37 2343 -31
rect 2211 -71 2223 -37
rect 2331 -71 2343 -37
rect 2211 -77 2343 -71
rect 2409 -37 2541 -31
rect 2409 -71 2421 -37
rect 2529 -71 2541 -37
rect 2409 -77 2541 -71
rect 2607 -37 2739 -31
rect 2607 -71 2619 -37
rect 2727 -71 2739 -37
rect 2607 -77 2739 -71
rect 2805 -37 2937 -31
rect 2805 -71 2817 -37
rect 2925 -71 2937 -37
rect 2805 -77 2937 -71
rect 3003 -37 3135 -31
rect 3003 -71 3015 -37
rect 3123 -71 3135 -37
rect 3003 -77 3135 -71
rect 3201 -37 3333 -31
rect 3201 -71 3213 -37
rect 3321 -71 3333 -37
rect 3201 -77 3333 -71
rect 3399 -37 3531 -31
rect 3399 -71 3411 -37
rect 3519 -71 3531 -37
rect 3399 -77 3531 -71
rect 3597 -37 3729 -31
rect 3597 -71 3609 -37
rect 3717 -71 3729 -37
rect 3597 -77 3729 -71
rect 3795 -37 3927 -31
rect 3795 -71 3807 -37
rect 3915 -71 3927 -37
rect 3795 -77 3927 -71
rect 3993 -37 4125 -31
rect 3993 -71 4005 -37
rect 4113 -71 4125 -37
rect 3993 -77 4125 -71
rect -4181 -130 -4135 -118
rect -4181 -1506 -4175 -130
rect -4141 -1506 -4135 -130
rect -4181 -1518 -4135 -1506
rect -3983 -130 -3937 -118
rect -3983 -1506 -3977 -130
rect -3943 -1506 -3937 -130
rect -3983 -1518 -3937 -1506
rect -3785 -130 -3739 -118
rect -3785 -1506 -3779 -130
rect -3745 -1506 -3739 -130
rect -3785 -1518 -3739 -1506
rect -3587 -130 -3541 -118
rect -3587 -1506 -3581 -130
rect -3547 -1506 -3541 -130
rect -3587 -1518 -3541 -1506
rect -3389 -130 -3343 -118
rect -3389 -1506 -3383 -130
rect -3349 -1506 -3343 -130
rect -3389 -1518 -3343 -1506
rect -3191 -130 -3145 -118
rect -3191 -1506 -3185 -130
rect -3151 -1506 -3145 -130
rect -3191 -1518 -3145 -1506
rect -2993 -130 -2947 -118
rect -2993 -1506 -2987 -130
rect -2953 -1506 -2947 -130
rect -2993 -1518 -2947 -1506
rect -2795 -130 -2749 -118
rect -2795 -1506 -2789 -130
rect -2755 -1506 -2749 -130
rect -2795 -1518 -2749 -1506
rect -2597 -130 -2551 -118
rect -2597 -1506 -2591 -130
rect -2557 -1506 -2551 -130
rect -2597 -1518 -2551 -1506
rect -2399 -130 -2353 -118
rect -2399 -1506 -2393 -130
rect -2359 -1506 -2353 -130
rect -2399 -1518 -2353 -1506
rect -2201 -130 -2155 -118
rect -2201 -1506 -2195 -130
rect -2161 -1506 -2155 -130
rect -2201 -1518 -2155 -1506
rect -2003 -130 -1957 -118
rect -2003 -1506 -1997 -130
rect -1963 -1506 -1957 -130
rect -2003 -1518 -1957 -1506
rect -1805 -130 -1759 -118
rect -1805 -1506 -1799 -130
rect -1765 -1506 -1759 -130
rect -1805 -1518 -1759 -1506
rect -1607 -130 -1561 -118
rect -1607 -1506 -1601 -130
rect -1567 -1506 -1561 -130
rect -1607 -1518 -1561 -1506
rect -1409 -130 -1363 -118
rect -1409 -1506 -1403 -130
rect -1369 -1506 -1363 -130
rect -1409 -1518 -1363 -1506
rect -1211 -130 -1165 -118
rect -1211 -1506 -1205 -130
rect -1171 -1506 -1165 -130
rect -1211 -1518 -1165 -1506
rect -1013 -130 -967 -118
rect -1013 -1506 -1007 -130
rect -973 -1506 -967 -130
rect -1013 -1518 -967 -1506
rect -815 -130 -769 -118
rect -815 -1506 -809 -130
rect -775 -1506 -769 -130
rect -815 -1518 -769 -1506
rect -617 -130 -571 -118
rect -617 -1506 -611 -130
rect -577 -1506 -571 -130
rect -617 -1518 -571 -1506
rect -419 -130 -373 -118
rect -419 -1506 -413 -130
rect -379 -1506 -373 -130
rect -419 -1518 -373 -1506
rect -221 -130 -175 -118
rect -221 -1506 -215 -130
rect -181 -1506 -175 -130
rect -221 -1518 -175 -1506
rect -23 -130 23 -118
rect -23 -1506 -17 -130
rect 17 -1506 23 -130
rect -23 -1518 23 -1506
rect 175 -130 221 -118
rect 175 -1506 181 -130
rect 215 -1506 221 -130
rect 175 -1518 221 -1506
rect 373 -130 419 -118
rect 373 -1506 379 -130
rect 413 -1506 419 -130
rect 373 -1518 419 -1506
rect 571 -130 617 -118
rect 571 -1506 577 -130
rect 611 -1506 617 -130
rect 571 -1518 617 -1506
rect 769 -130 815 -118
rect 769 -1506 775 -130
rect 809 -1506 815 -130
rect 769 -1518 815 -1506
rect 967 -130 1013 -118
rect 967 -1506 973 -130
rect 1007 -1506 1013 -130
rect 967 -1518 1013 -1506
rect 1165 -130 1211 -118
rect 1165 -1506 1171 -130
rect 1205 -1506 1211 -130
rect 1165 -1518 1211 -1506
rect 1363 -130 1409 -118
rect 1363 -1506 1369 -130
rect 1403 -1506 1409 -130
rect 1363 -1518 1409 -1506
rect 1561 -130 1607 -118
rect 1561 -1506 1567 -130
rect 1601 -1506 1607 -130
rect 1561 -1518 1607 -1506
rect 1759 -130 1805 -118
rect 1759 -1506 1765 -130
rect 1799 -1506 1805 -130
rect 1759 -1518 1805 -1506
rect 1957 -130 2003 -118
rect 1957 -1506 1963 -130
rect 1997 -1506 2003 -130
rect 1957 -1518 2003 -1506
rect 2155 -130 2201 -118
rect 2155 -1506 2161 -130
rect 2195 -1506 2201 -130
rect 2155 -1518 2201 -1506
rect 2353 -130 2399 -118
rect 2353 -1506 2359 -130
rect 2393 -1506 2399 -130
rect 2353 -1518 2399 -1506
rect 2551 -130 2597 -118
rect 2551 -1506 2557 -130
rect 2591 -1506 2597 -130
rect 2551 -1518 2597 -1506
rect 2749 -130 2795 -118
rect 2749 -1506 2755 -130
rect 2789 -1506 2795 -130
rect 2749 -1518 2795 -1506
rect 2947 -130 2993 -118
rect 2947 -1506 2953 -130
rect 2987 -1506 2993 -130
rect 2947 -1518 2993 -1506
rect 3145 -130 3191 -118
rect 3145 -1506 3151 -130
rect 3185 -1506 3191 -130
rect 3145 -1518 3191 -1506
rect 3343 -130 3389 -118
rect 3343 -1506 3349 -130
rect 3383 -1506 3389 -130
rect 3343 -1518 3389 -1506
rect 3541 -130 3587 -118
rect 3541 -1506 3547 -130
rect 3581 -1506 3587 -130
rect 3541 -1518 3587 -1506
rect 3739 -130 3785 -118
rect 3739 -1506 3745 -130
rect 3779 -1506 3785 -130
rect 3739 -1518 3785 -1506
rect 3937 -130 3983 -118
rect 3937 -1506 3943 -130
rect 3977 -1506 3983 -130
rect 3937 -1518 3983 -1506
rect 4135 -130 4181 -118
rect 4135 -1506 4141 -130
rect 4175 -1506 4181 -130
rect 4135 -1518 4181 -1506
rect -4125 -1565 -3993 -1559
rect -4125 -1599 -4113 -1565
rect -4005 -1599 -3993 -1565
rect -4125 -1605 -3993 -1599
rect -3927 -1565 -3795 -1559
rect -3927 -1599 -3915 -1565
rect -3807 -1599 -3795 -1565
rect -3927 -1605 -3795 -1599
rect -3729 -1565 -3597 -1559
rect -3729 -1599 -3717 -1565
rect -3609 -1599 -3597 -1565
rect -3729 -1605 -3597 -1599
rect -3531 -1565 -3399 -1559
rect -3531 -1599 -3519 -1565
rect -3411 -1599 -3399 -1565
rect -3531 -1605 -3399 -1599
rect -3333 -1565 -3201 -1559
rect -3333 -1599 -3321 -1565
rect -3213 -1599 -3201 -1565
rect -3333 -1605 -3201 -1599
rect -3135 -1565 -3003 -1559
rect -3135 -1599 -3123 -1565
rect -3015 -1599 -3003 -1565
rect -3135 -1605 -3003 -1599
rect -2937 -1565 -2805 -1559
rect -2937 -1599 -2925 -1565
rect -2817 -1599 -2805 -1565
rect -2937 -1605 -2805 -1599
rect -2739 -1565 -2607 -1559
rect -2739 -1599 -2727 -1565
rect -2619 -1599 -2607 -1565
rect -2739 -1605 -2607 -1599
rect -2541 -1565 -2409 -1559
rect -2541 -1599 -2529 -1565
rect -2421 -1599 -2409 -1565
rect -2541 -1605 -2409 -1599
rect -2343 -1565 -2211 -1559
rect -2343 -1599 -2331 -1565
rect -2223 -1599 -2211 -1565
rect -2343 -1605 -2211 -1599
rect -2145 -1565 -2013 -1559
rect -2145 -1599 -2133 -1565
rect -2025 -1599 -2013 -1565
rect -2145 -1605 -2013 -1599
rect -1947 -1565 -1815 -1559
rect -1947 -1599 -1935 -1565
rect -1827 -1599 -1815 -1565
rect -1947 -1605 -1815 -1599
rect -1749 -1565 -1617 -1559
rect -1749 -1599 -1737 -1565
rect -1629 -1599 -1617 -1565
rect -1749 -1605 -1617 -1599
rect -1551 -1565 -1419 -1559
rect -1551 -1599 -1539 -1565
rect -1431 -1599 -1419 -1565
rect -1551 -1605 -1419 -1599
rect -1353 -1565 -1221 -1559
rect -1353 -1599 -1341 -1565
rect -1233 -1599 -1221 -1565
rect -1353 -1605 -1221 -1599
rect -1155 -1565 -1023 -1559
rect -1155 -1599 -1143 -1565
rect -1035 -1599 -1023 -1565
rect -1155 -1605 -1023 -1599
rect -957 -1565 -825 -1559
rect -957 -1599 -945 -1565
rect -837 -1599 -825 -1565
rect -957 -1605 -825 -1599
rect -759 -1565 -627 -1559
rect -759 -1599 -747 -1565
rect -639 -1599 -627 -1565
rect -759 -1605 -627 -1599
rect -561 -1565 -429 -1559
rect -561 -1599 -549 -1565
rect -441 -1599 -429 -1565
rect -561 -1605 -429 -1599
rect -363 -1565 -231 -1559
rect -363 -1599 -351 -1565
rect -243 -1599 -231 -1565
rect -363 -1605 -231 -1599
rect -165 -1565 -33 -1559
rect -165 -1599 -153 -1565
rect -45 -1599 -33 -1565
rect -165 -1605 -33 -1599
rect 33 -1565 165 -1559
rect 33 -1599 45 -1565
rect 153 -1599 165 -1565
rect 33 -1605 165 -1599
rect 231 -1565 363 -1559
rect 231 -1599 243 -1565
rect 351 -1599 363 -1565
rect 231 -1605 363 -1599
rect 429 -1565 561 -1559
rect 429 -1599 441 -1565
rect 549 -1599 561 -1565
rect 429 -1605 561 -1599
rect 627 -1565 759 -1559
rect 627 -1599 639 -1565
rect 747 -1599 759 -1565
rect 627 -1605 759 -1599
rect 825 -1565 957 -1559
rect 825 -1599 837 -1565
rect 945 -1599 957 -1565
rect 825 -1605 957 -1599
rect 1023 -1565 1155 -1559
rect 1023 -1599 1035 -1565
rect 1143 -1599 1155 -1565
rect 1023 -1605 1155 -1599
rect 1221 -1565 1353 -1559
rect 1221 -1599 1233 -1565
rect 1341 -1599 1353 -1565
rect 1221 -1605 1353 -1599
rect 1419 -1565 1551 -1559
rect 1419 -1599 1431 -1565
rect 1539 -1599 1551 -1565
rect 1419 -1605 1551 -1599
rect 1617 -1565 1749 -1559
rect 1617 -1599 1629 -1565
rect 1737 -1599 1749 -1565
rect 1617 -1605 1749 -1599
rect 1815 -1565 1947 -1559
rect 1815 -1599 1827 -1565
rect 1935 -1599 1947 -1565
rect 1815 -1605 1947 -1599
rect 2013 -1565 2145 -1559
rect 2013 -1599 2025 -1565
rect 2133 -1599 2145 -1565
rect 2013 -1605 2145 -1599
rect 2211 -1565 2343 -1559
rect 2211 -1599 2223 -1565
rect 2331 -1599 2343 -1565
rect 2211 -1605 2343 -1599
rect 2409 -1565 2541 -1559
rect 2409 -1599 2421 -1565
rect 2529 -1599 2541 -1565
rect 2409 -1605 2541 -1599
rect 2607 -1565 2739 -1559
rect 2607 -1599 2619 -1565
rect 2727 -1599 2739 -1565
rect 2607 -1605 2739 -1599
rect 2805 -1565 2937 -1559
rect 2805 -1599 2817 -1565
rect 2925 -1599 2937 -1565
rect 2805 -1605 2937 -1599
rect 3003 -1565 3135 -1559
rect 3003 -1599 3015 -1565
rect 3123 -1599 3135 -1565
rect 3003 -1605 3135 -1599
rect 3201 -1565 3333 -1559
rect 3201 -1599 3213 -1565
rect 3321 -1599 3333 -1565
rect 3201 -1605 3333 -1599
rect 3399 -1565 3531 -1559
rect 3399 -1599 3411 -1565
rect 3519 -1599 3531 -1565
rect 3399 -1605 3531 -1599
rect 3597 -1565 3729 -1559
rect 3597 -1599 3609 -1565
rect 3717 -1599 3729 -1565
rect 3597 -1605 3729 -1599
rect 3795 -1565 3927 -1559
rect 3795 -1599 3807 -1565
rect 3915 -1599 3927 -1565
rect 3795 -1605 3927 -1599
rect 3993 -1565 4125 -1559
rect 3993 -1599 4005 -1565
rect 4113 -1599 4125 -1565
rect 3993 -1605 4125 -1599
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 7 l 0.7 m 2 nf 42 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
