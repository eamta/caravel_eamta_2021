magic
tech sky130A
magscale 1 2
timestamp 1615909117
<< error_p >>
rect -2920 -236 -2862 -230
rect -2802 -236 -2744 -230
rect -2684 -236 -2626 -230
rect -2566 -236 -2508 -230
rect -2448 -236 -2390 -230
rect -2330 -236 -2272 -230
rect -2212 -236 -2154 -230
rect -2094 -236 -2036 -230
rect -1976 -236 -1918 -230
rect -1858 -236 -1800 -230
rect -1740 -236 -1682 -230
rect -1622 -236 -1564 -230
rect -1504 -236 -1446 -230
rect -1386 -236 -1328 -230
rect -1268 -236 -1210 -230
rect -1150 -236 -1092 -230
rect -1032 -236 -974 -230
rect -914 -236 -856 -230
rect -796 -236 -738 -230
rect -678 -236 -620 -230
rect -560 -236 -502 -230
rect -442 -236 -384 -230
rect -324 -236 -266 -230
rect -206 -236 -148 -230
rect -88 -236 -30 -230
rect 30 -236 88 -230
rect 148 -236 206 -230
rect 266 -236 324 -230
rect 384 -236 442 -230
rect 502 -236 560 -230
rect 620 -236 678 -230
rect 738 -236 796 -230
rect 856 -236 914 -230
rect 974 -236 1032 -230
rect 1092 -236 1150 -230
rect 1210 -236 1268 -230
rect 1328 -236 1386 -230
rect 1446 -236 1504 -230
rect 1564 -236 1622 -230
rect 1682 -236 1740 -230
rect 1800 -236 1858 -230
rect 1918 -236 1976 -230
rect 2036 -236 2094 -230
rect 2154 -236 2212 -230
rect 2272 -236 2330 -230
rect 2390 -236 2448 -230
rect 2508 -236 2566 -230
rect 2626 -236 2684 -230
rect 2744 -236 2802 -230
rect 2862 -236 2920 -230
rect -2920 -270 -2908 -236
rect -2802 -270 -2790 -236
rect -2684 -270 -2672 -236
rect -2566 -270 -2554 -236
rect -2448 -270 -2436 -236
rect -2330 -270 -2318 -236
rect -2212 -270 -2200 -236
rect -2094 -270 -2082 -236
rect -1976 -270 -1964 -236
rect -1858 -270 -1846 -236
rect -1740 -270 -1728 -236
rect -1622 -270 -1610 -236
rect -1504 -270 -1492 -236
rect -1386 -270 -1374 -236
rect -1268 -270 -1256 -236
rect -1150 -270 -1138 -236
rect -1032 -270 -1020 -236
rect -914 -270 -902 -236
rect -796 -270 -784 -236
rect -678 -270 -666 -236
rect -560 -270 -548 -236
rect -442 -270 -430 -236
rect -324 -270 -312 -236
rect -206 -270 -194 -236
rect -88 -270 -76 -236
rect 30 -270 42 -236
rect 148 -270 160 -236
rect 266 -270 278 -236
rect 384 -270 396 -236
rect 502 -270 514 -236
rect 620 -270 632 -236
rect 738 -270 750 -236
rect 856 -270 868 -236
rect 974 -270 986 -236
rect 1092 -270 1104 -236
rect 1210 -270 1222 -236
rect 1328 -270 1340 -236
rect 1446 -270 1458 -236
rect 1564 -270 1576 -236
rect 1682 -270 1694 -236
rect 1800 -270 1812 -236
rect 1918 -270 1930 -236
rect 2036 -270 2048 -236
rect 2154 -270 2166 -236
rect 2272 -270 2284 -236
rect 2390 -270 2402 -236
rect 2508 -270 2520 -236
rect 2626 -270 2638 -236
rect 2744 -270 2756 -236
rect 2862 -270 2874 -236
rect -2920 -276 -2862 -270
rect -2802 -276 -2744 -270
rect -2684 -276 -2626 -270
rect -2566 -276 -2508 -270
rect -2448 -276 -2390 -270
rect -2330 -276 -2272 -270
rect -2212 -276 -2154 -270
rect -2094 -276 -2036 -270
rect -1976 -276 -1918 -270
rect -1858 -276 -1800 -270
rect -1740 -276 -1682 -270
rect -1622 -276 -1564 -270
rect -1504 -276 -1446 -270
rect -1386 -276 -1328 -270
rect -1268 -276 -1210 -270
rect -1150 -276 -1092 -270
rect -1032 -276 -974 -270
rect -914 -276 -856 -270
rect -796 -276 -738 -270
rect -678 -276 -620 -270
rect -560 -276 -502 -270
rect -442 -276 -384 -270
rect -324 -276 -266 -270
rect -206 -276 -148 -270
rect -88 -276 -30 -270
rect 30 -276 88 -270
rect 148 -276 206 -270
rect 266 -276 324 -270
rect 384 -276 442 -270
rect 502 -276 560 -270
rect 620 -276 678 -270
rect 738 -276 796 -270
rect 856 -276 914 -270
rect 974 -276 1032 -270
rect 1092 -276 1150 -270
rect 1210 -276 1268 -270
rect 1328 -276 1386 -270
rect 1446 -276 1504 -270
rect 1564 -276 1622 -270
rect 1682 -276 1740 -270
rect 1800 -276 1858 -270
rect 1918 -276 1976 -270
rect 2036 -276 2094 -270
rect 2154 -276 2212 -270
rect 2272 -276 2330 -270
rect 2390 -276 2448 -270
rect 2508 -276 2566 -270
rect 2626 -276 2684 -270
rect 2744 -276 2802 -270
rect 2862 -276 2920 -270
<< nwell >>
rect -3117 -409 3117 409
<< pmos >>
rect -2921 -189 -2861 261
rect -2803 -189 -2743 261
rect -2685 -189 -2625 261
rect -2567 -189 -2507 261
rect -2449 -189 -2389 261
rect -2331 -189 -2271 261
rect -2213 -189 -2153 261
rect -2095 -189 -2035 261
rect -1977 -189 -1917 261
rect -1859 -189 -1799 261
rect -1741 -189 -1681 261
rect -1623 -189 -1563 261
rect -1505 -189 -1445 261
rect -1387 -189 -1327 261
rect -1269 -189 -1209 261
rect -1151 -189 -1091 261
rect -1033 -189 -973 261
rect -915 -189 -855 261
rect -797 -189 -737 261
rect -679 -189 -619 261
rect -561 -189 -501 261
rect -443 -189 -383 261
rect -325 -189 -265 261
rect -207 -189 -147 261
rect -89 -189 -29 261
rect 29 -189 89 261
rect 147 -189 207 261
rect 265 -189 325 261
rect 383 -189 443 261
rect 501 -189 561 261
rect 619 -189 679 261
rect 737 -189 797 261
rect 855 -189 915 261
rect 973 -189 1033 261
rect 1091 -189 1151 261
rect 1209 -189 1269 261
rect 1327 -189 1387 261
rect 1445 -189 1505 261
rect 1563 -189 1623 261
rect 1681 -189 1741 261
rect 1799 -189 1859 261
rect 1917 -189 1977 261
rect 2035 -189 2095 261
rect 2153 -189 2213 261
rect 2271 -189 2331 261
rect 2389 -189 2449 261
rect 2507 -189 2567 261
rect 2625 -189 2685 261
rect 2743 -189 2803 261
rect 2861 -189 2921 261
<< pdiff >>
rect -2979 249 -2921 261
rect -2979 -177 -2967 249
rect -2933 -177 -2921 249
rect -2979 -189 -2921 -177
rect -2861 249 -2803 261
rect -2861 -177 -2849 249
rect -2815 -177 -2803 249
rect -2861 -189 -2803 -177
rect -2743 249 -2685 261
rect -2743 -177 -2731 249
rect -2697 -177 -2685 249
rect -2743 -189 -2685 -177
rect -2625 249 -2567 261
rect -2625 -177 -2613 249
rect -2579 -177 -2567 249
rect -2625 -189 -2567 -177
rect -2507 249 -2449 261
rect -2507 -177 -2495 249
rect -2461 -177 -2449 249
rect -2507 -189 -2449 -177
rect -2389 249 -2331 261
rect -2389 -177 -2377 249
rect -2343 -177 -2331 249
rect -2389 -189 -2331 -177
rect -2271 249 -2213 261
rect -2271 -177 -2259 249
rect -2225 -177 -2213 249
rect -2271 -189 -2213 -177
rect -2153 249 -2095 261
rect -2153 -177 -2141 249
rect -2107 -177 -2095 249
rect -2153 -189 -2095 -177
rect -2035 249 -1977 261
rect -2035 -177 -2023 249
rect -1989 -177 -1977 249
rect -2035 -189 -1977 -177
rect -1917 249 -1859 261
rect -1917 -177 -1905 249
rect -1871 -177 -1859 249
rect -1917 -189 -1859 -177
rect -1799 249 -1741 261
rect -1799 -177 -1787 249
rect -1753 -177 -1741 249
rect -1799 -189 -1741 -177
rect -1681 249 -1623 261
rect -1681 -177 -1669 249
rect -1635 -177 -1623 249
rect -1681 -189 -1623 -177
rect -1563 249 -1505 261
rect -1563 -177 -1551 249
rect -1517 -177 -1505 249
rect -1563 -189 -1505 -177
rect -1445 249 -1387 261
rect -1445 -177 -1433 249
rect -1399 -177 -1387 249
rect -1445 -189 -1387 -177
rect -1327 249 -1269 261
rect -1327 -177 -1315 249
rect -1281 -177 -1269 249
rect -1327 -189 -1269 -177
rect -1209 249 -1151 261
rect -1209 -177 -1197 249
rect -1163 -177 -1151 249
rect -1209 -189 -1151 -177
rect -1091 249 -1033 261
rect -1091 -177 -1079 249
rect -1045 -177 -1033 249
rect -1091 -189 -1033 -177
rect -973 249 -915 261
rect -973 -177 -961 249
rect -927 -177 -915 249
rect -973 -189 -915 -177
rect -855 249 -797 261
rect -855 -177 -843 249
rect -809 -177 -797 249
rect -855 -189 -797 -177
rect -737 249 -679 261
rect -737 -177 -725 249
rect -691 -177 -679 249
rect -737 -189 -679 -177
rect -619 249 -561 261
rect -619 -177 -607 249
rect -573 -177 -561 249
rect -619 -189 -561 -177
rect -501 249 -443 261
rect -501 -177 -489 249
rect -455 -177 -443 249
rect -501 -189 -443 -177
rect -383 249 -325 261
rect -383 -177 -371 249
rect -337 -177 -325 249
rect -383 -189 -325 -177
rect -265 249 -207 261
rect -265 -177 -253 249
rect -219 -177 -207 249
rect -265 -189 -207 -177
rect -147 249 -89 261
rect -147 -177 -135 249
rect -101 -177 -89 249
rect -147 -189 -89 -177
rect -29 249 29 261
rect -29 -177 -17 249
rect 17 -177 29 249
rect -29 -189 29 -177
rect 89 249 147 261
rect 89 -177 101 249
rect 135 -177 147 249
rect 89 -189 147 -177
rect 207 249 265 261
rect 207 -177 219 249
rect 253 -177 265 249
rect 207 -189 265 -177
rect 325 249 383 261
rect 325 -177 337 249
rect 371 -177 383 249
rect 325 -189 383 -177
rect 443 249 501 261
rect 443 -177 455 249
rect 489 -177 501 249
rect 443 -189 501 -177
rect 561 249 619 261
rect 561 -177 573 249
rect 607 -177 619 249
rect 561 -189 619 -177
rect 679 249 737 261
rect 679 -177 691 249
rect 725 -177 737 249
rect 679 -189 737 -177
rect 797 249 855 261
rect 797 -177 809 249
rect 843 -177 855 249
rect 797 -189 855 -177
rect 915 249 973 261
rect 915 -177 927 249
rect 961 -177 973 249
rect 915 -189 973 -177
rect 1033 249 1091 261
rect 1033 -177 1045 249
rect 1079 -177 1091 249
rect 1033 -189 1091 -177
rect 1151 249 1209 261
rect 1151 -177 1163 249
rect 1197 -177 1209 249
rect 1151 -189 1209 -177
rect 1269 249 1327 261
rect 1269 -177 1281 249
rect 1315 -177 1327 249
rect 1269 -189 1327 -177
rect 1387 249 1445 261
rect 1387 -177 1399 249
rect 1433 -177 1445 249
rect 1387 -189 1445 -177
rect 1505 249 1563 261
rect 1505 -177 1517 249
rect 1551 -177 1563 249
rect 1505 -189 1563 -177
rect 1623 249 1681 261
rect 1623 -177 1635 249
rect 1669 -177 1681 249
rect 1623 -189 1681 -177
rect 1741 249 1799 261
rect 1741 -177 1753 249
rect 1787 -177 1799 249
rect 1741 -189 1799 -177
rect 1859 249 1917 261
rect 1859 -177 1871 249
rect 1905 -177 1917 249
rect 1859 -189 1917 -177
rect 1977 249 2035 261
rect 1977 -177 1989 249
rect 2023 -177 2035 249
rect 1977 -189 2035 -177
rect 2095 249 2153 261
rect 2095 -177 2107 249
rect 2141 -177 2153 249
rect 2095 -189 2153 -177
rect 2213 249 2271 261
rect 2213 -177 2225 249
rect 2259 -177 2271 249
rect 2213 -189 2271 -177
rect 2331 249 2389 261
rect 2331 -177 2343 249
rect 2377 -177 2389 249
rect 2331 -189 2389 -177
rect 2449 249 2507 261
rect 2449 -177 2461 249
rect 2495 -177 2507 249
rect 2449 -189 2507 -177
rect 2567 249 2625 261
rect 2567 -177 2579 249
rect 2613 -177 2625 249
rect 2567 -189 2625 -177
rect 2685 249 2743 261
rect 2685 -177 2697 249
rect 2731 -177 2743 249
rect 2685 -189 2743 -177
rect 2803 249 2861 261
rect 2803 -177 2815 249
rect 2849 -177 2861 249
rect 2803 -189 2861 -177
rect 2921 249 2979 261
rect 2921 -177 2933 249
rect 2967 -177 2979 249
rect 2921 -189 2979 -177
<< pdiffc >>
rect -2967 -177 -2933 249
rect -2849 -177 -2815 249
rect -2731 -177 -2697 249
rect -2613 -177 -2579 249
rect -2495 -177 -2461 249
rect -2377 -177 -2343 249
rect -2259 -177 -2225 249
rect -2141 -177 -2107 249
rect -2023 -177 -1989 249
rect -1905 -177 -1871 249
rect -1787 -177 -1753 249
rect -1669 -177 -1635 249
rect -1551 -177 -1517 249
rect -1433 -177 -1399 249
rect -1315 -177 -1281 249
rect -1197 -177 -1163 249
rect -1079 -177 -1045 249
rect -961 -177 -927 249
rect -843 -177 -809 249
rect -725 -177 -691 249
rect -607 -177 -573 249
rect -489 -177 -455 249
rect -371 -177 -337 249
rect -253 -177 -219 249
rect -135 -177 -101 249
rect -17 -177 17 249
rect 101 -177 135 249
rect 219 -177 253 249
rect 337 -177 371 249
rect 455 -177 489 249
rect 573 -177 607 249
rect 691 -177 725 249
rect 809 -177 843 249
rect 927 -177 961 249
rect 1045 -177 1079 249
rect 1163 -177 1197 249
rect 1281 -177 1315 249
rect 1399 -177 1433 249
rect 1517 -177 1551 249
rect 1635 -177 1669 249
rect 1753 -177 1787 249
rect 1871 -177 1905 249
rect 1989 -177 2023 249
rect 2107 -177 2141 249
rect 2225 -177 2259 249
rect 2343 -177 2377 249
rect 2461 -177 2495 249
rect 2579 -177 2613 249
rect 2697 -177 2731 249
rect 2815 -177 2849 249
rect 2933 -177 2967 249
<< nsubdiff >>
rect -3081 339 -2985 373
rect 2985 339 3081 373
rect -3081 276 -3047 339
rect 3047 276 3081 339
rect -3081 -339 -3047 -276
rect 3047 -339 3081 -276
rect -3081 -373 -2985 -339
rect 2985 -373 3081 -339
<< nsubdiffcont >>
rect -2985 339 2985 373
rect -3081 -276 -3047 276
rect 3047 -276 3081 276
rect -2985 -373 2985 -339
<< poly >>
rect -2921 261 -2861 287
rect -2803 261 -2743 287
rect -2685 261 -2625 287
rect -2567 261 -2507 287
rect -2449 261 -2389 287
rect -2331 261 -2271 287
rect -2213 261 -2153 287
rect -2095 261 -2035 287
rect -1977 261 -1917 287
rect -1859 261 -1799 287
rect -1741 261 -1681 287
rect -1623 261 -1563 287
rect -1505 261 -1445 287
rect -1387 261 -1327 287
rect -1269 261 -1209 287
rect -1151 261 -1091 287
rect -1033 261 -973 287
rect -915 261 -855 287
rect -797 261 -737 287
rect -679 261 -619 287
rect -561 261 -501 287
rect -443 261 -383 287
rect -325 261 -265 287
rect -207 261 -147 287
rect -89 261 -29 287
rect 29 261 89 287
rect 147 261 207 287
rect 265 261 325 287
rect 383 261 443 287
rect 501 261 561 287
rect 619 261 679 287
rect 737 261 797 287
rect 855 261 915 287
rect 973 261 1033 287
rect 1091 261 1151 287
rect 1209 261 1269 287
rect 1327 261 1387 287
rect 1445 261 1505 287
rect 1563 261 1623 287
rect 1681 261 1741 287
rect 1799 261 1859 287
rect 1917 261 1977 287
rect 2035 261 2095 287
rect 2153 261 2213 287
rect 2271 261 2331 287
rect 2389 261 2449 287
rect 2507 261 2567 287
rect 2625 261 2685 287
rect 2743 261 2803 287
rect 2861 261 2921 287
rect -2921 -220 -2861 -189
rect -2803 -220 -2743 -189
rect -2685 -220 -2625 -189
rect -2567 -220 -2507 -189
rect -2449 -220 -2389 -189
rect -2331 -220 -2271 -189
rect -2213 -220 -2153 -189
rect -2095 -220 -2035 -189
rect -1977 -220 -1917 -189
rect -1859 -220 -1799 -189
rect -1741 -220 -1681 -189
rect -1623 -220 -1563 -189
rect -1505 -220 -1445 -189
rect -1387 -220 -1327 -189
rect -1269 -220 -1209 -189
rect -1151 -220 -1091 -189
rect -1033 -220 -973 -189
rect -915 -220 -855 -189
rect -797 -220 -737 -189
rect -679 -220 -619 -189
rect -561 -220 -501 -189
rect -443 -220 -383 -189
rect -325 -220 -265 -189
rect -207 -220 -147 -189
rect -89 -220 -29 -189
rect 29 -220 89 -189
rect 147 -220 207 -189
rect 265 -220 325 -189
rect 383 -220 443 -189
rect 501 -220 561 -189
rect 619 -220 679 -189
rect 737 -220 797 -189
rect 855 -220 915 -189
rect 973 -220 1033 -189
rect 1091 -220 1151 -189
rect 1209 -220 1269 -189
rect 1327 -220 1387 -189
rect 1445 -220 1505 -189
rect 1563 -220 1623 -189
rect 1681 -220 1741 -189
rect 1799 -220 1859 -189
rect 1917 -220 1977 -189
rect 2035 -220 2095 -189
rect 2153 -220 2213 -189
rect 2271 -220 2331 -189
rect 2389 -220 2449 -189
rect 2507 -220 2567 -189
rect 2625 -220 2685 -189
rect 2743 -220 2803 -189
rect 2861 -220 2921 -189
rect -2924 -236 -2858 -220
rect -2924 -270 -2908 -236
rect -2874 -270 -2858 -236
rect -2924 -286 -2858 -270
rect -2806 -236 -2740 -220
rect -2806 -270 -2790 -236
rect -2756 -270 -2740 -236
rect -2806 -286 -2740 -270
rect -2688 -236 -2622 -220
rect -2688 -270 -2672 -236
rect -2638 -270 -2622 -236
rect -2688 -286 -2622 -270
rect -2570 -236 -2504 -220
rect -2570 -270 -2554 -236
rect -2520 -270 -2504 -236
rect -2570 -286 -2504 -270
rect -2452 -236 -2386 -220
rect -2452 -270 -2436 -236
rect -2402 -270 -2386 -236
rect -2452 -286 -2386 -270
rect -2334 -236 -2268 -220
rect -2334 -270 -2318 -236
rect -2284 -270 -2268 -236
rect -2334 -286 -2268 -270
rect -2216 -236 -2150 -220
rect -2216 -270 -2200 -236
rect -2166 -270 -2150 -236
rect -2216 -286 -2150 -270
rect -2098 -236 -2032 -220
rect -2098 -270 -2082 -236
rect -2048 -270 -2032 -236
rect -2098 -286 -2032 -270
rect -1980 -236 -1914 -220
rect -1980 -270 -1964 -236
rect -1930 -270 -1914 -236
rect -1980 -286 -1914 -270
rect -1862 -236 -1796 -220
rect -1862 -270 -1846 -236
rect -1812 -270 -1796 -236
rect -1862 -286 -1796 -270
rect -1744 -236 -1678 -220
rect -1744 -270 -1728 -236
rect -1694 -270 -1678 -236
rect -1744 -286 -1678 -270
rect -1626 -236 -1560 -220
rect -1626 -270 -1610 -236
rect -1576 -270 -1560 -236
rect -1626 -286 -1560 -270
rect -1508 -236 -1442 -220
rect -1508 -270 -1492 -236
rect -1458 -270 -1442 -236
rect -1508 -286 -1442 -270
rect -1390 -236 -1324 -220
rect -1390 -270 -1374 -236
rect -1340 -270 -1324 -236
rect -1390 -286 -1324 -270
rect -1272 -236 -1206 -220
rect -1272 -270 -1256 -236
rect -1222 -270 -1206 -236
rect -1272 -286 -1206 -270
rect -1154 -236 -1088 -220
rect -1154 -270 -1138 -236
rect -1104 -270 -1088 -236
rect -1154 -286 -1088 -270
rect -1036 -236 -970 -220
rect -1036 -270 -1020 -236
rect -986 -270 -970 -236
rect -1036 -286 -970 -270
rect -918 -236 -852 -220
rect -918 -270 -902 -236
rect -868 -270 -852 -236
rect -918 -286 -852 -270
rect -800 -236 -734 -220
rect -800 -270 -784 -236
rect -750 -270 -734 -236
rect -800 -286 -734 -270
rect -682 -236 -616 -220
rect -682 -270 -666 -236
rect -632 -270 -616 -236
rect -682 -286 -616 -270
rect -564 -236 -498 -220
rect -564 -270 -548 -236
rect -514 -270 -498 -236
rect -564 -286 -498 -270
rect -446 -236 -380 -220
rect -446 -270 -430 -236
rect -396 -270 -380 -236
rect -446 -286 -380 -270
rect -328 -236 -262 -220
rect -328 -270 -312 -236
rect -278 -270 -262 -236
rect -328 -286 -262 -270
rect -210 -236 -144 -220
rect -210 -270 -194 -236
rect -160 -270 -144 -236
rect -210 -286 -144 -270
rect -92 -236 -26 -220
rect -92 -270 -76 -236
rect -42 -270 -26 -236
rect -92 -286 -26 -270
rect 26 -236 92 -220
rect 26 -270 42 -236
rect 76 -270 92 -236
rect 26 -286 92 -270
rect 144 -236 210 -220
rect 144 -270 160 -236
rect 194 -270 210 -236
rect 144 -286 210 -270
rect 262 -236 328 -220
rect 262 -270 278 -236
rect 312 -270 328 -236
rect 262 -286 328 -270
rect 380 -236 446 -220
rect 380 -270 396 -236
rect 430 -270 446 -236
rect 380 -286 446 -270
rect 498 -236 564 -220
rect 498 -270 514 -236
rect 548 -270 564 -236
rect 498 -286 564 -270
rect 616 -236 682 -220
rect 616 -270 632 -236
rect 666 -270 682 -236
rect 616 -286 682 -270
rect 734 -236 800 -220
rect 734 -270 750 -236
rect 784 -270 800 -236
rect 734 -286 800 -270
rect 852 -236 918 -220
rect 852 -270 868 -236
rect 902 -270 918 -236
rect 852 -286 918 -270
rect 970 -236 1036 -220
rect 970 -270 986 -236
rect 1020 -270 1036 -236
rect 970 -286 1036 -270
rect 1088 -236 1154 -220
rect 1088 -270 1104 -236
rect 1138 -270 1154 -236
rect 1088 -286 1154 -270
rect 1206 -236 1272 -220
rect 1206 -270 1222 -236
rect 1256 -270 1272 -236
rect 1206 -286 1272 -270
rect 1324 -236 1390 -220
rect 1324 -270 1340 -236
rect 1374 -270 1390 -236
rect 1324 -286 1390 -270
rect 1442 -236 1508 -220
rect 1442 -270 1458 -236
rect 1492 -270 1508 -236
rect 1442 -286 1508 -270
rect 1560 -236 1626 -220
rect 1560 -270 1576 -236
rect 1610 -270 1626 -236
rect 1560 -286 1626 -270
rect 1678 -236 1744 -220
rect 1678 -270 1694 -236
rect 1728 -270 1744 -236
rect 1678 -286 1744 -270
rect 1796 -236 1862 -220
rect 1796 -270 1812 -236
rect 1846 -270 1862 -236
rect 1796 -286 1862 -270
rect 1914 -236 1980 -220
rect 1914 -270 1930 -236
rect 1964 -270 1980 -236
rect 1914 -286 1980 -270
rect 2032 -236 2098 -220
rect 2032 -270 2048 -236
rect 2082 -270 2098 -236
rect 2032 -286 2098 -270
rect 2150 -236 2216 -220
rect 2150 -270 2166 -236
rect 2200 -270 2216 -236
rect 2150 -286 2216 -270
rect 2268 -236 2334 -220
rect 2268 -270 2284 -236
rect 2318 -270 2334 -236
rect 2268 -286 2334 -270
rect 2386 -236 2452 -220
rect 2386 -270 2402 -236
rect 2436 -270 2452 -236
rect 2386 -286 2452 -270
rect 2504 -236 2570 -220
rect 2504 -270 2520 -236
rect 2554 -270 2570 -236
rect 2504 -286 2570 -270
rect 2622 -236 2688 -220
rect 2622 -270 2638 -236
rect 2672 -270 2688 -236
rect 2622 -286 2688 -270
rect 2740 -236 2806 -220
rect 2740 -270 2756 -236
rect 2790 -270 2806 -236
rect 2740 -286 2806 -270
rect 2858 -236 2924 -220
rect 2858 -270 2874 -236
rect 2908 -270 2924 -236
rect 2858 -286 2924 -270
<< polycont >>
rect -2908 -270 -2874 -236
rect -2790 -270 -2756 -236
rect -2672 -270 -2638 -236
rect -2554 -270 -2520 -236
rect -2436 -270 -2402 -236
rect -2318 -270 -2284 -236
rect -2200 -270 -2166 -236
rect -2082 -270 -2048 -236
rect -1964 -270 -1930 -236
rect -1846 -270 -1812 -236
rect -1728 -270 -1694 -236
rect -1610 -270 -1576 -236
rect -1492 -270 -1458 -236
rect -1374 -270 -1340 -236
rect -1256 -270 -1222 -236
rect -1138 -270 -1104 -236
rect -1020 -270 -986 -236
rect -902 -270 -868 -236
rect -784 -270 -750 -236
rect -666 -270 -632 -236
rect -548 -270 -514 -236
rect -430 -270 -396 -236
rect -312 -270 -278 -236
rect -194 -270 -160 -236
rect -76 -270 -42 -236
rect 42 -270 76 -236
rect 160 -270 194 -236
rect 278 -270 312 -236
rect 396 -270 430 -236
rect 514 -270 548 -236
rect 632 -270 666 -236
rect 750 -270 784 -236
rect 868 -270 902 -236
rect 986 -270 1020 -236
rect 1104 -270 1138 -236
rect 1222 -270 1256 -236
rect 1340 -270 1374 -236
rect 1458 -270 1492 -236
rect 1576 -270 1610 -236
rect 1694 -270 1728 -236
rect 1812 -270 1846 -236
rect 1930 -270 1964 -236
rect 2048 -270 2082 -236
rect 2166 -270 2200 -236
rect 2284 -270 2318 -236
rect 2402 -270 2436 -236
rect 2520 -270 2554 -236
rect 2638 -270 2672 -236
rect 2756 -270 2790 -236
rect 2874 -270 2908 -236
<< locali >>
rect -3081 339 -2985 373
rect 2985 339 3081 373
rect -3081 276 -3047 339
rect 3047 276 3081 339
rect -2967 249 -2933 265
rect -2967 -193 -2933 -177
rect -2849 249 -2815 265
rect -2849 -193 -2815 -177
rect -2731 249 -2697 265
rect -2731 -193 -2697 -177
rect -2613 249 -2579 265
rect -2613 -193 -2579 -177
rect -2495 249 -2461 265
rect -2495 -193 -2461 -177
rect -2377 249 -2343 265
rect -2377 -193 -2343 -177
rect -2259 249 -2225 265
rect -2259 -193 -2225 -177
rect -2141 249 -2107 265
rect -2141 -193 -2107 -177
rect -2023 249 -1989 265
rect -2023 -193 -1989 -177
rect -1905 249 -1871 265
rect -1905 -193 -1871 -177
rect -1787 249 -1753 265
rect -1787 -193 -1753 -177
rect -1669 249 -1635 265
rect -1669 -193 -1635 -177
rect -1551 249 -1517 265
rect -1551 -193 -1517 -177
rect -1433 249 -1399 265
rect -1433 -193 -1399 -177
rect -1315 249 -1281 265
rect -1315 -193 -1281 -177
rect -1197 249 -1163 265
rect -1197 -193 -1163 -177
rect -1079 249 -1045 265
rect -1079 -193 -1045 -177
rect -961 249 -927 265
rect -961 -193 -927 -177
rect -843 249 -809 265
rect -843 -193 -809 -177
rect -725 249 -691 265
rect -725 -193 -691 -177
rect -607 249 -573 265
rect -607 -193 -573 -177
rect -489 249 -455 265
rect -489 -193 -455 -177
rect -371 249 -337 265
rect -371 -193 -337 -177
rect -253 249 -219 265
rect -253 -193 -219 -177
rect -135 249 -101 265
rect -135 -193 -101 -177
rect -17 249 17 265
rect -17 -193 17 -177
rect 101 249 135 265
rect 101 -193 135 -177
rect 219 249 253 265
rect 219 -193 253 -177
rect 337 249 371 265
rect 337 -193 371 -177
rect 455 249 489 265
rect 455 -193 489 -177
rect 573 249 607 265
rect 573 -193 607 -177
rect 691 249 725 265
rect 691 -193 725 -177
rect 809 249 843 265
rect 809 -193 843 -177
rect 927 249 961 265
rect 927 -193 961 -177
rect 1045 249 1079 265
rect 1045 -193 1079 -177
rect 1163 249 1197 265
rect 1163 -193 1197 -177
rect 1281 249 1315 265
rect 1281 -193 1315 -177
rect 1399 249 1433 265
rect 1399 -193 1433 -177
rect 1517 249 1551 265
rect 1517 -193 1551 -177
rect 1635 249 1669 265
rect 1635 -193 1669 -177
rect 1753 249 1787 265
rect 1753 -193 1787 -177
rect 1871 249 1905 265
rect 1871 -193 1905 -177
rect 1989 249 2023 265
rect 1989 -193 2023 -177
rect 2107 249 2141 265
rect 2107 -193 2141 -177
rect 2225 249 2259 265
rect 2225 -193 2259 -177
rect 2343 249 2377 265
rect 2343 -193 2377 -177
rect 2461 249 2495 265
rect 2461 -193 2495 -177
rect 2579 249 2613 265
rect 2579 -193 2613 -177
rect 2697 249 2731 265
rect 2697 -193 2731 -177
rect 2815 249 2849 265
rect 2815 -193 2849 -177
rect 2933 249 2967 265
rect 2933 -193 2967 -177
rect -2924 -270 -2908 -236
rect -2874 -270 -2858 -236
rect -2806 -270 -2790 -236
rect -2756 -270 -2740 -236
rect -2688 -270 -2672 -236
rect -2638 -270 -2622 -236
rect -2570 -270 -2554 -236
rect -2520 -270 -2504 -236
rect -2452 -270 -2436 -236
rect -2402 -270 -2386 -236
rect -2334 -270 -2318 -236
rect -2284 -270 -2268 -236
rect -2216 -270 -2200 -236
rect -2166 -270 -2150 -236
rect -2098 -270 -2082 -236
rect -2048 -270 -2032 -236
rect -1980 -270 -1964 -236
rect -1930 -270 -1914 -236
rect -1862 -270 -1846 -236
rect -1812 -270 -1796 -236
rect -1744 -270 -1728 -236
rect -1694 -270 -1678 -236
rect -1626 -270 -1610 -236
rect -1576 -270 -1560 -236
rect -1508 -270 -1492 -236
rect -1458 -270 -1442 -236
rect -1390 -270 -1374 -236
rect -1340 -270 -1324 -236
rect -1272 -270 -1256 -236
rect -1222 -270 -1206 -236
rect -1154 -270 -1138 -236
rect -1104 -270 -1088 -236
rect -1036 -270 -1020 -236
rect -986 -270 -970 -236
rect -918 -270 -902 -236
rect -868 -270 -852 -236
rect -800 -270 -784 -236
rect -750 -270 -734 -236
rect -682 -270 -666 -236
rect -632 -270 -616 -236
rect -564 -270 -548 -236
rect -514 -270 -498 -236
rect -446 -270 -430 -236
rect -396 -270 -380 -236
rect -328 -270 -312 -236
rect -278 -270 -262 -236
rect -210 -270 -194 -236
rect -160 -270 -144 -236
rect -92 -270 -76 -236
rect -42 -270 -26 -236
rect 26 -270 42 -236
rect 76 -270 92 -236
rect 144 -270 160 -236
rect 194 -270 210 -236
rect 262 -270 278 -236
rect 312 -270 328 -236
rect 380 -270 396 -236
rect 430 -270 446 -236
rect 498 -270 514 -236
rect 548 -270 564 -236
rect 616 -270 632 -236
rect 666 -270 682 -236
rect 734 -270 750 -236
rect 784 -270 800 -236
rect 852 -270 868 -236
rect 902 -270 918 -236
rect 970 -270 986 -236
rect 1020 -270 1036 -236
rect 1088 -270 1104 -236
rect 1138 -270 1154 -236
rect 1206 -270 1222 -236
rect 1256 -270 1272 -236
rect 1324 -270 1340 -236
rect 1374 -270 1390 -236
rect 1442 -270 1458 -236
rect 1492 -270 1508 -236
rect 1560 -270 1576 -236
rect 1610 -270 1626 -236
rect 1678 -270 1694 -236
rect 1728 -270 1744 -236
rect 1796 -270 1812 -236
rect 1846 -270 1862 -236
rect 1914 -270 1930 -236
rect 1964 -270 1980 -236
rect 2032 -270 2048 -236
rect 2082 -270 2098 -236
rect 2150 -270 2166 -236
rect 2200 -270 2216 -236
rect 2268 -270 2284 -236
rect 2318 -270 2334 -236
rect 2386 -270 2402 -236
rect 2436 -270 2452 -236
rect 2504 -270 2520 -236
rect 2554 -270 2570 -236
rect 2622 -270 2638 -236
rect 2672 -270 2688 -236
rect 2740 -270 2756 -236
rect 2790 -270 2806 -236
rect 2858 -270 2874 -236
rect 2908 -270 2924 -236
rect -3081 -339 -3047 -276
rect 3047 -339 3081 -276
rect -3081 -373 -2985 -339
rect 2985 -373 3081 -339
<< viali >>
rect -2967 -177 -2933 249
rect -2849 -177 -2815 249
rect -2731 -177 -2697 249
rect -2613 -177 -2579 249
rect -2495 -177 -2461 249
rect -2377 -177 -2343 249
rect -2259 -177 -2225 249
rect -2141 -177 -2107 249
rect -2023 -177 -1989 249
rect -1905 -177 -1871 249
rect -1787 -177 -1753 249
rect -1669 -177 -1635 249
rect -1551 -177 -1517 249
rect -1433 -177 -1399 249
rect -1315 -177 -1281 249
rect -1197 -177 -1163 249
rect -1079 -177 -1045 249
rect -961 -177 -927 249
rect -843 -177 -809 249
rect -725 -177 -691 249
rect -607 -177 -573 249
rect -489 -177 -455 249
rect -371 -177 -337 249
rect -253 -177 -219 249
rect -135 -177 -101 249
rect -17 -177 17 249
rect 101 -177 135 249
rect 219 -177 253 249
rect 337 -177 371 249
rect 455 -177 489 249
rect 573 -177 607 249
rect 691 -177 725 249
rect 809 -177 843 249
rect 927 -177 961 249
rect 1045 -177 1079 249
rect 1163 -177 1197 249
rect 1281 -177 1315 249
rect 1399 -177 1433 249
rect 1517 -177 1551 249
rect 1635 -177 1669 249
rect 1753 -177 1787 249
rect 1871 -177 1905 249
rect 1989 -177 2023 249
rect 2107 -177 2141 249
rect 2225 -177 2259 249
rect 2343 -177 2377 249
rect 2461 -177 2495 249
rect 2579 -177 2613 249
rect 2697 -177 2731 249
rect 2815 -177 2849 249
rect 2933 -177 2967 249
rect -2908 -270 -2874 -236
rect -2790 -270 -2756 -236
rect -2672 -270 -2638 -236
rect -2554 -270 -2520 -236
rect -2436 -270 -2402 -236
rect -2318 -270 -2284 -236
rect -2200 -270 -2166 -236
rect -2082 -270 -2048 -236
rect -1964 -270 -1930 -236
rect -1846 -270 -1812 -236
rect -1728 -270 -1694 -236
rect -1610 -270 -1576 -236
rect -1492 -270 -1458 -236
rect -1374 -270 -1340 -236
rect -1256 -270 -1222 -236
rect -1138 -270 -1104 -236
rect -1020 -270 -986 -236
rect -902 -270 -868 -236
rect -784 -270 -750 -236
rect -666 -270 -632 -236
rect -548 -270 -514 -236
rect -430 -270 -396 -236
rect -312 -270 -278 -236
rect -194 -270 -160 -236
rect -76 -270 -42 -236
rect 42 -270 76 -236
rect 160 -270 194 -236
rect 278 -270 312 -236
rect 396 -270 430 -236
rect 514 -270 548 -236
rect 632 -270 666 -236
rect 750 -270 784 -236
rect 868 -270 902 -236
rect 986 -270 1020 -236
rect 1104 -270 1138 -236
rect 1222 -270 1256 -236
rect 1340 -270 1374 -236
rect 1458 -270 1492 -236
rect 1576 -270 1610 -236
rect 1694 -270 1728 -236
rect 1812 -270 1846 -236
rect 1930 -270 1964 -236
rect 2048 -270 2082 -236
rect 2166 -270 2200 -236
rect 2284 -270 2318 -236
rect 2402 -270 2436 -236
rect 2520 -270 2554 -236
rect 2638 -270 2672 -236
rect 2756 -270 2790 -236
rect 2874 -270 2908 -236
<< metal1 >>
rect -2973 249 -2927 261
rect -2973 -177 -2967 249
rect -2933 -177 -2927 249
rect -2973 -189 -2927 -177
rect -2855 249 -2809 261
rect -2855 -177 -2849 249
rect -2815 -177 -2809 249
rect -2855 -189 -2809 -177
rect -2737 249 -2691 261
rect -2737 -177 -2731 249
rect -2697 -177 -2691 249
rect -2737 -189 -2691 -177
rect -2619 249 -2573 261
rect -2619 -177 -2613 249
rect -2579 -177 -2573 249
rect -2619 -189 -2573 -177
rect -2501 249 -2455 261
rect -2501 -177 -2495 249
rect -2461 -177 -2455 249
rect -2501 -189 -2455 -177
rect -2383 249 -2337 261
rect -2383 -177 -2377 249
rect -2343 -177 -2337 249
rect -2383 -189 -2337 -177
rect -2265 249 -2219 261
rect -2265 -177 -2259 249
rect -2225 -177 -2219 249
rect -2265 -189 -2219 -177
rect -2147 249 -2101 261
rect -2147 -177 -2141 249
rect -2107 -177 -2101 249
rect -2147 -189 -2101 -177
rect -2029 249 -1983 261
rect -2029 -177 -2023 249
rect -1989 -177 -1983 249
rect -2029 -189 -1983 -177
rect -1911 249 -1865 261
rect -1911 -177 -1905 249
rect -1871 -177 -1865 249
rect -1911 -189 -1865 -177
rect -1793 249 -1747 261
rect -1793 -177 -1787 249
rect -1753 -177 -1747 249
rect -1793 -189 -1747 -177
rect -1675 249 -1629 261
rect -1675 -177 -1669 249
rect -1635 -177 -1629 249
rect -1675 -189 -1629 -177
rect -1557 249 -1511 261
rect -1557 -177 -1551 249
rect -1517 -177 -1511 249
rect -1557 -189 -1511 -177
rect -1439 249 -1393 261
rect -1439 -177 -1433 249
rect -1399 -177 -1393 249
rect -1439 -189 -1393 -177
rect -1321 249 -1275 261
rect -1321 -177 -1315 249
rect -1281 -177 -1275 249
rect -1321 -189 -1275 -177
rect -1203 249 -1157 261
rect -1203 -177 -1197 249
rect -1163 -177 -1157 249
rect -1203 -189 -1157 -177
rect -1085 249 -1039 261
rect -1085 -177 -1079 249
rect -1045 -177 -1039 249
rect -1085 -189 -1039 -177
rect -967 249 -921 261
rect -967 -177 -961 249
rect -927 -177 -921 249
rect -967 -189 -921 -177
rect -849 249 -803 261
rect -849 -177 -843 249
rect -809 -177 -803 249
rect -849 -189 -803 -177
rect -731 249 -685 261
rect -731 -177 -725 249
rect -691 -177 -685 249
rect -731 -189 -685 -177
rect -613 249 -567 261
rect -613 -177 -607 249
rect -573 -177 -567 249
rect -613 -189 -567 -177
rect -495 249 -449 261
rect -495 -177 -489 249
rect -455 -177 -449 249
rect -495 -189 -449 -177
rect -377 249 -331 261
rect -377 -177 -371 249
rect -337 -177 -331 249
rect -377 -189 -331 -177
rect -259 249 -213 261
rect -259 -177 -253 249
rect -219 -177 -213 249
rect -259 -189 -213 -177
rect -141 249 -95 261
rect -141 -177 -135 249
rect -101 -177 -95 249
rect -141 -189 -95 -177
rect -23 249 23 261
rect -23 -177 -17 249
rect 17 -177 23 249
rect -23 -189 23 -177
rect 95 249 141 261
rect 95 -177 101 249
rect 135 -177 141 249
rect 95 -189 141 -177
rect 213 249 259 261
rect 213 -177 219 249
rect 253 -177 259 249
rect 213 -189 259 -177
rect 331 249 377 261
rect 331 -177 337 249
rect 371 -177 377 249
rect 331 -189 377 -177
rect 449 249 495 261
rect 449 -177 455 249
rect 489 -177 495 249
rect 449 -189 495 -177
rect 567 249 613 261
rect 567 -177 573 249
rect 607 -177 613 249
rect 567 -189 613 -177
rect 685 249 731 261
rect 685 -177 691 249
rect 725 -177 731 249
rect 685 -189 731 -177
rect 803 249 849 261
rect 803 -177 809 249
rect 843 -177 849 249
rect 803 -189 849 -177
rect 921 249 967 261
rect 921 -177 927 249
rect 961 -177 967 249
rect 921 -189 967 -177
rect 1039 249 1085 261
rect 1039 -177 1045 249
rect 1079 -177 1085 249
rect 1039 -189 1085 -177
rect 1157 249 1203 261
rect 1157 -177 1163 249
rect 1197 -177 1203 249
rect 1157 -189 1203 -177
rect 1275 249 1321 261
rect 1275 -177 1281 249
rect 1315 -177 1321 249
rect 1275 -189 1321 -177
rect 1393 249 1439 261
rect 1393 -177 1399 249
rect 1433 -177 1439 249
rect 1393 -189 1439 -177
rect 1511 249 1557 261
rect 1511 -177 1517 249
rect 1551 -177 1557 249
rect 1511 -189 1557 -177
rect 1629 249 1675 261
rect 1629 -177 1635 249
rect 1669 -177 1675 249
rect 1629 -189 1675 -177
rect 1747 249 1793 261
rect 1747 -177 1753 249
rect 1787 -177 1793 249
rect 1747 -189 1793 -177
rect 1865 249 1911 261
rect 1865 -177 1871 249
rect 1905 -177 1911 249
rect 1865 -189 1911 -177
rect 1983 249 2029 261
rect 1983 -177 1989 249
rect 2023 -177 2029 249
rect 1983 -189 2029 -177
rect 2101 249 2147 261
rect 2101 -177 2107 249
rect 2141 -177 2147 249
rect 2101 -189 2147 -177
rect 2219 249 2265 261
rect 2219 -177 2225 249
rect 2259 -177 2265 249
rect 2219 -189 2265 -177
rect 2337 249 2383 261
rect 2337 -177 2343 249
rect 2377 -177 2383 249
rect 2337 -189 2383 -177
rect 2455 249 2501 261
rect 2455 -177 2461 249
rect 2495 -177 2501 249
rect 2455 -189 2501 -177
rect 2573 249 2619 261
rect 2573 -177 2579 249
rect 2613 -177 2619 249
rect 2573 -189 2619 -177
rect 2691 249 2737 261
rect 2691 -177 2697 249
rect 2731 -177 2737 249
rect 2691 -189 2737 -177
rect 2809 249 2855 261
rect 2809 -177 2815 249
rect 2849 -177 2855 249
rect 2809 -189 2855 -177
rect 2927 249 2973 261
rect 2927 -177 2933 249
rect 2967 -177 2973 249
rect 2927 -189 2973 -177
rect -2920 -236 -2862 -230
rect -2920 -270 -2908 -236
rect -2874 -270 -2862 -236
rect -2920 -276 -2862 -270
rect -2802 -236 -2744 -230
rect -2802 -270 -2790 -236
rect -2756 -270 -2744 -236
rect -2802 -276 -2744 -270
rect -2684 -236 -2626 -230
rect -2684 -270 -2672 -236
rect -2638 -270 -2626 -236
rect -2684 -276 -2626 -270
rect -2566 -236 -2508 -230
rect -2566 -270 -2554 -236
rect -2520 -270 -2508 -236
rect -2566 -276 -2508 -270
rect -2448 -236 -2390 -230
rect -2448 -270 -2436 -236
rect -2402 -270 -2390 -236
rect -2448 -276 -2390 -270
rect -2330 -236 -2272 -230
rect -2330 -270 -2318 -236
rect -2284 -270 -2272 -236
rect -2330 -276 -2272 -270
rect -2212 -236 -2154 -230
rect -2212 -270 -2200 -236
rect -2166 -270 -2154 -236
rect -2212 -276 -2154 -270
rect -2094 -236 -2036 -230
rect -2094 -270 -2082 -236
rect -2048 -270 -2036 -236
rect -2094 -276 -2036 -270
rect -1976 -236 -1918 -230
rect -1976 -270 -1964 -236
rect -1930 -270 -1918 -236
rect -1976 -276 -1918 -270
rect -1858 -236 -1800 -230
rect -1858 -270 -1846 -236
rect -1812 -270 -1800 -236
rect -1858 -276 -1800 -270
rect -1740 -236 -1682 -230
rect -1740 -270 -1728 -236
rect -1694 -270 -1682 -236
rect -1740 -276 -1682 -270
rect -1622 -236 -1564 -230
rect -1622 -270 -1610 -236
rect -1576 -270 -1564 -236
rect -1622 -276 -1564 -270
rect -1504 -236 -1446 -230
rect -1504 -270 -1492 -236
rect -1458 -270 -1446 -236
rect -1504 -276 -1446 -270
rect -1386 -236 -1328 -230
rect -1386 -270 -1374 -236
rect -1340 -270 -1328 -236
rect -1386 -276 -1328 -270
rect -1268 -236 -1210 -230
rect -1268 -270 -1256 -236
rect -1222 -270 -1210 -236
rect -1268 -276 -1210 -270
rect -1150 -236 -1092 -230
rect -1150 -270 -1138 -236
rect -1104 -270 -1092 -236
rect -1150 -276 -1092 -270
rect -1032 -236 -974 -230
rect -1032 -270 -1020 -236
rect -986 -270 -974 -236
rect -1032 -276 -974 -270
rect -914 -236 -856 -230
rect -914 -270 -902 -236
rect -868 -270 -856 -236
rect -914 -276 -856 -270
rect -796 -236 -738 -230
rect -796 -270 -784 -236
rect -750 -270 -738 -236
rect -796 -276 -738 -270
rect -678 -236 -620 -230
rect -678 -270 -666 -236
rect -632 -270 -620 -236
rect -678 -276 -620 -270
rect -560 -236 -502 -230
rect -560 -270 -548 -236
rect -514 -270 -502 -236
rect -560 -276 -502 -270
rect -442 -236 -384 -230
rect -442 -270 -430 -236
rect -396 -270 -384 -236
rect -442 -276 -384 -270
rect -324 -236 -266 -230
rect -324 -270 -312 -236
rect -278 -270 -266 -236
rect -324 -276 -266 -270
rect -206 -236 -148 -230
rect -206 -270 -194 -236
rect -160 -270 -148 -236
rect -206 -276 -148 -270
rect -88 -236 -30 -230
rect -88 -270 -76 -236
rect -42 -270 -30 -236
rect -88 -276 -30 -270
rect 30 -236 88 -230
rect 30 -270 42 -236
rect 76 -270 88 -236
rect 30 -276 88 -270
rect 148 -236 206 -230
rect 148 -270 160 -236
rect 194 -270 206 -236
rect 148 -276 206 -270
rect 266 -236 324 -230
rect 266 -270 278 -236
rect 312 -270 324 -236
rect 266 -276 324 -270
rect 384 -236 442 -230
rect 384 -270 396 -236
rect 430 -270 442 -236
rect 384 -276 442 -270
rect 502 -236 560 -230
rect 502 -270 514 -236
rect 548 -270 560 -236
rect 502 -276 560 -270
rect 620 -236 678 -230
rect 620 -270 632 -236
rect 666 -270 678 -236
rect 620 -276 678 -270
rect 738 -236 796 -230
rect 738 -270 750 -236
rect 784 -270 796 -236
rect 738 -276 796 -270
rect 856 -236 914 -230
rect 856 -270 868 -236
rect 902 -270 914 -236
rect 856 -276 914 -270
rect 974 -236 1032 -230
rect 974 -270 986 -236
rect 1020 -270 1032 -236
rect 974 -276 1032 -270
rect 1092 -236 1150 -230
rect 1092 -270 1104 -236
rect 1138 -270 1150 -236
rect 1092 -276 1150 -270
rect 1210 -236 1268 -230
rect 1210 -270 1222 -236
rect 1256 -270 1268 -236
rect 1210 -276 1268 -270
rect 1328 -236 1386 -230
rect 1328 -270 1340 -236
rect 1374 -270 1386 -236
rect 1328 -276 1386 -270
rect 1446 -236 1504 -230
rect 1446 -270 1458 -236
rect 1492 -270 1504 -236
rect 1446 -276 1504 -270
rect 1564 -236 1622 -230
rect 1564 -270 1576 -236
rect 1610 -270 1622 -236
rect 1564 -276 1622 -270
rect 1682 -236 1740 -230
rect 1682 -270 1694 -236
rect 1728 -270 1740 -236
rect 1682 -276 1740 -270
rect 1800 -236 1858 -230
rect 1800 -270 1812 -236
rect 1846 -270 1858 -236
rect 1800 -276 1858 -270
rect 1918 -236 1976 -230
rect 1918 -270 1930 -236
rect 1964 -270 1976 -236
rect 1918 -276 1976 -270
rect 2036 -236 2094 -230
rect 2036 -270 2048 -236
rect 2082 -270 2094 -236
rect 2036 -276 2094 -270
rect 2154 -236 2212 -230
rect 2154 -270 2166 -236
rect 2200 -270 2212 -236
rect 2154 -276 2212 -270
rect 2272 -236 2330 -230
rect 2272 -270 2284 -236
rect 2318 -270 2330 -236
rect 2272 -276 2330 -270
rect 2390 -236 2448 -230
rect 2390 -270 2402 -236
rect 2436 -270 2448 -236
rect 2390 -276 2448 -270
rect 2508 -236 2566 -230
rect 2508 -270 2520 -236
rect 2554 -270 2566 -236
rect 2508 -276 2566 -270
rect 2626 -236 2684 -230
rect 2626 -270 2638 -236
rect 2672 -270 2684 -236
rect 2626 -276 2684 -270
rect 2744 -236 2802 -230
rect 2744 -270 2756 -236
rect 2790 -270 2802 -236
rect 2744 -276 2802 -270
rect 2862 -236 2920 -230
rect 2862 -270 2874 -236
rect 2908 -270 2920 -236
rect 2862 -276 2920 -270
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -3064 -356 3064 356
string parameters w 2.25 l 0.3 m 1 nf 50 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
