magic
tech sky130A
magscale 1 2
timestamp 1619566814
<< viali >>
rect -11340 2630 -7240 2670
rect -11340 -980 -11300 2630
rect -7270 2110 -7200 2480
rect -7270 1500 -7200 1870
rect -7270 900 -7200 1270
rect -7270 290 -7200 660
rect -7270 -320 -7200 50
rect -7270 -930 -7200 -560
rect -6930 -6460 -6880 -1350
rect -11330 -6500 -6880 -6460
<< metal1 >>
rect -11490 4140 -11480 4980
rect -11330 4860 -7320 4980
rect -11330 4140 -11240 4860
rect -11180 4140 -11040 4860
rect -10980 4140 -10860 4860
rect -10800 4140 -10660 4860
rect -10600 4140 -10480 4860
rect -10420 4140 -10280 4860
rect -10220 4140 -10080 4860
rect -10020 4140 -9900 4860
rect -9840 4140 -9700 4860
rect -9640 4140 -9520 4860
rect -9460 4140 -9320 4860
rect -9260 4140 -9120 4860
rect -9060 4140 -8940 4860
rect -8880 4140 -8740 4860
rect -8680 4140 -8540 4860
rect -8480 4140 -8360 4860
rect -8300 4140 -8160 4860
rect -8100 4140 -7980 4860
rect -7920 4140 -7780 4860
rect -7720 4140 -7580 4860
rect -7520 4140 -7380 4860
rect -7320 4140 -7310 4860
rect -11490 2630 -11480 2740
rect -11330 2670 -7270 2740
rect -11480 -980 -11340 2630
rect -11300 2624 -7270 2630
rect -11300 -980 -11294 2624
rect -7280 2620 -7270 2624
rect -7090 2620 -7080 2740
rect -6940 2570 -6930 2580
rect -11200 2530 -6930 2570
rect -6940 2520 -6930 2530
rect -6540 2520 -6530 2580
rect -7276 2480 -7194 2492
rect -11150 2400 -11140 2470
rect -11080 2400 -11070 2470
rect -10960 2400 -10950 2460
rect -10890 2400 -10880 2460
rect -10770 2400 -10760 2460
rect -10700 2400 -10690 2460
rect -10580 2410 -10570 2470
rect -10510 2410 -10500 2470
rect -10380 2410 -10370 2470
rect -10310 2410 -10300 2470
rect -10190 2410 -10180 2470
rect -10120 2410 -10110 2470
rect -10000 2410 -9990 2470
rect -9930 2410 -9920 2470
rect -9810 2410 -9800 2470
rect -9740 2410 -9730 2470
rect -9620 2410 -9610 2470
rect -9550 2410 -9540 2470
rect -9420 2410 -9410 2470
rect -9350 2410 -9340 2470
rect -9230 2410 -9220 2470
rect -9160 2410 -9150 2470
rect -9040 2410 -9030 2470
rect -8970 2410 -8960 2470
rect -8850 2410 -8840 2470
rect -8780 2410 -8770 2470
rect -8650 2410 -8640 2470
rect -8580 2410 -8570 2470
rect -8460 2400 -8450 2460
rect -8390 2400 -8380 2460
rect -8270 2400 -8260 2460
rect -8200 2400 -8190 2460
rect -8080 2400 -8070 2460
rect -8010 2400 -8000 2460
rect -7890 2400 -7880 2460
rect -7820 2400 -7810 2460
rect -7690 2400 -7680 2460
rect -7620 2400 -7610 2460
rect -7500 2400 -7490 2460
rect -7430 2400 -7420 2460
rect -11250 2300 -11240 2370
rect -11180 2300 -11170 2370
rect -11060 2310 -11050 2370
rect -10990 2310 -10980 2370
rect -10860 2310 -10850 2370
rect -10790 2310 -10780 2370
rect -10670 2310 -10660 2370
rect -10600 2310 -10590 2370
rect -10480 2310 -10470 2370
rect -10410 2310 -10400 2370
rect -10290 2310 -10280 2370
rect -10220 2310 -10210 2370
rect -10100 2310 -10090 2370
rect -10030 2310 -10020 2370
rect -9900 2310 -9890 2370
rect -9830 2310 -9820 2370
rect -9710 2310 -9700 2370
rect -9640 2310 -9630 2370
rect -9520 2310 -9510 2370
rect -9450 2310 -9440 2370
rect -9330 2310 -9320 2370
rect -9260 2310 -9250 2370
rect -9140 2310 -9130 2370
rect -9070 2310 -9060 2370
rect -8940 2310 -8930 2370
rect -8870 2310 -8860 2370
rect -8750 2310 -8740 2370
rect -8680 2310 -8670 2370
rect -8560 2310 -8550 2370
rect -8490 2310 -8480 2370
rect -8370 2310 -8360 2370
rect -8300 2310 -8290 2370
rect -8170 2310 -8160 2370
rect -8100 2310 -8090 2370
rect -7980 2310 -7970 2370
rect -7910 2310 -7900 2370
rect -7790 2310 -7780 2370
rect -7720 2310 -7710 2370
rect -7600 2310 -7590 2370
rect -7530 2310 -7520 2370
rect -7400 2310 -7390 2370
rect -7330 2310 -7320 2370
rect -11150 2210 -11140 2280
rect -11080 2210 -11070 2280
rect -10960 2210 -10950 2280
rect -10890 2210 -10880 2280
rect -10770 2200 -10760 2270
rect -10700 2200 -10690 2270
rect -10580 2200 -10570 2270
rect -10510 2200 -10500 2270
rect -10380 2200 -10370 2270
rect -10310 2200 -10300 2270
rect -10190 2200 -10180 2270
rect -10120 2200 -10110 2270
rect -10000 2200 -9990 2270
rect -9930 2200 -9920 2270
rect -9810 2200 -9800 2270
rect -9740 2200 -9730 2270
rect -9620 2200 -9610 2270
rect -9550 2200 -9540 2270
rect -9420 2200 -9410 2270
rect -9350 2200 -9340 2270
rect -9230 2200 -9220 2270
rect -9160 2200 -9150 2270
rect -9040 2200 -9030 2270
rect -8970 2200 -8960 2270
rect -8850 2200 -8840 2270
rect -8780 2200 -8770 2270
rect -8650 2200 -8640 2270
rect -8580 2200 -8570 2270
rect -8460 2200 -8450 2270
rect -8390 2200 -8380 2270
rect -8270 2200 -8260 2270
rect -8200 2200 -8190 2270
rect -8080 2200 -8070 2270
rect -8010 2200 -8000 2270
rect -7890 2200 -7880 2270
rect -7820 2200 -7810 2270
rect -7690 2200 -7680 2270
rect -7620 2200 -7610 2270
rect -7500 2200 -7490 2270
rect -7430 2200 -7420 2270
rect -11250 2100 -11240 2170
rect -11180 2100 -11170 2170
rect -11060 2100 -11050 2170
rect -10990 2100 -10980 2170
rect -10860 2100 -10850 2170
rect -10790 2100 -10780 2170
rect -10670 2100 -10660 2170
rect -10600 2100 -10590 2170
rect -10480 2100 -10470 2170
rect -10410 2100 -10400 2170
rect -10290 2100 -10280 2170
rect -10220 2100 -10210 2170
rect -10100 2100 -10090 2170
rect -10030 2100 -10020 2170
rect -9900 2100 -9890 2170
rect -9830 2100 -9820 2170
rect -9710 2100 -9700 2170
rect -9640 2100 -9630 2170
rect -9520 2100 -9510 2170
rect -9450 2100 -9440 2170
rect -9330 2100 -9320 2170
rect -9260 2100 -9250 2170
rect -9140 2100 -9130 2170
rect -9070 2100 -9060 2170
rect -8940 2100 -8930 2170
rect -8870 2100 -8860 2170
rect -8750 2100 -8740 2170
rect -8680 2100 -8670 2170
rect -8560 2100 -8550 2170
rect -8490 2100 -8480 2170
rect -8370 2100 -8360 2170
rect -8300 2100 -8290 2170
rect -8170 2100 -8160 2170
rect -8100 2100 -8090 2170
rect -7980 2100 -7970 2170
rect -7910 2100 -7900 2170
rect -7790 2100 -7780 2170
rect -7720 2100 -7710 2170
rect -7600 2100 -7590 2170
rect -7530 2100 -7520 2170
rect -7400 2100 -7390 2170
rect -7330 2100 -7320 2170
rect -7280 2110 -7270 2480
rect -7200 2110 -7190 2480
rect -7276 2098 -7194 2110
rect -11200 1910 -6930 2060
rect -6540 1910 -6530 2060
rect -7276 1870 -7194 1882
rect -11150 1790 -11140 1850
rect -11080 1790 -11070 1850
rect -10960 1790 -10950 1850
rect -10890 1790 -10880 1850
rect -10770 1790 -10760 1850
rect -10700 1790 -10690 1850
rect -10580 1790 -10570 1850
rect -10510 1790 -10500 1850
rect -10380 1790 -10370 1850
rect -10310 1790 -10300 1850
rect -10190 1790 -10180 1850
rect -10120 1790 -10110 1850
rect -10000 1790 -9990 1850
rect -9930 1790 -9920 1850
rect -9810 1790 -9800 1850
rect -9740 1790 -9730 1850
rect -9620 1790 -9610 1850
rect -9550 1790 -9540 1850
rect -9420 1790 -9410 1850
rect -9350 1790 -9340 1850
rect -9230 1790 -9220 1850
rect -9160 1790 -9150 1850
rect -9040 1790 -9030 1850
rect -8970 1790 -8960 1850
rect -8850 1790 -8840 1850
rect -8780 1790 -8770 1850
rect -8650 1790 -8640 1850
rect -8580 1790 -8570 1850
rect -8460 1790 -8450 1850
rect -8390 1790 -8380 1850
rect -8270 1790 -8260 1850
rect -8200 1790 -8190 1850
rect -8080 1790 -8070 1850
rect -8010 1790 -8000 1850
rect -7890 1790 -7880 1850
rect -7820 1790 -7810 1850
rect -7690 1790 -7680 1850
rect -7620 1790 -7610 1850
rect -7500 1790 -7490 1850
rect -7430 1790 -7420 1850
rect -11250 1650 -11240 1710
rect -11180 1650 -11170 1710
rect -11060 1670 -11050 1730
rect -10990 1670 -10980 1730
rect -10860 1670 -10850 1730
rect -10790 1670 -10780 1730
rect -10670 1670 -10660 1730
rect -10600 1670 -10590 1730
rect -10480 1670 -10470 1730
rect -10410 1670 -10400 1730
rect -10290 1670 -10280 1730
rect -10220 1670 -10210 1730
rect -10100 1670 -10090 1730
rect -10030 1670 -10020 1730
rect -9900 1670 -9890 1730
rect -9830 1670 -9820 1730
rect -9710 1670 -9700 1730
rect -9640 1670 -9630 1730
rect -9520 1670 -9510 1730
rect -9450 1670 -9440 1730
rect -9330 1670 -9320 1730
rect -9260 1670 -9250 1730
rect -9140 1670 -9130 1730
rect -9070 1670 -9060 1730
rect -8940 1670 -8930 1730
rect -8870 1670 -8860 1730
rect -8750 1670 -8740 1730
rect -8680 1670 -8670 1730
rect -8560 1670 -8550 1730
rect -8490 1670 -8480 1730
rect -8370 1670 -8360 1730
rect -8300 1670 -8290 1730
rect -8170 1670 -8160 1730
rect -8100 1670 -8090 1730
rect -7980 1670 -7970 1730
rect -7910 1670 -7900 1730
rect -7790 1670 -7780 1730
rect -7720 1670 -7710 1730
rect -7600 1670 -7590 1730
rect -7530 1670 -7520 1730
rect -7400 1670 -7390 1730
rect -7330 1670 -7320 1730
rect -11150 1570 -11140 1630
rect -11080 1570 -11070 1630
rect -10960 1580 -10950 1640
rect -10890 1580 -10880 1640
rect -10770 1580 -10760 1640
rect -10700 1580 -10690 1640
rect -10580 1580 -10570 1640
rect -10510 1580 -10500 1640
rect -10380 1580 -10370 1640
rect -10310 1580 -10300 1640
rect -10190 1580 -10180 1640
rect -10120 1580 -10110 1640
rect -10000 1580 -9990 1640
rect -9930 1580 -9920 1640
rect -9810 1580 -9800 1640
rect -9740 1580 -9730 1640
rect -9620 1580 -9610 1640
rect -9550 1580 -9540 1640
rect -9420 1580 -9410 1640
rect -9350 1580 -9340 1640
rect -9230 1580 -9220 1640
rect -9160 1580 -9150 1640
rect -9040 1580 -9030 1640
rect -8970 1580 -8960 1640
rect -8850 1580 -8840 1640
rect -8780 1580 -8770 1640
rect -8650 1580 -8640 1640
rect -8580 1580 -8570 1640
rect -8460 1580 -8450 1640
rect -8390 1580 -8380 1640
rect -8270 1580 -8260 1640
rect -8200 1580 -8190 1640
rect -8080 1580 -8070 1640
rect -8010 1580 -8000 1640
rect -7890 1580 -7880 1640
rect -7820 1580 -7810 1640
rect -7690 1580 -7680 1640
rect -7620 1580 -7610 1640
rect -7500 1580 -7490 1640
rect -7430 1580 -7420 1640
rect -11250 1490 -11240 1550
rect -11180 1490 -11170 1550
rect -11050 1490 -11040 1550
rect -10980 1490 -10970 1550
rect -10860 1490 -10850 1550
rect -10790 1490 -10780 1550
rect -10670 1490 -10660 1550
rect -10600 1490 -10590 1550
rect -10480 1490 -10470 1550
rect -10410 1490 -10400 1550
rect -10290 1490 -10280 1550
rect -10220 1490 -10210 1550
rect -10100 1490 -10090 1550
rect -10030 1490 -10020 1550
rect -9900 1490 -9890 1550
rect -9830 1490 -9820 1550
rect -9710 1490 -9700 1550
rect -9640 1490 -9630 1550
rect -9520 1490 -9510 1550
rect -9450 1490 -9440 1550
rect -9330 1490 -9320 1550
rect -9260 1490 -9250 1550
rect -9140 1490 -9130 1550
rect -9070 1490 -9060 1550
rect -8940 1490 -8930 1550
rect -8870 1490 -8860 1550
rect -8750 1490 -8740 1550
rect -8680 1490 -8670 1550
rect -8560 1490 -8550 1550
rect -8490 1490 -8480 1550
rect -8370 1490 -8360 1550
rect -8300 1490 -8290 1550
rect -8170 1490 -8160 1550
rect -8100 1490 -8090 1550
rect -7980 1490 -7970 1550
rect -7910 1490 -7900 1550
rect -7790 1490 -7780 1550
rect -7720 1490 -7710 1550
rect -7600 1490 -7590 1550
rect -7530 1490 -7520 1550
rect -7400 1490 -7390 1550
rect -7330 1490 -7320 1550
rect -7280 1500 -7270 1870
rect -7200 1500 -7190 1870
rect -7276 1488 -7194 1500
rect -11200 1310 -6930 1460
rect -6540 1310 -6530 1460
rect -7276 1270 -7194 1282
rect -11150 1160 -11140 1220
rect -11080 1160 -11070 1220
rect -10960 1160 -10950 1220
rect -10890 1160 -10880 1220
rect -10770 1160 -10760 1220
rect -10700 1160 -10690 1220
rect -10580 1160 -10570 1220
rect -10510 1160 -10500 1220
rect -10380 1160 -10370 1220
rect -10310 1160 -10300 1220
rect -10190 1160 -10180 1220
rect -10120 1160 -10110 1220
rect -10000 1160 -9990 1220
rect -9930 1160 -9920 1220
rect -9810 1160 -9800 1220
rect -9740 1160 -9730 1220
rect -9620 1160 -9610 1220
rect -9550 1160 -9540 1220
rect -9420 1160 -9410 1220
rect -9350 1160 -9340 1220
rect -9230 1160 -9220 1220
rect -9160 1160 -9150 1220
rect -9040 1160 -9030 1220
rect -8970 1160 -8960 1220
rect -8850 1160 -8840 1220
rect -8780 1160 -8770 1220
rect -8650 1160 -8640 1220
rect -8580 1160 -8570 1220
rect -8460 1160 -8450 1220
rect -8390 1160 -8380 1220
rect -8270 1160 -8260 1220
rect -8200 1160 -8190 1220
rect -8080 1160 -8070 1220
rect -8010 1160 -8000 1220
rect -7890 1160 -7880 1220
rect -7820 1160 -7810 1220
rect -7690 1160 -7680 1220
rect -7620 1160 -7610 1220
rect -7500 1160 -7490 1220
rect -7430 1160 -7420 1220
rect -11250 1070 -11240 1130
rect -11180 1070 -11170 1130
rect -11060 1070 -11050 1130
rect -10990 1070 -10980 1130
rect -10860 1070 -10850 1130
rect -10790 1070 -10780 1130
rect -10670 1070 -10660 1130
rect -10600 1070 -10590 1130
rect -10480 1070 -10470 1130
rect -10410 1070 -10400 1130
rect -10290 1070 -10280 1130
rect -10220 1070 -10210 1130
rect -10100 1070 -10090 1130
rect -10030 1070 -10020 1130
rect -9900 1070 -9890 1130
rect -9830 1070 -9820 1130
rect -9710 1070 -9700 1130
rect -9640 1070 -9630 1130
rect -9520 1070 -9510 1130
rect -9450 1070 -9440 1130
rect -9330 1070 -9320 1130
rect -9260 1070 -9250 1130
rect -9140 1070 -9130 1130
rect -9070 1070 -9060 1130
rect -8940 1070 -8930 1130
rect -8870 1070 -8860 1130
rect -8750 1070 -8740 1130
rect -8680 1070 -8670 1130
rect -8560 1070 -8550 1130
rect -8490 1070 -8480 1130
rect -8370 1070 -8360 1130
rect -8300 1070 -8290 1130
rect -8170 1070 -8160 1130
rect -8100 1070 -8090 1130
rect -7980 1070 -7970 1130
rect -7910 1070 -7900 1130
rect -7790 1070 -7780 1130
rect -7720 1070 -7710 1130
rect -7600 1070 -7590 1130
rect -7530 1070 -7520 1130
rect -7400 1070 -7390 1130
rect -7330 1070 -7320 1130
rect -11150 970 -11140 1030
rect -11080 970 -11070 1030
rect -10960 970 -10950 1030
rect -10890 970 -10880 1030
rect -10770 970 -10760 1030
rect -10700 970 -10690 1030
rect -10580 970 -10570 1030
rect -10510 970 -10500 1030
rect -10380 970 -10370 1030
rect -10310 970 -10300 1030
rect -10190 970 -10180 1030
rect -10120 970 -10110 1030
rect -10000 970 -9990 1030
rect -9930 970 -9920 1030
rect -9810 970 -9800 1030
rect -9740 970 -9730 1030
rect -9620 970 -9610 1030
rect -9550 970 -9540 1030
rect -9420 970 -9410 1030
rect -9350 970 -9340 1030
rect -9230 970 -9220 1030
rect -9160 970 -9150 1030
rect -9040 970 -9030 1030
rect -8970 970 -8960 1030
rect -8850 970 -8840 1030
rect -8780 970 -8770 1030
rect -8650 970 -8640 1030
rect -8580 970 -8570 1030
rect -8460 980 -8450 1040
rect -8390 980 -8380 1040
rect -8270 980 -8260 1040
rect -8200 980 -8190 1040
rect -8080 980 -8070 1040
rect -8010 980 -8000 1040
rect -7890 980 -7880 1040
rect -7820 980 -7810 1040
rect -7690 980 -7680 1040
rect -7620 980 -7610 1040
rect -7500 980 -7490 1040
rect -7430 980 -7420 1040
rect -11250 880 -11240 940
rect -11180 880 -11170 940
rect -11060 880 -11050 940
rect -10990 880 -10980 940
rect -10860 880 -10850 940
rect -10790 880 -10780 940
rect -10670 880 -10660 940
rect -10600 880 -10590 940
rect -10480 880 -10470 940
rect -10410 880 -10400 940
rect -10290 880 -10280 940
rect -10220 880 -10210 940
rect -10100 880 -10090 940
rect -10030 880 -10020 940
rect -9900 880 -9890 940
rect -9830 880 -9820 940
rect -9710 880 -9700 940
rect -9640 880 -9630 940
rect -9520 880 -9510 940
rect -9450 880 -9440 940
rect -9330 880 -9320 940
rect -9260 880 -9250 940
rect -9140 880 -9130 940
rect -9070 880 -9060 940
rect -8940 880 -8930 940
rect -8870 880 -8860 940
rect -8750 880 -8740 940
rect -8680 880 -8670 940
rect -8560 880 -8550 940
rect -8490 880 -8480 940
rect -8370 890 -8360 950
rect -8300 890 -8290 950
rect -8170 890 -8160 950
rect -8100 890 -8090 950
rect -7980 890 -7970 950
rect -7910 890 -7900 950
rect -7790 890 -7780 950
rect -7720 890 -7710 950
rect -7600 890 -7590 950
rect -7530 890 -7520 950
rect -7400 890 -7390 950
rect -7330 890 -7320 950
rect -7280 900 -7270 1270
rect -7200 900 -7190 1270
rect -7276 888 -7194 900
rect -11200 700 -6930 850
rect -6540 700 -6530 850
rect -7276 660 -7194 672
rect -11150 560 -11140 620
rect -11080 560 -11070 620
rect -10960 560 -10950 620
rect -10890 560 -10880 620
rect -10770 560 -10760 620
rect -10700 560 -10690 620
rect -10580 560 -10570 620
rect -10510 560 -10500 620
rect -10380 560 -10370 620
rect -10310 560 -10300 620
rect -10190 560 -10180 620
rect -10120 560 -10110 620
rect -10000 560 -9990 620
rect -9930 560 -9920 620
rect -9810 560 -9800 620
rect -9740 560 -9730 620
rect -9610 560 -9600 620
rect -9540 560 -9530 620
rect -9420 560 -9410 620
rect -9350 560 -9340 620
rect -9230 560 -9220 620
rect -9160 560 -9150 620
rect -9040 560 -9030 620
rect -8970 560 -8960 620
rect -8850 560 -8840 620
rect -8780 560 -8770 620
rect -8650 560 -8640 620
rect -8580 560 -8570 620
rect -8460 560 -8450 620
rect -8390 560 -8380 620
rect -8270 560 -8260 620
rect -8200 560 -8190 620
rect -8080 560 -8070 620
rect -8010 560 -8000 620
rect -7890 560 -7880 620
rect -7820 560 -7810 620
rect -7690 560 -7680 620
rect -7620 560 -7610 620
rect -7500 560 -7490 620
rect -7430 560 -7420 620
rect -11250 460 -11240 520
rect -11180 460 -11170 520
rect -11060 460 -11050 520
rect -10990 460 -10980 520
rect -10860 460 -10850 520
rect -10790 460 -10780 520
rect -10670 460 -10660 520
rect -10600 460 -10590 520
rect -10480 460 -10470 520
rect -10410 460 -10400 520
rect -10290 460 -10280 520
rect -10220 460 -10210 520
rect -10100 460 -10090 520
rect -10030 460 -10020 520
rect -9900 460 -9890 520
rect -9830 460 -9820 520
rect -9710 460 -9700 520
rect -9640 460 -9630 520
rect -9520 460 -9510 520
rect -9450 460 -9440 520
rect -9330 460 -9320 520
rect -9260 460 -9250 520
rect -9140 460 -9130 520
rect -9070 460 -9060 520
rect -8940 460 -8930 520
rect -8870 460 -8860 520
rect -8750 460 -8740 520
rect -8680 460 -8670 520
rect -8560 460 -8550 520
rect -8490 460 -8480 520
rect -8370 460 -8360 520
rect -8300 460 -8290 520
rect -8170 460 -8160 520
rect -8100 460 -8090 520
rect -7980 460 -7970 520
rect -7910 460 -7900 520
rect -7790 460 -7780 520
rect -7720 460 -7710 520
rect -7600 460 -7590 520
rect -7530 460 -7520 520
rect -7400 460 -7390 520
rect -7330 460 -7320 520
rect -11150 360 -11140 420
rect -11080 360 -11070 420
rect -10960 360 -10950 420
rect -10890 360 -10880 420
rect -10770 360 -10760 420
rect -10700 360 -10690 420
rect -10580 360 -10570 420
rect -10510 360 -10500 420
rect -10380 360 -10370 420
rect -10310 360 -10300 420
rect -10190 360 -10180 420
rect -10120 360 -10110 420
rect -10000 360 -9990 420
rect -9930 360 -9920 420
rect -9810 360 -9800 420
rect -9740 360 -9730 420
rect -9620 360 -9610 420
rect -9550 360 -9540 420
rect -9420 360 -9410 420
rect -9350 360 -9340 420
rect -9230 360 -9220 420
rect -9160 360 -9150 420
rect -9040 360 -9030 420
rect -8970 360 -8960 420
rect -8850 360 -8840 420
rect -8780 360 -8770 420
rect -8650 360 -8640 420
rect -8580 360 -8570 420
rect -8460 360 -8450 420
rect -8390 360 -8380 420
rect -8270 360 -8260 420
rect -8200 360 -8190 420
rect -8080 360 -8070 420
rect -8010 360 -8000 420
rect -7890 360 -7880 420
rect -7820 360 -7810 420
rect -7690 360 -7680 420
rect -7620 360 -7610 420
rect -7500 360 -7490 420
rect -7430 360 -7420 420
rect -11250 270 -11240 330
rect -11180 270 -11170 330
rect -11060 270 -11050 330
rect -10990 270 -10980 330
rect -10860 270 -10850 330
rect -10790 270 -10780 330
rect -10670 270 -10660 330
rect -10600 270 -10590 330
rect -10480 270 -10470 330
rect -10410 270 -10400 330
rect -10290 270 -10280 330
rect -10220 270 -10210 330
rect -10100 270 -10090 330
rect -10030 270 -10020 330
rect -9900 270 -9890 330
rect -9830 270 -9820 330
rect -9710 270 -9700 330
rect -9640 270 -9630 330
rect -9520 270 -9510 330
rect -9450 270 -9440 330
rect -9330 270 -9320 330
rect -9260 270 -9250 330
rect -9140 270 -9130 330
rect -9070 270 -9060 330
rect -8940 270 -8930 330
rect -8870 270 -8860 330
rect -8750 270 -8740 330
rect -8680 270 -8670 330
rect -8560 270 -8550 330
rect -8490 270 -8480 330
rect -8370 270 -8360 330
rect -8300 270 -8290 330
rect -8170 270 -8160 330
rect -8100 270 -8090 330
rect -7980 270 -7970 330
rect -7910 270 -7900 330
rect -7790 270 -7780 330
rect -7720 270 -7710 330
rect -7600 270 -7590 330
rect -7530 270 -7520 330
rect -7400 270 -7390 330
rect -7330 270 -7320 330
rect -7280 290 -7270 660
rect -7200 290 -7190 660
rect -7276 278 -7194 290
rect -11200 90 -6930 240
rect -6540 90 -6530 240
rect -7276 50 -7194 62
rect -11150 -40 -11140 20
rect -11080 -40 -11070 20
rect -10960 -40 -10950 20
rect -10890 -40 -10880 20
rect -10770 -40 -10760 20
rect -10700 -40 -10690 20
rect -10580 -40 -10570 20
rect -10510 -40 -10500 20
rect -10380 -40 -10370 20
rect -10310 -40 -10300 20
rect -10190 -40 -10180 20
rect -10120 -40 -10110 20
rect -10000 -40 -9990 20
rect -9930 -40 -9920 20
rect -9810 -40 -9800 20
rect -9740 -40 -9730 20
rect -9620 -40 -9610 20
rect -9550 -40 -9540 20
rect -9420 -40 -9410 20
rect -9350 -40 -9340 20
rect -9230 -40 -9220 20
rect -9160 -40 -9150 20
rect -9040 -50 -9030 10
rect -8970 -50 -8960 10
rect -8850 -50 -8840 10
rect -8780 -50 -8770 10
rect -8650 -50 -8640 10
rect -8580 -50 -8570 10
rect -8460 -50 -8450 10
rect -8390 -50 -8380 10
rect -8270 -50 -8260 10
rect -8200 -50 -8190 10
rect -8080 -50 -8070 10
rect -8010 -50 -8000 10
rect -7890 -50 -7880 10
rect -7820 -50 -7810 10
rect -7690 -50 -7680 10
rect -7620 -50 -7610 10
rect -7500 -50 -7490 10
rect -7430 -50 -7420 10
rect -11250 -140 -11240 -80
rect -11180 -140 -11170 -80
rect -11060 -140 -11050 -80
rect -10990 -140 -10980 -80
rect -10860 -130 -10850 -70
rect -10790 -130 -10780 -70
rect -10670 -130 -10660 -70
rect -10600 -130 -10590 -70
rect -10480 -130 -10470 -70
rect -10410 -130 -10400 -70
rect -10290 -130 -10280 -70
rect -10220 -130 -10210 -70
rect -10100 -130 -10090 -70
rect -10030 -130 -10020 -70
rect -9900 -130 -9890 -70
rect -9830 -130 -9820 -70
rect -9710 -130 -9700 -70
rect -9640 -130 -9630 -70
rect -9520 -130 -9510 -70
rect -9450 -130 -9440 -70
rect -9330 -130 -9320 -70
rect -9260 -130 -9250 -70
rect -9140 -130 -9130 -70
rect -9070 -130 -9060 -70
rect -8940 -140 -8930 -80
rect -8870 -140 -8860 -80
rect -8750 -140 -8740 -80
rect -8680 -140 -8670 -80
rect -8560 -140 -8550 -80
rect -8490 -140 -8480 -80
rect -8370 -140 -8360 -80
rect -8300 -140 -8290 -80
rect -8170 -140 -8160 -80
rect -8100 -140 -8090 -80
rect -7980 -140 -7970 -80
rect -7910 -140 -7900 -80
rect -7790 -140 -7780 -80
rect -7720 -140 -7710 -80
rect -7600 -140 -7590 -80
rect -7530 -140 -7520 -80
rect -7400 -140 -7390 -80
rect -7330 -140 -7320 -80
rect -11150 -230 -11140 -170
rect -11080 -230 -11070 -170
rect -10960 -230 -10950 -170
rect -10890 -230 -10880 -170
rect -10770 -230 -10760 -170
rect -10700 -230 -10690 -170
rect -10580 -230 -10570 -170
rect -10510 -230 -10500 -170
rect -10380 -230 -10370 -170
rect -10310 -230 -10300 -170
rect -10190 -230 -10180 -170
rect -10120 -230 -10110 -170
rect -10000 -230 -9990 -170
rect -9930 -230 -9920 -170
rect -9810 -230 -9800 -170
rect -9740 -230 -9730 -170
rect -9620 -230 -9610 -170
rect -9550 -230 -9540 -170
rect -9420 -230 -9410 -170
rect -9350 -230 -9340 -170
rect -9230 -230 -9220 -170
rect -9160 -230 -9150 -170
rect -9040 -230 -9030 -170
rect -8970 -230 -8960 -170
rect -8850 -230 -8840 -170
rect -8780 -230 -8770 -170
rect -8650 -230 -8640 -170
rect -8580 -230 -8570 -170
rect -8460 -230 -8450 -170
rect -8390 -230 -8380 -170
rect -8270 -230 -8260 -170
rect -8200 -230 -8190 -170
rect -8080 -230 -8070 -170
rect -8010 -230 -8000 -170
rect -7890 -230 -7880 -170
rect -7820 -230 -7810 -170
rect -7690 -230 -7680 -170
rect -7620 -230 -7610 -170
rect -7500 -230 -7490 -170
rect -7430 -230 -7420 -170
rect -11250 -320 -11240 -260
rect -11180 -320 -11170 -260
rect -11060 -320 -11050 -260
rect -10990 -320 -10980 -260
rect -10860 -320 -10850 -260
rect -10790 -320 -10780 -260
rect -10670 -320 -10660 -260
rect -10600 -320 -10590 -260
rect -10480 -320 -10470 -260
rect -10410 -320 -10400 -260
rect -10290 -320 -10280 -260
rect -10220 -320 -10210 -260
rect -10100 -320 -10090 -260
rect -10030 -320 -10020 -260
rect -9900 -320 -9890 -260
rect -9830 -320 -9820 -260
rect -9710 -320 -9700 -260
rect -9640 -320 -9630 -260
rect -9520 -320 -9510 -260
rect -9450 -320 -9440 -260
rect -9330 -320 -9320 -260
rect -9260 -320 -9250 -260
rect -9140 -320 -9130 -260
rect -9070 -320 -9060 -260
rect -8940 -320 -8930 -260
rect -8870 -320 -8860 -260
rect -8750 -320 -8740 -260
rect -8680 -320 -8670 -260
rect -8560 -320 -8550 -260
rect -8490 -320 -8480 -260
rect -8370 -320 -8360 -260
rect -8300 -320 -8290 -260
rect -8170 -320 -8160 -260
rect -8100 -320 -8090 -260
rect -7980 -320 -7970 -260
rect -7910 -320 -7900 -260
rect -7790 -320 -7780 -260
rect -7720 -320 -7710 -260
rect -7600 -320 -7590 -260
rect -7530 -320 -7520 -260
rect -7400 -320 -7390 -260
rect -7330 -320 -7320 -260
rect -7280 -320 -7270 50
rect -7200 -320 -7190 50
rect -7276 -332 -7194 -320
rect -11200 -520 -6930 -370
rect -6540 -520 -6530 -370
rect -7276 -560 -7194 -548
rect -11150 -640 -11140 -580
rect -11080 -640 -11070 -580
rect -10960 -640 -10950 -580
rect -10890 -640 -10880 -580
rect -10770 -640 -10760 -580
rect -10700 -640 -10690 -580
rect -10580 -640 -10570 -580
rect -10510 -640 -10500 -580
rect -10380 -640 -10370 -580
rect -10310 -640 -10300 -580
rect -10190 -640 -10180 -580
rect -10120 -640 -10110 -580
rect -10000 -640 -9990 -580
rect -9930 -640 -9920 -580
rect -9810 -640 -9800 -580
rect -9740 -640 -9730 -580
rect -9620 -640 -9610 -580
rect -9550 -640 -9540 -580
rect -9420 -640 -9410 -580
rect -9350 -640 -9340 -580
rect -9230 -640 -9220 -580
rect -9160 -640 -9150 -580
rect -9040 -640 -9030 -580
rect -8970 -640 -8960 -580
rect -8850 -640 -8840 -580
rect -8780 -640 -8770 -580
rect -8650 -640 -8640 -580
rect -8580 -640 -8570 -580
rect -8460 -640 -8450 -580
rect -8390 -640 -8380 -580
rect -8270 -640 -8260 -580
rect -8200 -640 -8190 -580
rect -8080 -640 -8070 -580
rect -8010 -640 -8000 -580
rect -7890 -640 -7880 -580
rect -7820 -640 -7810 -580
rect -7690 -640 -7680 -580
rect -7620 -640 -7610 -580
rect -7500 -640 -7490 -580
rect -7430 -640 -7420 -580
rect -11250 -740 -11240 -680
rect -11180 -740 -11170 -680
rect -11060 -740 -11050 -680
rect -10990 -740 -10980 -680
rect -10860 -740 -10850 -680
rect -10790 -740 -10780 -680
rect -10670 -740 -10660 -680
rect -10600 -740 -10590 -680
rect -10480 -740 -10470 -680
rect -10410 -740 -10400 -680
rect -10290 -740 -10280 -680
rect -10220 -740 -10210 -680
rect -10100 -740 -10090 -680
rect -10030 -740 -10020 -680
rect -9900 -740 -9890 -680
rect -9830 -740 -9820 -680
rect -9710 -740 -9700 -680
rect -9640 -740 -9630 -680
rect -9520 -740 -9510 -680
rect -9450 -740 -9440 -680
rect -9330 -740 -9320 -680
rect -9260 -740 -9250 -680
rect -9140 -740 -9130 -680
rect -9070 -740 -9060 -680
rect -8940 -740 -8930 -680
rect -8870 -740 -8860 -680
rect -8750 -740 -8740 -680
rect -8680 -740 -8670 -680
rect -8560 -740 -8550 -680
rect -8490 -740 -8480 -680
rect -8370 -740 -8360 -680
rect -8300 -740 -8290 -680
rect -8170 -740 -8160 -680
rect -8100 -740 -8090 -680
rect -7980 -740 -7970 -680
rect -7910 -740 -7900 -680
rect -7790 -740 -7780 -680
rect -7720 -740 -7710 -680
rect -7600 -740 -7590 -680
rect -7530 -740 -7520 -680
rect -7400 -740 -7390 -680
rect -7330 -740 -7320 -680
rect -11150 -830 -11140 -770
rect -11080 -830 -11070 -770
rect -10960 -830 -10950 -770
rect -10890 -830 -10880 -770
rect -10770 -830 -10760 -770
rect -10700 -830 -10690 -770
rect -10580 -830 -10570 -770
rect -10510 -830 -10500 -770
rect -10380 -830 -10370 -770
rect -10310 -830 -10300 -770
rect -10190 -830 -10180 -770
rect -10120 -830 -10110 -770
rect -10000 -830 -9990 -770
rect -9930 -830 -9920 -770
rect -9810 -830 -9800 -770
rect -9740 -830 -9730 -770
rect -9620 -830 -9610 -770
rect -9550 -830 -9540 -770
rect -9420 -830 -9410 -770
rect -9350 -830 -9340 -770
rect -9230 -830 -9220 -770
rect -9160 -830 -9150 -770
rect -9040 -830 -9030 -770
rect -8970 -830 -8960 -770
rect -8850 -830 -8840 -770
rect -8780 -830 -8770 -770
rect -8650 -830 -8640 -770
rect -8580 -830 -8570 -770
rect -8460 -830 -8450 -770
rect -8390 -830 -8380 -770
rect -8270 -830 -8260 -770
rect -8200 -830 -8190 -770
rect -8080 -830 -8070 -770
rect -8010 -830 -8000 -770
rect -7890 -830 -7880 -770
rect -7820 -830 -7810 -770
rect -7690 -830 -7680 -770
rect -7620 -830 -7610 -770
rect -7500 -830 -7490 -770
rect -7430 -830 -7420 -770
rect -11250 -920 -11240 -860
rect -11180 -920 -11170 -860
rect -11060 -920 -11050 -860
rect -10990 -920 -10980 -860
rect -10860 -920 -10850 -860
rect -10790 -920 -10780 -860
rect -10670 -920 -10660 -860
rect -10600 -920 -10590 -860
rect -10480 -920 -10470 -860
rect -10410 -920 -10400 -860
rect -10290 -920 -10280 -860
rect -10220 -920 -10210 -860
rect -10100 -920 -10090 -860
rect -10030 -920 -10020 -860
rect -9900 -920 -9890 -860
rect -9830 -920 -9820 -860
rect -9710 -920 -9700 -860
rect -9640 -920 -9630 -860
rect -9520 -920 -9510 -860
rect -9450 -920 -9440 -860
rect -9330 -920 -9320 -860
rect -9260 -920 -9250 -860
rect -9140 -920 -9130 -860
rect -9070 -920 -9060 -860
rect -8940 -920 -8930 -860
rect -8870 -920 -8860 -860
rect -8750 -920 -8740 -860
rect -8680 -920 -8670 -860
rect -8560 -920 -8550 -860
rect -8490 -920 -8480 -860
rect -8370 -920 -8360 -860
rect -8300 -920 -8290 -860
rect -8170 -920 -8160 -860
rect -8100 -920 -8090 -860
rect -7980 -920 -7970 -860
rect -7910 -920 -7900 -860
rect -7790 -920 -7780 -860
rect -7720 -920 -7710 -860
rect -7600 -920 -7590 -860
rect -7530 -920 -7520 -860
rect -7400 -920 -7390 -860
rect -7330 -920 -7320 -860
rect -7280 -930 -7270 -560
rect -7200 -930 -7190 -560
rect -7276 -942 -7194 -930
rect -6940 -980 -6930 -960
rect -11346 -992 -11294 -980
rect -11200 -1020 -6930 -980
rect -6540 -1020 -6530 -960
rect -11340 -1250 -11240 -1050
rect -11180 -1250 -10400 -1050
rect -10340 -1250 -9560 -1050
rect -9500 -1250 -8720 -1050
rect -8660 -1250 -7900 -1050
rect -7840 -1250 -7060 -1050
rect -7000 -1250 -6930 -1050
rect -6540 -1250 -6530 -1050
rect -11180 -1290 -7040 -1280
rect -11480 -1320 -7040 -1290
rect -6936 -1350 -6874 -1338
rect -11250 -1660 -11240 -1360
rect -11180 -1660 -11170 -1360
rect -10830 -1660 -10820 -1360
rect -10760 -1660 -10750 -1360
rect -10410 -1660 -10400 -1360
rect -10340 -1660 -10330 -1360
rect -9990 -1660 -9980 -1360
rect -9920 -1660 -9910 -1360
rect -9570 -1660 -9560 -1360
rect -9500 -1660 -9490 -1360
rect -9150 -1660 -9140 -1360
rect -9080 -1660 -9070 -1360
rect -8730 -1660 -8720 -1360
rect -8660 -1660 -8650 -1360
rect -8310 -1660 -8300 -1360
rect -8240 -1660 -8230 -1360
rect -7910 -1660 -7900 -1360
rect -7840 -1660 -7830 -1360
rect -7490 -1660 -7480 -1360
rect -7420 -1660 -7410 -1360
rect -7070 -1660 -7060 -1360
rect -7000 -1660 -6990 -1360
rect -11490 -1840 -11480 -1700
rect -11290 -1840 -7050 -1700
rect -11250 -2180 -11240 -1880
rect -11180 -2180 -11170 -1880
rect -10830 -2180 -10820 -1880
rect -10760 -2180 -10750 -1880
rect -10410 -2180 -10400 -1880
rect -10340 -2180 -10330 -1880
rect -9990 -2180 -9980 -1880
rect -9920 -2180 -9910 -1880
rect -9570 -2180 -9560 -1880
rect -9500 -2180 -9490 -1880
rect -9150 -2180 -9140 -1880
rect -9080 -2180 -9070 -1880
rect -8730 -2180 -8720 -1880
rect -8660 -2180 -8650 -1880
rect -8310 -2180 -8300 -1880
rect -8240 -2180 -8230 -1880
rect -7910 -2180 -7900 -1880
rect -7840 -2180 -7830 -1880
rect -7490 -2180 -7480 -1880
rect -7420 -2180 -7410 -1880
rect -7070 -2180 -7060 -1880
rect -7000 -2180 -6990 -1880
rect -11490 -2360 -11480 -2220
rect -11290 -2360 -7050 -2220
rect -11250 -2700 -11240 -2400
rect -11180 -2700 -11170 -2400
rect -10830 -2700 -10820 -2400
rect -10760 -2700 -10750 -2400
rect -10410 -2700 -10400 -2400
rect -10340 -2700 -10330 -2400
rect -9990 -2700 -9980 -2400
rect -9920 -2700 -9910 -2400
rect -9570 -2700 -9560 -2400
rect -9500 -2700 -9490 -2400
rect -9150 -2700 -9140 -2400
rect -9080 -2700 -9070 -2400
rect -8730 -2700 -8720 -2400
rect -8660 -2700 -8650 -2400
rect -8310 -2700 -8300 -2400
rect -8240 -2700 -8230 -2400
rect -7910 -2700 -7900 -2400
rect -7840 -2700 -7830 -2400
rect -7490 -2700 -7480 -2400
rect -7420 -2700 -7410 -2400
rect -7070 -2700 -7060 -2400
rect -7000 -2700 -6990 -2400
rect -11490 -2880 -11480 -2740
rect -11290 -2880 -7050 -2740
rect -11250 -3200 -11240 -2920
rect -11180 -3200 -11170 -2920
rect -10830 -3200 -10820 -2920
rect -10760 -3200 -10750 -2920
rect -10410 -3200 -10400 -2920
rect -10340 -3200 -10330 -2920
rect -9990 -3200 -9980 -2920
rect -9920 -3200 -9910 -2920
rect -9570 -3200 -9560 -2920
rect -9500 -3200 -9490 -2920
rect -9150 -3200 -9140 -2920
rect -9080 -3200 -9070 -2920
rect -8730 -3200 -8720 -2920
rect -8660 -3200 -8650 -2920
rect -8310 -3200 -8300 -2920
rect -8240 -3200 -8230 -2920
rect -7910 -3200 -7900 -2920
rect -7840 -3200 -7830 -2920
rect -7490 -3200 -7480 -2920
rect -7420 -3200 -7410 -2920
rect -7070 -3200 -7060 -2920
rect -7000 -3200 -6990 -2920
rect -11490 -3390 -11480 -3250
rect -11290 -3390 -7050 -3250
rect -11180 -3400 -7060 -3390
rect -11250 -3720 -11240 -3440
rect -11180 -3720 -11170 -3440
rect -10830 -3720 -10820 -3440
rect -10760 -3720 -10750 -3440
rect -10410 -3720 -10400 -3440
rect -10340 -3720 -10330 -3440
rect -9990 -3720 -9980 -3440
rect -9920 -3720 -9910 -3440
rect -9570 -3720 -9560 -3440
rect -9500 -3720 -9490 -3440
rect -9150 -3720 -9140 -3440
rect -9080 -3720 -9070 -3440
rect -8730 -3720 -8720 -3440
rect -8660 -3720 -8650 -3440
rect -8310 -3720 -8300 -3440
rect -8240 -3720 -8230 -3440
rect -7910 -3720 -7900 -3440
rect -7840 -3720 -7830 -3440
rect -7490 -3720 -7480 -3440
rect -7420 -3720 -7410 -3440
rect -7070 -3720 -7060 -3440
rect -7000 -3720 -6990 -3440
rect -11490 -3910 -11480 -3770
rect -11290 -3910 -7050 -3770
rect -11180 -3920 -7060 -3910
rect -11250 -4240 -11240 -3960
rect -11180 -4240 -11170 -3960
rect -10830 -4240 -10820 -3960
rect -10760 -4240 -10750 -3960
rect -10410 -4240 -10400 -3960
rect -10340 -4240 -10330 -3960
rect -9990 -4240 -9980 -3960
rect -9920 -4240 -9910 -3960
rect -9570 -4240 -9560 -3960
rect -9500 -4240 -9490 -3960
rect -9150 -4240 -9140 -3960
rect -9080 -4240 -9070 -3960
rect -8730 -4240 -8720 -3960
rect -8660 -4240 -8650 -3960
rect -8310 -4240 -8300 -3960
rect -8240 -4240 -8230 -3960
rect -7910 -4240 -7900 -3960
rect -7840 -4240 -7830 -3960
rect -7490 -4240 -7480 -3960
rect -7420 -4240 -7410 -3960
rect -7070 -4240 -7060 -3960
rect -7000 -4240 -6990 -3960
rect -11180 -4290 -7060 -4280
rect -11490 -4430 -11480 -4290
rect -11290 -4430 -7050 -4290
rect -11250 -4760 -11240 -4480
rect -11180 -4760 -11170 -4480
rect -10830 -4760 -10820 -4480
rect -10760 -4760 -10750 -4480
rect -10410 -4760 -10400 -4480
rect -10340 -4760 -10330 -4480
rect -9990 -4760 -9980 -4480
rect -9920 -4760 -9910 -4480
rect -9570 -4760 -9560 -4480
rect -9500 -4760 -9490 -4480
rect -9150 -4760 -9140 -4480
rect -9080 -4760 -9070 -4480
rect -8730 -4760 -8720 -4480
rect -8660 -4760 -8650 -4480
rect -8310 -4760 -8300 -4480
rect -8240 -4760 -8230 -4480
rect -7910 -4760 -7900 -4480
rect -7840 -4760 -7830 -4480
rect -7490 -4760 -7480 -4480
rect -7420 -4760 -7410 -4480
rect -7070 -4760 -7060 -4480
rect -7000 -4760 -6990 -4480
rect -11180 -4810 -7060 -4800
rect -11490 -4950 -11480 -4810
rect -11290 -4950 -7050 -4810
rect -11250 -5280 -11240 -5000
rect -11180 -5280 -11170 -5000
rect -10830 -5280 -10820 -5000
rect -10760 -5280 -10750 -5000
rect -10410 -5280 -10400 -5000
rect -10340 -5280 -10330 -5000
rect -9990 -5280 -9980 -5000
rect -9920 -5280 -9910 -5000
rect -9570 -5280 -9560 -5000
rect -9500 -5280 -9490 -5000
rect -9150 -5280 -9140 -5000
rect -9080 -5280 -9070 -5000
rect -8730 -5280 -8720 -5000
rect -8660 -5280 -8650 -5000
rect -8310 -5280 -8300 -5000
rect -8240 -5280 -8230 -5000
rect -7910 -5280 -7900 -5000
rect -7840 -5280 -7830 -5000
rect -7490 -5280 -7480 -5000
rect -7420 -5280 -7410 -5000
rect -7070 -5280 -7060 -5000
rect -7000 -5280 -6990 -5000
rect -11180 -5330 -7060 -5320
rect -11490 -5470 -11480 -5330
rect -11290 -5470 -7050 -5330
rect -11250 -5800 -11240 -5520
rect -11180 -5800 -11170 -5520
rect -10830 -5800 -10820 -5520
rect -10760 -5800 -10750 -5520
rect -10410 -5800 -10400 -5520
rect -10340 -5800 -10330 -5520
rect -9990 -5800 -9980 -5520
rect -9920 -5800 -9910 -5520
rect -9570 -5800 -9560 -5520
rect -9500 -5800 -9490 -5520
rect -9150 -5800 -9140 -5520
rect -9080 -5800 -9070 -5520
rect -8730 -5800 -8720 -5520
rect -8660 -5800 -8650 -5520
rect -8310 -5800 -8300 -5520
rect -8240 -5800 -8230 -5520
rect -7910 -5800 -7900 -5520
rect -7840 -5800 -7830 -5520
rect -7490 -5800 -7480 -5520
rect -7420 -5800 -7410 -5520
rect -7050 -5800 -7040 -5520
rect -6980 -5800 -6970 -5520
rect -11180 -5850 -7060 -5840
rect -11490 -5990 -11480 -5850
rect -11290 -5990 -7050 -5850
rect -11250 -6320 -11240 -6040
rect -11180 -6320 -11170 -6040
rect -10830 -6320 -10820 -6040
rect -10760 -6320 -10750 -6040
rect -10410 -6320 -10400 -6040
rect -10340 -6320 -10330 -6040
rect -9990 -6320 -9980 -6040
rect -9920 -6320 -9910 -6040
rect -9570 -6320 -9560 -6040
rect -9500 -6320 -9490 -6040
rect -9150 -6320 -9140 -6040
rect -9080 -6320 -9070 -6040
rect -8730 -6320 -8720 -6040
rect -8660 -6320 -8650 -6040
rect -8310 -6320 -8300 -6040
rect -8240 -6320 -8230 -6040
rect -7910 -6320 -7900 -6040
rect -7840 -6320 -7830 -6040
rect -7490 -6320 -7480 -6040
rect -7420 -6320 -7410 -6040
rect -7070 -6320 -7060 -6040
rect -7000 -6320 -6990 -6040
rect -11480 -6390 -7050 -6360
rect -11180 -6400 -7060 -6390
rect -6936 -6454 -6930 -1350
rect -11342 -6460 -6930 -6454
rect -11342 -6500 -11330 -6460
rect -6880 -6500 -6730 -1350
rect -11342 -6506 -6874 -6500
rect -6936 -6512 -6874 -6506
<< via1 >>
rect -11480 4140 -11330 4980
rect -11240 4140 -11180 4860
rect -11040 4140 -10980 4860
rect -10860 4140 -10800 4860
rect -10660 4140 -10600 4860
rect -10480 4140 -10420 4860
rect -10280 4140 -10220 4860
rect -10080 4140 -10020 4860
rect -9900 4140 -9840 4860
rect -9700 4140 -9640 4860
rect -9520 4140 -9460 4860
rect -9320 4140 -9260 4860
rect -9120 4140 -9060 4860
rect -8940 4140 -8880 4860
rect -8740 4140 -8680 4860
rect -8540 4140 -8480 4860
rect -8360 4140 -8300 4860
rect -8160 4140 -8100 4860
rect -7980 4140 -7920 4860
rect -7780 4140 -7720 4860
rect -7580 4140 -7520 4860
rect -7380 4140 -7320 4860
rect -11480 2670 -11330 2740
rect -7270 2670 -7090 2740
rect -11480 2630 -11340 2670
rect -11340 2630 -11330 2670
rect -7270 2630 -7240 2670
rect -7240 2630 -7090 2670
rect -7270 2620 -7090 2630
rect -6930 2520 -6540 2580
rect -11140 2400 -11080 2470
rect -10950 2400 -10890 2460
rect -10760 2400 -10700 2460
rect -10570 2410 -10510 2470
rect -10370 2410 -10310 2470
rect -10180 2410 -10120 2470
rect -9990 2410 -9930 2470
rect -9800 2410 -9740 2470
rect -9610 2410 -9550 2470
rect -9410 2410 -9350 2470
rect -9220 2410 -9160 2470
rect -9030 2410 -8970 2470
rect -8840 2410 -8780 2470
rect -8640 2410 -8580 2470
rect -8450 2400 -8390 2460
rect -8260 2400 -8200 2460
rect -8070 2400 -8010 2460
rect -7880 2400 -7820 2460
rect -7680 2400 -7620 2460
rect -7490 2400 -7430 2460
rect -11240 2300 -11180 2370
rect -11050 2310 -10990 2370
rect -10850 2310 -10790 2370
rect -10660 2310 -10600 2370
rect -10470 2310 -10410 2370
rect -10280 2310 -10220 2370
rect -10090 2310 -10030 2370
rect -9890 2310 -9830 2370
rect -9700 2310 -9640 2370
rect -9510 2310 -9450 2370
rect -9320 2310 -9260 2370
rect -9130 2310 -9070 2370
rect -8930 2310 -8870 2370
rect -8740 2310 -8680 2370
rect -8550 2310 -8490 2370
rect -8360 2310 -8300 2370
rect -8160 2310 -8100 2370
rect -7970 2310 -7910 2370
rect -7780 2310 -7720 2370
rect -7590 2310 -7530 2370
rect -7390 2310 -7330 2370
rect -11140 2210 -11080 2280
rect -10950 2210 -10890 2280
rect -10760 2200 -10700 2270
rect -10570 2200 -10510 2270
rect -10370 2200 -10310 2270
rect -10180 2200 -10120 2270
rect -9990 2200 -9930 2270
rect -9800 2200 -9740 2270
rect -9610 2200 -9550 2270
rect -9410 2200 -9350 2270
rect -9220 2200 -9160 2270
rect -9030 2200 -8970 2270
rect -8840 2200 -8780 2270
rect -8640 2200 -8580 2270
rect -8450 2200 -8390 2270
rect -8260 2200 -8200 2270
rect -8070 2200 -8010 2270
rect -7880 2200 -7820 2270
rect -7680 2200 -7620 2270
rect -7490 2200 -7430 2270
rect -11240 2100 -11180 2170
rect -11050 2100 -10990 2170
rect -10850 2100 -10790 2170
rect -10660 2100 -10600 2170
rect -10470 2100 -10410 2170
rect -10280 2100 -10220 2170
rect -10090 2100 -10030 2170
rect -9890 2100 -9830 2170
rect -9700 2100 -9640 2170
rect -9510 2100 -9450 2170
rect -9320 2100 -9260 2170
rect -9130 2100 -9070 2170
rect -8930 2100 -8870 2170
rect -8740 2100 -8680 2170
rect -8550 2100 -8490 2170
rect -8360 2100 -8300 2170
rect -8160 2100 -8100 2170
rect -7970 2100 -7910 2170
rect -7780 2100 -7720 2170
rect -7590 2100 -7530 2170
rect -7390 2100 -7330 2170
rect -7270 2110 -7200 2480
rect -6930 1910 -6540 2060
rect -11140 1790 -11080 1850
rect -10950 1790 -10890 1850
rect -10760 1790 -10700 1850
rect -10570 1790 -10510 1850
rect -10370 1790 -10310 1850
rect -10180 1790 -10120 1850
rect -9990 1790 -9930 1850
rect -9800 1790 -9740 1850
rect -9610 1790 -9550 1850
rect -9410 1790 -9350 1850
rect -9220 1790 -9160 1850
rect -9030 1790 -8970 1850
rect -8840 1790 -8780 1850
rect -8640 1790 -8580 1850
rect -8450 1790 -8390 1850
rect -8260 1790 -8200 1850
rect -8070 1790 -8010 1850
rect -7880 1790 -7820 1850
rect -7680 1790 -7620 1850
rect -7490 1790 -7430 1850
rect -11240 1650 -11180 1710
rect -11050 1670 -10990 1730
rect -10850 1670 -10790 1730
rect -10660 1670 -10600 1730
rect -10470 1670 -10410 1730
rect -10280 1670 -10220 1730
rect -10090 1670 -10030 1730
rect -9890 1670 -9830 1730
rect -9700 1670 -9640 1730
rect -9510 1670 -9450 1730
rect -9320 1670 -9260 1730
rect -9130 1670 -9070 1730
rect -8930 1670 -8870 1730
rect -8740 1670 -8680 1730
rect -8550 1670 -8490 1730
rect -8360 1670 -8300 1730
rect -8160 1670 -8100 1730
rect -7970 1670 -7910 1730
rect -7780 1670 -7720 1730
rect -7590 1670 -7530 1730
rect -7390 1670 -7330 1730
rect -11140 1570 -11080 1630
rect -10950 1580 -10890 1640
rect -10760 1580 -10700 1640
rect -10570 1580 -10510 1640
rect -10370 1580 -10310 1640
rect -10180 1580 -10120 1640
rect -9990 1580 -9930 1640
rect -9800 1580 -9740 1640
rect -9610 1580 -9550 1640
rect -9410 1580 -9350 1640
rect -9220 1580 -9160 1640
rect -9030 1580 -8970 1640
rect -8840 1580 -8780 1640
rect -8640 1580 -8580 1640
rect -8450 1580 -8390 1640
rect -8260 1580 -8200 1640
rect -8070 1580 -8010 1640
rect -7880 1580 -7820 1640
rect -7680 1580 -7620 1640
rect -7490 1580 -7430 1640
rect -11240 1490 -11180 1550
rect -11040 1490 -10980 1550
rect -10850 1490 -10790 1550
rect -10660 1490 -10600 1550
rect -10470 1490 -10410 1550
rect -10280 1490 -10220 1550
rect -10090 1490 -10030 1550
rect -9890 1490 -9830 1550
rect -9700 1490 -9640 1550
rect -9510 1490 -9450 1550
rect -9320 1490 -9260 1550
rect -9130 1490 -9070 1550
rect -8930 1490 -8870 1550
rect -8740 1490 -8680 1550
rect -8550 1490 -8490 1550
rect -8360 1490 -8300 1550
rect -8160 1490 -8100 1550
rect -7970 1490 -7910 1550
rect -7780 1490 -7720 1550
rect -7590 1490 -7530 1550
rect -7390 1490 -7330 1550
rect -7270 1500 -7200 1870
rect -6930 1310 -6540 1460
rect -11140 1160 -11080 1220
rect -10950 1160 -10890 1220
rect -10760 1160 -10700 1220
rect -10570 1160 -10510 1220
rect -10370 1160 -10310 1220
rect -10180 1160 -10120 1220
rect -9990 1160 -9930 1220
rect -9800 1160 -9740 1220
rect -9610 1160 -9550 1220
rect -9410 1160 -9350 1220
rect -9220 1160 -9160 1220
rect -9030 1160 -8970 1220
rect -8840 1160 -8780 1220
rect -8640 1160 -8580 1220
rect -8450 1160 -8390 1220
rect -8260 1160 -8200 1220
rect -8070 1160 -8010 1220
rect -7880 1160 -7820 1220
rect -7680 1160 -7620 1220
rect -7490 1160 -7430 1220
rect -11240 1070 -11180 1130
rect -11050 1070 -10990 1130
rect -10850 1070 -10790 1130
rect -10660 1070 -10600 1130
rect -10470 1070 -10410 1130
rect -10280 1070 -10220 1130
rect -10090 1070 -10030 1130
rect -9890 1070 -9830 1130
rect -9700 1070 -9640 1130
rect -9510 1070 -9450 1130
rect -9320 1070 -9260 1130
rect -9130 1070 -9070 1130
rect -8930 1070 -8870 1130
rect -8740 1070 -8680 1130
rect -8550 1070 -8490 1130
rect -8360 1070 -8300 1130
rect -8160 1070 -8100 1130
rect -7970 1070 -7910 1130
rect -7780 1070 -7720 1130
rect -7590 1070 -7530 1130
rect -7390 1070 -7330 1130
rect -11140 970 -11080 1030
rect -10950 970 -10890 1030
rect -10760 970 -10700 1030
rect -10570 970 -10510 1030
rect -10370 970 -10310 1030
rect -10180 970 -10120 1030
rect -9990 970 -9930 1030
rect -9800 970 -9740 1030
rect -9610 970 -9550 1030
rect -9410 970 -9350 1030
rect -9220 970 -9160 1030
rect -9030 970 -8970 1030
rect -8840 970 -8780 1030
rect -8640 970 -8580 1030
rect -8450 980 -8390 1040
rect -8260 980 -8200 1040
rect -8070 980 -8010 1040
rect -7880 980 -7820 1040
rect -7680 980 -7620 1040
rect -7490 980 -7430 1040
rect -11240 880 -11180 940
rect -11050 880 -10990 940
rect -10850 880 -10790 940
rect -10660 880 -10600 940
rect -10470 880 -10410 940
rect -10280 880 -10220 940
rect -10090 880 -10030 940
rect -9890 880 -9830 940
rect -9700 880 -9640 940
rect -9510 880 -9450 940
rect -9320 880 -9260 940
rect -9130 880 -9070 940
rect -8930 880 -8870 940
rect -8740 880 -8680 940
rect -8550 880 -8490 940
rect -8360 890 -8300 950
rect -8160 890 -8100 950
rect -7970 890 -7910 950
rect -7780 890 -7720 950
rect -7590 890 -7530 950
rect -7390 890 -7330 950
rect -7270 900 -7200 1270
rect -6930 700 -6540 850
rect -11140 560 -11080 620
rect -10950 560 -10890 620
rect -10760 560 -10700 620
rect -10570 560 -10510 620
rect -10370 560 -10310 620
rect -10180 560 -10120 620
rect -9990 560 -9930 620
rect -9800 560 -9740 620
rect -9600 560 -9540 620
rect -9410 560 -9350 620
rect -9220 560 -9160 620
rect -9030 560 -8970 620
rect -8840 560 -8780 620
rect -8640 560 -8580 620
rect -8450 560 -8390 620
rect -8260 560 -8200 620
rect -8070 560 -8010 620
rect -7880 560 -7820 620
rect -7680 560 -7620 620
rect -7490 560 -7430 620
rect -11240 460 -11180 520
rect -11050 460 -10990 520
rect -10850 460 -10790 520
rect -10660 460 -10600 520
rect -10470 460 -10410 520
rect -10280 460 -10220 520
rect -10090 460 -10030 520
rect -9890 460 -9830 520
rect -9700 460 -9640 520
rect -9510 460 -9450 520
rect -9320 460 -9260 520
rect -9130 460 -9070 520
rect -8930 460 -8870 520
rect -8740 460 -8680 520
rect -8550 460 -8490 520
rect -8360 460 -8300 520
rect -8160 460 -8100 520
rect -7970 460 -7910 520
rect -7780 460 -7720 520
rect -7590 460 -7530 520
rect -7390 460 -7330 520
rect -11140 360 -11080 420
rect -10950 360 -10890 420
rect -10760 360 -10700 420
rect -10570 360 -10510 420
rect -10370 360 -10310 420
rect -10180 360 -10120 420
rect -9990 360 -9930 420
rect -9800 360 -9740 420
rect -9610 360 -9550 420
rect -9410 360 -9350 420
rect -9220 360 -9160 420
rect -9030 360 -8970 420
rect -8840 360 -8780 420
rect -8640 360 -8580 420
rect -8450 360 -8390 420
rect -8260 360 -8200 420
rect -8070 360 -8010 420
rect -7880 360 -7820 420
rect -7680 360 -7620 420
rect -7490 360 -7430 420
rect -11240 270 -11180 330
rect -11050 270 -10990 330
rect -10850 270 -10790 330
rect -10660 270 -10600 330
rect -10470 270 -10410 330
rect -10280 270 -10220 330
rect -10090 270 -10030 330
rect -9890 270 -9830 330
rect -9700 270 -9640 330
rect -9510 270 -9450 330
rect -9320 270 -9260 330
rect -9130 270 -9070 330
rect -8930 270 -8870 330
rect -8740 270 -8680 330
rect -8550 270 -8490 330
rect -8360 270 -8300 330
rect -8160 270 -8100 330
rect -7970 270 -7910 330
rect -7780 270 -7720 330
rect -7590 270 -7530 330
rect -7390 270 -7330 330
rect -7270 290 -7200 660
rect -6930 90 -6540 240
rect -11140 -40 -11080 20
rect -10950 -40 -10890 20
rect -10760 -40 -10700 20
rect -10570 -40 -10510 20
rect -10370 -40 -10310 20
rect -10180 -40 -10120 20
rect -9990 -40 -9930 20
rect -9800 -40 -9740 20
rect -9610 -40 -9550 20
rect -9410 -40 -9350 20
rect -9220 -40 -9160 20
rect -9030 -50 -8970 10
rect -8840 -50 -8780 10
rect -8640 -50 -8580 10
rect -8450 -50 -8390 10
rect -8260 -50 -8200 10
rect -8070 -50 -8010 10
rect -7880 -50 -7820 10
rect -7680 -50 -7620 10
rect -7490 -50 -7430 10
rect -11240 -140 -11180 -80
rect -11050 -140 -10990 -80
rect -10850 -130 -10790 -70
rect -10660 -130 -10600 -70
rect -10470 -130 -10410 -70
rect -10280 -130 -10220 -70
rect -10090 -130 -10030 -70
rect -9890 -130 -9830 -70
rect -9700 -130 -9640 -70
rect -9510 -130 -9450 -70
rect -9320 -130 -9260 -70
rect -9130 -130 -9070 -70
rect -8930 -140 -8870 -80
rect -8740 -140 -8680 -80
rect -8550 -140 -8490 -80
rect -8360 -140 -8300 -80
rect -8160 -140 -8100 -80
rect -7970 -140 -7910 -80
rect -7780 -140 -7720 -80
rect -7590 -140 -7530 -80
rect -7390 -140 -7330 -80
rect -11140 -230 -11080 -170
rect -10950 -230 -10890 -170
rect -10760 -230 -10700 -170
rect -10570 -230 -10510 -170
rect -10370 -230 -10310 -170
rect -10180 -230 -10120 -170
rect -9990 -230 -9930 -170
rect -9800 -230 -9740 -170
rect -9610 -230 -9550 -170
rect -9410 -230 -9350 -170
rect -9220 -230 -9160 -170
rect -9030 -230 -8970 -170
rect -8840 -230 -8780 -170
rect -8640 -230 -8580 -170
rect -8450 -230 -8390 -170
rect -8260 -230 -8200 -170
rect -8070 -230 -8010 -170
rect -7880 -230 -7820 -170
rect -7680 -230 -7620 -170
rect -7490 -230 -7430 -170
rect -11240 -320 -11180 -260
rect -11050 -320 -10990 -260
rect -10850 -320 -10790 -260
rect -10660 -320 -10600 -260
rect -10470 -320 -10410 -260
rect -10280 -320 -10220 -260
rect -10090 -320 -10030 -260
rect -9890 -320 -9830 -260
rect -9700 -320 -9640 -260
rect -9510 -320 -9450 -260
rect -9320 -320 -9260 -260
rect -9130 -320 -9070 -260
rect -8930 -320 -8870 -260
rect -8740 -320 -8680 -260
rect -8550 -320 -8490 -260
rect -8360 -320 -8300 -260
rect -8160 -320 -8100 -260
rect -7970 -320 -7910 -260
rect -7780 -320 -7720 -260
rect -7590 -320 -7530 -260
rect -7390 -320 -7330 -260
rect -7270 -320 -7200 50
rect -6930 -520 -6540 -370
rect -11140 -640 -11080 -580
rect -10950 -640 -10890 -580
rect -10760 -640 -10700 -580
rect -10570 -640 -10510 -580
rect -10370 -640 -10310 -580
rect -10180 -640 -10120 -580
rect -9990 -640 -9930 -580
rect -9800 -640 -9740 -580
rect -9610 -640 -9550 -580
rect -9410 -640 -9350 -580
rect -9220 -640 -9160 -580
rect -9030 -640 -8970 -580
rect -8840 -640 -8780 -580
rect -8640 -640 -8580 -580
rect -8450 -640 -8390 -580
rect -8260 -640 -8200 -580
rect -8070 -640 -8010 -580
rect -7880 -640 -7820 -580
rect -7680 -640 -7620 -580
rect -7490 -640 -7430 -580
rect -11240 -740 -11180 -680
rect -11050 -740 -10990 -680
rect -10850 -740 -10790 -680
rect -10660 -740 -10600 -680
rect -10470 -740 -10410 -680
rect -10280 -740 -10220 -680
rect -10090 -740 -10030 -680
rect -9890 -740 -9830 -680
rect -9700 -740 -9640 -680
rect -9510 -740 -9450 -680
rect -9320 -740 -9260 -680
rect -9130 -740 -9070 -680
rect -8930 -740 -8870 -680
rect -8740 -740 -8680 -680
rect -8550 -740 -8490 -680
rect -8360 -740 -8300 -680
rect -8160 -740 -8100 -680
rect -7970 -740 -7910 -680
rect -7780 -740 -7720 -680
rect -7590 -740 -7530 -680
rect -7390 -740 -7330 -680
rect -11140 -830 -11080 -770
rect -10950 -830 -10890 -770
rect -10760 -830 -10700 -770
rect -10570 -830 -10510 -770
rect -10370 -830 -10310 -770
rect -10180 -830 -10120 -770
rect -9990 -830 -9930 -770
rect -9800 -830 -9740 -770
rect -9610 -830 -9550 -770
rect -9410 -830 -9350 -770
rect -9220 -830 -9160 -770
rect -9030 -830 -8970 -770
rect -8840 -830 -8780 -770
rect -8640 -830 -8580 -770
rect -8450 -830 -8390 -770
rect -8260 -830 -8200 -770
rect -8070 -830 -8010 -770
rect -7880 -830 -7820 -770
rect -7680 -830 -7620 -770
rect -7490 -830 -7430 -770
rect -11240 -920 -11180 -860
rect -11050 -920 -10990 -860
rect -10850 -920 -10790 -860
rect -10660 -920 -10600 -860
rect -10470 -920 -10410 -860
rect -10280 -920 -10220 -860
rect -10090 -920 -10030 -860
rect -9890 -920 -9830 -860
rect -9700 -920 -9640 -860
rect -9510 -920 -9450 -860
rect -9320 -920 -9260 -860
rect -9130 -920 -9070 -860
rect -8930 -920 -8870 -860
rect -8740 -920 -8680 -860
rect -8550 -920 -8490 -860
rect -8360 -920 -8300 -860
rect -8160 -920 -8100 -860
rect -7970 -920 -7910 -860
rect -7780 -920 -7720 -860
rect -7590 -920 -7530 -860
rect -7390 -920 -7330 -860
rect -7270 -930 -7200 -560
rect -6930 -1020 -6540 -960
rect -11240 -1250 -11180 -1050
rect -10400 -1250 -10340 -1050
rect -9560 -1250 -9500 -1050
rect -8720 -1250 -8660 -1050
rect -7900 -1250 -7840 -1050
rect -7060 -1250 -7000 -1050
rect -6930 -1250 -6540 -1050
rect -11240 -1660 -11180 -1360
rect -10820 -1660 -10760 -1360
rect -10400 -1660 -10340 -1360
rect -9980 -1660 -9920 -1360
rect -9560 -1660 -9500 -1360
rect -9140 -1660 -9080 -1360
rect -8720 -1660 -8660 -1360
rect -8300 -1660 -8240 -1360
rect -7900 -1660 -7840 -1360
rect -7480 -1660 -7420 -1360
rect -7060 -1660 -7000 -1360
rect -11480 -1840 -11290 -1700
rect -11240 -2180 -11180 -1880
rect -10820 -2180 -10760 -1880
rect -10400 -2180 -10340 -1880
rect -9980 -2180 -9920 -1880
rect -9560 -2180 -9500 -1880
rect -9140 -2180 -9080 -1880
rect -8720 -2180 -8660 -1880
rect -8300 -2180 -8240 -1880
rect -7900 -2180 -7840 -1880
rect -7480 -2180 -7420 -1880
rect -7060 -2180 -7000 -1880
rect -11480 -2360 -11290 -2220
rect -11240 -2700 -11180 -2400
rect -10820 -2700 -10760 -2400
rect -10400 -2700 -10340 -2400
rect -9980 -2700 -9920 -2400
rect -9560 -2700 -9500 -2400
rect -9140 -2700 -9080 -2400
rect -8720 -2700 -8660 -2400
rect -8300 -2700 -8240 -2400
rect -7900 -2700 -7840 -2400
rect -7480 -2700 -7420 -2400
rect -7060 -2700 -7000 -2400
rect -11480 -2880 -11290 -2740
rect -11240 -3200 -11180 -2920
rect -10820 -3200 -10760 -2920
rect -10400 -3200 -10340 -2920
rect -9980 -3200 -9920 -2920
rect -9560 -3200 -9500 -2920
rect -9140 -3200 -9080 -2920
rect -8720 -3200 -8660 -2920
rect -8300 -3200 -8240 -2920
rect -7900 -3200 -7840 -2920
rect -7480 -3200 -7420 -2920
rect -7060 -3200 -7000 -2920
rect -11480 -3390 -11290 -3250
rect -11240 -3720 -11180 -3440
rect -10820 -3720 -10760 -3440
rect -10400 -3720 -10340 -3440
rect -9980 -3720 -9920 -3440
rect -9560 -3720 -9500 -3440
rect -9140 -3720 -9080 -3440
rect -8720 -3720 -8660 -3440
rect -8300 -3720 -8240 -3440
rect -7900 -3720 -7840 -3440
rect -7480 -3720 -7420 -3440
rect -7060 -3720 -7000 -3440
rect -11480 -3910 -11290 -3770
rect -11240 -4240 -11180 -3960
rect -10820 -4240 -10760 -3960
rect -10400 -4240 -10340 -3960
rect -9980 -4240 -9920 -3960
rect -9560 -4240 -9500 -3960
rect -9140 -4240 -9080 -3960
rect -8720 -4240 -8660 -3960
rect -8300 -4240 -8240 -3960
rect -7900 -4240 -7840 -3960
rect -7480 -4240 -7420 -3960
rect -7060 -4240 -7000 -3960
rect -11480 -4430 -11290 -4290
rect -11240 -4760 -11180 -4480
rect -10820 -4760 -10760 -4480
rect -10400 -4760 -10340 -4480
rect -9980 -4760 -9920 -4480
rect -9560 -4760 -9500 -4480
rect -9140 -4760 -9080 -4480
rect -8720 -4760 -8660 -4480
rect -8300 -4760 -8240 -4480
rect -7900 -4760 -7840 -4480
rect -7480 -4760 -7420 -4480
rect -7060 -4760 -7000 -4480
rect -11480 -4950 -11290 -4810
rect -11240 -5280 -11180 -5000
rect -10820 -5280 -10760 -5000
rect -10400 -5280 -10340 -5000
rect -9980 -5280 -9920 -5000
rect -9560 -5280 -9500 -5000
rect -9140 -5280 -9080 -5000
rect -8720 -5280 -8660 -5000
rect -8300 -5280 -8240 -5000
rect -7900 -5280 -7840 -5000
rect -7480 -5280 -7420 -5000
rect -7060 -5280 -7000 -5000
rect -11480 -5470 -11290 -5330
rect -11240 -5800 -11180 -5520
rect -10820 -5800 -10760 -5520
rect -10400 -5800 -10340 -5520
rect -9980 -5800 -9920 -5520
rect -9560 -5800 -9500 -5520
rect -9140 -5800 -9080 -5520
rect -8720 -5800 -8660 -5520
rect -8300 -5800 -8240 -5520
rect -7900 -5800 -7840 -5520
rect -7480 -5800 -7420 -5520
rect -7040 -5800 -6980 -5520
rect -11480 -5990 -11290 -5850
rect -11240 -6320 -11180 -6040
rect -10820 -6320 -10760 -6040
rect -10400 -6320 -10340 -6040
rect -9980 -6320 -9920 -6040
rect -9560 -6320 -9500 -6040
rect -9140 -6320 -9080 -6040
rect -8720 -6320 -8660 -6040
rect -8300 -6320 -8240 -6040
rect -7900 -6320 -7840 -6040
rect -7480 -6320 -7420 -6040
rect -7060 -6320 -7000 -6040
<< metal2 >>
rect -11480 4980 -11330 4990
rect -11480 2740 -11330 4140
rect -11480 2620 -11330 2630
rect -11240 4860 -11180 4980
rect -11240 2370 -11180 4140
rect -11240 2170 -11180 2300
rect -11240 1710 -11180 2100
rect -11240 1550 -11180 1650
rect -11240 1130 -11180 1490
rect -11240 940 -11180 1070
rect -11240 520 -11180 880
rect -11240 330 -11180 460
rect -11240 -80 -11180 270
rect -11240 -260 -11180 -140
rect -11240 -680 -11180 -320
rect -11240 -860 -11180 -740
rect -11240 -940 -11180 -920
rect -11140 3980 -11080 4980
rect -11140 2470 -11080 3160
rect -11140 2280 -11080 2400
rect -11140 1850 -11080 2210
rect -11140 1630 -11080 1790
rect -11140 1220 -11080 1570
rect -11140 1030 -11080 1160
rect -11140 620 -11080 970
rect -11140 420 -11080 560
rect -11140 20 -11080 360
rect -11140 -170 -11080 -40
rect -11140 -580 -11080 -230
rect -11140 -770 -11080 -640
rect -11140 -940 -11080 -830
rect -11050 4860 -10980 4980
rect -11050 4140 -11040 4860
rect -11050 4130 -10980 4140
rect -11050 2370 -10990 4130
rect -10950 3990 -10890 4980
rect -10860 4860 -10790 4980
rect -10800 4140 -10790 4860
rect -10860 4130 -10790 4140
rect -10960 3980 -10890 3990
rect -10900 3160 -10890 3980
rect -10960 3150 -10890 3160
rect -11050 2170 -10990 2310
rect -11050 1730 -10990 2100
rect -11050 1560 -10990 1670
rect -10950 2460 -10890 3150
rect -10950 2280 -10890 2400
rect -10950 1850 -10890 2210
rect -10950 1640 -10890 1790
rect -11050 1550 -10980 1560
rect -11050 1490 -11040 1550
rect -11050 1480 -10980 1490
rect -11050 1130 -10990 1480
rect -11050 940 -10990 1070
rect -11050 520 -10990 880
rect -11050 330 -10990 460
rect -11050 -80 -10990 270
rect -11050 -260 -10990 -140
rect -11050 -680 -10990 -320
rect -11050 -860 -10990 -740
rect -11050 -940 -10990 -920
rect -10950 1220 -10890 1580
rect -10950 1030 -10890 1160
rect -10950 620 -10890 970
rect -10950 420 -10890 560
rect -10950 20 -10890 360
rect -10950 -170 -10890 -40
rect -10950 -580 -10890 -230
rect -10950 -770 -10890 -640
rect -10950 -940 -10890 -830
rect -10850 2370 -10790 4130
rect -10850 2170 -10790 2310
rect -10850 1730 -10790 2100
rect -10850 1550 -10790 1670
rect -10850 1130 -10790 1490
rect -10850 940 -10790 1070
rect -10850 520 -10790 880
rect -10850 330 -10790 460
rect -10850 -70 -10790 270
rect -10850 -260 -10790 -130
rect -10850 -680 -10790 -320
rect -10850 -860 -10790 -740
rect -10850 -940 -10790 -920
rect -10760 3980 -10700 4980
rect -10760 2460 -10700 3160
rect -10760 2270 -10700 2400
rect -10760 1850 -10700 2200
rect -10760 1640 -10700 1790
rect -10760 1220 -10700 1580
rect -10760 1030 -10700 1160
rect -10760 620 -10700 970
rect -10760 420 -10700 560
rect -10760 20 -10700 360
rect -10760 -170 -10700 -40
rect -10760 -580 -10700 -230
rect -10760 -770 -10700 -640
rect -10760 -940 -10700 -830
rect -10660 4860 -10600 4980
rect -10660 2370 -10600 4140
rect -10660 2170 -10600 2310
rect -10660 1730 -10600 2100
rect -10660 1550 -10600 1670
rect -10660 1130 -10600 1490
rect -10660 940 -10600 1070
rect -10660 520 -10600 880
rect -10660 330 -10600 460
rect -10660 -70 -10600 270
rect -10660 -260 -10600 -130
rect -10660 -680 -10600 -320
rect -10660 -860 -10600 -740
rect -10660 -940 -10600 -920
rect -10570 3990 -10510 4980
rect -10480 4860 -10410 4980
rect -10420 4140 -10410 4860
rect -10480 4130 -10410 4140
rect -10570 3980 -10500 3990
rect -10570 3160 -10560 3980
rect -10570 3150 -10500 3160
rect -10570 2470 -10510 3150
rect -10570 2270 -10510 2410
rect -10570 1850 -10510 2200
rect -10570 1640 -10510 1790
rect -10570 1220 -10510 1580
rect -10570 1030 -10510 1160
rect -10570 620 -10510 970
rect -10570 420 -10510 560
rect -10570 20 -10510 360
rect -10570 -170 -10510 -40
rect -10570 -580 -10510 -230
rect -10570 -770 -10510 -640
rect -10570 -940 -10510 -830
rect -10470 2370 -10410 4130
rect -10370 3990 -10310 4980
rect -10380 3980 -10310 3990
rect -10320 3160 -10310 3980
rect -10380 3150 -10310 3160
rect -10470 2170 -10410 2310
rect -10470 1730 -10410 2100
rect -10470 1550 -10410 1670
rect -10470 1130 -10410 1490
rect -10470 940 -10410 1070
rect -10470 520 -10410 880
rect -10470 330 -10410 460
rect -10470 -70 -10410 270
rect -10470 -260 -10410 -130
rect -10470 -680 -10410 -320
rect -10470 -860 -10410 -740
rect -10470 -940 -10410 -920
rect -10370 2470 -10310 3150
rect -10370 2270 -10310 2410
rect -10370 1850 -10310 2200
rect -10370 1640 -10310 1790
rect -10370 1220 -10310 1580
rect -10370 1030 -10310 1160
rect -10370 620 -10310 970
rect -10370 420 -10310 560
rect -10370 20 -10310 360
rect -10370 -170 -10310 -40
rect -10370 -580 -10310 -230
rect -10370 -770 -10310 -640
rect -10370 -940 -10310 -830
rect -10280 4860 -10220 4980
rect -10280 2370 -10220 4140
rect -10280 2170 -10220 2310
rect -10280 1730 -10220 2100
rect -10280 1550 -10220 1670
rect -10280 1130 -10220 1490
rect -10280 940 -10220 1070
rect -10280 520 -10220 880
rect -10280 330 -10220 460
rect -10280 -70 -10220 270
rect -10280 -260 -10220 -130
rect -10280 -680 -10220 -320
rect -10280 -860 -10220 -740
rect -10280 -940 -10220 -920
rect -10180 3980 -10120 4980
rect -10180 2470 -10120 3160
rect -10180 2270 -10120 2410
rect -10180 1850 -10120 2200
rect -10180 1640 -10120 1790
rect -10180 1220 -10120 1580
rect -10180 1030 -10120 1160
rect -10180 620 -10120 970
rect -10180 420 -10120 560
rect -10180 20 -10120 360
rect -10180 -170 -10120 -40
rect -10180 -580 -10120 -230
rect -10180 -770 -10120 -640
rect -10180 -940 -10120 -830
rect -10090 4860 -10020 4980
rect -10090 4140 -10080 4860
rect -10090 4130 -10020 4140
rect -10090 2370 -10030 4130
rect -9990 3990 -9930 4980
rect -9900 4860 -9830 4980
rect -9840 4140 -9830 4860
rect -9900 4130 -9830 4140
rect -10000 3980 -9930 3990
rect -9940 3160 -9930 3980
rect -10000 3150 -9930 3160
rect -10090 2170 -10030 2310
rect -10090 1730 -10030 2100
rect -10090 1550 -10030 1670
rect -10090 1130 -10030 1490
rect -10090 940 -10030 1070
rect -10090 520 -10030 880
rect -10090 330 -10030 460
rect -10090 -70 -10030 270
rect -10090 -260 -10030 -130
rect -10090 -680 -10030 -320
rect -10090 -860 -10030 -740
rect -10090 -940 -10030 -920
rect -9990 2470 -9930 3150
rect -9990 2270 -9930 2410
rect -9990 1850 -9930 2200
rect -9990 1640 -9930 1790
rect -9990 1220 -9930 1580
rect -9990 1030 -9930 1160
rect -9990 620 -9930 970
rect -9990 420 -9930 560
rect -9990 20 -9930 360
rect -9990 -170 -9930 -40
rect -9990 -580 -9930 -230
rect -9990 -770 -9930 -640
rect -9990 -940 -9930 -830
rect -9890 2370 -9830 4130
rect -9890 2170 -9830 2310
rect -9890 1730 -9830 2100
rect -9890 1550 -9830 1670
rect -9890 1130 -9830 1490
rect -9890 940 -9830 1070
rect -9890 520 -9830 880
rect -9890 330 -9830 460
rect -9890 -70 -9830 270
rect -9890 -260 -9830 -130
rect -9890 -680 -9830 -320
rect -9890 -860 -9830 -740
rect -9890 -940 -9830 -920
rect -9800 3980 -9740 4980
rect -9800 2470 -9740 3160
rect -9800 2270 -9740 2410
rect -9800 1850 -9740 2200
rect -9800 1640 -9740 1790
rect -9800 1220 -9740 1580
rect -9800 1030 -9740 1160
rect -9800 620 -9740 970
rect -9800 420 -9740 560
rect -9800 20 -9740 360
rect -9800 -170 -9740 -40
rect -9800 -580 -9740 -230
rect -9800 -770 -9740 -640
rect -9800 -940 -9740 -830
rect -9700 4860 -9640 4980
rect -9700 2370 -9640 4140
rect -9700 2170 -9640 2310
rect -9700 1730 -9640 2100
rect -9700 1550 -9640 1670
rect -9700 1130 -9640 1490
rect -9700 940 -9640 1070
rect -9700 520 -9640 880
rect -9700 330 -9640 460
rect -9700 -70 -9640 270
rect -9700 -260 -9640 -130
rect -9700 -680 -9640 -320
rect -9700 -860 -9640 -740
rect -9700 -940 -9640 -920
rect -9610 3990 -9550 4980
rect -9520 4860 -9450 4980
rect -9460 4140 -9450 4860
rect -9520 4130 -9450 4140
rect -9610 3980 -9540 3990
rect -9610 3160 -9600 3980
rect -9610 3150 -9540 3160
rect -9610 2470 -9550 3150
rect -9610 2270 -9550 2410
rect -9610 1850 -9550 2200
rect -9610 1640 -9550 1790
rect -9610 1220 -9550 1580
rect -9610 1030 -9550 1160
rect -9610 630 -9550 970
rect -9510 2370 -9450 4130
rect -9410 3990 -9350 4980
rect -9420 3980 -9350 3990
rect -9360 3160 -9350 3980
rect -9420 3150 -9350 3160
rect -9510 2170 -9450 2310
rect -9510 1730 -9450 2100
rect -9510 1550 -9450 1670
rect -9510 1130 -9450 1490
rect -9510 940 -9450 1070
rect -9610 620 -9540 630
rect -9610 560 -9600 620
rect -9610 550 -9540 560
rect -9610 420 -9550 550
rect -9610 20 -9550 360
rect -9610 -170 -9550 -40
rect -9610 -580 -9550 -230
rect -9610 -770 -9550 -640
rect -9610 -940 -9550 -830
rect -9510 520 -9450 880
rect -9510 330 -9450 460
rect -9510 -70 -9450 270
rect -9510 -260 -9450 -130
rect -9510 -680 -9450 -320
rect -9510 -860 -9450 -740
rect -9510 -940 -9450 -920
rect -9410 2470 -9350 3150
rect -9410 2270 -9350 2410
rect -9410 1850 -9350 2200
rect -9410 1640 -9350 1790
rect -9410 1220 -9350 1580
rect -9410 1030 -9350 1160
rect -9410 620 -9350 970
rect -9410 420 -9350 560
rect -9410 20 -9350 360
rect -9410 -170 -9350 -40
rect -9410 -580 -9350 -230
rect -9410 -770 -9350 -640
rect -9410 -940 -9350 -830
rect -9320 4860 -9260 4980
rect -9320 2370 -9260 4140
rect -9320 2170 -9260 2310
rect -9320 1730 -9260 2100
rect -9320 1550 -9260 1670
rect -9320 1130 -9260 1490
rect -9320 940 -9260 1070
rect -9320 520 -9260 880
rect -9320 330 -9260 460
rect -9320 -70 -9260 270
rect -9320 -260 -9260 -130
rect -9320 -680 -9260 -320
rect -9320 -860 -9260 -740
rect -9320 -940 -9260 -920
rect -9220 3980 -9160 4980
rect -9220 2470 -9160 3160
rect -9220 2270 -9160 2410
rect -9220 1850 -9160 2200
rect -9220 1640 -9160 1790
rect -9220 1220 -9160 1580
rect -9220 1030 -9160 1160
rect -9220 620 -9160 970
rect -9220 420 -9160 560
rect -9220 20 -9160 360
rect -9220 -170 -9160 -40
rect -9220 -580 -9160 -230
rect -9220 -770 -9160 -640
rect -9220 -940 -9160 -830
rect -9130 4860 -9060 4980
rect -9130 4140 -9120 4860
rect -9130 4130 -9060 4140
rect -9130 2370 -9070 4130
rect -9030 3990 -8970 4980
rect -8940 4860 -8870 4980
rect -8880 4140 -8870 4860
rect -8940 4130 -8870 4140
rect -9040 3980 -8970 3990
rect -8980 3160 -8970 3980
rect -9040 3150 -8970 3160
rect -9130 2170 -9070 2310
rect -9130 1730 -9070 2100
rect -9130 1550 -9070 1670
rect -9130 1130 -9070 1490
rect -9130 940 -9070 1070
rect -9130 520 -9070 880
rect -9130 330 -9070 460
rect -9130 -70 -9070 270
rect -9130 -260 -9070 -130
rect -9130 -680 -9070 -320
rect -9130 -860 -9070 -740
rect -9130 -940 -9070 -920
rect -9030 2470 -8970 3150
rect -9030 2270 -8970 2410
rect -9030 1850 -8970 2200
rect -9030 1640 -8970 1790
rect -9030 1220 -8970 1580
rect -9030 1030 -8970 1160
rect -9030 620 -8970 970
rect -9030 420 -8970 560
rect -9030 10 -8970 360
rect -9030 -170 -8970 -50
rect -9030 -580 -8970 -230
rect -9030 -770 -8970 -640
rect -9030 -940 -8970 -830
rect -8930 2370 -8870 4130
rect -8930 2170 -8870 2310
rect -8930 1730 -8870 2100
rect -8930 1550 -8870 1670
rect -8930 1130 -8870 1490
rect -8930 940 -8870 1070
rect -8930 520 -8870 880
rect -8930 330 -8870 460
rect -8930 -80 -8870 270
rect -8930 -260 -8870 -140
rect -8930 -680 -8870 -320
rect -8930 -860 -8870 -740
rect -8930 -940 -8870 -920
rect -8840 3980 -8780 4980
rect -8840 2470 -8780 3160
rect -8840 2270 -8780 2410
rect -8840 1850 -8780 2200
rect -8840 1640 -8780 1790
rect -8840 1220 -8780 1580
rect -8840 1030 -8780 1160
rect -8840 620 -8780 970
rect -8840 420 -8780 560
rect -8840 10 -8780 360
rect -8840 -170 -8780 -50
rect -8840 -580 -8780 -230
rect -8840 -770 -8780 -640
rect -8840 -940 -8780 -830
rect -8740 4860 -8680 4980
rect -8740 2370 -8680 4140
rect -8740 2170 -8680 2310
rect -8740 1730 -8680 2100
rect -8740 1550 -8680 1670
rect -8740 1130 -8680 1490
rect -8740 940 -8680 1070
rect -8740 520 -8680 880
rect -8740 330 -8680 460
rect -8740 -80 -8680 270
rect -8740 -260 -8680 -140
rect -8740 -680 -8680 -320
rect -8740 -860 -8680 -740
rect -8740 -940 -8680 -920
rect -8640 3980 -8580 4980
rect -8640 2470 -8580 3160
rect -8640 2270 -8580 2410
rect -8640 1850 -8580 2200
rect -8640 1640 -8580 1790
rect -8640 1220 -8580 1580
rect -8640 1030 -8580 1160
rect -8640 620 -8580 970
rect -8640 420 -8580 560
rect -8640 10 -8580 360
rect -8640 -170 -8580 -50
rect -8640 -580 -8580 -230
rect -8640 -770 -8580 -640
rect -8640 -940 -8580 -830
rect -8550 4860 -8480 4980
rect -8550 4140 -8540 4860
rect -8550 4130 -8480 4140
rect -8550 2370 -8490 4130
rect -8450 3990 -8390 4980
rect -8460 3980 -8390 3990
rect -8400 3160 -8390 3980
rect -8460 3150 -8390 3160
rect -8550 2170 -8490 2310
rect -8550 1730 -8490 2100
rect -8550 1550 -8490 1670
rect -8550 1130 -8490 1490
rect -8550 940 -8490 1070
rect -8550 520 -8490 880
rect -8550 330 -8490 460
rect -8550 -80 -8490 270
rect -8550 -260 -8490 -140
rect -8550 -680 -8490 -320
rect -8550 -860 -8490 -740
rect -8550 -940 -8490 -920
rect -8450 2460 -8390 3150
rect -8450 2270 -8390 2400
rect -8450 1850 -8390 2200
rect -8450 1640 -8390 1790
rect -8450 1220 -8390 1580
rect -8450 1040 -8390 1160
rect -8450 620 -8390 980
rect -8450 420 -8390 560
rect -8450 10 -8390 360
rect -8450 -170 -8390 -50
rect -8450 -580 -8390 -230
rect -8450 -770 -8390 -640
rect -8450 -940 -8390 -830
rect -8360 4860 -8300 4980
rect -8360 2370 -8300 4140
rect -8360 2170 -8300 2310
rect -8360 1730 -8300 2100
rect -8360 1550 -8300 1670
rect -8360 1130 -8300 1490
rect -8360 950 -8300 1070
rect -8360 520 -8300 890
rect -8360 330 -8300 460
rect -8360 -80 -8300 270
rect -8360 -260 -8300 -140
rect -8360 -680 -8300 -320
rect -8360 -860 -8300 -740
rect -8360 -940 -8300 -920
rect -8260 3980 -8200 4980
rect -8260 2460 -8200 3160
rect -8260 2270 -8200 2400
rect -8260 1850 -8200 2200
rect -8260 1640 -8200 1790
rect -8260 1220 -8200 1580
rect -8260 1040 -8200 1160
rect -8260 620 -8200 980
rect -8260 420 -8200 560
rect -8260 10 -8200 360
rect -8260 -170 -8200 -50
rect -8260 -580 -8200 -230
rect -8260 -770 -8200 -640
rect -8260 -940 -8200 -830
rect -8160 4860 -8100 4980
rect -8160 2370 -8100 4140
rect -8160 2170 -8100 2310
rect -8160 1730 -8100 2100
rect -8160 1550 -8100 1670
rect -8160 1130 -8100 1490
rect -8160 950 -8100 1070
rect -8160 520 -8100 890
rect -8160 330 -8100 460
rect -8160 -80 -8100 270
rect -8160 -260 -8100 -140
rect -8160 -680 -8100 -320
rect -8160 -860 -8100 -740
rect -8160 -940 -8100 -920
rect -8070 3990 -8010 4980
rect -7980 4860 -7910 4980
rect -7920 4140 -7910 4860
rect -7980 4130 -7910 4140
rect -8070 3980 -8000 3990
rect -8070 3160 -8060 3980
rect -8070 3150 -8000 3160
rect -8070 2460 -8010 3150
rect -8070 2270 -8010 2400
rect -8070 1850 -8010 2200
rect -8070 1640 -8010 1790
rect -8070 1220 -8010 1580
rect -8070 1040 -8010 1160
rect -8070 620 -8010 980
rect -8070 420 -8010 560
rect -8070 10 -8010 360
rect -8070 -170 -8010 -50
rect -8070 -580 -8010 -230
rect -8070 -770 -8010 -640
rect -8070 -940 -8010 -830
rect -7970 2370 -7910 4130
rect -7970 2170 -7910 2310
rect -7970 1730 -7910 2100
rect -7970 1550 -7910 1670
rect -7970 1130 -7910 1490
rect -7970 950 -7910 1070
rect -7970 520 -7910 890
rect -7970 330 -7910 460
rect -7970 -80 -7910 270
rect -7970 -260 -7910 -140
rect -7970 -680 -7910 -320
rect -7970 -860 -7910 -740
rect -7970 -940 -7910 -920
rect -7880 3980 -7820 4980
rect -7880 2460 -7820 3160
rect -7880 2270 -7820 2400
rect -7880 1850 -7820 2200
rect -7880 1640 -7820 1790
rect -7880 1220 -7820 1580
rect -7880 1040 -7820 1160
rect -7880 620 -7820 980
rect -7880 420 -7820 560
rect -7880 10 -7820 360
rect -7880 -170 -7820 -50
rect -7880 -580 -7820 -230
rect -7880 -770 -7820 -640
rect -7880 -940 -7820 -830
rect -7780 4860 -7720 4980
rect -7780 2370 -7720 4140
rect -7780 2170 -7720 2310
rect -7780 1730 -7720 2100
rect -7780 1550 -7720 1670
rect -7780 1130 -7720 1490
rect -7780 950 -7720 1070
rect -7780 520 -7720 890
rect -7780 330 -7720 460
rect -7780 -80 -7720 270
rect -7780 -260 -7720 -140
rect -7780 -680 -7720 -320
rect -7780 -860 -7720 -740
rect -7780 -940 -7720 -920
rect -7680 3980 -7620 4980
rect -7680 2460 -7620 3160
rect -7680 2270 -7620 2400
rect -7680 1850 -7620 2200
rect -7680 1640 -7620 1790
rect -7680 1220 -7620 1580
rect -7680 1040 -7620 1160
rect -7680 620 -7620 980
rect -7680 420 -7620 560
rect -7680 10 -7620 360
rect -7680 -170 -7620 -50
rect -7680 -580 -7620 -230
rect -7680 -770 -7620 -640
rect -7680 -940 -7620 -830
rect -7590 4860 -7520 4980
rect -7590 4140 -7580 4860
rect -7590 4130 -7520 4140
rect -7590 2370 -7530 4130
rect -7490 3980 -7420 4980
rect -7590 2170 -7530 2310
rect -7590 1730 -7530 2100
rect -7590 1550 -7530 1670
rect -7590 1130 -7530 1490
rect -7590 950 -7530 1070
rect -7590 520 -7530 890
rect -7590 330 -7530 460
rect -7590 -80 -7530 270
rect -7590 -260 -7530 -140
rect -7590 -680 -7530 -320
rect -7590 -860 -7530 -740
rect -7590 -940 -7530 -920
rect -7490 3160 -7480 3480
rect -7490 3150 -7420 3160
rect -7390 4860 -7320 4980
rect -7390 4140 -7380 4860
rect -7390 4130 -7320 4140
rect -7490 2460 -7430 3150
rect -7490 2270 -7430 2400
rect -7490 1850 -7430 2200
rect -7490 1640 -7430 1790
rect -7490 1220 -7430 1580
rect -7490 1040 -7430 1160
rect -7490 620 -7430 980
rect -7490 420 -7430 560
rect -7490 10 -7430 360
rect -7490 -170 -7430 -50
rect -7490 -580 -7430 -230
rect -7490 -770 -7430 -640
rect -7490 -940 -7430 -830
rect -7390 2370 -7330 4130
rect -7390 2170 -7330 2310
rect -7390 1730 -7330 2100
rect -7390 1550 -7330 1670
rect -7390 1130 -7330 1490
rect -7390 950 -7330 1070
rect -7390 520 -7330 890
rect -7390 330 -7330 460
rect -7390 -80 -7330 270
rect -7390 -260 -7330 -140
rect -7390 -680 -7330 -320
rect -7390 -860 -7330 -740
rect -7390 -940 -7330 -920
rect -7270 2740 -7090 2750
rect -7270 2480 -7090 2620
rect -7200 2110 -7090 2480
rect -7270 1870 -7090 2110
rect -7200 1500 -7090 1870
rect -7270 1270 -7090 1500
rect -7200 900 -7090 1270
rect -7270 660 -7090 900
rect -7200 290 -7090 660
rect -7270 50 -7090 290
rect -7200 -320 -7090 50
rect -7270 -560 -7090 -320
rect -7200 -930 -7090 -560
rect -7270 -960 -7090 -930
rect -6930 2580 -6540 2590
rect -6930 2060 -6540 2520
rect -6930 1460 -6540 1910
rect -6930 850 -6540 1310
rect -6930 240 -6540 700
rect -6930 -370 -6540 90
rect -6930 -960 -6540 -520
rect -11240 -1050 -11180 -1040
rect -10400 -1050 -10340 -1040
rect -11480 -1700 -11290 -1290
rect -11480 -2220 -11290 -1840
rect -11480 -2740 -11290 -2360
rect -11480 -3250 -11290 -2880
rect -11480 -3770 -11290 -3390
rect -11480 -4290 -11290 -3910
rect -11480 -4810 -11290 -4430
rect -11480 -5330 -11290 -4950
rect -11480 -5850 -11290 -5470
rect -11480 -6390 -11290 -5990
rect -11240 -1360 -11180 -1250
rect -11240 -1880 -11180 -1660
rect -11240 -2400 -11180 -2180
rect -11240 -2920 -11180 -2700
rect -11240 -3440 -11180 -3200
rect -11240 -3960 -11180 -3720
rect -11240 -4480 -11180 -4240
rect -11240 -5000 -11180 -4760
rect -11240 -5520 -11180 -5280
rect -11240 -6040 -11180 -5800
rect -11240 -6640 -11180 -6320
rect -10820 -1360 -10760 -1200
rect -10820 -1880 -10760 -1660
rect -10820 -2400 -10760 -2180
rect -10820 -2920 -10760 -2700
rect -10820 -3440 -10760 -3200
rect -10820 -3960 -10760 -3720
rect -10820 -4480 -10760 -4240
rect -10820 -5000 -10760 -4760
rect -10820 -5520 -10760 -5280
rect -10820 -6040 -10760 -5800
rect -10820 -6450 -10760 -6320
rect -9560 -1050 -9500 -1040
rect -10400 -1360 -10340 -1250
rect -10400 -1880 -10340 -1660
rect -10400 -2400 -10340 -2180
rect -10400 -2920 -10340 -2700
rect -10400 -3440 -10340 -3200
rect -10400 -3960 -10340 -3720
rect -10400 -4480 -10340 -4240
rect -10400 -5000 -10340 -4760
rect -10400 -5520 -10340 -5280
rect -10400 -6040 -10340 -5800
rect -10400 -6640 -10340 -6320
rect -9980 -1360 -9920 -1180
rect -9980 -1880 -9920 -1660
rect -9980 -2400 -9920 -2180
rect -9980 -2920 -9920 -2700
rect -9980 -3440 -9920 -3200
rect -9980 -3960 -9920 -3720
rect -9980 -4480 -9920 -4240
rect -9980 -5000 -9920 -4760
rect -9980 -5520 -9920 -5280
rect -9980 -6040 -9920 -5800
rect -9980 -6450 -9920 -6320
rect -10820 -6780 -10760 -6770
rect -8720 -1050 -8660 -1040
rect -9560 -1360 -9500 -1250
rect -9560 -1880 -9500 -1660
rect -9560 -2400 -9500 -2180
rect -9560 -2920 -9500 -2700
rect -9560 -3440 -9500 -3200
rect -9560 -3960 -9500 -3720
rect -9560 -4480 -9500 -4240
rect -9560 -5000 -9500 -4760
rect -9560 -5520 -9500 -5280
rect -9560 -6040 -9500 -5800
rect -9560 -6640 -9500 -6320
rect -9140 -1360 -9080 -1180
rect -9140 -1880 -9080 -1660
rect -9140 -2400 -9080 -2180
rect -9140 -2920 -9080 -2700
rect -9140 -3440 -9080 -3200
rect -9140 -3960 -9080 -3720
rect -9140 -4480 -9080 -4240
rect -9140 -5000 -9080 -4760
rect -9140 -5520 -9080 -5280
rect -9140 -6040 -9080 -5800
rect -9140 -6450 -9080 -6320
rect -9980 -6780 -9920 -6770
rect -7900 -1050 -7840 -1040
rect -8720 -1360 -8660 -1250
rect -8720 -1880 -8660 -1660
rect -8720 -2400 -8660 -2180
rect -8720 -2920 -8660 -2700
rect -8720 -3440 -8660 -3200
rect -8720 -3960 -8660 -3720
rect -8720 -4480 -8660 -4240
rect -8720 -5000 -8660 -4760
rect -8720 -5520 -8660 -5280
rect -8720 -6040 -8660 -5800
rect -8720 -6640 -8660 -6320
rect -8300 -1360 -8240 -1180
rect -8300 -1880 -8240 -1660
rect -8300 -2400 -8240 -2180
rect -8300 -2920 -8240 -2700
rect -8300 -3440 -8240 -3200
rect -8300 -3960 -8240 -3720
rect -8300 -4480 -8240 -4240
rect -8300 -5000 -8240 -4760
rect -8300 -5520 -8240 -5280
rect -8300 -6040 -8240 -5800
rect -8300 -6460 -8240 -6320
rect -9140 -6780 -9080 -6770
rect -7060 -1050 -7000 -1040
rect -7900 -1360 -7840 -1250
rect -7900 -1880 -7840 -1660
rect -7900 -2400 -7840 -2180
rect -7900 -2920 -7840 -2700
rect -7900 -3440 -7840 -3200
rect -7900 -3960 -7840 -3720
rect -7900 -4480 -7840 -4240
rect -7900 -5000 -7840 -4760
rect -7900 -5520 -7840 -5280
rect -7900 -6040 -7840 -5800
rect -7900 -6640 -7840 -6320
rect -7480 -1360 -7420 -1180
rect -7480 -1880 -7420 -1660
rect -7480 -2400 -7420 -2180
rect -7480 -2920 -7420 -2700
rect -7480 -3440 -7420 -3200
rect -7480 -3960 -7420 -3720
rect -7480 -4480 -7420 -4240
rect -7480 -5000 -7420 -4760
rect -7480 -5520 -7420 -5280
rect -7480 -6040 -7420 -5800
rect -7480 -6450 -7420 -6320
rect -7060 -1360 -7000 -1250
rect -6930 -1050 -6540 -1020
rect -6930 -1260 -6540 -1250
rect -7060 -1880 -7000 -1660
rect -7060 -2400 -7000 -2180
rect -7060 -2920 -7000 -2700
rect -7060 -3440 -7000 -3200
rect -7060 -3960 -7000 -3720
rect -7060 -4480 -7000 -4240
rect -7060 -5000 -7000 -4760
rect -7060 -5510 -7000 -5280
rect -7060 -5520 -6980 -5510
rect -7060 -5800 -7040 -5520
rect -7060 -5810 -6980 -5800
rect -7060 -6040 -7000 -5810
rect -7060 -6640 -7000 -6320
rect -7480 -6780 -7420 -6770
rect -8300 -6790 -8240 -6780
<< via2 >>
rect -11140 3160 -11080 3980
rect -10960 3160 -10900 3980
rect -10760 3160 -10700 3980
rect -10560 3160 -10500 3980
rect -10380 3160 -10320 3980
rect -10180 3160 -10120 3980
rect -10000 3160 -9940 3980
rect -9800 3160 -9740 3980
rect -9600 3160 -9540 3980
rect -9420 3160 -9360 3980
rect -9220 3160 -9160 3980
rect -9040 3160 -8980 3980
rect -8840 3160 -8780 3980
rect -8640 3160 -8580 3980
rect -8460 3160 -8400 3980
rect -8260 3160 -8200 3980
rect -8060 3160 -8000 3980
rect -7880 3160 -7820 3980
rect -7680 3160 -7620 3980
rect -7480 3160 -7420 3980
rect -10820 -6770 -10760 -6450
rect -9980 -6770 -9920 -6450
rect -9140 -6770 -9080 -6450
rect -8300 -6780 -8240 -6460
rect -7480 -6770 -7420 -6450
<< metal3 >>
rect -11150 3980 -11070 3985
rect -10970 3980 -10890 3985
rect -10770 3980 -10690 3985
rect -10570 3980 -10490 3985
rect -10390 3980 -10310 3985
rect -10190 3980 -10110 3985
rect -10010 3980 -9930 3985
rect -9810 3980 -9730 3985
rect -9610 3980 -9530 3985
rect -9430 3980 -9350 3985
rect -9230 3980 -9150 3985
rect -9050 3980 -8970 3985
rect -8850 3980 -8770 3985
rect -8650 3980 -8570 3985
rect -8470 3980 -8390 3985
rect -8270 3980 -8190 3985
rect -8070 3980 -7990 3985
rect -7890 3980 -7810 3985
rect -7690 3980 -7610 3985
rect -7490 3980 -7410 3985
rect -11240 3160 -11140 3980
rect -11080 3160 -10960 3980
rect -10900 3160 -10760 3980
rect -10700 3160 -10560 3980
rect -10500 3160 -10380 3980
rect -10320 3160 -10180 3980
rect -10120 3160 -10000 3980
rect -9940 3160 -9800 3980
rect -9740 3160 -9600 3980
rect -9540 3160 -9420 3980
rect -9360 3160 -9220 3980
rect -9160 3160 -9040 3980
rect -8980 3160 -8840 3980
rect -8780 3160 -8640 3980
rect -8580 3160 -8460 3980
rect -8400 3160 -8260 3980
rect -8200 3160 -8060 3980
rect -8000 3160 -7880 3980
rect -7820 3160 -7680 3980
rect -7620 3160 -7480 3980
rect -7420 3160 -7390 3980
rect -11240 3150 -7390 3160
rect -6740 3150 -6730 3980
rect -3470 3120 -3260 3200
rect -140 3120 70 3200
rect -10830 -6450 -10750 -6445
rect -10830 -6490 -10820 -6450
rect -11240 -6770 -10820 -6490
rect -10760 -6490 -10750 -6450
rect -9990 -6450 -9910 -6445
rect -9990 -6490 -9980 -6450
rect -10760 -6770 -9980 -6490
rect -9920 -6490 -9910 -6450
rect -9150 -6450 -9070 -6445
rect -9150 -6490 -9140 -6450
rect -9920 -6770 -9140 -6490
rect -9080 -6490 -9070 -6450
rect -7490 -6450 -7410 -6445
rect -8310 -6460 -8230 -6455
rect -8310 -6490 -8300 -6460
rect -9080 -6770 -8300 -6490
rect -10830 -6775 -10750 -6770
rect -9990 -6775 -9910 -6770
rect -9150 -6775 -9070 -6770
rect -8310 -6780 -8300 -6770
rect -8240 -6490 -8230 -6460
rect -7490 -6490 -7480 -6450
rect -8240 -6770 -7480 -6490
rect -7420 -6490 -7410 -6450
rect -3400 -6490 -3260 3120
rect -80 -6490 60 3120
rect -7420 -6500 -6890 -6490
rect -6610 -6500 3280 -6490
rect -7420 -6770 3280 -6500
rect -8240 -6780 -8230 -6770
rect -7490 -6775 -7410 -6770
rect -8310 -6785 -8230 -6780
<< via3 >>
rect -7390 3150 -6740 3980
<< metal4 >>
rect -7391 3980 -6739 3981
rect -7391 3150 -7390 3980
rect -6740 3430 2580 3980
rect -6740 3310 -6650 3430
rect -6740 3150 -6640 3310
rect -5110 3180 -4960 3430
rect -1780 3220 -1650 3430
rect 1530 3210 1670 3430
rect -7391 3149 -6739 3150
use sky130_fd_pr__nfet_01v8_RE4H9G  sky130_fd_pr__nfet_01v8_RE4H9G_0
timestamp 1619113446
transform 1 0 -9287 0 1 773
box -2087 -1925 2087 1925
use sky130_fd_pr__cap_mim_m3_1_6BP6N2  sky130_fd_pr__cap_mim_m3_1_6BP6N2_0
timestamp 1619113446
transform 1 0 -1669 0 1 -1700
box -4969 -4950 4968 4950
use sky130_fd_pr__nfet_01v8_B8HNLY  sky130_fd_pr__nfet_01v8_B8HNLY_0
timestamp 1619113446
transform 1 0 -9116 0 1 -3842
box -2257 -2691 2257 2691
<< labels >>
rlabel metal4 -6740 3430 2580 3980 1 vout
rlabel metal1 -11340 -1250 -11240 -1050 1 vin
rlabel metal1 -11330 4140 -11240 4980 1 vss
rlabel metal2 -11480 -1700 -11290 -1290 1 vdd
rlabel metal3 -7420 -6770 3280 -6500 1 net1
<< end >>
