magic
tech sky130A
magscale 1 2
timestamp 1624053917
<< error_s >>
rect 5348 2621 5383 2655
rect 9312 2621 9347 2655
rect 13276 2621 13311 2655
rect 17240 2621 17275 2655
rect 5349 2602 5383 2621
rect 5735 2602 5788 2603
rect 9313 2602 9347 2621
rect 9699 2602 9752 2603
rect 13277 2602 13311 2621
rect 13663 2602 13716 2603
rect 17241 2602 17275 2621
rect 17627 2602 17680 2603
rect 5179 2553 5237 2559
rect 5179 2519 5191 2553
rect 5179 2513 5237 2519
rect 3556 2397 3591 2431
rect 2086 2363 2121 2381
rect 2050 2348 2121 2363
rect 2401 2348 2436 2382
rect 3557 2378 3591 2397
rect 2050 2110 2120 2348
rect 2402 2329 2436 2348
rect 3576 2335 3591 2378
rect 2421 2286 2436 2329
rect 2232 2280 2290 2286
rect 2232 2246 2244 2280
rect 2232 2240 2290 2246
rect 1668 2072 2120 2110
rect 2200 2072 2234 2106
rect 2288 2072 2322 2106
rect 2402 2072 2436 2286
rect 2455 2295 2490 2329
rect 2455 2072 2489 2295
rect 2601 2227 2659 2233
rect 2601 2193 2613 2227
rect 2771 2204 2805 2233
rect 2601 2187 2659 2193
rect 2771 2168 2841 2204
rect 2771 2134 2859 2168
rect 3139 2134 3174 2168
rect 2771 2110 2858 2134
rect 3140 2115 3174 2134
rect 3205 2151 3210 2204
rect 3241 2151 3275 2335
rect 3387 2329 3445 2335
rect 3387 2295 3399 2329
rect 3387 2289 3445 2295
rect 3557 2169 3591 2335
rect 3610 2344 3645 2378
rect 3925 2344 3960 2378
rect 3557 2151 3597 2169
rect 3205 2136 3597 2151
rect 3205 2115 3596 2136
rect 3159 2110 3174 2115
rect 3193 2110 3596 2115
rect 2569 2072 2603 2106
rect 2657 2072 2691 2106
rect 2771 2072 3596 2110
rect 3610 2072 3644 2344
rect 3926 2325 3960 2344
rect 3945 2297 3960 2325
rect 3979 2297 4014 2325
rect 4075 2297 4233 2325
rect 4027 2291 4233 2297
rect 4294 2291 4329 2325
rect 3756 2276 3814 2282
rect 3756 2242 3768 2276
rect 3926 2263 3960 2282
rect 4027 2263 4185 2291
rect 3756 2236 3814 2242
rect 3724 2170 3758 2199
rect 3658 2136 3678 2170
rect 3712 2136 3858 2170
rect 3892 2136 3912 2170
rect 3712 2102 3801 2115
rect 3844 2106 3846 2136
rect 3853 2106 3858 2136
rect 3686 2072 3801 2102
rect 3812 2072 3874 2106
rect 334 2021 369 2055
rect 335 2002 369 2021
rect 1668 2038 3874 2072
rect 3878 2072 3912 2136
rect 3926 2091 3965 2263
rect 3979 2091 4013 2263
rect 4105 2211 4121 2223
rect 4105 2201 4125 2211
rect 4105 2195 4121 2201
rect 4089 2180 4091 2189
rect 4099 2180 4123 2195
rect 4137 2189 4161 2223
rect 4261 2201 4281 2291
rect 4073 2161 4139 2180
rect 4077 2155 4135 2161
rect 4093 2142 4127 2146
rect 4139 2142 4163 2145
rect 4181 2142 4201 2146
rect 4081 2130 4139 2142
rect 4175 2130 4201 2142
rect 4081 2127 4136 2130
rect 4045 2114 4047 2118
rect 4059 2114 4079 2118
rect 4033 2110 4085 2114
rect 4087 2110 4127 2127
rect 4033 2091 4079 2110
rect 4093 2091 4127 2110
rect 4133 2114 4167 2118
rect 4133 2110 4173 2114
rect 4175 2110 4205 2130
rect 4133 2091 4167 2110
rect 4181 2106 4205 2110
rect 4213 2106 4215 2146
rect 4181 2091 4215 2106
rect 4222 2091 4227 2142
rect 4247 2091 4281 2201
rect 4295 2244 4329 2291
rect 4348 2244 4383 2272
rect 4444 2244 4602 2272
rect 5179 2263 5237 2269
rect 4295 2210 4335 2244
rect 4396 2238 4602 2244
rect 4663 2238 4698 2255
rect 4396 2210 4554 2238
rect 4295 2091 4334 2210
rect 4348 2091 4382 2210
rect 4474 2158 4490 2170
rect 4474 2148 4494 2158
rect 4474 2142 4490 2148
rect 4458 2127 4460 2136
rect 4468 2127 4492 2142
rect 4506 2138 4530 2170
rect 4630 2148 4650 2238
rect 4504 2130 4552 2138
rect 4442 2110 4508 2127
rect 4442 2108 4580 2110
rect 4504 2106 4580 2108
rect 3926 2083 4382 2091
rect 4462 2089 4496 2106
rect 4504 2102 4584 2106
rect 4508 2089 4532 2092
rect 4450 2083 4508 2089
rect 4550 2083 4584 2102
rect 3926 2072 4584 2083
rect 4591 2072 4596 2089
rect 4616 2072 4650 2148
rect 4664 2237 4698 2238
rect 4664 2201 4734 2237
rect 5179 2229 5191 2263
rect 5179 2223 5237 2229
rect 4664 2167 4752 2201
rect 4664 2110 4751 2167
rect 5129 2148 5287 2161
rect 5368 2148 5383 2602
rect 5402 2568 5437 2602
rect 5717 2568 5788 2602
rect 5402 2148 5436 2568
rect 5718 2567 5788 2568
rect 5735 2533 5806 2567
rect 6086 2533 6121 2567
rect 5548 2500 5606 2506
rect 5548 2466 5560 2500
rect 5548 2460 5606 2466
rect 5627 2327 5650 2381
rect 5735 2363 5805 2533
rect 6087 2514 6121 2533
rect 9143 2553 9201 2559
rect 9143 2519 9155 2553
rect 5917 2465 5975 2471
rect 5917 2431 5929 2465
rect 5917 2425 5975 2431
rect 5885 2363 5919 2388
rect 5996 2382 6019 2384
rect 6106 2382 6121 2514
rect 6140 2480 6175 2514
rect 6455 2480 6490 2514
rect 9143 2513 9201 2519
rect 6140 2382 6174 2480
rect 6456 2461 6490 2480
rect 6475 2418 6490 2461
rect 6286 2412 6344 2418
rect 6286 2382 6298 2412
rect 6050 2381 6073 2382
rect 6050 2363 6085 2381
rect 5735 2348 6085 2363
rect 6140 2348 6400 2382
rect 5681 2293 5704 2327
rect 5735 2293 6084 2348
rect 5681 2248 5715 2293
rect 5684 2231 5715 2248
rect 5548 2210 5606 2216
rect 5548 2176 5560 2210
rect 5548 2170 5606 2176
rect 5129 2127 5340 2148
rect 5052 2110 5067 2127
rect 5086 2126 5121 2127
rect 5182 2126 5340 2127
rect 5086 2114 5402 2126
rect 5086 2110 5120 2114
rect 5681 2110 5715 2231
rect 5718 2110 6084 2293
rect 4664 2078 6084 2110
rect 6087 2078 6121 2348
rect 6140 2221 6174 2348
rect 6366 2335 6400 2348
rect 6254 2331 6288 2335
rect 6342 2331 6400 2335
rect 6242 2323 6300 2331
rect 6330 2323 6400 2331
rect 6242 2280 6289 2323
rect 6342 2314 6400 2323
rect 6192 2246 6212 2280
rect 6216 2246 6289 2280
rect 6130 2199 6174 2221
rect 6242 2199 6288 2246
rect 6130 2187 6175 2199
rect 6254 2187 6288 2199
rect 6140 2078 6208 2187
rect 6252 2163 6288 2187
rect 6252 2151 6286 2163
rect 6252 2106 6298 2151
rect 6252 2104 6332 2106
rect 4664 2072 6210 2078
rect 6252 2072 6324 2104
rect 6332 2072 6348 2104
rect 6366 2072 6400 2314
rect 6419 2295 6454 2329
rect 6419 2072 6453 2295
rect 6456 2072 6490 2418
rect 6509 2427 6544 2461
rect 6509 2329 6543 2427
rect 7520 2397 7555 2431
rect 7521 2378 7555 2397
rect 6655 2359 6713 2365
rect 6655 2329 6667 2359
rect 6825 2336 6859 2365
rect 6509 2295 6753 2329
rect 6509 2168 6543 2295
rect 6735 2282 6753 2295
rect 6623 2278 6657 2282
rect 6711 2278 6753 2282
rect 6825 2300 6895 2336
rect 6611 2270 6669 2278
rect 6699 2270 6757 2278
rect 6611 2227 6658 2270
rect 6711 2261 6757 2270
rect 6561 2193 6581 2227
rect 6585 2193 6658 2227
rect 6735 2222 6757 2261
rect 6825 2266 6913 2300
rect 6734 2204 6769 2222
rect 6825 2204 6912 2266
rect 6499 2146 6543 2168
rect 6611 2146 6657 2193
rect 6734 2168 6912 2204
rect 7024 2198 7082 2204
rect 7024 2168 7036 2198
rect 6499 2134 6544 2146
rect 6623 2134 6657 2146
rect 6509 2072 6577 2134
rect 6621 2110 6657 2134
rect 6735 2134 7138 2168
rect 6735 2126 6912 2134
rect 7104 2130 7138 2134
rect 6992 2126 7026 2130
rect 7080 2126 7138 2130
rect 6621 2106 6655 2110
rect 6621 2098 6657 2106
rect 6667 2098 6669 2126
rect 6699 2110 6912 2126
rect 6980 2110 7038 2126
rect 7068 2110 7138 2126
rect 7169 2151 7264 2336
rect 7540 2335 7555 2378
rect 7351 2329 7409 2335
rect 7351 2295 7363 2329
rect 7351 2289 7409 2295
rect 7521 2169 7555 2335
rect 7574 2344 7609 2378
rect 7889 2344 7924 2378
rect 7521 2151 7561 2169
rect 7169 2136 7561 2151
rect 7169 2115 7560 2136
rect 7157 2110 7560 2115
rect 6699 2098 7560 2110
rect 6621 2085 6667 2098
rect 6711 2094 7560 2098
rect 6735 2085 7560 2094
rect 6621 2072 7560 2085
rect 7574 2072 7608 2344
rect 7890 2325 7924 2344
rect 7909 2297 7924 2325
rect 7943 2297 7978 2325
rect 8039 2297 8197 2325
rect 7991 2291 8197 2297
rect 8258 2291 8293 2325
rect 7720 2276 7778 2282
rect 7720 2242 7732 2276
rect 7890 2263 7924 2282
rect 7991 2263 8149 2291
rect 7720 2236 7778 2242
rect 7688 2170 7722 2199
rect 7622 2136 7642 2170
rect 7676 2136 7822 2170
rect 7856 2136 7876 2170
rect 7676 2102 7765 2115
rect 7808 2106 7810 2136
rect 7817 2106 7822 2136
rect 7650 2072 7765 2102
rect 7776 2072 7838 2106
rect 3878 2038 3880 2072
rect 3892 2038 3916 2072
rect 721 2002 774 2003
rect -17 1814 281 1867
rect 354 1814 369 2002
rect 388 1968 423 2002
rect 703 1968 774 2002
rect 388 1814 422 1968
rect 704 1967 774 1968
rect 721 1933 792 1967
rect 1072 1933 1107 1967
rect 534 1900 592 1906
rect 534 1866 546 1900
rect 534 1860 592 1866
rect -17 1761 650 1814
rect 721 1761 791 1933
rect 1073 1914 1107 1933
rect 1668 1966 2120 2038
rect 2188 2019 2228 2038
rect 2266 2019 2334 2038
rect 2204 2000 2318 2006
rect 2244 1984 2288 1990
rect 2213 1972 2325 1984
rect 2132 1966 2148 1972
rect 2213 1969 2328 1972
rect 1668 1956 2158 1966
rect 1668 1946 2164 1956
rect 1668 1940 2120 1946
rect 1668 1932 2112 1940
rect 1092 1871 1107 1914
rect 903 1865 961 1871
rect 903 1831 915 1865
rect 903 1825 961 1831
rect -17 1725 791 1761
rect -17 1706 983 1725
rect -17 1691 993 1706
rect -17 1629 791 1691
rect 859 1657 872 1670
rect -17 1623 837 1629
rect -17 1589 791 1623
rect 837 1589 841 1623
rect 859 1604 875 1657
rect 871 1600 875 1604
rect 949 1600 993 1691
rect 1073 1672 1107 1871
rect 1126 1880 1161 1914
rect 1441 1880 1476 1914
rect 1668 1897 2103 1932
rect 1126 1672 1160 1880
rect 1442 1861 1476 1880
rect 1272 1812 1330 1818
rect 1272 1778 1284 1812
rect 1272 1772 1330 1778
rect 1002 1604 1027 1672
rect 1073 1638 1352 1672
rect -17 1583 837 1589
rect -17 1564 791 1583
rect -17 1517 815 1564
rect 949 1563 983 1600
rect 903 1557 983 1563
rect -17 1472 791 1517
rect 865 1506 869 1546
rect 899 1538 928 1557
rect 949 1538 983 1557
rect 899 1523 983 1538
rect 903 1517 983 1523
rect 949 1510 983 1517
rect 835 1472 869 1506
rect 875 1489 989 1510
rect 949 1472 983 1489
rect 1002 1472 1036 1604
rect 1073 1472 1107 1638
rect 1126 1576 1160 1638
rect 1318 1637 1352 1638
rect 1461 1637 1476 1861
rect 1495 1827 1530 1861
rect 1681 1853 2103 1897
rect 2114 1870 2120 1940
rect 2138 1940 2164 1946
rect 2138 1922 2158 1940
rect 2228 1938 2328 1969
rect 2333 1956 2354 1984
rect 2402 1966 2436 2038
rect 2455 1984 2489 2038
rect 2594 2010 2603 2038
rect 2540 1990 2569 1996
rect 2586 1990 2615 2010
rect 2540 1984 2615 1990
rect 2370 1956 2436 1966
rect 2364 1946 2436 1956
rect 2364 1940 2401 1946
rect 2228 1932 2290 1938
rect 2228 1922 2266 1932
rect 2308 1906 2328 1938
rect 2380 1922 2401 1940
rect 2402 1940 2436 1946
rect 2402 1932 2414 1940
rect 2415 1932 2436 1940
rect 2402 1922 2436 1932
rect 2402 1870 2414 1922
rect 2114 1859 2159 1870
rect 1704 1827 1845 1853
rect 2086 1836 2090 1853
rect 2114 1847 2148 1859
rect 2103 1836 2159 1847
rect 2208 1836 2354 1870
rect 2369 1859 2414 1870
rect 2380 1847 2414 1859
rect 2415 1847 2436 1922
rect 2369 1836 2436 1847
rect 2440 1836 2490 1984
rect 2540 1978 2603 1984
rect 2540 1972 2569 1978
rect 2594 1962 2603 1978
rect 2628 1967 2637 2038
rect 2678 1990 2703 2038
rect 2657 1984 2703 1990
rect 2771 1984 3596 2038
rect 3610 2015 3644 2038
rect 3712 2034 3788 2038
rect 3712 2015 3770 2034
rect 3798 2015 3858 2038
rect 3610 2002 3832 2015
rect 3844 2011 3846 2015
rect 3840 2002 3842 2010
rect 3610 2000 3842 2002
rect 2657 1978 2691 1984
rect 2617 1966 2645 1967
rect 2732 1966 2757 1984
rect 2563 1906 2574 1953
rect 2616 1925 2674 1966
rect 2601 1919 2674 1925
rect 2597 1885 2674 1919
rect 2601 1879 2663 1885
rect 2616 1869 2663 1879
rect 1495 1637 1529 1827
rect 1668 1800 1734 1808
rect 1716 1780 1737 1793
rect 1668 1772 1737 1780
rect 1716 1763 1737 1772
rect 1811 1763 1845 1827
rect 2032 1825 2090 1836
rect 1953 1804 2090 1825
rect 2208 1804 2266 1836
rect 2296 1804 2354 1836
rect 2440 1817 2489 1836
rect 2771 1817 3608 1984
rect 3610 1966 3644 2000
rect 3676 1987 3678 1991
rect 3690 1987 3710 1991
rect 3734 1987 3798 2000
rect 3840 1987 3842 2000
rect 3664 1966 3717 1987
rect 3734 1984 3810 1987
rect 3734 1972 3849 1984
rect 3610 1956 3717 1966
rect 3718 1968 3849 1972
rect 3718 1956 3740 1968
rect 3610 1946 3740 1956
rect 3610 1922 3655 1946
rect 3664 1922 3740 1946
rect 3752 1956 3849 1968
rect 3752 1934 3818 1956
rect 3610 1866 3644 1922
rect 3664 1866 3670 1922
rect 3676 1900 3710 1922
rect 3718 1906 3740 1922
rect 3764 1922 3828 1934
rect 3764 1918 3818 1922
rect 3672 1866 3710 1900
rect 3764 1866 3798 1918
rect 3878 1906 3916 2038
rect 3926 2038 7838 2072
rect 7842 2072 7876 2136
rect 7890 2091 7929 2263
rect 7943 2091 7977 2263
rect 8069 2211 8085 2223
rect 8069 2201 8089 2211
rect 8069 2195 8085 2201
rect 8053 2180 8055 2189
rect 8063 2180 8087 2195
rect 8101 2189 8125 2223
rect 8225 2201 8245 2291
rect 8037 2161 8103 2180
rect 8041 2155 8099 2161
rect 8057 2142 8091 2146
rect 8103 2142 8127 2145
rect 8145 2142 8165 2146
rect 8045 2130 8103 2142
rect 8139 2130 8165 2142
rect 8045 2127 8100 2130
rect 8009 2114 8011 2118
rect 8023 2114 8043 2118
rect 7997 2110 8049 2114
rect 8051 2110 8091 2127
rect 7997 2091 8043 2110
rect 8057 2091 8091 2110
rect 8097 2114 8131 2118
rect 8097 2110 8137 2114
rect 8139 2110 8169 2130
rect 8097 2091 8131 2110
rect 8145 2106 8169 2110
rect 8177 2106 8179 2146
rect 8145 2091 8179 2106
rect 8186 2091 8191 2142
rect 8211 2091 8245 2201
rect 8259 2244 8293 2291
rect 8312 2244 8347 2272
rect 8408 2244 8566 2272
rect 9143 2263 9201 2269
rect 8259 2210 8299 2244
rect 8360 2238 8566 2244
rect 8627 2238 8662 2255
rect 8360 2210 8518 2238
rect 8259 2091 8298 2210
rect 8312 2091 8346 2210
rect 8438 2158 8454 2170
rect 8438 2148 8458 2158
rect 8438 2142 8454 2148
rect 8422 2127 8424 2136
rect 8432 2127 8456 2142
rect 8470 2138 8494 2170
rect 8594 2148 8614 2238
rect 8468 2130 8516 2138
rect 8406 2110 8472 2127
rect 8406 2108 8544 2110
rect 8468 2106 8544 2108
rect 7890 2083 8346 2091
rect 8426 2089 8460 2106
rect 8468 2102 8548 2106
rect 8472 2089 8496 2092
rect 8414 2083 8472 2089
rect 8514 2083 8548 2102
rect 7890 2072 8548 2083
rect 8555 2072 8560 2089
rect 8580 2072 8614 2148
rect 8628 2237 8662 2238
rect 8628 2201 8698 2237
rect 9143 2229 9155 2263
rect 9143 2223 9201 2229
rect 8628 2167 8716 2201
rect 8628 2110 8715 2167
rect 9093 2148 9251 2161
rect 9332 2148 9347 2602
rect 9366 2568 9401 2602
rect 9681 2568 9752 2602
rect 9366 2148 9400 2568
rect 9682 2567 9752 2568
rect 9699 2533 9770 2567
rect 10050 2533 10085 2567
rect 9512 2500 9570 2506
rect 9512 2466 9524 2500
rect 9512 2460 9570 2466
rect 9591 2327 9614 2381
rect 9699 2363 9769 2533
rect 10051 2514 10085 2533
rect 13107 2553 13165 2559
rect 13107 2519 13119 2553
rect 9881 2465 9939 2471
rect 9881 2431 9893 2465
rect 9881 2425 9939 2431
rect 9849 2363 9883 2388
rect 9960 2382 9983 2384
rect 10070 2382 10085 2514
rect 10104 2480 10139 2514
rect 10419 2480 10454 2514
rect 13107 2513 13165 2519
rect 10104 2382 10138 2480
rect 10420 2461 10454 2480
rect 10439 2418 10454 2461
rect 10250 2412 10308 2418
rect 10250 2382 10262 2412
rect 10014 2381 10037 2382
rect 10014 2363 10049 2381
rect 9699 2348 10049 2363
rect 10104 2348 10364 2382
rect 9645 2293 9668 2327
rect 9699 2293 10048 2348
rect 9645 2248 9679 2293
rect 9648 2231 9679 2248
rect 9512 2210 9570 2216
rect 9512 2176 9524 2210
rect 9512 2170 9570 2176
rect 9093 2127 9304 2148
rect 9016 2110 9031 2127
rect 9050 2126 9085 2127
rect 9146 2126 9304 2127
rect 9050 2114 9366 2126
rect 9050 2110 9084 2114
rect 9645 2110 9679 2231
rect 9682 2110 10048 2293
rect 8628 2078 10048 2110
rect 10051 2078 10085 2348
rect 10104 2221 10138 2348
rect 10330 2335 10364 2348
rect 10218 2331 10252 2335
rect 10306 2331 10364 2335
rect 10206 2323 10264 2331
rect 10294 2323 10364 2331
rect 10206 2280 10253 2323
rect 10306 2314 10364 2323
rect 10156 2246 10176 2280
rect 10180 2246 10253 2280
rect 10094 2199 10138 2221
rect 10206 2199 10252 2246
rect 10094 2187 10139 2199
rect 10218 2187 10252 2199
rect 10104 2078 10172 2187
rect 10216 2163 10252 2187
rect 10216 2151 10250 2163
rect 10216 2106 10262 2151
rect 10216 2104 10296 2106
rect 8628 2072 10174 2078
rect 10216 2072 10288 2104
rect 10296 2072 10312 2104
rect 10330 2072 10364 2314
rect 10383 2295 10418 2329
rect 10383 2072 10417 2295
rect 10420 2072 10454 2418
rect 10473 2427 10508 2461
rect 10473 2329 10507 2427
rect 11484 2397 11519 2431
rect 11485 2378 11519 2397
rect 10619 2359 10677 2365
rect 10619 2329 10631 2359
rect 10789 2336 10823 2365
rect 10473 2295 10717 2329
rect 10473 2168 10507 2295
rect 10699 2282 10717 2295
rect 10587 2278 10621 2282
rect 10675 2278 10717 2282
rect 10789 2300 10859 2336
rect 10575 2270 10633 2278
rect 10663 2270 10721 2278
rect 10575 2227 10622 2270
rect 10675 2261 10721 2270
rect 10525 2193 10545 2227
rect 10549 2193 10622 2227
rect 10699 2222 10721 2261
rect 10789 2266 10877 2300
rect 10698 2204 10733 2222
rect 10789 2204 10876 2266
rect 10463 2146 10507 2168
rect 10575 2146 10621 2193
rect 10698 2168 10876 2204
rect 10988 2198 11046 2204
rect 10988 2168 11000 2198
rect 10463 2134 10508 2146
rect 10587 2134 10621 2146
rect 10473 2072 10541 2134
rect 10585 2110 10621 2134
rect 10699 2134 11102 2168
rect 10699 2126 10876 2134
rect 11068 2130 11102 2134
rect 10956 2126 10990 2130
rect 11044 2126 11102 2130
rect 10585 2106 10619 2110
rect 10585 2098 10621 2106
rect 10631 2098 10633 2126
rect 10663 2110 10876 2126
rect 10944 2110 11002 2126
rect 11032 2110 11102 2126
rect 11133 2151 11228 2336
rect 11504 2335 11519 2378
rect 11315 2329 11373 2335
rect 11315 2295 11327 2329
rect 11315 2289 11373 2295
rect 11485 2169 11519 2335
rect 11538 2344 11573 2378
rect 11853 2344 11888 2378
rect 11485 2151 11525 2169
rect 11133 2136 11525 2151
rect 11133 2115 11524 2136
rect 11121 2110 11524 2115
rect 10663 2098 11524 2110
rect 10585 2085 10631 2098
rect 10675 2094 11524 2098
rect 10699 2085 11524 2094
rect 10585 2072 11524 2085
rect 11538 2072 11572 2344
rect 11854 2325 11888 2344
rect 11873 2297 11888 2325
rect 11907 2297 11942 2325
rect 12003 2297 12161 2325
rect 11955 2291 12161 2297
rect 12222 2291 12257 2325
rect 11684 2276 11742 2282
rect 11684 2242 11696 2276
rect 11854 2263 11888 2282
rect 11955 2263 12113 2291
rect 11684 2236 11742 2242
rect 11652 2170 11686 2199
rect 11586 2136 11606 2170
rect 11640 2136 11786 2170
rect 11820 2136 11840 2170
rect 11640 2102 11729 2115
rect 11772 2106 11774 2136
rect 11781 2106 11786 2136
rect 11614 2072 11729 2102
rect 11740 2072 11802 2106
rect 7842 2038 7844 2072
rect 7856 2038 7880 2072
rect 3926 2007 6210 2038
rect 6252 2025 6298 2038
rect 6240 2019 6298 2025
rect 6252 2015 6286 2019
rect 6366 2007 6400 2038
rect 6419 2007 6453 2038
rect 6456 2007 6490 2038
rect 6509 2011 6577 2038
rect 6509 2010 6544 2011
rect 6558 2010 6567 2011
rect 6509 2007 6543 2010
rect 3926 2004 6456 2007
rect 3926 1984 6453 2004
rect 6462 1984 6509 2007
rect 6521 1990 6543 2007
rect 6550 1990 6579 2010
rect 6521 1984 6579 1990
rect 3926 1973 6567 1984
rect 3926 1956 6400 1973
rect 6404 1968 6495 1973
rect 6509 1972 6567 1973
rect 3926 1948 6335 1956
rect 6344 1948 6400 1956
rect 3926 1945 6400 1948
rect 6401 1945 6495 1968
rect 3926 1938 6306 1945
rect 6344 1939 6365 1945
rect 6366 1939 6400 1945
rect 6404 1939 6454 1945
rect 3926 1932 6254 1938
rect 3926 1922 6230 1932
rect 6272 1922 6306 1938
rect 3926 1914 6227 1922
rect 6272 1914 6292 1922
rect 6317 1921 6454 1939
rect 6317 1914 6453 1921
rect 6461 1914 6495 1945
rect 3878 1866 3912 1906
rect 3926 1880 6495 1914
rect 6504 1966 6567 1972
rect 6592 1967 6601 2038
rect 6629 2031 6693 2038
rect 6629 2017 6701 2031
rect 6629 1990 6667 2017
rect 6621 1978 6667 1990
rect 6735 1984 7560 2038
rect 7574 2015 7608 2038
rect 7676 2034 7752 2038
rect 7676 2015 7734 2034
rect 7762 2015 7822 2038
rect 7574 2002 7796 2015
rect 7808 2011 7810 2015
rect 7804 2002 7806 2010
rect 7574 2000 7806 2002
rect 6581 1966 6609 1967
rect 6626 1966 6667 1978
rect 6696 1966 6721 1984
rect 6504 1962 6655 1966
rect 6504 1954 6638 1962
rect 6735 1954 7572 1984
rect 6504 1906 7572 1954
rect 3926 1870 6227 1880
rect 6287 1877 6318 1880
rect 6319 1877 6335 1880
rect 6287 1871 6337 1877
rect 6351 1871 6401 1880
rect 6404 1871 6453 1880
rect 6287 1870 6353 1871
rect 6366 1870 6400 1871
rect 3926 1866 6400 1870
rect 3610 1836 6400 1866
rect 6404 1855 6416 1871
rect 6419 1855 6453 1871
rect 6404 1836 6454 1855
rect 3610 1832 6230 1836
rect 2440 1812 2674 1817
rect 2732 1812 3608 1817
rect 2440 1804 3608 1812
rect 3664 1812 3694 1832
rect 3764 1819 3782 1832
rect 3878 1831 3928 1832
rect 3931 1831 6230 1832
rect 3664 1807 3710 1812
rect 2032 1788 2034 1794
rect 1990 1778 2002 1788
rect 2032 1778 2044 1788
rect 2440 1783 3596 1804
rect 3676 1803 3710 1807
rect 3722 1794 3752 1807
rect 3764 1803 3798 1812
rect 3859 1804 6230 1831
rect 6260 1828 6282 1836
rect 6287 1828 6318 1836
rect 6419 1828 6453 1836
rect 6260 1824 6341 1828
rect 6395 1824 6453 1828
rect 6260 1812 6354 1824
rect 6383 1817 6453 1824
rect 6456 1817 6495 1880
rect 6509 1892 7572 1906
rect 6509 1861 6548 1892
rect 6561 1885 6638 1892
rect 6735 1886 7572 1892
rect 6562 1869 6627 1885
rect 6562 1861 6596 1869
rect 6686 1861 7572 1886
rect 6509 1832 7572 1861
rect 7574 1966 7608 2000
rect 7640 1987 7642 1991
rect 7654 1987 7674 1991
rect 7698 1987 7762 2000
rect 7804 1987 7806 2000
rect 7628 1966 7681 1987
rect 7698 1984 7774 1987
rect 7698 1972 7813 1984
rect 7574 1956 7681 1966
rect 7682 1968 7813 1972
rect 7682 1956 7704 1968
rect 7574 1946 7704 1956
rect 7574 1922 7619 1946
rect 7628 1922 7704 1946
rect 7716 1956 7813 1968
rect 7716 1934 7782 1956
rect 7574 1866 7608 1922
rect 7628 1866 7634 1922
rect 7640 1900 7674 1922
rect 7682 1906 7704 1922
rect 7728 1922 7792 1934
rect 7728 1918 7782 1922
rect 7636 1866 7674 1900
rect 7728 1866 7762 1918
rect 7842 1906 7880 2038
rect 7890 2038 11802 2072
rect 11806 2072 11840 2136
rect 11854 2091 11893 2263
rect 11907 2091 11941 2263
rect 12033 2211 12049 2223
rect 12033 2201 12053 2211
rect 12033 2195 12049 2201
rect 12017 2180 12019 2189
rect 12027 2180 12051 2195
rect 12065 2189 12089 2223
rect 12189 2201 12209 2291
rect 12001 2161 12067 2180
rect 12005 2155 12063 2161
rect 12021 2142 12055 2146
rect 12067 2142 12091 2145
rect 12109 2142 12129 2146
rect 12009 2130 12067 2142
rect 12103 2130 12129 2142
rect 12009 2127 12064 2130
rect 11973 2114 11975 2118
rect 11987 2114 12007 2118
rect 11961 2110 12013 2114
rect 12015 2110 12055 2127
rect 11961 2091 12007 2110
rect 12021 2091 12055 2110
rect 12061 2114 12095 2118
rect 12061 2110 12101 2114
rect 12103 2110 12133 2130
rect 12061 2091 12095 2110
rect 12109 2106 12133 2110
rect 12141 2106 12143 2146
rect 12109 2091 12143 2106
rect 12150 2091 12155 2142
rect 12175 2091 12209 2201
rect 12223 2244 12257 2291
rect 12276 2244 12311 2272
rect 12372 2244 12530 2272
rect 13107 2263 13165 2269
rect 12223 2210 12263 2244
rect 12324 2238 12530 2244
rect 12591 2238 12626 2255
rect 12324 2210 12482 2238
rect 12223 2091 12262 2210
rect 12276 2091 12310 2210
rect 12402 2158 12418 2170
rect 12402 2148 12422 2158
rect 12402 2142 12418 2148
rect 12386 2127 12388 2136
rect 12396 2127 12420 2142
rect 12434 2138 12458 2170
rect 12558 2148 12578 2238
rect 12432 2130 12480 2138
rect 12370 2110 12436 2127
rect 12370 2108 12508 2110
rect 12432 2106 12508 2108
rect 11854 2083 12310 2091
rect 12390 2089 12424 2106
rect 12432 2102 12512 2106
rect 12436 2089 12460 2092
rect 12378 2083 12436 2089
rect 12478 2083 12512 2102
rect 11854 2072 12512 2083
rect 12519 2072 12524 2089
rect 12544 2072 12578 2148
rect 12592 2237 12626 2238
rect 12592 2201 12662 2237
rect 13107 2229 13119 2263
rect 13107 2223 13165 2229
rect 12592 2167 12680 2201
rect 12592 2110 12679 2167
rect 13057 2148 13215 2161
rect 13296 2148 13311 2602
rect 13330 2568 13365 2602
rect 13645 2568 13716 2602
rect 13330 2148 13364 2568
rect 13646 2567 13716 2568
rect 13663 2533 13734 2567
rect 14014 2533 14049 2567
rect 13476 2500 13534 2506
rect 13476 2466 13488 2500
rect 13476 2460 13534 2466
rect 13555 2327 13578 2381
rect 13663 2363 13733 2533
rect 14015 2514 14049 2533
rect 17071 2553 17129 2559
rect 17071 2519 17083 2553
rect 13845 2465 13903 2471
rect 13845 2431 13857 2465
rect 13845 2425 13903 2431
rect 13813 2363 13847 2388
rect 13924 2382 13947 2384
rect 14034 2382 14049 2514
rect 14068 2480 14103 2514
rect 14383 2480 14418 2514
rect 17071 2513 17129 2519
rect 14068 2382 14102 2480
rect 14384 2461 14418 2480
rect 14403 2418 14418 2461
rect 14214 2412 14272 2418
rect 14214 2382 14226 2412
rect 13978 2381 14001 2382
rect 13978 2363 14013 2381
rect 13663 2348 14013 2363
rect 14068 2348 14328 2382
rect 13609 2293 13632 2327
rect 13663 2293 14012 2348
rect 13609 2248 13643 2293
rect 13612 2231 13643 2248
rect 13476 2210 13534 2216
rect 13476 2176 13488 2210
rect 13476 2170 13534 2176
rect 13057 2127 13268 2148
rect 12980 2110 12995 2127
rect 13014 2126 13049 2127
rect 13110 2126 13268 2127
rect 13014 2114 13330 2126
rect 13014 2110 13048 2114
rect 13609 2110 13643 2231
rect 13646 2110 14012 2293
rect 12592 2078 14012 2110
rect 14015 2078 14049 2348
rect 14068 2221 14102 2348
rect 14294 2335 14328 2348
rect 14182 2331 14216 2335
rect 14270 2331 14328 2335
rect 14170 2323 14228 2331
rect 14258 2323 14328 2331
rect 14170 2280 14217 2323
rect 14270 2314 14328 2323
rect 14120 2246 14140 2280
rect 14144 2246 14217 2280
rect 14058 2199 14102 2221
rect 14170 2199 14216 2246
rect 14058 2187 14103 2199
rect 14182 2187 14216 2199
rect 14068 2078 14136 2187
rect 14180 2163 14216 2187
rect 14180 2151 14214 2163
rect 14180 2106 14226 2151
rect 14180 2104 14260 2106
rect 12592 2072 14138 2078
rect 14180 2072 14252 2104
rect 14260 2072 14276 2104
rect 14294 2072 14328 2314
rect 14347 2295 14382 2329
rect 14347 2072 14381 2295
rect 14384 2072 14418 2418
rect 14437 2427 14472 2461
rect 14437 2329 14471 2427
rect 15448 2397 15483 2431
rect 15449 2378 15483 2397
rect 14583 2359 14641 2365
rect 14583 2329 14595 2359
rect 14753 2336 14787 2365
rect 14437 2295 14681 2329
rect 14437 2168 14471 2295
rect 14663 2282 14681 2295
rect 14551 2278 14585 2282
rect 14639 2278 14681 2282
rect 14753 2300 14823 2336
rect 14539 2270 14597 2278
rect 14627 2270 14685 2278
rect 14539 2227 14586 2270
rect 14639 2261 14685 2270
rect 14489 2193 14509 2227
rect 14513 2193 14586 2227
rect 14663 2222 14685 2261
rect 14753 2266 14841 2300
rect 14662 2204 14697 2222
rect 14753 2204 14840 2266
rect 14427 2146 14471 2168
rect 14539 2146 14585 2193
rect 14662 2168 14840 2204
rect 14952 2198 15010 2204
rect 14952 2168 14964 2198
rect 14427 2134 14472 2146
rect 14551 2134 14585 2146
rect 14437 2072 14505 2134
rect 14549 2110 14585 2134
rect 14663 2134 15066 2168
rect 14663 2126 14840 2134
rect 15032 2130 15066 2134
rect 14920 2126 14954 2130
rect 15008 2126 15066 2130
rect 14549 2106 14583 2110
rect 14549 2098 14585 2106
rect 14595 2098 14597 2126
rect 14627 2110 14840 2126
rect 14908 2110 14966 2126
rect 14996 2110 15066 2126
rect 15097 2151 15192 2336
rect 15468 2335 15483 2378
rect 15279 2329 15337 2335
rect 15279 2295 15291 2329
rect 15279 2289 15337 2295
rect 15449 2169 15483 2335
rect 15502 2344 15537 2378
rect 15817 2344 15852 2378
rect 15449 2151 15489 2169
rect 15097 2136 15489 2151
rect 15097 2115 15488 2136
rect 15085 2110 15488 2115
rect 14627 2098 15488 2110
rect 14549 2085 14595 2098
rect 14639 2094 15488 2098
rect 14663 2085 15488 2094
rect 14549 2072 15488 2085
rect 15502 2072 15536 2344
rect 15818 2325 15852 2344
rect 15837 2297 15852 2325
rect 15871 2297 15906 2325
rect 15967 2297 16125 2325
rect 15919 2291 16125 2297
rect 16186 2291 16221 2325
rect 15648 2276 15706 2282
rect 15648 2242 15660 2276
rect 15818 2263 15852 2282
rect 15919 2263 16077 2291
rect 15648 2236 15706 2242
rect 15616 2170 15650 2199
rect 15550 2136 15570 2170
rect 15604 2136 15750 2170
rect 15784 2136 15804 2170
rect 15604 2102 15693 2115
rect 15736 2106 15738 2136
rect 15745 2106 15750 2136
rect 15578 2072 15693 2102
rect 15704 2072 15766 2106
rect 11806 2038 11808 2072
rect 11820 2038 11844 2072
rect 7890 2007 10174 2038
rect 10216 2025 10262 2038
rect 10204 2019 10262 2025
rect 10216 2015 10250 2019
rect 10330 2007 10364 2038
rect 10383 2007 10417 2038
rect 10420 2007 10454 2038
rect 10473 2011 10541 2038
rect 10473 2010 10508 2011
rect 10522 2010 10531 2011
rect 10473 2007 10507 2010
rect 7890 2004 10420 2007
rect 7890 1984 10417 2004
rect 10426 1984 10473 2007
rect 10485 1990 10507 2007
rect 10514 1990 10543 2010
rect 10485 1984 10543 1990
rect 7890 1973 10531 1984
rect 7890 1956 10364 1973
rect 7890 1945 10282 1956
rect 7890 1938 10256 1945
rect 10270 1939 10282 1945
rect 10308 1945 10364 1956
rect 10308 1939 10329 1945
rect 10330 1939 10364 1945
rect 10368 1945 10459 1973
rect 10473 1972 10531 1973
rect 10368 1939 10418 1945
rect 7890 1932 10218 1938
rect 7890 1922 10194 1932
rect 7842 1866 7876 1906
rect 7890 1870 10191 1922
rect 10236 1911 10256 1938
rect 10265 1921 10418 1939
rect 10265 1911 10417 1921
rect 10236 1906 10417 1911
rect 10267 1893 10282 1906
rect 10330 1905 10364 1906
rect 10251 1877 10282 1893
rect 10283 1877 10365 1905
rect 10251 1872 10365 1877
rect 10251 1871 10301 1872
rect 10315 1871 10365 1872
rect 10368 1871 10417 1906
rect 10251 1870 10317 1871
rect 10330 1870 10364 1871
rect 7890 1866 10364 1870
rect 7574 1836 10364 1866
rect 10368 1855 10380 1871
rect 10383 1855 10417 1871
rect 10368 1836 10418 1855
rect 7574 1832 10194 1836
rect 6509 1827 7560 1832
rect 6509 1817 6548 1827
rect 6562 1817 6596 1827
rect 6625 1824 6638 1827
rect 6688 1824 7560 1827
rect 6656 1817 7560 1824
rect 6260 1804 6366 1812
rect 6383 1811 7560 1817
rect 3859 1797 6227 1804
rect 6282 1800 6366 1804
rect 1984 1774 2012 1778
rect 2022 1774 2050 1778
rect 1984 1763 2050 1774
rect 2086 1771 2159 1782
rect 2208 1779 2354 1782
rect 2191 1778 2221 1779
rect 2086 1763 2148 1771
rect 1681 1759 2148 1763
rect 2190 1759 2222 1778
rect 2255 1771 2307 1779
rect 2369 1778 2436 1782
rect 2440 1778 2490 1783
rect 2788 1778 3596 1783
rect 3686 1791 3788 1794
rect 3686 1778 3801 1791
rect 3859 1778 3928 1797
rect 3931 1782 6227 1797
rect 6259 1796 6261 1800
rect 6271 1796 6381 1800
rect 6247 1782 6387 1796
rect 6389 1783 7560 1811
rect 7628 1822 7634 1832
rect 7628 1807 7649 1822
rect 7728 1819 7746 1832
rect 7842 1831 7892 1832
rect 7895 1831 10194 1832
rect 7686 1794 7716 1807
rect 6389 1782 6419 1783
rect 3931 1778 6419 1782
rect 6422 1778 6429 1783
rect 6456 1778 6495 1783
rect 6509 1778 6548 1783
rect 6562 1778 6596 1783
rect 6620 1778 6638 1783
rect 6752 1778 7560 1783
rect 2369 1771 3596 1778
rect 2266 1759 2296 1771
rect 2380 1759 2414 1771
rect 1670 1754 2159 1759
rect 2190 1754 2233 1759
rect 1670 1748 2233 1754
rect 2255 1748 2307 1759
rect 2369 1748 2414 1759
rect 1670 1736 2120 1748
rect 2190 1744 2201 1748
rect 2211 1744 2232 1748
rect 2221 1738 2232 1744
rect 2191 1736 2232 1738
rect 1670 1727 2250 1736
rect 1681 1700 2250 1727
rect 2296 1710 2298 1716
rect 2254 1700 2266 1710
rect 2296 1700 2308 1710
rect 1640 1637 1649 1678
rect 1668 1637 1677 1700
rect 1681 1684 2314 1700
rect 2402 1686 2414 1748
rect 2415 1744 3596 1771
rect 2415 1686 2436 1744
rect 1681 1666 2308 1684
rect 1681 1660 2278 1666
rect 2294 1660 2308 1666
rect 1681 1656 2308 1660
rect 1681 1650 2298 1656
rect 1681 1640 2294 1650
rect 1681 1637 2263 1640
rect 1318 1618 2263 1637
rect 2276 1630 2294 1640
rect 1228 1604 1241 1617
rect 1126 1570 1206 1576
rect 1126 1538 1160 1570
rect 1206 1538 1210 1570
rect 1228 1551 1244 1604
rect 1240 1547 1244 1551
rect 1318 1586 2250 1618
rect 1318 1576 1918 1586
rect 2010 1582 2022 1586
rect 2033 1582 2250 1586
rect 1318 1557 1932 1576
rect 2006 1564 2250 1582
rect 2010 1558 2250 1564
rect 1318 1553 1952 1557
rect 1318 1548 1959 1553
rect 2033 1548 2250 1558
rect 1126 1536 1210 1538
rect 1318 1542 1965 1548
rect 1972 1542 2250 1548
rect 1318 1541 2250 1542
rect 1126 1530 1206 1536
rect 1126 1511 1160 1530
rect 1318 1526 1965 1541
rect 1972 1531 2250 1541
rect 2276 1584 2311 1599
rect 2276 1531 2296 1584
rect 2402 1531 2436 1686
rect 2440 1729 2490 1744
rect 2788 1729 3596 1744
rect 2440 1710 3596 1729
rect 2440 1695 2674 1710
rect 2440 1655 2490 1695
rect 2788 1694 3596 1710
rect 2440 1624 2577 1655
rect 2647 1643 2674 1674
rect 2616 1633 2674 1643
rect 2601 1624 2674 1633
rect 2455 1618 2489 1624
rect 2528 1618 2530 1624
rect 2455 1608 2498 1618
rect 2528 1608 2540 1618
rect 2455 1592 2546 1608
rect 2601 1593 2613 1624
rect 2616 1593 2663 1624
rect 2790 1622 2805 1694
rect 3056 1676 3066 1694
rect 3076 1690 3104 1694
rect 3078 1684 3104 1690
rect 3078 1676 3098 1684
rect 3056 1666 3098 1676
rect 3072 1656 3098 1666
rect 3157 1658 3596 1694
rect 3610 1769 6419 1778
rect 3610 1767 3681 1769
rect 3610 1755 3670 1767
rect 3610 1744 3681 1755
rect 3682 1748 6419 1769
rect 3682 1744 6299 1748
rect 3610 1658 3644 1744
rect 3704 1726 3801 1744
rect 3704 1720 3766 1726
rect 3704 1710 3752 1720
rect 3802 1692 3849 1723
rect 3782 1682 3849 1692
rect 3756 1658 3849 1682
rect 3859 1658 3912 1744
rect 3925 1725 6227 1744
rect 6247 1731 6299 1744
rect 3072 1650 3088 1656
rect 3157 1655 3681 1658
rect 3157 1642 3591 1655
rect 3610 1649 3681 1655
rect 3694 1649 3912 1658
rect 3610 1642 3912 1649
rect 3157 1641 3912 1642
rect 2771 1604 2805 1622
rect 2455 1531 2489 1592
rect 2496 1584 2540 1592
rect 2601 1587 2659 1593
rect 2496 1574 2725 1584
rect 2771 1574 3210 1604
rect 2528 1564 2542 1574
rect 2771 1568 2841 1574
rect 2528 1558 2530 1564
rect 2535 1562 2542 1564
rect 2569 1546 2603 1550
rect 2563 1540 2615 1546
rect 2657 1540 2691 1550
rect 2788 1540 3174 1568
rect 3205 1551 3210 1574
rect 3241 1551 3275 1641
rect 3355 1636 3370 1641
rect 3385 1636 3401 1641
rect 3389 1633 3401 1636
rect 3400 1551 3401 1633
rect 3431 1636 3449 1641
rect 3431 1633 3443 1636
rect 3431 1551 3434 1633
rect 3557 1624 3912 1641
rect 3926 1710 6227 1725
rect 3926 1700 6230 1710
rect 6242 1700 6299 1731
rect 3926 1646 6299 1700
rect 3557 1608 3591 1624
rect 3610 1608 3644 1624
rect 3796 1608 3800 1624
rect 3840 1616 3842 1624
rect 3828 1608 3842 1616
rect 3859 1608 3893 1624
rect 3557 1606 3893 1608
rect 3557 1590 3872 1606
rect 3557 1574 3724 1590
rect 3737 1580 3812 1590
rect 3752 1574 3812 1580
rect 3838 1574 3872 1590
rect 3892 1574 3893 1606
rect 3557 1570 3591 1574
rect 3610 1570 3644 1574
rect 3752 1570 3770 1574
rect 3825 1570 3858 1574
rect 3859 1570 3893 1574
rect 3926 1621 6227 1646
rect 6240 1630 6299 1646
rect 3557 1551 3912 1570
rect 3205 1540 3912 1551
rect 2563 1534 2570 1540
rect 2571 1531 2615 1540
rect 1972 1530 2495 1531
rect 2002 1526 2495 1530
rect 1318 1514 2495 1526
rect 1126 1510 1184 1511
rect 1318 1510 1898 1514
rect 1907 1510 1918 1514
rect 1919 1510 1959 1514
rect 1966 1510 2024 1514
rect 2033 1510 2495 1514
rect 1120 1506 1234 1510
rect 1318 1506 2495 1510
rect 2586 1506 2615 1531
rect 2788 1534 2869 1540
rect 2893 1534 2949 1540
rect 3045 1534 3097 1540
rect 2788 1510 2858 1534
rect 2924 1510 2938 1524
rect 3056 1510 3074 1524
rect 3170 1510 3174 1540
rect 3194 1515 3591 1540
rect 3193 1510 3591 1515
rect 2788 1506 3591 1510
rect 3610 1536 3681 1540
rect 3712 1536 3912 1540
rect 1116 1502 1238 1506
rect 1284 1504 2495 1506
rect 1116 1472 1184 1502
rect 1204 1472 1238 1502
rect 1268 1472 1272 1504
rect 1284 1472 1297 1504
rect 1318 1478 2495 1504
rect 2569 1478 2615 1506
rect 2657 1478 2691 1506
rect 2771 1484 3596 1506
rect 3610 1484 3644 1536
rect 3662 1484 3670 1526
rect 3752 1506 3858 1536
rect 3859 1506 3912 1536
rect 3752 1502 3770 1506
rect 3686 1484 3788 1502
rect 2771 1478 3788 1484
rect 1318 1472 3788 1478
rect 3812 1484 3912 1506
rect 3926 1557 6232 1621
rect 6242 1616 6299 1630
rect 6300 1744 6419 1748
rect 6429 1776 7560 1778
rect 7658 1776 7716 1794
rect 6429 1766 7716 1776
rect 7718 1766 7765 1807
rect 6429 1749 7765 1766
rect 6429 1744 6628 1749
rect 6300 1644 6341 1744
rect 6344 1735 6419 1744
rect 6242 1599 6293 1616
rect 3926 1531 6227 1557
rect 6240 1538 6293 1599
rect 6300 1551 6304 1644
rect 6307 1640 6341 1644
rect 6342 1729 6419 1735
rect 6422 1729 6429 1744
rect 6456 1729 6495 1744
rect 6509 1729 6548 1744
rect 6562 1729 6596 1744
rect 6628 1731 6630 1744
rect 6636 1743 6638 1749
rect 6640 1743 6655 1747
rect 6664 1744 6735 1749
rect 6750 1744 7765 1749
rect 6664 1743 6750 1744
rect 6752 1743 7765 1744
rect 6636 1731 7765 1743
rect 6628 1729 7765 1731
rect 6342 1726 7765 1729
rect 7823 1804 10194 1831
rect 10224 1828 10282 1836
rect 10383 1828 10417 1836
rect 10224 1827 10305 1828
rect 10224 1804 10259 1827
rect 10269 1824 10305 1827
rect 10308 1824 10341 1827
rect 10359 1824 10417 1828
rect 10265 1809 10317 1824
rect 10347 1817 10417 1824
rect 10425 1817 10459 1945
rect 10468 1966 10531 1972
rect 10556 1967 10565 2038
rect 10593 2031 10657 2038
rect 10593 2017 10665 2031
rect 10593 1990 10631 2017
rect 10585 1978 10631 1990
rect 10699 1984 11524 2038
rect 11538 2015 11572 2038
rect 11640 2034 11716 2038
rect 11640 2015 11698 2034
rect 11726 2015 11786 2038
rect 11538 2002 11760 2015
rect 11772 2011 11774 2015
rect 11768 2002 11770 2010
rect 11538 2000 11770 2002
rect 10545 1966 10573 1967
rect 10590 1966 10631 1978
rect 10660 1966 10685 1984
rect 10468 1962 10619 1966
rect 10468 1954 10602 1962
rect 10699 1954 11536 1984
rect 10468 1906 11536 1954
rect 10473 1892 11536 1906
rect 10473 1817 10512 1892
rect 10525 1885 10602 1892
rect 10526 1869 10591 1885
rect 10699 1871 11536 1892
rect 10526 1817 10560 1869
rect 10589 1825 10602 1869
rect 10668 1855 11536 1871
rect 10660 1852 11536 1855
rect 10574 1817 10602 1825
rect 10652 1832 11536 1852
rect 11538 1966 11572 2000
rect 11604 1987 11606 1991
rect 11618 1987 11638 1991
rect 11662 1987 11726 2000
rect 11768 1987 11770 2000
rect 11592 1966 11645 1987
rect 11662 1984 11738 1987
rect 11662 1972 11777 1984
rect 11538 1956 11645 1966
rect 11646 1968 11777 1972
rect 11646 1956 11668 1968
rect 11538 1946 11668 1956
rect 11538 1922 11583 1946
rect 11592 1922 11668 1946
rect 11680 1956 11777 1968
rect 11680 1934 11746 1956
rect 11538 1866 11572 1922
rect 11592 1866 11598 1922
rect 11604 1900 11638 1922
rect 11646 1906 11668 1922
rect 11692 1922 11756 1934
rect 11692 1918 11746 1922
rect 11600 1866 11638 1900
rect 11692 1866 11726 1918
rect 11806 1906 11844 2038
rect 11854 2038 15766 2072
rect 15770 2072 15804 2136
rect 15770 2038 15772 2072
rect 15784 2038 15808 2072
rect 11854 2007 14138 2038
rect 14180 2025 14226 2038
rect 14168 2019 14226 2025
rect 14180 2015 14214 2019
rect 14294 2007 14328 2038
rect 14347 2007 14381 2038
rect 14384 2007 14418 2038
rect 14437 2011 14505 2038
rect 14437 2010 14472 2011
rect 14486 2010 14495 2011
rect 14437 2007 14471 2010
rect 11854 2004 14384 2007
rect 11854 1984 14381 2004
rect 14390 1984 14437 2007
rect 14449 1990 14471 2007
rect 14478 1990 14507 2010
rect 14449 1984 14507 1990
rect 11854 1973 14495 1984
rect 11854 1956 14328 1973
rect 11854 1945 14246 1956
rect 11854 1938 14220 1945
rect 14234 1939 14246 1945
rect 14272 1945 14328 1956
rect 14272 1939 14293 1945
rect 14294 1939 14328 1945
rect 14332 1945 14423 1973
rect 14437 1972 14495 1973
rect 14332 1939 14382 1945
rect 11854 1932 14182 1938
rect 11854 1922 14158 1932
rect 11806 1866 11840 1906
rect 11854 1870 14155 1922
rect 14200 1911 14220 1938
rect 14229 1921 14382 1939
rect 14229 1911 14381 1921
rect 14200 1906 14381 1911
rect 14231 1893 14246 1906
rect 14294 1905 14328 1906
rect 14215 1877 14246 1893
rect 14247 1877 14329 1905
rect 14215 1872 14329 1877
rect 14215 1871 14265 1872
rect 14279 1871 14329 1872
rect 14332 1871 14381 1906
rect 14215 1870 14281 1871
rect 14294 1870 14328 1871
rect 11854 1866 14328 1870
rect 11538 1836 14328 1866
rect 14332 1855 14344 1871
rect 14347 1855 14381 1871
rect 14332 1836 14382 1855
rect 11538 1832 14158 1836
rect 10652 1824 11524 1832
rect 10636 1817 11524 1824
rect 10347 1811 11524 1817
rect 7823 1798 10191 1804
rect 6342 1720 7730 1726
rect 6342 1710 7716 1720
rect 6342 1695 7704 1710
rect 6342 1656 6453 1695
rect 6342 1644 6415 1656
rect 6419 1644 6453 1656
rect 6342 1613 6400 1644
rect 6404 1642 6454 1644
rect 6456 1642 6495 1695
rect 6509 1661 6548 1695
rect 6562 1661 6596 1695
rect 6628 1674 6668 1695
rect 6509 1643 6596 1661
rect 6611 1643 6668 1674
rect 6509 1642 6668 1643
rect 6404 1627 6668 1642
rect 6404 1624 6548 1627
rect 6335 1597 6400 1613
rect 6419 1608 6548 1624
rect 6561 1608 6668 1627
rect 6335 1563 6401 1597
rect 6335 1551 6400 1563
rect 6300 1540 6305 1551
rect 6332 1540 6400 1551
rect 6419 1540 6453 1608
rect 6300 1538 6453 1540
rect 6240 1531 6453 1538
rect 6456 1584 6548 1608
rect 6562 1593 6668 1608
rect 6562 1584 6596 1593
rect 6611 1584 6668 1593
rect 6456 1574 6668 1584
rect 6456 1531 6495 1574
rect 6499 1568 6506 1574
rect 6509 1568 6548 1574
rect 6499 1550 6548 1568
rect 6562 1568 6596 1574
rect 6562 1550 6601 1568
rect 6499 1534 6601 1550
rect 6611 1563 6668 1574
rect 6669 1603 6710 1695
rect 6716 1694 7704 1695
rect 6716 1666 6788 1694
rect 6711 1622 6788 1666
rect 6791 1622 6798 1666
rect 6800 1622 6810 1694
rect 6711 1604 6810 1622
rect 6825 1658 7704 1694
rect 7823 1658 7892 1798
rect 6825 1624 7892 1658
rect 7895 1782 10191 1798
rect 10223 1796 10257 1800
rect 10211 1782 10263 1796
rect 10265 1782 10305 1809
rect 10308 1800 10317 1809
rect 10308 1796 10345 1800
rect 10308 1782 10351 1796
rect 10353 1783 11524 1811
rect 11592 1822 11598 1832
rect 11592 1807 11613 1822
rect 11692 1819 11710 1832
rect 11806 1831 11856 1832
rect 11859 1831 14158 1832
rect 11650 1794 11680 1807
rect 10353 1782 10383 1783
rect 7895 1748 10383 1782
rect 10391 1778 10393 1783
rect 10425 1778 10459 1783
rect 10473 1778 10512 1783
rect 10526 1778 10560 1783
rect 10574 1778 10602 1783
rect 10716 1778 11524 1783
rect 7895 1710 10191 1748
rect 7895 1700 10194 1710
rect 10211 1700 10263 1748
rect 7895 1646 10263 1700
rect 6825 1608 7686 1624
rect 7792 1608 7804 1616
rect 7823 1608 7857 1624
rect 6825 1604 7857 1608
rect 6669 1591 6696 1603
rect 6669 1578 6673 1591
rect 6711 1590 7857 1604
rect 6711 1586 7686 1590
rect 7802 1587 7812 1590
rect 7823 1587 7857 1590
rect 7895 1621 10191 1646
rect 10204 1630 10222 1646
rect 10223 1630 10263 1646
rect 10265 1644 10305 1748
rect 10271 1640 10305 1644
rect 10308 1729 10383 1748
rect 10393 1776 11524 1778
rect 11622 1776 11680 1794
rect 10393 1766 11680 1776
rect 11682 1766 11729 1807
rect 10393 1749 11729 1766
rect 10393 1744 10592 1749
rect 10626 1744 10680 1749
rect 10714 1744 11729 1749
rect 10391 1729 10393 1744
rect 10425 1729 10459 1744
rect 10473 1729 10512 1744
rect 10526 1729 10560 1744
rect 10592 1729 10594 1744
rect 10606 1743 10626 1744
rect 10628 1743 10674 1744
rect 10606 1731 10632 1743
rect 10602 1729 10632 1731
rect 10634 1729 10674 1743
rect 10680 1743 10714 1744
rect 10716 1743 11729 1744
rect 10680 1729 11729 1743
rect 10308 1726 11729 1729
rect 11787 1804 14158 1831
rect 14188 1828 14246 1836
rect 14347 1828 14381 1836
rect 14188 1827 14269 1828
rect 14188 1804 14223 1827
rect 14233 1824 14269 1827
rect 14272 1824 14305 1827
rect 14323 1824 14381 1828
rect 14229 1809 14281 1824
rect 14311 1817 14381 1824
rect 14389 1817 14423 1945
rect 14432 1966 14495 1972
rect 14520 1967 14529 2038
rect 14557 2031 14621 2038
rect 14557 2017 14629 2031
rect 14557 1990 14595 2017
rect 14549 1978 14595 1990
rect 14663 1984 15488 2038
rect 15502 2015 15536 2038
rect 15604 2034 15680 2038
rect 15604 2015 15662 2034
rect 15690 2015 15750 2038
rect 15502 2002 15724 2015
rect 15736 2011 15738 2015
rect 15732 2002 15734 2010
rect 15502 2000 15734 2002
rect 14509 1966 14537 1967
rect 14554 1966 14595 1978
rect 14624 1966 14649 1984
rect 14432 1962 14583 1966
rect 14432 1954 14566 1962
rect 14663 1954 15500 1984
rect 14432 1906 15500 1954
rect 14437 1892 15500 1906
rect 14437 1817 14476 1892
rect 14489 1885 14566 1892
rect 14490 1869 14555 1885
rect 14663 1871 15500 1892
rect 14490 1817 14524 1869
rect 14553 1825 14566 1869
rect 14632 1855 15500 1871
rect 14624 1852 15500 1855
rect 14538 1817 14566 1825
rect 14616 1832 15500 1852
rect 15502 1966 15536 2000
rect 15568 1987 15570 1991
rect 15582 1987 15602 1991
rect 15626 1987 15690 2000
rect 15732 1987 15734 2000
rect 15556 1966 15609 1987
rect 15626 1984 15702 1987
rect 15626 1972 15741 1984
rect 15502 1956 15609 1966
rect 15610 1968 15741 1972
rect 15610 1956 15632 1968
rect 15502 1946 15632 1956
rect 15502 1922 15547 1946
rect 15556 1922 15632 1946
rect 15644 1956 15741 1968
rect 15644 1934 15710 1956
rect 15502 1866 15536 1922
rect 15556 1866 15562 1922
rect 15568 1900 15602 1922
rect 15610 1906 15632 1922
rect 15656 1922 15720 1934
rect 15656 1918 15710 1922
rect 15564 1866 15602 1900
rect 15656 1866 15690 1918
rect 15770 1906 15808 2038
rect 15770 1866 15804 1906
rect 15818 1866 15857 2263
rect 15502 1832 15820 1866
rect 14616 1824 15488 1832
rect 14600 1817 15488 1824
rect 14311 1811 15488 1817
rect 11787 1798 14155 1804
rect 10308 1720 11694 1726
rect 10308 1710 11680 1720
rect 10308 1695 11668 1710
rect 10308 1656 10417 1695
rect 10308 1644 10379 1656
rect 10383 1655 10417 1656
rect 10425 1655 10459 1695
rect 10473 1661 10512 1695
rect 10526 1661 10560 1695
rect 10592 1674 10632 1695
rect 10383 1644 10472 1655
rect 10308 1631 10364 1644
rect 6711 1585 6965 1586
rect 7033 1585 7104 1586
rect 7134 1585 7168 1586
rect 7169 1585 7179 1586
rect 7194 1585 7228 1586
rect 6711 1578 7228 1585
rect 6669 1574 7228 1578
rect 6611 1546 6662 1563
rect 6621 1540 6662 1546
rect 6623 1534 6662 1540
rect 3926 1529 6495 1531
rect 6509 1529 6601 1534
rect 3926 1506 6601 1529
rect 3926 1495 6495 1506
rect 6509 1504 6601 1506
rect 6509 1495 6596 1504
rect 3926 1491 6596 1495
rect 3926 1484 3966 1491
rect 3812 1472 3966 1484
rect -17 1470 1250 1472
rect 1257 1470 3966 1472
rect -17 1468 3966 1470
rect 3973 1480 4127 1491
rect 3973 1472 4013 1480
rect 4023 1472 4088 1480
rect 4093 1472 4127 1480
rect 4133 1472 4167 1491
rect 4175 1472 4227 1491
rect 4228 1472 4281 1491
rect 4295 1478 6596 1491
rect 6621 1485 6662 1534
rect 6669 1498 6673 1574
rect 6711 1560 7233 1574
rect 6704 1551 7233 1560
rect 6704 1540 7179 1551
rect 7194 1540 7233 1551
rect 6704 1534 7233 1540
rect 6704 1510 6965 1534
rect 7033 1530 7091 1534
rect 7104 1530 7233 1534
rect 6992 1526 7026 1530
rect 7033 1529 7233 1530
rect 7247 1532 7281 1586
rect 7045 1526 7079 1529
rect 7080 1526 7138 1529
rect 6980 1510 7038 1526
rect 7045 1525 7138 1526
rect 7158 1525 7228 1529
rect 7055 1517 7228 1525
rect 7055 1515 7178 1517
rect 7194 1515 7228 1517
rect 7247 1526 7293 1532
rect 7300 1526 7334 1586
rect 7380 1574 7686 1586
rect 7705 1576 7757 1587
rect 7490 1570 7686 1574
rect 7716 1574 7746 1576
rect 7802 1574 7875 1587
rect 7716 1570 7875 1574
rect 7402 1532 7413 1566
rect 7414 1540 7448 1570
rect 7490 1553 7875 1570
rect 7895 1557 10196 1621
rect 10211 1616 10263 1630
rect 10211 1599 10257 1616
rect 7490 1540 7780 1553
rect 7804 1547 7857 1553
rect 7490 1532 7686 1540
rect 7348 1526 7686 1532
rect 7247 1515 7686 1526
rect 7055 1510 7228 1515
rect 7233 1510 7686 1515
rect 6704 1502 7686 1510
rect 7716 1536 7761 1540
rect 7793 1536 7857 1547
rect 7716 1519 7760 1536
rect 7716 1506 7766 1519
rect 7823 1506 7857 1536
rect 7721 1502 7760 1506
rect 6669 1485 6674 1498
rect 6704 1496 7760 1502
rect 7779 1501 7857 1506
rect 6704 1494 7752 1496
rect 6621 1478 6678 1485
rect 6716 1484 7752 1494
rect 7763 1485 7857 1501
rect 7763 1484 7800 1485
rect 7813 1484 7857 1485
rect 6716 1478 7800 1484
rect 4295 1472 7800 1478
rect 7804 1474 7857 1484
rect 7861 1484 7876 1553
rect 7895 1531 10191 1557
rect 10204 1531 10257 1599
rect 10281 1597 10364 1631
rect 10368 1642 10472 1644
rect 10473 1643 10560 1661
rect 10575 1643 10632 1674
rect 10473 1642 10632 1643
rect 10368 1627 10632 1642
rect 10368 1624 10512 1627
rect 10383 1620 10417 1624
rect 10425 1620 10512 1624
rect 10299 1563 10365 1597
rect 10383 1592 10512 1620
rect 10525 1608 10632 1627
rect 10299 1547 10364 1563
rect 10308 1540 10364 1547
rect 10383 1540 10417 1592
rect 10424 1584 10512 1592
rect 10526 1593 10632 1608
rect 10526 1584 10560 1593
rect 10580 1584 10591 1593
rect 10592 1584 10632 1593
rect 10634 1603 10674 1695
rect 10680 1694 11668 1695
rect 10680 1622 10752 1694
rect 10760 1622 10762 1666
rect 10769 1622 10774 1694
rect 10680 1604 10774 1622
rect 10794 1621 10828 1694
rect 10842 1658 11668 1694
rect 11787 1658 11856 1798
rect 10842 1624 11856 1658
rect 11859 1782 14155 1798
rect 14187 1796 14221 1800
rect 14175 1782 14227 1796
rect 14229 1782 14269 1809
rect 14272 1800 14281 1809
rect 14272 1796 14309 1800
rect 14272 1782 14315 1796
rect 14317 1783 15488 1811
rect 15556 1822 15562 1832
rect 15556 1807 15577 1822
rect 15656 1819 15674 1832
rect 15614 1794 15644 1807
rect 14317 1782 14347 1783
rect 11859 1748 14347 1782
rect 14355 1778 14357 1783
rect 14389 1778 14423 1783
rect 14437 1778 14476 1783
rect 14490 1778 14524 1783
rect 14538 1778 14566 1783
rect 14680 1778 15488 1783
rect 11859 1710 14155 1748
rect 11859 1700 14158 1710
rect 14175 1700 14227 1748
rect 11859 1646 14227 1700
rect 10842 1621 11650 1624
rect 10794 1608 11650 1621
rect 11756 1608 11768 1616
rect 11787 1608 11821 1624
rect 10794 1604 11821 1608
rect 10634 1591 10660 1603
rect 10424 1574 10632 1584
rect 10680 1590 11821 1604
rect 10680 1586 11650 1590
rect 11766 1587 11776 1590
rect 11787 1587 11821 1590
rect 11859 1621 14155 1646
rect 14168 1630 14186 1646
rect 14187 1630 14227 1646
rect 14229 1644 14269 1748
rect 14235 1640 14269 1644
rect 14272 1729 14347 1748
rect 14357 1776 15488 1778
rect 15586 1776 15644 1794
rect 14357 1766 15644 1776
rect 15646 1766 15693 1807
rect 14357 1749 15693 1766
rect 14357 1744 14556 1749
rect 14590 1744 14644 1749
rect 14678 1744 15693 1749
rect 14355 1729 14357 1744
rect 14389 1729 14423 1744
rect 14437 1729 14476 1744
rect 14490 1729 14524 1744
rect 14556 1729 14558 1744
rect 14570 1743 14590 1744
rect 14592 1743 14638 1744
rect 14570 1731 14596 1743
rect 14566 1729 14596 1731
rect 14598 1729 14638 1743
rect 14644 1743 14678 1744
rect 14680 1743 15693 1744
rect 14644 1729 15693 1743
rect 14272 1726 15693 1729
rect 14272 1720 15658 1726
rect 14272 1710 15644 1720
rect 14272 1695 15632 1710
rect 14272 1656 14381 1695
rect 14272 1644 14343 1656
rect 14347 1655 14381 1656
rect 14389 1655 14423 1695
rect 14437 1661 14476 1695
rect 14490 1661 14524 1695
rect 14556 1674 14596 1695
rect 14347 1644 14436 1655
rect 14272 1631 14328 1644
rect 10680 1585 10929 1586
rect 10997 1585 11014 1586
rect 11098 1585 11132 1586
rect 10680 1578 11179 1585
rect 10634 1575 11179 1578
rect 10634 1574 10929 1575
rect 10265 1531 10417 1540
rect 7895 1529 10423 1531
rect 10425 1529 10459 1574
rect 10463 1568 10470 1574
rect 10473 1568 10512 1574
rect 10463 1550 10512 1568
rect 10526 1568 10560 1574
rect 10526 1550 10565 1568
rect 10463 1534 10565 1550
rect 10580 1563 10632 1574
rect 10650 1568 10929 1574
rect 10943 1574 11179 1575
rect 10943 1568 11197 1574
rect 10650 1565 11197 1568
rect 10580 1562 10626 1563
rect 10580 1550 10588 1562
rect 10592 1550 10626 1562
rect 10580 1546 10626 1550
rect 10585 1540 10626 1546
rect 10650 1560 10680 1565
rect 10686 1560 11197 1565
rect 10650 1551 11197 1560
rect 10650 1544 11143 1551
rect 10592 1534 10626 1540
rect 10473 1529 10565 1534
rect 7895 1506 10565 1529
rect 7895 1495 10423 1506
rect 10425 1495 10459 1506
rect 10473 1504 10565 1506
rect 10473 1495 10560 1504
rect 7895 1491 10473 1495
rect 7895 1484 7930 1491
rect 7937 1484 7971 1491
rect 7861 1474 7971 1484
rect 7804 1472 7971 1474
rect 7976 1480 8059 1491
rect 7976 1472 8052 1480
rect 8097 1472 8131 1491
rect 8139 1472 8173 1491
rect 8192 1472 8245 1491
rect 8264 1478 10473 1491
rect 10478 1478 10560 1495
rect 10585 1478 10626 1534
rect 10668 1540 11143 1544
rect 11163 1540 11197 1551
rect 10668 1534 11197 1540
rect 10668 1510 10929 1534
rect 10997 1529 11049 1534
rect 11068 1529 11197 1534
rect 11211 1532 11245 1586
rect 10995 1524 11014 1529
rect 11034 1525 11043 1529
rect 10984 1510 11014 1524
rect 11055 1510 11056 1529
rect 11068 1525 11102 1529
rect 11122 1525 11179 1529
rect 11068 1517 11179 1525
rect 11068 1515 11142 1517
rect 11163 1515 11179 1517
rect 11211 1526 11257 1532
rect 11264 1526 11298 1586
rect 11344 1574 11650 1586
rect 11669 1576 11721 1587
rect 11454 1570 11650 1574
rect 11680 1574 11710 1576
rect 11766 1574 11839 1587
rect 11680 1570 11839 1574
rect 11366 1532 11377 1566
rect 11378 1540 11412 1570
rect 11454 1553 11839 1570
rect 11859 1557 14160 1621
rect 14175 1616 14227 1630
rect 14175 1599 14221 1616
rect 11454 1540 11744 1553
rect 11768 1547 11821 1553
rect 11454 1532 11650 1540
rect 11312 1526 11650 1532
rect 11211 1515 11650 1526
rect 11068 1510 11179 1515
rect 11197 1510 11650 1515
rect 10668 1502 11650 1510
rect 11680 1536 11725 1540
rect 11757 1536 11821 1547
rect 11680 1519 11724 1536
rect 11680 1506 11730 1519
rect 11787 1506 11821 1536
rect 11685 1502 11724 1506
rect 10668 1496 11724 1502
rect 11743 1501 11821 1506
rect 10668 1494 11716 1496
rect 10680 1484 11716 1494
rect 11727 1485 11821 1501
rect 11727 1484 11764 1485
rect 11777 1484 11821 1485
rect 10680 1478 11764 1484
rect 8264 1472 11764 1478
rect 11768 1474 11821 1484
rect 11825 1484 11840 1553
rect 11859 1531 14155 1557
rect 14168 1531 14221 1599
rect 14245 1597 14328 1631
rect 14332 1642 14436 1644
rect 14437 1643 14524 1661
rect 14539 1643 14596 1674
rect 14437 1642 14596 1643
rect 14332 1627 14596 1642
rect 14332 1624 14476 1627
rect 14347 1620 14381 1624
rect 14389 1620 14476 1624
rect 14263 1563 14329 1597
rect 14347 1592 14476 1620
rect 14489 1608 14596 1627
rect 14263 1547 14328 1563
rect 14272 1540 14328 1547
rect 14347 1540 14381 1592
rect 14388 1584 14476 1592
rect 14490 1593 14596 1608
rect 14490 1584 14524 1593
rect 14544 1584 14555 1593
rect 14556 1584 14596 1593
rect 14598 1603 14638 1695
rect 14644 1694 15632 1695
rect 14644 1622 14716 1694
rect 14724 1622 14726 1666
rect 14733 1622 14738 1694
rect 14644 1604 14738 1622
rect 14758 1621 14792 1694
rect 14806 1658 15632 1694
rect 15770 1658 15820 1832
rect 14806 1624 15820 1658
rect 15823 1697 15857 1866
rect 15871 1948 15905 2263
rect 15997 2211 16013 2223
rect 15997 2201 16017 2211
rect 15997 2195 16013 2201
rect 15981 2180 15983 2189
rect 15991 2180 16015 2195
rect 16029 2189 16053 2223
rect 16153 2201 16173 2291
rect 15965 2161 16031 2180
rect 15969 2155 16027 2161
rect 15985 2142 16019 2146
rect 16031 2142 16055 2145
rect 16073 2142 16093 2146
rect 15973 2130 16031 2142
rect 16067 2130 16093 2142
rect 15973 2127 16028 2130
rect 15937 2114 15939 2118
rect 15951 2114 15971 2118
rect 15925 2110 15977 2114
rect 15979 2110 16019 2127
rect 15925 2072 15971 2110
rect 15985 2072 16019 2110
rect 16025 2114 16059 2118
rect 16025 2110 16065 2114
rect 16067 2110 16097 2130
rect 16025 2072 16059 2110
rect 16073 2106 16097 2110
rect 16105 2106 16107 2146
rect 16073 2072 16107 2106
rect 16114 2072 16119 2142
rect 16139 2072 16173 2201
rect 16187 2244 16221 2291
rect 16240 2244 16275 2272
rect 16336 2244 16494 2272
rect 17071 2263 17129 2269
rect 16187 2210 16227 2244
rect 16288 2238 16494 2244
rect 16555 2238 16590 2255
rect 16288 2210 16446 2238
rect 16187 2072 16226 2210
rect 16240 2083 16274 2210
rect 16366 2158 16382 2170
rect 16366 2148 16386 2158
rect 16366 2142 16382 2148
rect 16350 2127 16352 2136
rect 16360 2127 16384 2142
rect 16398 2138 16422 2170
rect 16522 2148 16542 2238
rect 16396 2130 16444 2138
rect 16334 2110 16400 2127
rect 16334 2108 16472 2110
rect 16396 2106 16472 2108
rect 16354 2089 16388 2106
rect 16396 2102 16476 2106
rect 16400 2089 16424 2092
rect 16342 2083 16400 2089
rect 16442 2083 16476 2102
rect 16240 2072 16476 2083
rect 16483 2072 16488 2089
rect 16508 2072 16542 2148
rect 16556 2237 16590 2238
rect 16556 2201 16626 2237
rect 17071 2229 17083 2263
rect 17071 2223 17129 2229
rect 16556 2167 16644 2201
rect 16556 2110 16643 2167
rect 17021 2148 17179 2161
rect 17260 2148 17275 2602
rect 17294 2568 17329 2602
rect 17609 2568 17680 2602
rect 17294 2148 17328 2568
rect 17610 2567 17680 2568
rect 17627 2533 17698 2567
rect 17978 2533 18013 2567
rect 17440 2500 17498 2506
rect 17440 2466 17452 2500
rect 17440 2460 17498 2466
rect 17440 2210 17498 2216
rect 17440 2176 17452 2210
rect 17440 2170 17498 2176
rect 17021 2127 17232 2148
rect 16944 2110 16959 2127
rect 16978 2126 17013 2127
rect 17074 2126 17232 2127
rect 17627 2131 17697 2533
rect 17979 2514 18013 2533
rect 17809 2465 17867 2471
rect 17809 2431 17821 2465
rect 17809 2425 17867 2431
rect 17809 2157 17867 2163
rect 16978 2114 17294 2126
rect 16978 2110 17012 2114
rect 16556 2108 17524 2110
rect 16556 2095 17548 2108
rect 16556 2072 17601 2095
rect 15912 2061 17601 2072
rect 17627 2078 17733 2131
rect 17809 2123 17821 2157
rect 17809 2117 17867 2123
rect 17998 2078 18013 2514
rect 18032 2480 18067 2514
rect 18347 2480 18382 2514
rect 18032 2078 18066 2480
rect 18348 2461 18382 2480
rect 18178 2412 18236 2418
rect 18178 2378 18190 2412
rect 18178 2372 18236 2378
rect 18178 2104 18236 2110
rect 15912 2038 17524 2061
rect 15925 2000 15971 2038
rect 15985 2000 16019 2038
rect 15925 1974 15977 2000
rect 15979 1974 16019 2000
rect 16025 2002 16059 2038
rect 16073 2002 16097 2038
rect 16105 2002 16107 2038
rect 16114 2002 16119 2038
rect 15925 1962 16005 1974
rect 15925 1948 15980 1962
rect 15985 1958 16005 1962
rect 15992 1949 16005 1958
rect 16025 1962 16119 2002
rect 16025 1949 16071 1962
rect 16073 1958 16107 1962
rect 15992 1948 16071 1949
rect 15871 1920 15911 1948
rect 15937 1934 15977 1948
rect 15937 1920 15971 1934
rect 15871 1886 15971 1920
rect 15871 1813 15911 1886
rect 15937 1847 15971 1886
rect 15933 1813 15971 1847
rect 15983 1915 16071 1948
rect 16092 1936 16125 1948
rect 16092 1915 16138 1936
rect 15983 1881 16138 1915
rect 15983 1865 16071 1881
rect 15983 1813 16013 1865
rect 16056 1850 16071 1865
rect 16092 1865 16094 1881
rect 16104 1865 16138 1881
rect 16025 1813 16059 1847
rect 16092 1836 16138 1865
rect 16092 1813 16125 1836
rect 16139 1813 16173 2038
rect 16187 1813 16226 2038
rect 15871 1779 16071 1813
rect 16092 1779 16226 1813
rect 15892 1768 15911 1779
rect 15950 1769 15971 1779
rect 15983 1769 16013 1779
rect 15937 1768 15971 1769
rect 15980 1768 16013 1769
rect 16092 1768 16125 1779
rect 15937 1766 15983 1768
rect 15935 1754 15983 1766
rect 15983 1731 16013 1754
rect 15981 1713 16015 1731
rect 16139 1716 16173 1779
rect 15969 1707 16027 1713
rect 15969 1697 15981 1707
rect 16139 1697 16190 1716
rect 15823 1663 15874 1697
rect 15939 1686 16042 1697
rect 16109 1686 16190 1697
rect 15950 1674 16031 1686
rect 16120 1682 16190 1686
rect 15939 1663 16042 1674
rect 16120 1666 16173 1682
rect 15823 1624 15857 1663
rect 14806 1621 15614 1624
rect 14758 1608 15614 1621
rect 15762 1616 15764 1622
rect 15720 1608 15732 1616
rect 15762 1608 15774 1616
rect 14758 1604 15780 1608
rect 14598 1591 14624 1603
rect 14388 1574 14596 1584
rect 14644 1590 15780 1604
rect 15823 1590 15838 1624
rect 15939 1594 16042 1605
rect 15950 1590 16031 1594
rect 14644 1586 15614 1590
rect 15730 1587 15740 1590
rect 15754 1587 15774 1590
rect 14644 1585 14893 1586
rect 14961 1585 14978 1586
rect 15062 1585 15096 1586
rect 14644 1578 15143 1585
rect 14598 1575 15143 1578
rect 14598 1574 14893 1575
rect 14229 1531 14381 1540
rect 11859 1529 14387 1531
rect 14389 1529 14423 1574
rect 14427 1568 14434 1574
rect 14437 1568 14476 1574
rect 14427 1550 14476 1568
rect 14490 1568 14524 1574
rect 14490 1550 14529 1568
rect 14427 1534 14529 1550
rect 14544 1563 14596 1574
rect 14614 1568 14893 1574
rect 14907 1574 15143 1575
rect 14907 1568 15161 1574
rect 14614 1565 15161 1568
rect 14544 1562 14590 1563
rect 14544 1550 14552 1562
rect 14556 1550 14590 1562
rect 14544 1546 14590 1550
rect 14549 1540 14590 1546
rect 14614 1560 14644 1565
rect 14650 1560 15161 1565
rect 14614 1551 15161 1560
rect 14614 1544 15107 1551
rect 14556 1534 14590 1540
rect 14437 1529 14529 1534
rect 11859 1506 14529 1529
rect 11859 1495 14387 1506
rect 14389 1495 14423 1506
rect 14437 1504 14529 1506
rect 14437 1495 14524 1504
rect 11859 1491 14437 1495
rect 11859 1484 11894 1491
rect 11901 1484 11935 1491
rect 11825 1474 11935 1484
rect 11768 1472 11935 1474
rect 11940 1480 12023 1491
rect 11940 1472 12016 1480
rect 12061 1472 12095 1491
rect 12103 1472 12137 1491
rect 12156 1472 12209 1491
rect 12228 1478 14437 1491
rect 14442 1478 14524 1495
rect 14549 1478 14590 1534
rect 14632 1540 15107 1544
rect 15127 1540 15161 1551
rect 14632 1534 15161 1540
rect 14632 1510 14893 1534
rect 14961 1529 15013 1534
rect 15032 1529 15161 1534
rect 15175 1532 15209 1586
rect 14959 1524 14978 1529
rect 14998 1525 15007 1529
rect 14948 1510 14978 1524
rect 15019 1510 15020 1529
rect 15032 1525 15066 1529
rect 15086 1525 15143 1529
rect 15032 1517 15143 1525
rect 15032 1515 15106 1517
rect 15127 1515 15143 1517
rect 15175 1526 15221 1532
rect 15228 1526 15262 1586
rect 15308 1574 15614 1586
rect 15633 1576 15685 1587
rect 15730 1576 15775 1587
rect 15418 1570 15614 1574
rect 15644 1574 15674 1576
rect 15730 1574 15764 1576
rect 15644 1570 15803 1574
rect 15330 1532 15341 1566
rect 15342 1540 15376 1570
rect 15418 1553 15803 1570
rect 15823 1553 15837 1590
rect 15950 1582 16072 1590
rect 15939 1576 16083 1582
rect 16150 1576 16173 1666
rect 16192 1644 16226 1779
rect 16240 1814 16274 2038
rect 16294 2000 16340 2038
rect 16354 2000 16388 2038
rect 16294 1967 16346 2000
rect 16348 1967 16388 2000
rect 16394 2004 16428 2038
rect 16394 2000 16430 2004
rect 16442 2000 16466 2038
rect 16474 2004 16476 2038
rect 16394 1967 16434 2000
rect 16436 1967 16466 2000
rect 16483 1989 16488 2038
rect 16477 1970 16488 1989
rect 16294 1954 16466 1967
rect 16474 1954 16488 1970
rect 16294 1948 16488 1954
rect 16306 1936 16480 1948
rect 16280 1921 16480 1936
rect 16280 1909 16462 1921
rect 16474 1909 16480 1921
rect 16280 1881 16352 1909
rect 16354 1905 16480 1909
rect 16280 1836 16340 1881
rect 16346 1868 16352 1881
rect 16362 1881 16480 1905
rect 16362 1878 16430 1881
rect 16432 1878 16480 1881
rect 16362 1870 16480 1878
rect 16508 1939 16542 2038
rect 16556 1999 17524 2038
rect 16556 1983 17551 1999
rect 17627 1985 18102 2078
rect 18178 2070 18190 2104
rect 18178 2064 18236 2070
rect 18367 2007 18382 2461
rect 18401 2427 18436 2461
rect 18401 2007 18435 2427
rect 18547 2359 18605 2365
rect 18547 2325 18559 2359
rect 18717 2336 18751 2354
rect 18547 2319 18605 2325
rect 18717 2300 18787 2336
rect 18734 2266 18805 2300
rect 18547 2051 18605 2057
rect 18547 2017 18559 2051
rect 18547 2011 18605 2017
rect 18181 2002 18339 2007
rect 16556 1959 17535 1983
rect 16556 1953 17551 1959
rect 16556 1939 17524 1953
rect 16364 1862 16479 1870
rect 16240 1768 16294 1814
rect 16306 1794 16340 1836
rect 16302 1768 16340 1794
rect 16240 1760 16274 1768
rect 16294 1760 16340 1768
rect 16382 1828 16479 1862
rect 16382 1814 16448 1828
rect 16382 1812 16492 1814
rect 16382 1794 16396 1812
rect 16382 1760 16428 1794
rect 16440 1768 16492 1812
rect 16508 1797 17524 1939
rect 17682 1888 17697 1985
rect 17716 1888 17750 1985
rect 17862 1940 17920 1946
rect 17996 1945 18102 1985
rect 18128 1973 18339 2002
rect 18400 1973 18435 2007
rect 18128 1968 18291 1973
rect 18133 1945 18291 1968
rect 17862 1906 17874 1940
rect 17996 1932 18119 1945
rect 17862 1900 17920 1906
rect 18001 1888 18119 1932
rect 17632 1797 18119 1888
rect 18211 1893 18227 1905
rect 18211 1883 18231 1893
rect 18211 1877 18227 1883
rect 18195 1862 18197 1871
rect 18205 1862 18229 1877
rect 18243 1871 18267 1905
rect 18367 1878 18387 1973
rect 18179 1843 18245 1862
rect 18183 1837 18241 1843
rect 18199 1824 18233 1828
rect 18245 1824 18269 1827
rect 18287 1824 18307 1828
rect 18187 1812 18245 1824
rect 18281 1812 18307 1824
rect 18187 1809 18242 1812
rect 16508 1763 17595 1797
rect 17629 1763 18119 1797
rect 18151 1796 18153 1800
rect 18165 1796 18185 1800
rect 16508 1760 17524 1763
rect 16240 1743 17524 1760
rect 16240 1726 16280 1743
rect 16294 1741 17524 1743
rect 16294 1732 16911 1741
rect 16294 1729 16643 1732
rect 16671 1729 16709 1732
rect 16763 1729 16800 1732
rect 16294 1726 16629 1729
rect 16382 1716 16396 1726
rect 16508 1716 16629 1726
rect 16382 1701 16411 1716
rect 16472 1692 16626 1716
rect 16638 1707 16643 1729
rect 16663 1714 16721 1729
rect 16751 1716 16809 1729
rect 16663 1707 16709 1714
rect 16716 1707 16721 1714
rect 16732 1707 16809 1716
rect 16824 1707 16831 1732
rect 16843 1707 16858 1732
rect 16877 1707 16911 1732
rect 16925 1707 16964 1741
rect 16472 1682 16488 1692
rect 16508 1690 16626 1692
rect 16663 1696 16823 1707
rect 16334 1660 16338 1670
rect 16350 1660 16384 1678
rect 16508 1666 16595 1690
rect 16609 1684 16610 1690
rect 16663 1684 16812 1696
rect 16609 1682 16621 1684
rect 16609 1678 16629 1682
rect 16663 1678 16823 1684
rect 16609 1673 16824 1678
rect 16877 1673 16897 1707
rect 16716 1666 16721 1673
rect 16751 1666 16809 1673
rect 16334 1654 16396 1660
rect 16334 1644 16350 1654
rect 16508 1644 16522 1666
rect 16192 1633 16318 1644
rect 16323 1633 16411 1644
rect 16481 1633 16522 1644
rect 16192 1621 16226 1633
rect 16230 1621 16318 1633
rect 16334 1621 16400 1633
rect 16492 1621 16522 1633
rect 16192 1614 16318 1621
rect 16192 1576 16207 1614
rect 16219 1610 16318 1614
rect 16323 1610 16411 1621
rect 16481 1610 16522 1621
rect 16219 1583 16226 1610
rect 16334 1604 16338 1610
rect 16508 1576 16522 1610
rect 15939 1571 16139 1576
rect 15870 1553 15899 1571
rect 15418 1540 15708 1553
rect 15732 1547 15762 1553
rect 15418 1532 15614 1540
rect 15276 1526 15614 1532
rect 15175 1515 15614 1526
rect 15032 1510 15143 1515
rect 15161 1510 15614 1515
rect 14632 1502 15614 1510
rect 15644 1536 15689 1540
rect 15721 1536 15773 1547
rect 15644 1519 15688 1536
rect 15770 1523 15773 1536
rect 15770 1519 15779 1523
rect 15789 1519 15804 1553
rect 15644 1506 15694 1519
rect 15649 1502 15688 1506
rect 14632 1496 15688 1502
rect 15707 1501 15766 1506
rect 14632 1494 15680 1496
rect 14644 1484 15680 1494
rect 15691 1485 15766 1501
rect 15691 1484 15728 1485
rect 15736 1484 15766 1485
rect 15770 1484 15804 1519
rect 15823 1484 15857 1553
rect 15865 1488 15899 1553
rect 15904 1527 15938 1571
rect 15965 1561 15981 1571
rect 16024 1561 16139 1571
rect 15969 1555 16139 1561
rect 16024 1552 16139 1555
rect 16004 1540 16139 1552
rect 15904 1514 15933 1527
rect 15983 1514 16013 1524
rect 16024 1514 16139 1540
rect 15904 1499 15983 1514
rect 16013 1509 16139 1514
rect 16024 1508 16139 1509
rect 16150 1574 16207 1576
rect 16150 1548 16192 1574
rect 16150 1508 16207 1548
rect 16226 1508 16522 1576
rect 16525 1644 16595 1666
rect 16782 1654 16809 1666
rect 16767 1644 16809 1654
rect 16824 1644 16831 1673
rect 16525 1639 16675 1644
rect 16709 1639 16763 1644
rect 16767 1639 16824 1644
rect 16525 1546 16595 1639
rect 16782 1635 16811 1639
rect 16669 1610 16811 1635
rect 16707 1601 16765 1607
rect 16703 1576 16769 1601
rect 16707 1567 16719 1576
rect 16707 1561 16765 1567
rect 16612 1546 16614 1561
rect 16782 1551 16811 1610
rect 16525 1540 16614 1546
rect 16525 1508 16595 1540
rect 16025 1506 16059 1508
rect 15904 1488 15980 1499
rect 15865 1484 15980 1488
rect 14644 1478 15728 1484
rect 12228 1472 15728 1478
rect 15732 1472 15980 1484
rect -17 1438 3965 1468
rect 3973 1464 15779 1472
rect -17 1421 1036 1438
rect 1082 1421 1107 1438
rect -17 1367 774 1421
rect 835 1374 869 1401
rect 949 1367 988 1421
rect 1002 1367 1036 1421
rect 1116 1402 1160 1438
rect 1188 1402 1238 1436
rect 1318 1434 3788 1438
rect 1318 1416 3770 1434
rect 3812 1416 3965 1438
rect 1318 1402 3596 1416
rect 1116 1384 3596 1402
rect 3602 1404 3676 1416
rect 3694 1415 3858 1416
rect 3682 1411 3846 1415
rect 3682 1404 3832 1411
rect 3602 1402 3832 1404
rect 3602 1400 3842 1402
rect 3602 1388 3676 1400
rect 3608 1387 3680 1388
rect 3694 1387 3708 1400
rect 3718 1387 3752 1400
rect 3782 1391 3828 1400
rect 3764 1387 3828 1391
rect 3608 1384 3828 1387
rect 3859 1384 3916 1416
rect 3926 1384 3965 1416
rect 1116 1368 3608 1384
rect 1116 1367 1141 1368
rect -17 1362 1036 1367
rect -17 1353 823 1362
rect 853 1353 1036 1362
rect -17 1348 1036 1353
rect 1082 1348 1158 1367
rect -17 1334 1158 1348
rect -17 1333 1162 1334
rect -17 1331 791 1333
rect 793 1331 800 1333
rect -17 1321 800 1331
rect -17 1315 837 1321
rect -17 1299 841 1315
rect -17 1281 800 1299
rect 832 1281 841 1299
rect 854 1281 875 1333
rect 949 1312 988 1333
rect 949 1281 996 1312
rect -17 1275 837 1281
rect -17 1250 800 1275
rect 854 1250 856 1281
rect -17 1213 791 1250
rect 866 1247 875 1281
rect 899 1271 912 1281
rect 942 1271 996 1281
rect 899 1231 996 1271
rect 899 1225 983 1231
rect 899 1215 912 1225
rect 942 1222 983 1225
rect 1002 1222 1036 1333
rect 1042 1305 1070 1333
rect 1073 1314 1162 1333
rect 1204 1321 1238 1354
rect 1239 1348 1250 1368
rect 1318 1348 3608 1368
rect 1250 1343 1254 1348
rect 1284 1343 3608 1348
rect 1318 1336 3608 1343
rect 1296 1334 3608 1336
rect 1318 1314 3608 1334
rect 3610 1328 3965 1384
rect 3636 1326 3965 1328
rect 1073 1309 3608 1314
rect 1073 1305 1107 1309
rect 1042 1286 1107 1305
rect 1112 1298 3608 1309
rect 3610 1322 3740 1326
rect 3610 1298 3644 1322
rect 1112 1286 3644 1298
rect 1042 1236 1070 1286
rect 942 1215 1036 1222
rect 942 1213 947 1215
rect 949 1214 1036 1215
rect 1073 1214 1107 1286
rect 1124 1280 3644 1286
rect 1124 1270 1160 1280
rect 949 1213 1107 1214
rect -17 1202 1107 1213
rect -17 1179 993 1202
rect 1002 1183 1107 1202
rect -17 1168 800 1179
rect 854 1168 859 1179
rect 912 1168 916 1179
rect -17 1125 791 1168
rect 912 1163 917 1168
rect 968 1163 993 1179
rect 905 1132 993 1163
rect 882 1125 993 1132
rect -17 1091 993 1125
rect 1000 1168 1107 1183
rect 1000 1137 1030 1168
rect 1073 1160 1107 1168
rect 1126 1268 1160 1270
rect 1196 1270 1242 1280
rect 1318 1272 3644 1280
rect 3664 1272 3670 1322
rect 3676 1300 3710 1322
rect 3718 1310 3740 1322
rect 3764 1322 3828 1326
rect 3764 1318 3818 1322
rect 3718 1306 3758 1310
rect 3728 1300 3758 1306
rect 3764 1300 3798 1318
rect 3825 1310 3828 1322
rect 3859 1319 3916 1326
rect 3926 1319 3965 1326
rect 3979 1451 15779 1464
rect 15789 1462 15980 1472
rect 16092 1462 16125 1508
rect 16139 1462 16173 1508
rect 16192 1462 16226 1508
rect 16298 1502 16396 1508
rect 16298 1462 16394 1502
rect 15789 1461 16394 1462
rect 16434 1461 16435 1508
rect 16508 1499 16595 1508
rect 16843 1499 16858 1673
rect 16877 1499 16892 1673
rect 16508 1482 16668 1499
rect 16771 1488 16823 1499
rect 16782 1482 16812 1488
rect 16896 1482 16911 1673
rect 16508 1465 16911 1482
rect 16930 1506 16964 1707
rect 16978 1654 17012 1741
rect 17042 1731 17046 1741
rect 17098 1739 17122 1741
rect 17136 1739 17160 1741
rect 17093 1706 17186 1739
rect 17200 1706 17228 1741
rect 17093 1698 17138 1706
rect 17093 1697 17120 1698
rect 17151 1697 17200 1698
rect 17135 1688 17201 1697
rect 17260 1688 17280 1741
rect 17040 1676 17078 1688
rect 17132 1681 17200 1688
rect 17132 1676 17162 1681
rect 17032 1664 17078 1676
rect 17032 1654 17046 1664
rect 17120 1661 17178 1676
rect 17132 1654 17178 1661
rect 17185 1654 17200 1681
rect 17246 1654 17280 1688
rect 17294 1654 17333 1741
rect 16978 1643 17241 1654
rect 16978 1631 17230 1643
rect 16978 1620 17178 1631
rect 17189 1620 17241 1631
rect 17246 1620 17266 1654
rect 17299 1648 17333 1654
rect 17280 1620 17333 1648
rect 17032 1611 17118 1620
rect 17265 1614 17280 1620
rect 17299 1614 17333 1620
rect 17030 1586 17118 1611
rect 17280 1586 17333 1614
rect 17046 1561 17090 1586
rect 17096 1548 17106 1579
rect 17088 1544 17118 1548
rect 17072 1514 17138 1544
rect 17042 1506 17076 1510
rect 16930 1465 16965 1506
rect 17042 1494 17088 1506
rect 17142 1494 17153 1506
rect 17154 1494 17172 1510
rect 17042 1480 17172 1494
rect 17246 1506 17280 1560
rect 3979 1449 15770 1451
rect 3979 1438 15773 1449
rect 3979 1420 4013 1438
rect 4033 1424 4092 1438
rect 4017 1420 4092 1424
rect 4093 1420 4127 1438
rect 4133 1420 4167 1438
rect 3979 1400 4167 1420
rect 4175 1411 4227 1438
rect 4228 1411 4281 1438
rect 4295 1415 4536 1438
rect 4295 1411 4334 1415
rect 4342 1411 4382 1415
rect 4388 1411 4536 1415
rect 4175 1406 4536 1411
rect 4542 1406 4596 1438
rect 4175 1404 4596 1406
rect 4175 1400 4538 1404
rect 4542 1400 4596 1404
rect 3979 1362 4173 1400
rect 4175 1383 4281 1400
rect 4295 1383 4346 1400
rect 4175 1362 4346 1383
rect 3979 1348 4346 1362
rect 4348 1377 4596 1400
rect 4348 1367 4460 1377
rect 4462 1367 4596 1377
rect 4348 1348 4596 1367
rect 4597 1434 7693 1438
rect 7701 1434 7788 1438
rect 4597 1429 7689 1434
rect 4597 1348 4650 1429
rect 4664 1416 7689 1429
rect 7701 1425 7704 1434
rect 7694 1416 7704 1425
rect 7716 1416 7788 1434
rect 7804 1416 8542 1438
rect 4664 1415 7716 1416
rect 4664 1404 7729 1415
rect 7766 1408 7804 1416
rect 7735 1404 7804 1408
rect 7823 1404 7880 1416
rect 4664 1400 7880 1404
rect 4664 1387 7716 1400
rect 7723 1387 7880 1400
rect 4664 1384 7880 1387
rect 7892 1409 8542 1416
rect 8561 1434 11657 1438
rect 11665 1434 11752 1438
rect 8561 1429 11653 1434
rect 8561 1409 8614 1429
rect 8663 1428 8964 1429
rect 8966 1428 11653 1429
rect 8663 1424 11653 1428
rect 11665 1425 11668 1434
rect 8660 1421 11653 1424
rect 8660 1420 8809 1421
rect 8824 1420 11653 1421
rect 8660 1416 11653 1420
rect 11658 1416 11668 1425
rect 11680 1416 11752 1434
rect 11768 1416 12506 1438
rect 8660 1415 11680 1416
rect 8660 1409 11693 1415
rect 7892 1404 11693 1409
rect 11730 1408 11768 1416
rect 11699 1404 11768 1408
rect 11787 1404 11844 1416
rect 7892 1400 11844 1404
rect 7892 1394 11680 1400
rect 7892 1384 8831 1394
rect 4664 1348 7892 1384
rect 3979 1330 7892 1348
rect 3979 1319 4085 1330
rect 4091 1328 7892 1330
rect 4091 1319 4281 1328
rect 3804 1300 3842 1310
rect 3676 1272 3840 1300
rect 3859 1285 3928 1319
rect 3931 1285 4281 1319
rect 3878 1272 3912 1285
rect 1196 1268 1241 1270
rect 1126 1259 1241 1268
rect 1318 1259 3608 1272
rect 1126 1247 3608 1259
rect 3610 1266 3912 1272
rect 3926 1266 3965 1285
rect 3610 1247 3928 1266
rect 3931 1247 3965 1266
rect 1126 1246 3965 1247
rect 1126 1228 1160 1246
rect 1174 1238 3965 1246
rect 1174 1236 3608 1238
rect 1196 1229 3608 1236
rect 3610 1232 3965 1238
rect 3664 1229 3710 1232
rect 3764 1229 3798 1232
rect 3878 1229 3928 1232
rect 3931 1229 3965 1232
rect 3979 1272 4079 1285
rect 4091 1281 4281 1285
rect 4091 1272 4179 1281
rect 4187 1272 4202 1281
rect 4212 1272 4281 1281
rect 4295 1272 4334 1328
rect 4348 1318 4588 1328
rect 4348 1310 4382 1318
rect 4388 1310 4588 1318
rect 4346 1300 4448 1310
rect 4348 1272 4382 1300
rect 4388 1272 4448 1300
rect 4454 1309 4588 1310
rect 4454 1272 4460 1309
rect 4462 1305 4588 1309
rect 4470 1286 4588 1305
rect 4470 1272 4482 1286
rect 4490 1272 4588 1286
rect 4597 1326 7892 1328
rect 4597 1322 7704 1326
rect 4597 1272 7689 1322
rect 7694 1306 7704 1322
rect 7728 1322 7792 1326
rect 7728 1272 7769 1322
rect 7789 1272 7792 1322
rect 7823 1272 7892 1326
rect 3979 1238 4019 1272
rect 4020 1238 7892 1272
rect 1196 1228 3971 1229
rect 1126 1222 1210 1228
rect 1126 1160 1160 1222
rect 1196 1214 1210 1222
rect 1237 1214 3971 1228
rect 1196 1212 3971 1214
rect 1196 1168 1254 1212
rect 1284 1194 3971 1212
rect 1268 1178 3971 1194
rect 3979 1215 4079 1238
rect 3979 1213 4019 1215
rect 4045 1213 4079 1215
rect 4091 1215 4167 1238
rect 4091 1213 4121 1215
rect 4133 1213 4167 1215
rect 4200 1236 4587 1238
rect 4597 1236 7689 1238
rect 4200 1232 7689 1236
rect 4200 1215 4246 1232
rect 4200 1213 4233 1215
rect 4247 1213 4281 1232
rect 4295 1213 4334 1232
rect 3979 1204 4334 1213
rect 3979 1201 4179 1204
rect 4200 1201 4334 1204
rect 4348 1214 4382 1232
rect 4412 1215 4448 1232
rect 4348 1201 4402 1214
rect 4414 1202 4448 1215
rect 3979 1200 4408 1201
rect 3979 1199 4179 1200
rect 4200 1199 4334 1200
rect 3979 1179 4334 1199
rect 1284 1176 3971 1178
rect 4000 1176 4085 1179
rect 4088 1176 4179 1179
rect 4200 1176 4281 1179
rect 4288 1176 4334 1179
rect 1284 1173 4340 1176
rect 4348 1173 4402 1200
rect 4412 1199 4448 1202
rect 4458 1203 4459 1232
rect 4490 1229 7689 1232
rect 7728 1236 7769 1238
rect 7823 1236 7892 1238
rect 7728 1229 7762 1236
rect 7842 1229 7892 1236
rect 7895 1319 7929 1384
rect 7937 1362 8831 1384
rect 7937 1349 8762 1362
rect 8763 1358 8831 1362
rect 7937 1348 8787 1349
rect 8796 1348 8831 1358
rect 8840 1356 8854 1374
rect 8836 1348 8854 1356
rect 8877 1364 8911 1394
rect 8930 1374 8964 1394
rect 8966 1387 11680 1394
rect 11687 1387 11844 1400
rect 8966 1384 11844 1387
rect 11856 1409 12506 1416
rect 12525 1434 15621 1438
rect 15629 1434 15716 1438
rect 12525 1429 15617 1434
rect 12525 1409 12578 1429
rect 12627 1428 12928 1429
rect 12930 1428 15617 1429
rect 12627 1424 15617 1428
rect 15629 1425 15632 1434
rect 12624 1421 15617 1424
rect 12624 1420 12773 1421
rect 12788 1420 15617 1421
rect 12624 1416 15617 1420
rect 15622 1416 15632 1425
rect 15644 1416 15716 1434
rect 15732 1416 15773 1438
rect 15789 1439 16326 1461
rect 16382 1446 16411 1461
rect 16382 1439 16396 1446
rect 16434 1439 16440 1461
rect 15789 1416 16440 1439
rect 12624 1415 15644 1416
rect 12624 1409 15657 1415
rect 11856 1404 15657 1409
rect 15694 1408 15732 1416
rect 15770 1408 15808 1416
rect 15663 1404 15732 1408
rect 15751 1404 15808 1408
rect 11856 1400 15808 1404
rect 11856 1394 15644 1400
rect 11856 1384 12795 1394
rect 8966 1376 11856 1384
rect 8928 1364 8964 1374
rect 8877 1360 8916 1364
rect 8920 1360 8964 1364
rect 8877 1348 8964 1360
rect 9014 1356 9018 1376
rect 9032 1372 11856 1376
rect 8986 1348 9018 1356
rect 7937 1339 8967 1348
rect 9014 1339 9016 1348
rect 9026 1341 11856 1372
rect 7937 1327 9019 1339
rect 9026 1338 9182 1341
rect 9190 1338 11856 1341
rect 9026 1327 9166 1338
rect 7937 1326 9166 1327
rect 9214 1326 11856 1338
rect 7937 1319 9019 1326
rect 7895 1286 9019 1319
rect 9026 1309 9090 1326
rect 9097 1309 9131 1326
rect 9132 1321 9166 1326
rect 9132 1309 9165 1321
rect 9026 1306 9038 1309
rect 9044 1306 9086 1309
rect 9026 1296 9086 1306
rect 9097 1306 9169 1309
rect 9224 1306 9226 1326
rect 9246 1322 11668 1326
rect 9246 1306 11653 1322
rect 11658 1306 11668 1322
rect 11692 1322 11756 1326
rect 9097 1296 9170 1306
rect 9026 1286 9170 1296
rect 9224 1286 11653 1306
rect 7895 1285 11653 1286
rect 7895 1229 7929 1285
rect 7937 1272 11653 1285
rect 11692 1272 11733 1322
rect 11753 1272 11756 1322
rect 11787 1272 11856 1326
rect 7937 1238 11856 1272
rect 7937 1229 11653 1238
rect 11692 1236 11733 1238
rect 11787 1236 11856 1238
rect 11692 1229 11726 1236
rect 11806 1229 11856 1236
rect 11859 1319 11893 1384
rect 11901 1362 12795 1384
rect 11901 1349 12726 1362
rect 12727 1358 12795 1362
rect 11901 1348 12751 1349
rect 12760 1348 12795 1358
rect 12804 1356 12818 1374
rect 12800 1348 12818 1356
rect 12841 1364 12875 1394
rect 12894 1374 12928 1394
rect 12930 1387 15644 1394
rect 15651 1387 15808 1400
rect 12930 1384 15808 1387
rect 15820 1409 16440 1416
rect 16508 1429 16578 1465
rect 16930 1464 16964 1465
rect 16620 1446 17042 1464
rect 17246 1446 17288 1506
rect 16620 1429 17088 1446
rect 17142 1429 17288 1446
rect 16508 1409 16542 1429
rect 16578 1424 16832 1429
rect 16578 1409 16892 1424
rect 15820 1384 16578 1409
rect 12930 1376 15820 1384
rect 12892 1364 12928 1374
rect 12841 1360 12880 1364
rect 12884 1360 12928 1364
rect 12841 1348 12928 1360
rect 12978 1356 12982 1376
rect 12996 1372 15820 1376
rect 12950 1348 12982 1356
rect 11901 1339 12931 1348
rect 12978 1339 12980 1348
rect 12990 1341 15820 1372
rect 15823 1356 15857 1384
rect 15831 1354 15857 1356
rect 11901 1327 12983 1339
rect 12990 1338 13146 1341
rect 13154 1338 15820 1341
rect 12990 1327 13130 1338
rect 11901 1326 13130 1327
rect 13178 1326 15820 1338
rect 11901 1319 12983 1326
rect 11859 1286 12983 1319
rect 12990 1309 13054 1326
rect 13061 1309 13095 1326
rect 13096 1321 13130 1326
rect 13096 1309 13129 1321
rect 12990 1306 13002 1309
rect 13008 1306 13050 1309
rect 12990 1296 13050 1306
rect 13061 1306 13133 1309
rect 13188 1306 13190 1326
rect 13210 1322 15632 1326
rect 13210 1306 15617 1322
rect 15622 1306 15632 1322
rect 15656 1322 15720 1326
rect 13061 1296 13134 1306
rect 12990 1286 13134 1296
rect 13188 1286 15617 1306
rect 11859 1285 15617 1286
rect 11859 1229 11893 1285
rect 11901 1272 15617 1285
rect 15656 1272 15697 1322
rect 15717 1272 15720 1322
rect 15751 1310 15762 1326
rect 15770 1310 15820 1326
rect 15751 1272 15820 1310
rect 11901 1238 15820 1272
rect 11901 1229 15617 1238
rect 15656 1236 15697 1238
rect 15751 1236 15820 1238
rect 15656 1229 15690 1236
rect 15770 1229 15820 1236
rect 15823 1229 15857 1354
rect 15865 1373 16578 1384
rect 16620 1373 16673 1409
rect 15865 1339 16673 1373
rect 16724 1394 16892 1409
rect 16894 1412 17288 1429
rect 16894 1411 17042 1412
rect 17265 1411 17288 1412
rect 17299 1411 17333 1586
rect 17347 1614 17381 1741
rect 17400 1711 17430 1741
rect 17581 1737 17583 1763
rect 17590 1741 17595 1763
rect 17615 1741 18119 1763
rect 17455 1711 17476 1737
rect 17441 1703 17476 1711
rect 17615 1703 17617 1741
rect 17441 1695 17529 1703
rect 17441 1661 17491 1695
rect 17505 1669 17529 1695
rect 17441 1645 17476 1661
rect 17409 1623 17447 1635
rect 17459 1623 17476 1645
rect 17629 1635 18119 1741
rect 17401 1614 17453 1623
rect 17347 1601 17453 1614
rect 17467 1610 17476 1623
rect 17464 1601 17481 1610
rect 17501 1601 17535 1635
rect 17347 1567 17547 1601
rect 17615 1567 18119 1635
rect 17353 1564 17453 1567
rect 17379 1548 17453 1564
rect 17464 1564 17535 1567
rect 17464 1552 17481 1564
rect 17401 1533 17453 1548
rect 17467 1533 17476 1552
rect 17400 1529 17438 1533
rect 17400 1511 17430 1529
rect 17459 1511 17476 1533
rect 17501 1545 17535 1564
rect 17501 1529 17510 1545
rect 17441 1501 17476 1511
rect 17441 1495 17503 1501
rect 17632 1495 18119 1567
rect 18139 1616 18191 1796
rect 18193 1644 18233 1809
rect 18199 1640 18233 1644
rect 18239 1796 18273 1800
rect 18239 1644 18279 1796
rect 18281 1656 18311 1812
rect 18281 1644 18307 1656
rect 18239 1631 18285 1644
rect 18287 1640 18307 1644
rect 18319 1640 18321 1828
rect 18328 1644 18333 1824
rect 18353 1644 18387 1878
rect 18139 1606 18185 1616
rect 18139 1495 18173 1606
rect 18209 1597 18285 1631
rect 18353 1606 18355 1644
rect 18227 1563 18307 1597
rect 18227 1547 18285 1563
rect 18270 1532 18285 1547
rect 18367 1529 18387 1644
rect 18239 1495 18273 1529
rect 18353 1495 18387 1529
rect 18401 1949 18435 1973
rect 18734 1990 18804 2266
rect 18916 2198 18974 2204
rect 18916 2164 18928 2198
rect 18916 2158 18974 2164
rect 18916 1998 18974 2004
rect 18454 1949 18489 1954
rect 18550 1949 18708 1954
rect 18401 1892 18441 1949
rect 18497 1920 18708 1949
rect 18497 1915 18660 1920
rect 18502 1892 18660 1915
rect 18401 1495 18440 1892
rect 17441 1461 17472 1495
rect 17632 1478 18125 1495
rect 17441 1455 17503 1461
rect 17441 1445 17472 1455
rect 17354 1416 17367 1420
rect 17342 1411 17387 1416
rect 16894 1394 17411 1411
rect 16724 1357 16744 1394
rect 16870 1393 17411 1394
rect 16870 1376 17488 1393
rect 16870 1364 16938 1376
rect 16782 1357 16938 1364
rect 16724 1339 16938 1357
rect 16942 1357 16943 1376
rect 16972 1366 17006 1376
rect 17088 1375 17156 1376
rect 17263 1375 17488 1376
rect 16954 1357 17006 1366
rect 16942 1339 17006 1357
rect 15865 1328 16580 1339
rect 16603 1338 17006 1339
rect 16603 1328 16965 1338
rect 15865 1303 16578 1328
rect 16603 1303 16610 1328
rect 15865 1302 16610 1303
rect 16620 1327 16965 1328
rect 16972 1327 17006 1338
rect 17025 1341 17088 1375
rect 17142 1359 17488 1375
rect 17632 1359 17702 1478
rect 17814 1442 17872 1448
rect 17814 1408 17826 1442
rect 17814 1402 17872 1408
rect 17142 1341 17411 1359
rect 17025 1327 17059 1341
rect 17088 1327 17156 1341
rect 17200 1327 17230 1331
rect 17242 1327 17411 1341
rect 16620 1326 17411 1327
rect 15865 1272 16596 1302
rect 16620 1286 16947 1326
rect 16972 1306 17006 1326
rect 16965 1298 17006 1306
rect 17025 1306 17040 1326
rect 17200 1306 17230 1326
rect 17242 1323 17411 1326
rect 17242 1322 17276 1323
rect 17442 1322 17476 1359
rect 17632 1323 17685 1359
rect 17025 1298 17059 1306
rect 17183 1300 17230 1306
rect 16965 1286 17167 1298
rect 17183 1286 17217 1300
rect 17341 1298 17375 1306
rect 17233 1286 17411 1298
rect 16620 1277 17411 1286
rect 16603 1272 17411 1277
rect 15865 1268 17375 1272
rect 17411 1268 17437 1272
rect 15865 1238 17483 1268
rect 17632 1250 17665 1323
rect 18003 1306 18018 1478
rect 18037 1379 18071 1478
rect 18085 1461 18125 1478
rect 18139 1461 18285 1495
rect 18353 1461 18373 1495
rect 18195 1395 18229 1413
rect 18183 1389 18241 1395
rect 18183 1379 18195 1389
rect 18037 1345 18072 1379
rect 18168 1368 18256 1379
rect 18179 1356 18245 1368
rect 18168 1345 18256 1356
rect 18037 1287 18071 1345
rect 18037 1253 18072 1287
rect 18168 1276 18256 1287
rect 18179 1264 18245 1276
rect 18168 1253 18256 1264
rect 17702 1250 17798 1252
rect 4490 1228 7935 1229
rect 4490 1214 4556 1228
rect 4578 1214 7935 1228
rect 4490 1212 7935 1214
rect 4458 1201 4460 1203
rect 4490 1201 4536 1212
rect 4548 1201 7935 1212
rect 4454 1200 4536 1201
rect 4542 1200 7935 1201
rect 1284 1172 4408 1173
rect 1284 1168 4340 1172
rect 1318 1162 1334 1168
rect 1335 1162 4340 1168
rect 1286 1160 1316 1162
rect 1318 1160 4340 1162
rect 1036 1159 1329 1160
rect 1335 1159 4340 1160
rect 1036 1143 4340 1159
rect 1073 1141 4340 1143
rect 1000 1126 1041 1137
rect 1073 1131 1328 1141
rect 1335 1131 4340 1141
rect 1073 1126 4340 1131
rect 4348 1168 4402 1172
rect 4414 1168 4448 1199
rect 4458 1173 4460 1200
rect 4490 1173 4536 1200
rect 4548 1179 7935 1200
rect 4548 1173 4600 1179
rect 4616 1176 7935 1179
rect 7937 1176 11899 1229
rect 11901 1176 15863 1229
rect 15865 1176 16595 1238
rect 4616 1173 16595 1176
rect 4454 1172 4536 1173
rect 4542 1172 16595 1173
rect 4348 1160 4382 1168
rect 4402 1160 4448 1168
rect 4458 1160 4460 1172
rect 4490 1160 4536 1172
rect 4548 1168 4600 1172
rect 4616 1160 16595 1172
rect 4348 1143 16595 1160
rect 4348 1126 4388 1143
rect 4402 1132 16595 1143
rect 4402 1129 4751 1132
rect 4783 1129 4785 1132
rect 4898 1129 4905 1132
rect 4402 1126 4737 1129
rect 1000 1091 1005 1126
rect -17 1057 791 1091
rect 882 1082 1005 1091
rect 859 1066 871 1070
rect 882 1066 917 1082
rect 947 1072 1005 1082
rect 1073 1072 1107 1126
rect 1126 1072 1160 1126
rect 1216 1116 4340 1126
rect 1234 1094 4340 1116
rect 4408 1116 4448 1126
rect 4458 1116 4460 1126
rect 4408 1101 4460 1116
rect 4490 1113 4536 1126
rect 4580 1116 4737 1126
rect 4490 1109 4519 1113
rect 4490 1101 4542 1109
rect 1234 1082 2881 1094
rect 1234 1072 1286 1082
rect 1294 1072 1300 1082
rect 1322 1072 2881 1082
rect 947 1066 2881 1072
rect 859 1057 872 1066
rect -17 1047 875 1057
rect -17 1029 791 1047
rect -17 1023 837 1029
rect -17 1019 841 1023
rect -17 1008 791 1019
rect 837 1008 841 1019
rect -17 989 841 1008
rect 859 1008 875 1047
rect 912 1019 917 1066
rect 897 1008 917 1019
rect 859 1004 917 1008
rect 949 1044 2881 1066
rect 2949 1044 2953 1094
rect 2980 1059 3007 1094
rect 3056 1066 3095 1094
rect 2965 1044 3007 1059
rect 3157 1044 4340 1094
rect 4380 1081 4420 1099
rect 4580 1092 4734 1116
rect 4746 1107 4751 1129
rect 4771 1114 4829 1129
rect 4859 1116 4917 1129
rect 4771 1113 4823 1114
rect 4771 1107 4817 1113
rect 4824 1107 4829 1114
rect 4840 1107 4917 1116
rect 4930 1108 5352 1132
rect 5368 1116 5388 1132
rect 4930 1107 5354 1108
rect 4580 1082 4596 1092
rect 4616 1090 4734 1092
rect 4771 1096 5354 1107
rect 5373 1107 5388 1116
rect 5402 1107 5441 1132
rect 5455 1107 5489 1132
rect 5507 1111 5538 1132
rect 5549 1107 5580 1111
rect 5632 1107 8667 1132
rect 5373 1101 5402 1107
rect 4380 1073 4570 1081
rect 4442 1047 4446 1070
rect 4616 1066 4703 1090
rect 4717 1084 4718 1090
rect 4771 1084 4920 1096
rect 4930 1091 5354 1096
rect 4927 1090 5354 1091
rect 4927 1084 5005 1090
rect 4717 1082 4729 1084
rect 4717 1078 4737 1082
rect 4771 1078 5005 1084
rect 5038 1078 5072 1090
rect 4717 1073 5005 1078
rect 5019 1073 5072 1078
rect 4418 1044 4420 1047
rect 4442 1044 4448 1047
rect 4458 1044 4492 1054
rect 4616 1044 4630 1066
rect 949 1019 983 1044
rect 992 1038 2881 1044
rect 2961 1040 2995 1042
rect 3049 1040 3083 1042
rect 3157 1041 4426 1044
rect 992 1019 1036 1038
rect 949 1004 1036 1019
rect 1042 1010 1044 1038
rect 871 1000 905 1004
rect 949 1000 993 1004
rect -17 983 837 989
rect -17 974 791 983
rect 949 976 983 1000
rect 1002 976 1036 1004
rect 1073 976 1107 1038
rect 881 974 899 976
rect 912 974 942 976
rect -17 966 942 974
rect -17 957 875 966
rect 881 957 899 966
rect 912 963 942 966
rect 949 963 1107 976
rect 903 957 1107 963
rect -17 955 1107 957
rect -17 942 815 955
rect 823 942 1107 955
rect -17 940 1107 942
rect -17 917 815 940
rect 823 927 849 940
rect 823 924 834 927
rect -17 891 791 917
rect 862 908 1107 940
rect 1126 976 1160 1038
rect 1228 976 1241 1017
rect 1254 976 1284 1038
rect 1318 1010 2881 1038
rect 1126 966 1284 976
rect 1305 1004 2881 1010
rect 2927 1006 3117 1008
rect 3163 1004 3197 1041
rect 1305 986 3210 1004
rect 1305 975 1918 986
rect 2006 982 2022 986
rect 2033 982 3210 986
rect 1126 962 1286 966
rect 1305 963 1987 975
rect 2006 964 3210 982
rect 1126 951 1308 962
rect 1126 910 1284 951
rect 1286 920 1316 951
rect 1318 948 1987 963
rect 2010 958 3210 964
rect 2033 951 3210 958
rect 3216 978 3231 1041
rect 3318 1002 3333 1041
rect 3316 991 3333 1002
rect 3406 1006 3434 1041
rect 3532 1036 4426 1041
rect 4431 1036 4519 1044
rect 3532 1033 4519 1036
rect 4589 1033 4630 1044
rect 3532 1021 4508 1033
rect 4600 1032 4630 1033
rect 3532 1016 4519 1021
rect 3532 1010 4532 1016
rect 4534 1010 4630 1032
rect 3406 991 3449 1006
rect 3216 951 3242 978
rect 3316 960 3318 991
rect 3324 974 3458 978
rect 3532 976 4340 1010
rect 4394 976 4418 994
rect 4516 986 4532 1010
rect 4534 976 4568 998
rect 4616 976 4630 1010
rect 3358 951 3360 960
rect 3532 951 4630 976
rect 2033 948 4630 951
rect 1318 942 1965 948
rect 1972 942 4630 948
rect 1318 941 4630 942
rect 1318 926 1965 941
rect 1972 930 4630 941
rect 2002 926 4630 930
rect 1318 914 4630 926
rect 1318 910 1899 914
rect 1907 910 1918 914
rect 1919 910 1959 914
rect 1966 910 2024 914
rect 2033 910 4630 914
rect 854 906 989 908
rect 14 872 165 891
rect 182 872 298 891
rect 344 872 791 891
rect 835 889 989 906
rect 835 872 881 889
rect 949 872 983 889
rect 1002 872 1036 908
rect 1073 872 1107 908
rect 1120 908 1284 910
rect 1298 908 4630 910
rect 4633 1044 4703 1066
rect 4783 1051 4817 1073
rect 4824 1066 4829 1073
rect 4859 1066 4920 1073
rect 4871 1060 4920 1066
rect 4871 1054 4917 1060
rect 4861 1044 4917 1054
rect 4932 1044 4939 1073
rect 4951 1044 4966 1073
rect 4985 1060 5000 1073
rect 5004 1060 5019 1073
rect 4985 1044 5019 1060
rect 5038 1044 5072 1073
rect 5086 1054 5120 1090
rect 5198 1088 5328 1090
rect 5335 1088 5354 1090
rect 5198 1082 5248 1088
rect 5259 1082 5308 1088
rect 5309 1082 5374 1088
rect 5259 1081 5309 1082
rect 5152 1076 5154 1080
rect 5140 1064 5154 1076
rect 5164 1064 5186 1080
rect 5240 1076 5286 1081
rect 5140 1054 5186 1064
rect 5228 1054 5286 1076
rect 5293 1054 5309 1081
rect 5335 1073 5374 1082
rect 5388 1073 5402 1101
rect 5407 1096 8667 1107
rect 5407 1084 5538 1096
rect 5549 1094 8667 1096
rect 5549 1084 6864 1094
rect 5407 1073 6864 1084
rect 5354 1054 5388 1073
rect 5402 1054 5441 1073
rect 4633 1039 4783 1044
rect 4817 1039 4932 1044
rect 4633 946 4703 1039
rect 4876 1035 4901 1039
rect 4777 1010 4911 1035
rect 4956 1010 4962 1044
rect 4966 1039 5053 1044
rect 4811 1007 4840 1010
rect 4811 1001 4873 1007
rect 4811 976 4877 1001
rect 4720 946 4722 961
rect 4633 940 4722 946
rect 4750 946 4754 974
rect 4780 946 4784 974
rect 4811 967 4840 976
rect 4951 974 4966 1010
rect 4985 994 5019 1039
rect 4985 974 5000 994
rect 5004 974 5019 994
rect 5038 994 5053 1039
rect 5086 1043 5350 1054
rect 5086 1042 5138 1043
rect 5140 1042 5350 1043
rect 5086 1039 5350 1042
rect 5086 1031 5338 1039
rect 5086 1021 5286 1031
rect 5295 1021 5349 1031
rect 5354 1021 5374 1054
rect 5388 1039 5402 1054
rect 5407 1044 5441 1054
rect 5455 1044 5489 1073
rect 5549 1061 5599 1073
rect 5613 1069 6864 1073
rect 5549 1045 5584 1061
rect 5407 1039 5550 1044
rect 5086 1020 5385 1021
rect 4811 961 4873 967
rect 4811 951 4840 961
rect 4750 940 4784 946
rect 4985 940 4994 974
rect 5038 944 5072 994
rect 5140 986 5226 1020
rect 5228 1018 5274 1020
rect 5228 1012 5280 1018
rect 5228 986 5286 1012
rect 5154 961 5198 986
rect 5240 982 5274 986
rect 5290 974 5308 990
rect 5206 948 5308 974
rect 5196 946 5226 948
rect 5196 945 5230 946
rect 5168 944 5230 945
rect 5306 944 5336 946
rect 5038 940 5336 944
rect 5338 940 5340 974
rect 5354 948 5385 1020
rect 5354 940 5388 948
rect 4633 908 4703 940
rect 1120 906 1246 908
rect 1116 902 1246 906
rect 1116 889 1184 902
rect 1109 874 1184 889
rect 1116 872 1184 874
rect 1196 889 1246 902
rect 1196 872 1250 889
rect 1268 872 1272 904
rect 1284 872 4340 908
rect 4427 902 4504 908
rect 4427 877 4502 902
rect 14 864 4340 872
rect 36 837 37 864
rect 41 838 4340 864
rect 4434 861 4502 877
rect 4542 861 4543 908
rect 4616 899 4703 908
rect 4818 899 4830 908
rect 4906 899 4935 908
rect 4951 899 4966 940
rect 4985 908 5000 940
rect 5004 908 5019 940
rect 4985 899 5019 908
rect 4616 865 4776 899
rect 4818 865 5019 899
rect 5038 910 5072 940
rect 5168 914 5246 940
rect 5354 928 5365 940
rect 5373 928 5388 940
rect 5168 910 5218 914
rect 5038 908 5096 910
rect 5038 906 5053 908
rect 5072 906 5096 908
rect 48 837 85 838
rect 87 837 125 838
rect 36 787 125 837
rect 36 783 94 787
rect 136 783 137 838
rect 182 783 298 838
rect 344 815 404 838
rect 466 827 614 838
rect 494 816 614 827
rect 436 815 512 816
rect 344 783 370 815
rect 378 811 454 815
rect 382 784 454 811
rect 382 783 472 784
rect 546 783 570 816
rect 580 783 614 816
rect 36 753 182 783
rect 211 781 382 783
rect 36 738 211 753
rect 36 726 182 738
rect 214 726 382 781
rect 436 771 614 783
rect 436 738 582 771
rect 599 738 614 771
rect 436 726 614 738
rect 48 719 82 726
rect 211 719 298 726
rect 36 698 298 719
rect 436 718 472 726
rect 436 706 451 718
rect 546 710 570 726
rect 36 685 245 698
rect 55 672 82 685
rect 136 672 170 685
rect 182 672 236 685
rect 248 672 298 698
rect 336 700 370 706
rect 436 703 482 706
rect 448 700 482 703
rect 536 700 570 710
rect 336 672 570 700
rect 55 666 577 672
rect 580 666 614 726
rect 55 651 582 666
rect 55 639 182 651
rect 214 639 582 651
rect 55 638 582 639
rect 55 615 82 638
rect 264 632 382 638
rect 436 632 582 638
rect 599 632 614 666
rect 633 820 742 838
rect 757 821 1250 838
rect 633 770 668 820
rect 633 748 700 770
rect 735 762 800 820
rect 793 748 800 762
rect 633 730 800 748
rect 633 686 700 730
rect 775 710 800 730
rect 854 806 881 821
rect 949 806 988 821
rect 854 787 900 806
rect 854 762 881 787
rect 854 748 855 762
rect 866 748 875 749
rect 949 748 1000 806
rect 1002 748 1036 821
rect 1088 806 1250 821
rect 1042 802 1250 806
rect 1318 802 4340 838
rect 1042 787 4340 802
rect 4402 839 4434 861
rect 4443 849 4460 861
rect 4448 846 4460 849
rect 4458 839 4460 846
rect 4490 846 4519 861
rect 4490 839 4504 846
rect 4402 816 4504 839
rect 4520 816 4536 824
rect 4542 816 4548 861
rect 4402 790 4548 816
rect 4616 829 4688 865
rect 1042 770 1070 787
rect 1088 770 4340 787
rect 1042 768 4340 770
rect 1042 756 1250 768
rect 1042 748 1162 756
rect 854 740 1162 748
rect 1170 740 1174 756
rect 1196 748 1250 756
rect 1318 748 4340 768
rect 4388 756 4548 790
rect 4554 756 4570 790
rect 854 728 1088 740
rect 775 706 825 710
rect 832 706 841 715
rect 754 698 841 706
rect 854 706 875 728
rect 854 698 900 706
rect 754 686 900 698
rect 633 632 668 686
rect 775 681 875 686
rect 775 672 800 681
rect 841 672 856 681
rect 866 672 875 681
rect 949 672 988 728
rect 1002 672 1036 728
rect 1042 686 1076 728
rect 1077 720 1088 728
rect 1104 734 1158 740
rect 1104 709 1162 734
rect 1196 728 4340 748
rect 4402 729 4548 756
rect 4582 740 4588 806
rect 4616 757 4650 829
rect 4676 820 4754 829
rect 4686 790 4754 820
rect 4818 790 4830 865
rect 4906 820 4920 865
rect 5038 846 5072 906
rect 5073 891 5108 906
rect 5088 846 5108 891
rect 5150 898 5218 910
rect 5262 906 5296 910
rect 5354 908 5388 928
rect 5336 906 5353 908
rect 5150 894 5184 898
rect 5262 894 5280 906
rect 5150 880 5280 894
rect 5306 846 5307 905
rect 5338 894 5353 906
rect 5354 906 5394 908
rect 5354 894 5396 906
rect 5338 893 5396 894
rect 5350 846 5396 893
rect 5038 812 5396 846
rect 5054 806 5184 812
rect 4876 790 4878 801
rect 4907 790 4920 801
rect 4964 790 4966 801
rect 4686 757 4764 790
rect 4616 739 4776 757
rect 4616 729 4688 739
rect 4346 728 4400 729
rect 4402 728 4688 729
rect 4718 728 4776 739
rect 4818 756 4878 790
rect 4918 757 4966 790
rect 5006 790 5184 806
rect 5006 778 5206 790
rect 4906 756 4966 757
rect 4994 756 5040 757
rect 5062 756 5206 778
rect 4818 728 4876 756
rect 4906 728 4964 756
rect 4994 738 5062 756
rect 5072 740 5108 756
rect 5150 738 5184 756
rect 5306 741 5307 812
rect 5350 806 5396 812
rect 5337 790 5338 801
rect 5348 759 5396 806
rect 5407 793 5441 1039
rect 5455 1010 5489 1039
rect 5515 1035 5550 1039
rect 5512 1027 5550 1035
rect 5512 1023 5521 1027
rect 5567 1023 5584 1045
rect 5509 1010 5561 1023
rect 5575 1010 5584 1023
rect 5609 1011 5618 1027
rect 5632 1021 6864 1069
rect 6878 1021 8667 1094
rect 5632 1011 8667 1021
rect 5455 1001 5561 1010
rect 5572 1001 5589 1010
rect 5609 1001 8667 1011
rect 5455 986 8667 1001
rect 5455 967 5655 986
rect 5461 964 5561 967
rect 5487 948 5561 964
rect 5572 964 5643 967
rect 5572 952 5589 964
rect 5509 933 5561 948
rect 5575 933 5589 952
rect 5508 929 5546 933
rect 5508 911 5538 929
rect 5567 911 5589 933
rect 5609 945 5643 964
rect 5609 929 5618 945
rect 5549 905 5589 911
rect 5549 895 5584 905
rect 5549 845 5580 895
rect 5450 804 5495 820
rect 5450 793 5496 804
rect 5668 793 5673 805
rect 5689 793 5714 967
rect 5723 932 7583 986
rect 7585 969 8667 986
rect 8675 1111 9502 1132
rect 9514 1111 9534 1132
rect 8675 1107 9500 1111
rect 9513 1107 9544 1111
rect 9596 1107 12631 1132
rect 8675 1094 12631 1107
rect 8675 1073 10828 1094
rect 8675 1044 9500 1073
rect 9513 1061 9579 1073
rect 9513 1055 9575 1061
rect 9513 1045 9548 1055
rect 9514 1044 9548 1045
rect 9596 1044 10828 1073
rect 10877 1044 10882 1094
rect 10908 1059 10935 1094
rect 10984 1066 11023 1094
rect 10893 1044 10935 1059
rect 8675 1027 9514 1044
rect 8675 1023 9500 1027
rect 9531 1023 9548 1044
rect 9580 1040 10828 1044
rect 10889 1040 10923 1042
rect 10977 1040 11011 1042
rect 11085 1041 12631 1094
rect 9568 1023 10828 1040
rect 8675 1011 9517 1023
rect 8675 969 9534 1011
rect 7585 945 9534 969
rect 9539 973 9548 1023
rect 9573 1021 10828 1023
rect 11091 1021 11125 1041
rect 11144 1021 11159 1041
rect 9573 986 11233 1021
rect 11246 1002 11261 1041
rect 7585 935 9517 945
rect 5723 931 7570 932
rect 5723 929 6227 931
rect 6247 929 6293 931
rect 6301 929 7570 931
rect 5723 906 7570 929
rect 7585 910 8007 935
rect 8020 922 8066 935
rect 7585 906 8010 910
rect 8020 906 8098 922
rect 5723 895 6227 906
rect 6247 895 6293 906
rect 6344 895 6381 906
rect 6406 898 7570 906
rect 7582 898 8010 906
rect 6406 895 8010 898
rect 5723 878 8010 895
rect 5723 858 5918 878
rect 5723 848 5924 858
rect 5968 848 6126 878
rect 5723 842 6126 848
rect 5723 838 5966 842
rect 5968 838 6126 842
rect 5723 816 6126 838
rect 5723 793 5882 816
rect 5894 804 5898 816
rect 5908 808 6006 816
rect 5908 804 5980 808
rect 5407 759 5596 793
rect 5646 788 5661 793
rect 5668 788 5882 793
rect 5884 802 5980 804
rect 5884 792 5966 802
rect 5884 788 5954 792
rect 5668 759 5810 788
rect 5348 756 5384 759
rect 5296 738 5307 741
rect 5350 738 5384 756
rect 5462 738 5496 759
rect 4994 728 5073 738
rect 5291 728 5306 738
rect 1198 721 1202 728
rect 1204 721 1238 728
rect 1318 726 4546 728
rect 1318 719 4340 726
rect 1042 672 1070 686
rect 1088 672 1108 698
rect 1112 696 1162 709
rect 1196 706 1207 709
rect 1318 706 3596 719
rect 1196 705 1242 706
rect 1196 696 1207 705
rect 1208 696 1242 705
rect 1112 686 1242 696
rect 1296 686 3596 706
rect 1112 685 1228 686
rect 1112 684 1241 685
rect 1126 672 1241 684
rect 1318 672 3596 686
rect 3608 672 3636 698
rect 3664 672 3670 719
rect 3676 672 3710 719
rect 3730 706 3740 719
rect 3764 672 3798 719
rect 3878 698 4340 719
rect 4432 718 4448 726
rect 4458 700 4460 726
rect 4616 703 4686 728
rect 5050 726 5073 728
rect 5250 726 5263 728
rect 5291 726 5308 728
rect 5373 725 5384 738
rect 5550 722 5584 759
rect 5740 740 5810 759
rect 5814 774 5954 788
rect 5814 744 5892 774
rect 5908 754 5954 774
rect 6008 774 6018 804
rect 6040 788 6126 816
rect 6008 754 6042 774
rect 6054 754 6126 788
rect 6145 861 6492 878
rect 6145 816 6305 861
rect 6336 851 6492 861
rect 6335 838 6492 851
rect 6495 872 6596 878
rect 6616 872 6662 878
rect 6712 872 6762 878
rect 6495 861 6529 872
rect 6539 861 6674 872
rect 6495 842 6674 861
rect 6678 842 6762 872
rect 6811 861 8010 878
rect 8032 905 8098 906
rect 8120 911 8154 935
rect 8032 888 8108 905
rect 8120 888 8132 911
rect 8142 894 8154 911
rect 8176 888 8188 910
rect 8032 872 8044 888
rect 8064 876 8108 888
rect 8126 876 8164 880
rect 6495 838 6795 842
rect 6830 838 8010 861
rect 6335 836 6602 838
rect 6336 816 6602 836
rect 6616 826 8007 838
rect 8036 826 8040 860
rect 8064 854 8110 876
rect 8060 844 8110 854
rect 8060 838 8122 844
rect 8060 826 8110 838
rect 8200 832 8210 910
rect 8228 906 8667 935
rect 8228 884 8304 906
rect 8310 899 8667 906
rect 8692 933 9517 935
rect 9519 933 9525 945
rect 9539 933 9553 973
rect 8692 911 9502 933
rect 9531 929 9553 933
rect 9573 962 9614 986
rect 9573 950 9607 962
rect 9610 950 9614 962
rect 9573 946 9619 950
rect 9644 946 9648 986
rect 9687 984 11233 986
rect 9573 942 9678 946
rect 9573 933 9619 942
rect 9573 929 9607 933
rect 9514 911 9553 929
rect 8310 884 8378 899
rect 8597 888 8681 899
rect 8514 884 8670 888
rect 8228 882 8670 884
rect 8692 882 9500 911
rect 8234 832 8268 882
rect 8200 826 8268 832
rect 8599 831 8628 882
rect 8633 876 8670 882
rect 8674 876 9500 882
rect 8633 865 9500 876
rect 8692 829 9500 865
rect 9513 905 9553 911
rect 9608 918 9621 928
rect 9644 918 9648 942
rect 9653 918 9678 942
rect 9608 914 9678 918
rect 9608 912 9641 914
rect 9644 912 9648 914
rect 9608 907 9645 912
rect 9513 895 9548 905
rect 9608 895 9641 907
rect 9513 845 9544 895
rect 9574 861 9579 895
rect 9608 862 9621 895
rect 8692 828 8796 829
rect 8966 828 9500 829
rect 6616 825 8137 826
rect 6616 816 6965 825
rect 6145 779 6180 816
rect 6265 804 6318 816
rect 6344 805 6377 816
rect 6404 804 6416 816
rect 6265 798 6416 804
rect 6265 795 6318 798
rect 6265 789 6349 795
rect 6184 779 6213 788
rect 6287 779 6337 789
rect 6404 788 6416 798
rect 6427 788 6450 816
rect 6344 779 6388 788
rect 6404 779 6450 788
rect 6461 779 6495 816
rect 6514 804 6548 816
rect 6562 808 6971 816
rect 6145 768 6389 779
rect 6145 754 6378 768
rect 5814 740 5882 744
rect 5740 726 5814 740
rect 5872 738 5882 740
rect 5908 740 5909 754
rect 6054 740 6122 754
rect 6145 745 6364 754
rect 6404 745 6495 779
rect 6145 741 6180 745
rect 6287 741 6318 745
rect 5908 726 6054 740
rect 6145 739 6318 741
rect 6404 741 6405 745
rect 6427 741 6450 745
rect 6461 741 6495 745
rect 6111 726 6126 738
rect 5740 723 6126 726
rect 5776 706 6126 723
rect 6145 727 6287 739
rect 6303 727 6386 739
rect 6145 726 6386 727
rect 6404 727 6495 741
rect 6504 727 6548 804
rect 6594 795 6662 808
rect 6594 783 6660 795
rect 6696 783 6762 808
rect 6830 804 6971 808
rect 6997 804 6999 815
rect 7028 810 7031 815
rect 7050 811 7088 816
rect 7144 815 8137 825
rect 6796 789 6971 804
rect 7020 799 7031 810
rect 6997 789 7031 799
rect 7062 789 7065 804
rect 7073 801 7088 811
rect 7119 799 7131 811
rect 7085 789 7131 799
rect 7144 804 8132 815
rect 7144 803 8126 804
rect 7144 792 8137 803
rect 8164 792 8340 826
rect 8692 820 9500 828
rect 7144 789 8024 792
rect 6594 760 6626 783
rect 6628 779 6706 783
rect 6592 750 6626 760
rect 6638 774 6706 779
rect 6708 774 6716 783
rect 6796 778 8024 789
rect 6796 774 7131 778
rect 6638 754 6742 774
rect 6830 772 7131 774
rect 6830 760 6917 772
rect 6634 750 6744 754
rect 6592 738 6754 750
rect 6796 738 6917 760
rect 6931 755 7131 772
rect 7134 772 8024 778
rect 7134 766 7168 772
rect 7134 755 7179 766
rect 7194 755 7286 772
rect 6610 727 6754 738
rect 6830 727 6917 738
rect 6404 726 6550 727
rect 6580 726 6754 727
rect 6784 726 6917 727
rect 6962 726 6971 755
rect 6974 754 7031 755
rect 6997 741 7031 754
rect 7062 754 7119 755
rect 7134 754 7178 755
rect 7194 754 7240 755
rect 6997 738 7043 741
rect 7062 738 7065 754
rect 7085 738 7119 754
rect 7152 744 7178 754
rect 7152 738 7168 744
rect 7199 738 7240 754
rect 6991 726 7043 738
rect 4616 702 4630 703
rect 4633 702 4729 703
rect 4616 698 4704 702
rect 3878 672 4402 698
rect 4548 672 4704 698
rect 4718 692 4729 702
rect 4765 693 4931 703
rect 4953 702 5005 703
rect 4765 672 4923 693
rect 4953 692 4964 702
rect 4994 692 5005 702
rect 6145 698 6179 726
rect 6245 706 6260 726
rect 5740 672 6179 698
rect 6241 687 6303 706
rect 6337 687 6399 706
rect 6241 672 6399 687
rect 6461 698 6495 726
rect 6504 698 6917 726
rect 6985 721 7043 726
rect 7079 726 7125 738
rect 7079 721 7131 726
rect 7020 710 7043 721
rect 6461 696 6917 698
rect 6461 672 6830 696
rect 6847 672 6917 696
rect 6963 693 7153 710
rect 7041 683 7075 693
rect 7199 672 7233 738
rect 7252 672 7286 755
rect 7294 770 7340 772
rect 7364 770 7408 772
rect 7412 770 7488 772
rect 7294 762 7488 770
rect 7526 770 7542 772
rect 7549 770 8024 772
rect 8036 770 8040 792
rect 8060 788 8110 792
rect 8095 773 8110 788
rect 8200 770 8210 792
rect 7294 754 7472 762
rect 7294 746 7454 754
rect 7484 746 7488 757
rect 7526 755 8024 770
rect 7526 754 7560 755
rect 7294 738 7488 746
rect 7300 736 7334 738
rect 7354 736 7400 738
rect 7454 736 7488 738
rect 7534 736 7560 754
rect 7568 736 8024 755
rect 8064 762 8210 770
rect 8064 738 8220 762
rect 8164 736 8220 738
rect 8234 736 8268 792
rect 7300 719 8268 736
rect 8272 722 8298 792
rect 8305 773 8340 792
rect 8364 773 8394 816
rect 8728 810 9500 820
rect 9514 810 9534 845
rect 9550 810 9560 820
rect 9653 810 9678 914
rect 9687 904 9852 984
rect 9854 904 9884 984
rect 9930 904 9960 984
rect 10001 968 11233 984
rect 11244 991 11261 1002
rect 11334 1006 11362 1041
rect 11334 991 11377 1006
rect 11244 968 11246 991
rect 11460 986 12631 1041
rect 11252 974 11386 978
rect 11460 968 11547 986
rect 10001 932 11547 968
rect 11549 969 12631 986
rect 12639 1111 13466 1132
rect 13478 1111 13498 1132
rect 12639 1107 13464 1111
rect 13477 1107 13508 1111
rect 13560 1107 16595 1132
rect 12639 1094 16595 1107
rect 12639 1073 14792 1094
rect 12639 1044 13464 1073
rect 13477 1061 13543 1073
rect 13477 1055 13539 1061
rect 13477 1045 13512 1055
rect 13478 1044 13512 1045
rect 13560 1044 14792 1073
rect 14841 1044 14846 1094
rect 14872 1059 14899 1094
rect 14948 1066 14987 1094
rect 14857 1044 14899 1059
rect 12639 1027 13478 1044
rect 12639 1023 13464 1027
rect 13495 1023 13512 1044
rect 13544 1040 14792 1044
rect 14853 1040 14887 1042
rect 14941 1040 14975 1042
rect 15049 1041 16595 1094
rect 13532 1023 14792 1040
rect 12639 1011 13481 1023
rect 12639 969 13498 1011
rect 11549 945 13498 969
rect 13503 973 13512 1023
rect 13537 1021 14792 1023
rect 15055 1021 15089 1041
rect 15108 1021 15123 1041
rect 13537 986 15197 1021
rect 15210 1002 15225 1041
rect 11549 935 13481 945
rect 10001 931 11530 932
rect 10026 906 10052 931
rect 10056 906 10076 931
rect 9687 892 9880 904
rect 9687 889 9861 892
rect 9930 889 9975 904
rect 9687 884 9852 889
rect 10056 884 10090 906
rect 9687 858 9882 884
rect 9687 848 9888 858
rect 9932 848 10090 884
rect 9687 842 10090 848
rect 9687 838 9930 842
rect 9932 838 10090 842
rect 9687 816 10090 838
rect 9687 810 9852 816
rect 8728 809 9560 810
rect 8692 794 9560 809
rect 8692 773 8816 794
rect 8966 793 9560 794
rect 9562 804 9852 810
rect 9858 804 9862 816
rect 9872 808 9970 816
rect 9872 804 9944 808
rect 9562 802 9944 804
rect 9562 793 9930 802
rect 8966 792 9930 793
rect 8966 776 9918 792
rect 7300 702 7686 719
rect 7366 680 7400 702
rect 7454 685 7500 702
rect 7454 680 7488 685
rect 7534 672 7560 702
rect 7568 698 7686 702
rect 7723 706 7746 719
rect 7723 698 7769 706
rect 7568 685 7769 698
rect 7568 672 7723 685
rect 7735 672 7769 685
rect 7789 672 7792 719
rect 7811 710 7834 719
rect 7811 700 7842 710
rect 7823 672 7842 700
rect 7882 702 8268 719
rect 7882 672 8024 702
rect 8132 690 8198 702
rect 8222 700 8240 702
rect 8070 672 8260 674
rect 8306 672 8340 773
rect 8359 739 8510 773
rect 8582 739 8816 773
rect 8359 726 8394 739
rect 8359 672 8393 726
rect 8464 722 8498 739
rect 8675 730 8816 739
rect 8675 693 8681 730
rect 8692 698 8762 730
rect 8782 729 8816 730
rect 8848 729 8958 764
rect 9016 729 9084 776
rect 9124 775 9125 776
rect 9312 775 9625 776
rect 8782 728 9084 729
rect 9097 759 9625 775
rect 9632 774 9918 776
rect 9632 759 9856 774
rect 9097 756 9483 759
rect 9097 740 9102 756
rect 9124 741 9483 756
rect 9124 740 9131 741
rect 9097 729 9132 740
rect 9270 729 9300 731
rect 9335 729 9483 741
rect 9514 740 9548 759
rect 9704 744 9856 759
rect 9872 754 9918 774
rect 9972 774 9982 804
rect 10004 788 10090 816
rect 9972 754 10006 774
rect 10018 754 10090 788
rect 10109 884 10143 931
rect 10211 884 10224 931
rect 10308 884 10342 931
rect 10370 898 11530 931
rect 11549 910 11971 935
rect 11984 922 12030 935
rect 10370 884 11548 898
rect 10109 816 10269 884
rect 10300 878 11548 884
rect 10300 872 10624 878
rect 10676 872 11548 878
rect 10300 851 10456 872
rect 10299 838 10456 851
rect 10459 838 10638 872
rect 10642 838 11548 872
rect 10299 836 10624 838
rect 10300 816 10624 836
rect 10718 835 11548 838
rect 11549 838 11974 910
rect 11984 906 12062 922
rect 11996 905 12062 906
rect 12084 911 12118 935
rect 11996 888 12072 905
rect 12084 888 12096 911
rect 12106 894 12118 911
rect 12140 888 12152 910
rect 11996 872 12008 888
rect 12028 876 12072 888
rect 12090 876 12128 880
rect 11549 835 11971 838
rect 10718 826 11971 835
rect 12000 826 12004 860
rect 12028 854 12074 876
rect 12024 844 12074 854
rect 12024 838 12086 844
rect 12024 826 12074 838
rect 12164 832 12174 910
rect 12192 906 12631 935
rect 12192 884 12268 906
rect 12274 899 12631 906
rect 12656 933 13481 935
rect 13483 933 13489 945
rect 13503 933 13517 973
rect 12656 911 13466 933
rect 13495 929 13517 933
rect 13537 962 13578 986
rect 13537 950 13571 962
rect 13574 950 13578 962
rect 13537 946 13583 950
rect 13608 946 13612 986
rect 13651 984 15197 986
rect 13537 942 13642 946
rect 13537 933 13583 942
rect 13537 929 13571 933
rect 13478 911 13517 929
rect 12274 884 12342 899
rect 12561 888 12645 899
rect 12478 884 12634 888
rect 12192 882 12634 884
rect 12656 882 13464 911
rect 12198 832 12232 882
rect 12164 826 12232 832
rect 12563 831 12592 882
rect 12597 876 12634 882
rect 12638 876 13464 882
rect 12597 865 13464 876
rect 12656 829 13464 865
rect 13477 905 13517 911
rect 13572 918 13585 928
rect 13608 918 13612 942
rect 13617 918 13642 942
rect 13572 914 13642 918
rect 13572 912 13605 914
rect 13608 912 13612 914
rect 13572 907 13609 912
rect 13477 895 13512 905
rect 13572 895 13605 907
rect 13477 845 13508 895
rect 13538 861 13543 895
rect 13572 862 13585 895
rect 12656 828 12760 829
rect 12930 828 13464 829
rect 10718 825 12101 826
rect 10680 816 10714 822
rect 10718 816 10881 825
rect 9704 740 9852 744
rect 9872 740 9873 754
rect 10018 740 10086 754
rect 10109 741 10144 816
rect 10229 804 10282 816
rect 10308 805 10341 816
rect 10368 804 10380 816
rect 10229 798 10380 804
rect 10229 795 10282 798
rect 10229 789 10313 795
rect 10251 788 10301 789
rect 10148 754 10177 788
rect 10251 755 10282 788
rect 10308 755 10352 788
rect 10251 754 10352 755
rect 10251 749 10313 754
rect 10251 741 10282 749
rect 9097 728 9483 729
rect 8794 698 8796 728
rect 8870 726 8928 728
rect 8870 698 8936 726
rect 9044 698 9078 728
rect 9097 698 9131 728
rect 9197 702 9212 728
rect 9270 706 9300 728
rect 9335 723 9483 728
rect 9704 726 9778 740
rect 9836 738 9846 740
rect 9872 726 10018 740
rect 10109 739 10282 741
rect 10326 744 10352 754
rect 10368 754 10380 798
rect 10326 739 10342 744
rect 10368 741 10369 754
rect 10391 741 10414 816
rect 10425 741 10459 816
rect 10478 804 10512 816
rect 10075 726 10090 738
rect 9704 723 10090 726
rect 9255 702 9300 706
rect 8692 692 9239 698
rect 8692 677 8888 692
rect 8675 672 8888 677
rect 8918 672 9239 692
rect 9255 673 9289 702
rect 9312 698 9339 707
rect 9413 698 9447 706
rect 9704 698 9737 723
rect 9740 706 10090 723
rect 10109 726 10350 739
rect 10368 727 10459 741
rect 10468 727 10512 804
rect 10558 783 10624 816
rect 10660 783 10726 816
rect 10558 745 10590 783
rect 10592 779 10670 783
rect 10602 774 10670 779
rect 10602 754 10706 774
rect 10586 738 10590 745
rect 10598 736 10708 754
rect 10602 727 10708 736
rect 10794 727 10881 816
rect 10368 726 10881 727
rect 10926 726 10935 816
rect 10992 810 10995 815
rect 11014 811 11052 816
rect 10984 799 10995 810
rect 11026 799 11029 804
rect 11037 801 11052 811
rect 11060 811 11072 816
rect 11108 815 12101 825
rect 11060 799 11095 811
rect 10961 788 10995 799
rect 11015 788 11037 799
rect 11049 788 11095 799
rect 11108 804 12096 815
rect 11108 803 12090 804
rect 11108 792 12101 803
rect 12128 792 12304 826
rect 12656 820 13464 828
rect 11108 788 11988 792
rect 10938 754 10995 788
rect 10961 741 10995 754
rect 11026 754 11083 788
rect 11098 772 11988 788
rect 11098 754 11142 772
rect 11158 754 11204 772
rect 10961 738 11007 741
rect 11026 738 11029 754
rect 11049 738 11083 754
rect 11116 744 11142 754
rect 11116 738 11132 744
rect 11163 738 11204 754
rect 10955 726 11007 738
rect 10109 706 10143 726
rect 10109 698 10124 706
rect 9305 673 9483 698
rect 9278 672 9483 673
rect 9704 672 10124 698
rect 10205 672 10363 706
rect 10425 704 10459 726
rect 10426 700 10459 704
rect 10434 698 10459 700
rect 10468 698 10512 726
rect 10620 706 10624 726
rect 10636 706 10670 719
rect 10620 702 10672 706
rect 10718 700 10728 726
rect 10794 698 10881 726
rect 10949 721 11007 726
rect 11043 726 11089 738
rect 11043 721 11095 726
rect 10984 710 11007 721
rect 10434 696 10881 698
rect 10434 672 10794 696
rect 10811 672 10881 696
rect 10927 693 11117 710
rect 11005 683 11039 693
rect 11163 672 11197 738
rect 11216 672 11250 772
rect 11258 758 11304 772
rect 11328 758 11372 772
rect 11376 762 11452 772
rect 11376 758 11436 762
rect 11258 738 11284 758
rect 11318 754 11400 758
rect 11402 754 11436 758
rect 11318 743 11376 754
rect 11318 726 11364 743
rect 11448 726 11452 757
rect 11513 755 11988 772
rect 12000 770 12004 792
rect 12024 788 12074 792
rect 12059 773 12074 788
rect 12164 770 12174 792
rect 11330 716 11364 726
rect 11438 710 11464 726
rect 11330 680 11364 710
rect 11418 685 11464 710
rect 11418 680 11452 685
rect 11498 672 11524 755
rect 11532 736 11988 755
rect 12028 762 12174 770
rect 12028 738 12184 762
rect 12128 736 12184 738
rect 12198 736 12232 792
rect 11532 719 12232 736
rect 12236 722 12262 792
rect 12269 773 12304 792
rect 12328 773 12358 816
rect 12692 810 13464 820
rect 13478 810 13498 845
rect 13514 810 13524 820
rect 13617 810 13642 914
rect 13651 904 13816 984
rect 13818 904 13848 984
rect 13894 904 13924 984
rect 13965 968 15197 984
rect 15208 991 15225 1002
rect 15298 1006 15326 1041
rect 15298 991 15341 1006
rect 15208 968 15210 991
rect 15424 986 16595 1041
rect 15216 974 15350 978
rect 15424 968 15511 986
rect 13965 932 15511 968
rect 15513 969 16595 986
rect 16603 1233 17316 1238
rect 17341 1233 17411 1238
rect 16603 1214 17411 1233
rect 17632 1218 17798 1250
rect 17632 1214 17780 1218
rect 16603 1204 17780 1214
rect 16603 1197 17429 1204
rect 17490 1197 17780 1204
rect 16603 1180 17780 1197
rect 16603 1163 17553 1180
rect 16603 1023 17428 1163
rect 17632 1159 17780 1180
rect 17536 1118 17549 1128
rect 17536 1112 17598 1118
rect 17445 1095 17503 1101
rect 17441 1078 17475 1095
rect 17502 1078 17507 1095
rect 17441 1061 17507 1078
rect 17536 1078 17552 1112
rect 17581 1078 17602 1112
rect 17536 1072 17598 1078
rect 17536 1062 17549 1072
rect 17615 1069 17780 1159
rect 17814 1150 17872 1156
rect 17814 1116 17826 1150
rect 17814 1110 17872 1116
rect 17445 1055 17503 1061
rect 17508 1040 17541 1044
rect 17496 1028 17541 1040
rect 17496 1027 17542 1028
rect 17496 1023 17504 1027
rect 16603 1011 17429 1023
rect 17508 1011 17542 1027
rect 16603 969 17462 1011
rect 15513 952 16578 969
rect 16620 953 17462 969
rect 15513 935 16232 952
rect 13965 931 15494 932
rect 13990 906 14016 931
rect 14020 906 14040 931
rect 13651 892 13844 904
rect 13651 889 13825 892
rect 13894 889 13939 904
rect 13651 884 13816 889
rect 14020 884 14054 906
rect 13651 858 13846 884
rect 13651 848 13852 858
rect 13896 848 14054 884
rect 13651 842 14054 848
rect 13651 838 13894 842
rect 13896 838 14054 842
rect 13651 816 14054 838
rect 13651 810 13816 816
rect 12692 809 13524 810
rect 12656 794 13524 809
rect 12656 773 12780 794
rect 12930 793 13524 794
rect 13526 804 13816 810
rect 13822 804 13826 816
rect 13836 808 13934 816
rect 13836 804 13908 808
rect 13526 802 13908 804
rect 13526 793 13894 802
rect 12930 792 13894 793
rect 12930 776 13882 792
rect 11532 698 11619 719
rect 11687 706 11710 719
rect 11687 698 11733 706
rect 11532 685 11733 698
rect 11532 672 11687 685
rect 11699 672 11733 685
rect 11753 672 11756 719
rect 11775 710 11798 719
rect 11775 700 11806 710
rect 11787 672 11806 700
rect 11846 702 12232 719
rect 11846 672 11988 702
rect 12096 690 12162 702
rect 12186 700 12204 702
rect 12034 672 12224 674
rect 12270 672 12304 773
rect 12323 739 12474 773
rect 12546 739 12780 773
rect 12323 726 12358 739
rect 12323 672 12357 726
rect 12428 722 12462 739
rect 12639 730 12780 739
rect 12639 693 12645 730
rect 12656 698 12726 730
rect 12746 729 12780 730
rect 12812 729 12922 764
rect 12980 729 13048 776
rect 13088 775 13089 776
rect 13276 775 13589 776
rect 12746 728 13048 729
rect 13061 759 13589 775
rect 13596 774 13882 776
rect 13596 759 13820 774
rect 13061 756 13447 759
rect 13061 740 13066 756
rect 13088 741 13447 756
rect 13088 740 13095 741
rect 13061 729 13096 740
rect 13234 729 13264 731
rect 13299 729 13447 741
rect 13478 740 13512 759
rect 13668 744 13820 759
rect 13836 754 13882 774
rect 13936 774 13946 804
rect 13968 788 14054 816
rect 13936 754 13970 774
rect 13982 754 14054 788
rect 14073 884 14107 931
rect 14175 884 14188 931
rect 14272 884 14306 931
rect 14334 898 15494 931
rect 14334 884 15512 898
rect 14073 816 14233 884
rect 14264 878 15512 884
rect 14264 872 14588 878
rect 14640 872 15512 878
rect 14264 851 14420 872
rect 14263 838 14420 851
rect 14423 838 14602 872
rect 14606 838 15512 872
rect 14263 836 14588 838
rect 14264 816 14588 836
rect 14682 835 15512 838
rect 15513 835 15935 935
rect 15948 880 15953 935
rect 16156 882 16232 935
rect 16251 935 16578 952
rect 16595 945 17462 953
rect 17501 962 17542 1011
rect 17501 950 17535 962
rect 17501 945 17547 950
rect 16595 935 17429 945
rect 16251 918 16595 935
rect 16620 933 17429 935
rect 17502 933 17547 945
rect 16251 899 16578 918
rect 16525 882 16578 899
rect 16620 882 17428 933
rect 17502 929 17535 933
rect 17536 918 17549 928
rect 17536 912 17598 918
rect 17536 907 17573 912
rect 17445 895 17503 901
rect 17536 895 17569 907
rect 15948 876 15988 880
rect 16054 876 16094 880
rect 14682 826 15935 835
rect 15980 844 16038 860
rect 15980 838 16050 844
rect 15980 826 16004 838
rect 16162 832 16196 882
rect 16602 865 17428 882
rect 16138 826 16196 832
rect 16620 829 17428 865
rect 17441 861 17475 895
rect 17502 861 17507 895
rect 17536 878 17552 895
rect 17581 878 17602 912
rect 17615 889 17798 1069
rect 17536 872 17598 878
rect 17536 862 17549 872
rect 17445 855 17503 861
rect 17615 844 17780 889
rect 16894 827 17428 829
rect 14682 825 15953 826
rect 14644 816 14678 822
rect 14682 816 14845 825
rect 13668 740 13816 744
rect 13836 740 13837 754
rect 13982 740 14050 754
rect 14073 741 14108 816
rect 14193 804 14246 816
rect 14272 805 14305 816
rect 14332 804 14344 816
rect 14193 798 14344 804
rect 14193 795 14246 798
rect 14193 789 14277 795
rect 14215 788 14265 789
rect 14112 754 14141 788
rect 14215 755 14246 788
rect 14272 755 14316 788
rect 14215 754 14316 755
rect 14215 749 14277 754
rect 14215 741 14246 749
rect 13061 728 13447 729
rect 12758 698 12760 728
rect 12834 726 12892 728
rect 12834 698 12900 726
rect 13008 698 13042 728
rect 13061 698 13095 728
rect 13161 702 13176 728
rect 13234 706 13264 728
rect 13299 723 13447 728
rect 13668 726 13742 740
rect 13800 738 13810 740
rect 13836 726 13982 740
rect 14073 739 14246 741
rect 14290 744 14316 754
rect 14332 754 14344 798
rect 14290 739 14306 744
rect 14332 741 14333 754
rect 14355 741 14378 816
rect 14389 741 14423 816
rect 14442 804 14476 816
rect 14039 726 14054 738
rect 13668 723 14054 726
rect 13219 702 13264 706
rect 12656 692 13203 698
rect 12656 677 12852 692
rect 12639 672 12852 677
rect 12882 672 13203 692
rect 13219 673 13253 702
rect 13276 698 13303 707
rect 13377 698 13411 706
rect 13668 698 13701 723
rect 13704 706 14054 723
rect 14073 726 14314 739
rect 14332 727 14423 741
rect 14432 727 14476 804
rect 14522 783 14588 816
rect 14624 783 14690 816
rect 14522 745 14554 783
rect 14556 779 14634 783
rect 14566 774 14634 779
rect 14566 754 14670 774
rect 14550 738 14554 745
rect 14562 736 14672 754
rect 14566 727 14672 736
rect 14758 727 14845 816
rect 14332 726 14845 727
rect 14890 726 14899 816
rect 14956 810 14959 815
rect 14978 811 15016 816
rect 14948 799 14959 810
rect 14990 799 14993 804
rect 15001 801 15016 811
rect 15024 811 15036 816
rect 15024 799 15059 811
rect 14925 788 14959 799
rect 14979 788 15001 799
rect 15013 788 15059 799
rect 15072 792 15953 825
rect 15977 815 16196 826
rect 15988 803 16196 815
rect 15977 798 16196 803
rect 15977 792 16172 798
rect 16233 792 16268 826
rect 16656 809 16691 827
rect 15072 788 15952 792
rect 14902 754 14959 788
rect 14925 741 14959 754
rect 14990 754 15047 788
rect 15062 772 15952 788
rect 15062 754 15106 772
rect 15122 754 15168 772
rect 14925 738 14971 741
rect 14990 738 14993 754
rect 15013 738 15047 754
rect 15080 744 15106 754
rect 15080 738 15096 744
rect 15127 738 15168 754
rect 14919 726 14971 738
rect 14073 706 14107 726
rect 14073 698 14088 706
rect 13269 673 13447 698
rect 13242 672 13447 673
rect 13668 672 14088 698
rect 14169 672 14327 706
rect 14389 704 14423 726
rect 14390 700 14423 704
rect 14398 698 14423 700
rect 14432 698 14476 726
rect 14584 706 14588 726
rect 14600 706 14634 719
rect 14584 702 14636 706
rect 14682 700 14692 726
rect 14758 698 14845 726
rect 14913 721 14971 726
rect 15007 726 15053 738
rect 15007 721 15059 726
rect 14948 710 14971 721
rect 14398 696 14845 698
rect 14398 672 14758 696
rect 14775 672 14845 696
rect 14891 693 15081 710
rect 14969 683 15003 693
rect 15127 672 15161 738
rect 15180 672 15214 772
rect 15222 758 15268 772
rect 15292 758 15336 772
rect 15340 762 15416 772
rect 15340 758 15400 762
rect 15222 738 15248 758
rect 15282 754 15364 758
rect 15366 754 15400 758
rect 15282 743 15340 754
rect 15282 726 15328 743
rect 15412 726 15416 757
rect 15477 755 15952 772
rect 15294 716 15328 726
rect 15402 710 15428 726
rect 15294 680 15328 710
rect 15382 685 15428 710
rect 15382 680 15416 685
rect 15462 672 15488 755
rect 15496 736 15952 755
rect 16234 773 16268 792
rect 16620 794 16691 809
rect 15496 719 16157 736
rect 15496 698 15583 719
rect 15651 706 15674 719
rect 15651 698 15697 706
rect 15496 685 15697 698
rect 15496 672 15651 685
rect 15663 672 15697 685
rect 15717 672 15720 719
rect 15739 710 15762 719
rect 15739 700 15770 710
rect 15751 672 15770 700
rect 15810 706 16157 719
rect 15810 702 16196 706
rect 16234 702 16250 773
rect 674 671 4551 672
rect 674 670 1088 671
rect 1097 670 4551 671
rect 674 666 4551 670
rect 674 638 3928 666
rect 949 636 983 638
rect 1002 636 1036 638
rect 1042 636 1070 638
rect 1196 636 1241 638
rect 448 601 482 632
rect 536 615 562 632
rect 633 601 648 632
rect 654 613 667 632
rect 900 614 1042 636
rect 1076 614 1144 636
rect 900 613 1144 614
rect 654 604 1144 613
rect 1196 614 1296 636
rect 1318 629 3608 638
rect 3664 629 3694 638
rect 3764 629 3782 638
rect 3878 629 3928 638
rect 3931 629 3965 666
rect 4020 639 4281 666
rect 4300 639 4551 666
rect 4616 651 5567 672
rect 5838 652 6064 672
rect 6111 666 7686 672
rect 6111 653 7655 666
rect 6111 652 6179 653
rect 5776 651 6179 652
rect 4616 639 5591 651
rect 4020 638 5591 639
rect 5712 639 6179 651
rect 6287 650 6353 653
rect 6427 650 7655 653
rect 6193 639 7655 650
rect 7701 639 7852 672
rect 7882 671 8505 672
rect 7882 666 8531 671
rect 5712 638 7852 639
rect 7942 661 8531 666
rect 7942 653 8497 661
rect 8501 653 8531 661
rect 7942 638 8531 653
rect 1318 614 3971 629
rect 1196 604 3971 614
rect 654 601 800 604
rect 854 601 983 604
rect 1002 601 1088 604
rect 1196 602 1254 604
rect 1284 602 3971 604
rect 1196 601 3971 602
rect 236 600 3971 601
rect 448 599 482 600
rect 633 598 648 600
rect 654 579 800 600
rect 854 579 983 600
rect 1002 573 1088 600
rect 1196 574 1254 600
rect 1284 576 3971 600
rect 4033 576 4091 594
rect 4121 576 4179 594
rect 4266 576 4281 638
rect 4300 576 4334 638
rect 1284 574 4340 576
rect 1196 573 4340 574
rect 236 572 4340 573
rect 1002 568 1088 572
rect 1196 568 1254 572
rect 1284 568 4340 572
rect 1002 537 1030 568
rect 1318 560 4340 568
rect 1036 543 1088 560
rect 1113 549 1169 560
rect 1196 554 1318 560
rect 1196 550 1322 554
rect 1335 550 4340 560
rect 1124 537 1158 549
rect 1196 543 4340 550
rect 1002 526 1041 537
rect 1113 526 1169 537
rect 1200 532 4340 543
rect 1200 526 1388 532
rect 1335 516 1388 526
rect 932 482 936 516
rect 1234 492 1388 516
rect 1467 496 1585 507
rect 1335 490 1388 492
rect 1371 484 1372 490
rect 1478 484 1574 496
rect 1668 494 4340 532
rect 1371 478 1383 484
rect 1467 478 1585 484
rect 1371 473 1586 478
rect 1042 410 1044 444
rect 1337 439 1586 444
rect 1668 437 2881 494
rect 2949 444 2953 494
rect 2980 459 3007 494
rect 3056 466 3095 494
rect 2965 444 3007 459
rect 2961 440 2995 442
rect 3049 440 3083 442
rect 3157 441 4340 494
rect 1704 386 2881 437
rect 2927 406 3117 408
rect 816 340 820 374
rect 1374 346 1376 374
rect 1342 340 1376 346
rect 1884 342 1894 376
rect 1908 342 1928 376
rect 2109 374 2195 386
rect 2266 378 2296 386
rect 2380 378 2414 386
rect 2255 374 2307 378
rect 2369 374 2425 378
rect 2444 374 2459 386
rect 2109 367 2459 374
rect 2478 382 2512 386
rect 2520 384 2540 386
rect 2518 382 2540 384
rect 2586 382 2720 386
rect 2794 382 2881 386
rect 2478 374 2881 382
rect 2478 348 2512 374
rect 2528 364 2540 374
rect 2528 358 2530 364
rect 2794 348 2881 374
rect 2993 397 3051 403
rect 2993 363 3005 397
rect 2993 357 3051 363
rect 1640 235 1650 342
rect 1086 192 1088 230
rect 1668 207 1678 342
rect 2478 340 2881 348
rect 3056 347 3086 386
rect 3170 378 3197 441
rect 3163 340 3197 378
rect 3216 378 3231 441
rect 3318 402 3333 441
rect 3316 391 3333 402
rect 3406 406 3434 441
rect 3406 391 3449 406
rect 2098 337 2539 340
rect 2575 337 2627 340
rect 2779 337 2881 340
rect 2098 333 2528 337
rect 2114 306 2124 333
rect 2138 306 2158 333
rect 2478 325 2528 333
rect 2586 325 2616 337
rect 2478 314 2539 325
rect 2575 314 2627 325
rect 2788 319 2881 337
rect 2667 314 2881 319
rect 2788 306 2800 314
rect 2810 310 2872 314
rect 2810 306 2881 310
rect 3154 306 3163 329
rect 3170 306 3214 340
rect 3216 306 3242 378
rect 3316 360 3318 391
rect 3532 386 4340 441
rect 4446 454 4504 460
rect 4446 420 4458 454
rect 4446 414 4504 420
rect 3324 374 3458 378
rect 3358 344 3360 360
rect 3358 340 3424 344
rect 2811 295 2881 306
rect 3170 301 3197 306
rect 3216 301 3231 306
rect 3358 301 3360 340
rect 3532 301 3619 386
rect 3665 305 3670 386
rect 3693 333 3698 386
rect 3775 359 3782 386
rect 3786 359 3824 378
rect 3838 374 3888 386
rect 3768 345 3824 359
rect 3752 333 3824 345
rect 3825 333 3833 374
rect 3870 364 3882 374
rect 3870 358 3872 364
rect 3895 335 4340 386
rect 3693 329 3739 333
rect 3752 329 3833 333
rect 3752 325 3755 329
rect 3776 325 3796 329
rect 3693 306 3802 325
rect 3665 301 3855 305
rect 2951 295 3619 301
rect 2732 282 2748 288
rect 2714 272 2758 282
rect 2714 262 2764 272
rect 2738 256 2764 262
rect 2738 254 2758 256
rect 2714 238 2758 254
rect 2732 228 2758 238
rect 2732 222 2748 228
rect 2811 225 3619 295
rect 3727 272 3793 291
rect 3920 270 3935 335
rect 1124 156 1126 192
rect 1846 188 1850 216
rect 1884 164 1894 188
rect 1908 164 1928 188
rect 1884 154 1928 164
rect 1944 154 1956 216
rect 2076 188 2090 216
rect 2342 188 2354 216
rect 2114 164 2128 188
rect 2138 164 2158 188
rect 2114 154 2158 164
rect 2380 164 2392 188
rect 2404 164 2424 188
rect 2380 154 2424 164
rect 2440 154 2452 216
rect 2866 188 2878 216
rect 3132 188 3144 216
rect 3180 189 3619 225
rect 3636 189 3653 204
rect 3694 189 3708 216
rect 3901 189 3935 270
rect 3180 188 3935 189
rect 2904 164 2916 188
rect 2928 164 2948 188
rect 2904 154 2948 164
rect 3170 172 3608 188
rect 3625 178 3935 188
rect 3170 164 3182 172
rect 3194 164 3214 172
rect 3170 154 3214 164
rect 3230 154 3242 172
rect 3400 164 3414 172
rect 3424 164 3444 172
rect 3400 154 3444 164
rect 3462 154 3472 172
rect 3585 155 3608 172
rect 3636 155 3935 178
rect 3954 155 3988 335
rect 4264 282 4340 335
rect 4633 318 4703 638
rect 4827 600 4861 601
rect 4815 401 4873 407
rect 4815 367 4827 401
rect 4815 361 4873 367
rect 4633 282 4686 318
rect 5004 289 5019 638
rect 4979 265 5019 289
rect 5038 616 5073 638
rect 5134 616 5292 638
rect 5353 616 5388 638
rect 5776 633 5811 638
rect 5038 265 5072 616
rect 5354 597 5388 616
rect 5740 618 5811 633
rect 5038 235 5053 265
rect 5134 235 5292 246
rect 5373 236 5388 597
rect 5033 231 5053 235
rect 5129 212 5292 235
rect 5348 212 5388 236
rect 5407 563 5442 597
rect 5407 212 5441 563
rect 5553 495 5611 501
rect 5553 461 5565 495
rect 5553 455 5611 461
rect 5553 295 5611 301
rect 5553 261 5565 295
rect 5604 261 5611 295
rect 5553 255 5611 261
rect 5632 227 5639 329
rect 5129 201 5287 212
rect 5348 201 5383 212
rect 5349 182 5383 201
rect 5407 182 5437 212
rect 5740 201 5810 618
rect 5894 482 5898 584
rect 5922 550 5980 556
rect 5922 516 5934 550
rect 5922 510 5980 516
rect 5723 193 5810 201
rect 5503 182 5661 193
rect 3636 154 3680 155
rect 3694 154 3708 155
rect 1902 144 1928 154
rect 2132 144 2158 154
rect 2398 144 2424 154
rect 2922 144 2948 154
rect 3188 144 3214 154
rect 3418 144 3444 154
rect 3654 144 3680 154
rect 1902 138 1918 144
rect 2132 138 2148 144
rect 2398 138 2414 144
rect 2922 138 2938 144
rect 3188 138 3204 144
rect 3418 138 3434 144
rect 3654 138 3670 144
rect 3954 126 3982 155
rect 3954 121 3969 126
rect 3179 47 3653 72
rect 3187 38 3653 47
rect 3241 4 3591 11
rect 2050 -38 2086 -12
rect 2436 -38 2472 -12
rect 3205 -38 3241 -12
rect 3275 -38 3557 4
rect 3591 -38 3914 -12
rect 2086 -39 2867 -38
rect 1748 -72 2867 -39
rect 3241 -51 3591 -38
rect 3888 -42 3914 -38
rect 3610 -51 3888 -42
rect 3207 -57 3888 -51
rect 3207 -58 3309 -57
rect 3349 -58 3483 -57
rect 3523 -58 3888 -57
rect 3925 -58 3960 -42
rect 3205 -66 3960 -58
rect 2050 -93 2120 -72
rect 1717 -106 1804 -93
rect 1838 -106 2120 -93
rect 1762 -126 1792 -106
rect 1850 -107 2032 -106
rect 1837 -120 2032 -107
rect 1813 -126 2032 -120
rect 2050 -126 2120 -106
rect 2140 -106 2228 -72
rect 2266 -91 2455 -72
rect 2489 -91 2771 -72
rect 2805 -91 2841 -72
rect 2266 -106 2771 -91
rect 2778 -106 2841 -91
rect 2140 -110 2771 -106
rect 2140 -126 2228 -110
rect 2266 -120 2771 -110
rect 2244 -126 2771 -120
rect 2790 -126 2841 -106
rect 3205 -126 4340 -66
rect 1717 -127 2103 -126
rect 1086 -156 1088 -128
rect 1717 -155 1751 -127
rect 1846 -154 1850 -127
rect 1944 -138 1956 -127
rect 2033 -134 2103 -127
rect 1884 -144 1990 -138
rect 1874 -154 1990 -144
rect 1124 -192 1126 -156
rect 1716 -188 1751 -155
rect 1837 -161 1850 -157
rect 1304 -308 1412 -302
rect 83 -376 201 -365
rect 283 -376 369 -365
rect 94 -388 190 -376
rect 294 -388 324 -376
rect 334 -384 369 -376
rect 447 -384 482 -371
rect 816 -374 820 -340
rect 1374 -374 1376 -340
rect 1640 -342 1650 -235
rect 1668 -342 1678 -207
rect 1717 -216 1751 -188
rect 1825 -195 1850 -161
rect 1868 -161 1990 -154
rect 2033 -143 2112 -134
rect 2208 -138 2316 -126
rect 2033 -144 2120 -143
rect 2132 -144 2148 -138
rect 2208 -140 2328 -138
rect 2033 -154 2158 -144
rect 1868 -170 1934 -161
rect 1884 -179 1928 -170
rect 1884 -188 1918 -179
rect 1944 -188 1956 -161
rect 2033 -164 2164 -154
rect 2033 -170 2120 -164
rect 2033 -188 2112 -170
rect 1825 -204 1838 -195
rect 1844 -213 1850 -195
rect 1792 -216 1850 -213
rect 1859 -229 1872 -195
rect 1875 -216 1888 -195
rect 1944 -213 1947 -188
rect 1944 -216 2002 -213
rect 2033 -216 2103 -188
rect 2114 -216 2120 -170
rect 2138 -170 2164 -164
rect 2208 -167 2209 -140
rect 2213 -141 2328 -140
rect 2228 -167 2328 -141
rect 2342 -154 2436 -126
rect 2354 -167 2436 -154
rect 2138 -188 2158 -170
rect 2208 -183 2436 -167
rect 2166 -204 2436 -183
rect 2208 -216 2436 -204
rect 2440 -215 2490 -126
rect 2628 -155 2662 -138
rect 2674 -155 2742 -126
rect 2563 -204 2574 -159
rect 2628 -177 2742 -155
rect 2616 -187 2742 -177
rect 2601 -193 2742 -187
rect 2597 -200 2742 -193
rect 2771 -198 2805 -126
rect 2832 -198 2839 -138
rect 2841 -198 2878 -126
rect 2922 -144 2938 -138
rect 2894 -154 2948 -144
rect 2888 -164 2954 -154
rect 2888 -170 2916 -164
rect 2904 -188 2916 -170
rect 2928 -170 2954 -164
rect 2928 -188 2948 -170
rect 3112 -172 3144 -126
rect 3188 -144 3204 -138
rect 3205 -144 3212 -126
rect 3160 -154 3214 -144
rect 3154 -164 3220 -154
rect 3154 -170 3182 -164
rect 3194 -170 3220 -164
rect 3170 -174 3214 -170
rect 3230 -174 3275 -126
rect 3362 -138 3449 -126
rect 3462 -138 3472 -126
rect 3349 -150 3483 -138
rect 3321 -159 3511 -150
rect 3321 -172 3364 -159
rect 3376 -170 3450 -159
rect 3376 -172 3444 -170
rect 3462 -172 3472 -159
rect 3474 -172 3511 -159
rect 3321 -174 3376 -172
rect 3400 -174 3511 -172
rect 3170 -188 3276 -174
rect 3321 -184 3511 -174
rect 2771 -200 2878 -198
rect 2597 -215 2878 -200
rect 2440 -216 2878 -215
rect 2998 -216 3056 -198
rect 3086 -216 3144 -198
rect 3180 -204 3276 -188
rect 3330 -188 3511 -184
rect 3330 -204 3508 -188
rect 3180 -216 3212 -204
rect 3230 -208 3231 -204
rect 3241 -208 3275 -204
rect 3343 -208 3389 -204
rect 3400 -208 3401 -204
rect 3431 -208 3434 -204
rect 3443 -208 3504 -204
rect 3549 -208 4340 -126
rect 4348 -176 4383 -148
rect 4444 -176 4602 -148
rect 1907 -282 1933 -267
rect 1850 -304 1865 -292
rect 1907 -304 1918 -282
rect 1846 -310 1918 -304
rect 1919 -304 1952 -292
rect 1919 -310 1953 -304
rect 2033 -310 2043 -216
rect 2050 -310 2120 -216
rect 2200 -238 2234 -217
rect 2288 -221 2322 -217
rect 2276 -238 2322 -221
rect 1681 -314 2120 -310
rect 2138 -314 2158 -306
rect 2188 -314 2195 -259
rect 2276 -314 2296 -238
rect 2402 -314 2436 -216
rect 2452 -272 2489 -216
rect 2597 -227 2663 -216
rect 2601 -233 2659 -227
rect 2732 -228 2748 -222
rect 2771 -225 2841 -216
rect 3180 -225 3210 -216
rect 2714 -238 2758 -228
rect 2563 -261 2628 -238
rect 2662 -270 2691 -238
rect 2455 -278 2489 -272
rect 2664 -274 2691 -270
rect 2698 -254 2764 -238
rect 2698 -272 2758 -254
rect 2571 -275 2615 -274
rect 2563 -278 2615 -275
rect 2645 -278 2703 -274
rect 2732 -278 2758 -272
rect 2771 -269 3210 -225
rect 3216 -238 4340 -208
rect 4396 -182 4602 -176
rect 4663 -182 4698 -165
rect 5191 -178 5225 -165
rect 4396 -210 4554 -182
rect 3216 -268 3231 -238
rect 3241 -268 3275 -238
rect 3277 -242 3504 -238
rect 3509 -242 4340 -238
rect 3216 -269 3275 -268
rect 3400 -269 3401 -242
rect 3431 -269 3434 -242
rect 3532 -269 4340 -242
rect 2771 -278 4340 -269
rect 2442 -314 4340 -278
rect 1681 -348 4340 -314
rect 4348 -337 4382 -210
rect 4630 -229 4650 -182
rect 4664 -183 4698 -182
rect 4664 -219 4734 -183
rect 5175 -191 5241 -178
rect 5368 -212 5383 182
rect 5402 148 5437 182
rect 5498 159 5661 182
rect 5717 159 5810 193
rect 5894 174 5898 276
rect 5922 242 5980 248
rect 5922 208 5934 242
rect 5922 202 5980 208
rect 5498 148 5656 159
rect 5717 148 5806 159
rect 5402 -159 5436 148
rect 5718 147 5806 148
rect 6111 147 6126 638
rect 5735 106 5806 147
rect 5867 140 6025 147
rect 5867 113 6030 140
rect 5872 106 6030 113
rect 6086 106 6126 147
rect 6145 106 6179 638
rect 6225 600 6415 624
rect 6253 572 6299 596
rect 6341 572 6387 596
rect 6291 189 6349 195
rect 6291 155 6303 189
rect 6291 149 6349 155
rect 5548 80 5606 86
rect 5548 46 5560 80
rect 5548 40 5606 46
rect 5735 -106 5805 106
rect 6087 94 6121 106
rect 6145 94 6175 106
rect 6480 94 6495 638
rect 5889 -23 5898 79
rect 5917 45 5975 51
rect 5917 11 5929 45
rect 5917 5 5975 11
rect 6106 0 6121 94
rect 5885 -106 5919 -72
rect 5973 -106 6007 -72
rect 6087 -106 6121 0
rect 6140 53 6175 94
rect 6236 87 6394 94
rect 6236 60 6399 87
rect 6241 53 6399 60
rect 6455 53 6495 94
rect 6514 634 6548 638
rect 6514 604 6830 634
rect 6514 600 6549 604
rect 6645 600 6733 604
rect 6514 53 6548 600
rect 6847 581 6917 638
rect 6847 547 6918 581
rect 7218 547 7233 638
rect 7252 547 7286 638
rect 7394 604 7460 630
rect 7410 600 7444 604
rect 7568 590 7655 638
rect 7823 636 7842 638
rect 7739 600 7853 611
rect 7942 604 8024 638
rect 6847 511 6900 547
rect 7252 513 7267 547
rect 7585 494 7655 590
rect 7767 572 7825 583
rect 7767 543 7779 572
rect 7767 537 7825 543
rect 7585 458 7638 494
rect 6830 421 6864 439
rect 7954 422 8024 604
rect 8158 558 8164 600
rect 8186 562 8192 600
rect 8108 544 8164 558
rect 8136 524 8194 530
rect 8136 516 8192 524
rect 8136 490 8148 516
rect 8136 484 8194 490
rect 8306 484 8340 638
rect 6830 385 6900 421
rect 7954 388 8025 422
rect 8325 388 8340 484
rect 8359 388 8393 638
rect 8501 637 8531 638
rect 8560 637 8567 671
rect 8594 638 8601 672
rect 8626 653 8762 672
rect 8836 671 8970 672
rect 8602 639 8762 653
rect 8804 639 9002 671
rect 9010 639 9131 672
rect 9228 661 9316 672
rect 9379 668 9447 672
rect 9483 668 9509 672
rect 9704 670 9737 672
rect 9239 649 9305 661
rect 9228 646 9316 649
rect 9379 646 9542 668
rect 9145 639 9542 646
rect 8602 638 9542 639
rect 9676 653 9870 668
rect 10109 653 11619 672
rect 9676 639 11619 653
rect 11665 639 11816 672
rect 11846 671 12469 672
rect 11846 666 12495 671
rect 9676 638 11816 639
rect 11906 661 12495 666
rect 11906 653 12461 661
rect 12465 653 12495 661
rect 11906 638 12495 653
rect 8439 600 8629 627
rect 8467 572 8513 599
rect 8555 572 8601 599
rect 8505 471 8563 477
rect 8505 437 8517 471
rect 8505 431 8563 437
rect 8675 431 8762 638
rect 8842 600 8876 633
rect 8930 600 8964 633
rect 6847 351 6918 385
rect 7198 351 7233 385
rect 7621 368 7656 386
rect 6660 136 6718 142
rect 6660 102 6672 136
rect 6660 96 6718 102
rect 6847 53 6917 351
rect 7199 332 7233 351
rect 7585 353 7656 368
rect 7029 283 7087 289
rect 7029 249 7041 283
rect 7029 243 7087 249
rect 7029 83 7087 89
rect 7029 53 7041 83
rect 6140 -53 6174 53
rect 6456 41 6490 53
rect 6514 41 6544 53
rect 6475 -2 6490 41
rect 6286 -8 6344 -2
rect 6286 -19 6298 -8
rect 6282 -42 6348 -19
rect 6286 -48 6344 -42
rect 6456 -53 6490 -2
rect 6509 0 6544 41
rect 6605 34 6763 41
rect 6847 35 6918 53
rect 7014 42 7102 53
rect 7025 35 7091 42
rect 6605 7 6768 34
rect 6610 0 6768 7
rect 6847 19 7199 35
rect 6509 -34 6549 0
rect 6847 -19 6917 19
rect 7007 -19 7109 -15
rect 6629 -27 6739 -23
rect 6617 -34 6751 -27
rect 6140 -87 6180 -53
rect 6188 -87 6442 -53
rect 5516 -159 5550 -125
rect 5604 -159 5638 -125
rect 5735 -140 5811 -106
rect 5872 -140 6019 -106
rect 6030 -140 6041 -106
rect 5402 -193 5442 -159
rect 5504 -172 5650 -159
rect 5661 -160 5672 -159
rect 5513 -176 5641 -172
rect 5510 -193 5644 -176
rect 5033 -219 5349 -212
rect 4664 -229 5349 -219
rect 4630 -246 5349 -229
rect 4474 -262 4490 -250
rect 4474 -272 4494 -262
rect 4474 -278 4490 -272
rect 4468 -284 4492 -278
rect 4506 -282 4530 -250
rect 4630 -253 5072 -246
rect 4630 -265 4751 -253
rect 5033 -259 5072 -253
rect 4630 -272 4734 -265
rect 4538 -282 4540 -280
rect 4504 -284 4552 -282
rect 4442 -290 4552 -284
rect 4442 -309 4508 -290
rect 4616 -299 4734 -272
rect 4751 -287 5019 -265
rect 4765 -294 4785 -287
rect 4825 -294 4959 -287
rect 4999 -294 5019 -287
rect 4751 -299 5019 -294
rect 4442 -310 4554 -309
rect 4616 -310 4751 -299
rect 4985 -310 5019 -299
rect 5033 -280 5349 -259
rect 5368 -272 5388 -212
rect 5402 -272 5441 -193
rect 5632 -200 5634 -193
rect 5548 -210 5606 -204
rect 5544 -244 5610 -210
rect 5735 -221 5810 -140
rect 5896 -186 5919 -170
rect 5968 -186 6015 -161
rect 5896 -204 6015 -186
rect 5903 -208 6015 -204
rect 5903 -216 5931 -208
rect 5548 -250 5606 -244
rect 5718 -250 5810 -221
rect 5881 -229 5931 -216
rect 5934 -216 6015 -208
rect 5934 -229 6011 -216
rect 5881 -242 6011 -229
rect 5553 -261 5611 -255
rect 5033 -293 5073 -280
rect 5129 -293 5340 -280
rect 5033 -310 5072 -293
rect 5086 -294 5126 -293
rect 5146 -294 5340 -293
rect 5086 -306 5354 -294
rect 5388 -306 5402 -294
rect 5407 -306 5422 -274
rect 5549 -295 5615 -261
rect 5735 -289 5810 -250
rect 5889 -263 5898 -242
rect 5922 -248 5980 -242
rect 5917 -263 5975 -257
rect 5886 -276 6016 -263
rect 5886 -289 5963 -276
rect 5966 -289 6016 -276
rect 5735 -291 5841 -289
rect 5553 -301 5611 -295
rect 5086 -310 5120 -306
rect 5368 -310 5388 -306
rect 5402 -310 5441 -306
rect 4442 -312 4580 -310
rect 4428 -314 4580 -312
rect 4616 -312 5632 -310
rect 4428 -318 4584 -314
rect 4396 -331 4584 -318
rect 4616 -325 5656 -312
rect 4396 -337 4596 -331
rect 4348 -348 4596 -337
rect 4616 -348 5709 -325
rect 1681 -359 5709 -348
rect 5723 -342 5841 -291
rect 5898 -297 6010 -289
rect 5898 -301 5936 -297
rect 5891 -313 5936 -301
rect 5966 -301 5994 -297
rect 5966 -313 6001 -301
rect 6087 -303 6126 -106
rect 5891 -335 5924 -313
rect 5978 -335 6001 -313
rect 6092 -342 6126 -303
rect 6140 -342 6179 -87
rect 6242 -112 6300 -89
rect 6330 -112 6388 -89
rect 6254 -139 6288 -112
rect 6337 -139 6384 -112
rect 6254 -205 6300 -139
rect 6330 -155 6384 -139
rect 6303 -189 6384 -155
rect 6330 -205 6376 -189
rect 6254 -232 6288 -205
rect 6254 -257 6293 -232
rect 6330 -236 6335 -205
rect 6342 -232 6376 -205
rect 6259 -300 6293 -257
rect 6300 -269 6304 -237
rect 6342 -257 6381 -232
rect 6347 -269 6381 -257
rect 6300 -300 6305 -269
rect 6259 -316 6305 -300
rect 6332 -316 6381 -269
rect 5723 -359 6210 -342
rect 1681 -382 5632 -359
rect 334 -388 498 -384
rect 83 -397 201 -388
rect 283 -397 498 -388
rect 83 -399 498 -397
rect 570 -398 604 -384
rect 119 -411 190 -409
rect 119 -451 124 -411
rect 335 -414 498 -399
rect 335 -418 370 -414
rect 721 -418 774 -417
rect 229 -433 295 -431
rect 161 -497 166 -451
rect 195 -497 227 -467
rect 229 -497 269 -433
rect 161 -501 227 -497
rect 161 -517 166 -501
rect 136 -535 261 -531
rect 121 -541 139 -539
rect 354 -541 370 -418
rect 388 -429 535 -418
rect 388 -441 532 -429
rect 570 -432 638 -418
rect 701 -429 774 -418
rect 1042 -419 1044 -410
rect 388 -448 535 -441
rect 703 -448 774 -429
rect 992 -444 1141 -419
rect 1681 -437 4340 -382
rect 1337 -444 1586 -439
rect 388 -452 423 -448
rect 483 -452 535 -448
rect 700 -452 774 -448
rect 388 -541 422 -452
rect 494 -504 524 -462
rect 670 -482 700 -452
rect 704 -482 774 -452
rect 901 -464 953 -453
rect 912 -466 942 -464
rect 882 -476 950 -466
rect 958 -476 1107 -453
rect 700 -486 704 -482
rect 530 -541 566 -504
rect 712 -514 774 -482
rect 871 -478 1107 -476
rect 871 -487 961 -478
rect 989 -487 1073 -478
rect 712 -516 791 -514
rect 670 -532 700 -516
rect 704 -532 791 -516
rect 882 -532 912 -497
rect 932 -516 936 -487
rect 942 -532 950 -497
rect 1000 -526 1007 -497
rect 1092 -526 1107 -478
rect 1335 -473 1512 -470
rect 1335 -478 1586 -473
rect 1335 -484 1585 -478
rect 1335 -496 1574 -484
rect 1335 -505 1585 -496
rect 1668 -505 4340 -437
rect 1335 -506 4340 -505
rect 1126 -514 1169 -506
rect 1222 -514 1311 -506
rect 1331 -507 4340 -506
rect 1331 -514 1514 -507
rect 1126 -516 1514 -514
rect 1126 -523 1512 -516
rect 1668 -523 4340 -507
rect 1126 -526 4340 -523
rect 618 -541 791 -532
rect 0 -553 791 -541
rect -17 -579 791 -553
rect 1000 -537 4340 -526
rect 1000 -568 1030 -537
rect 1036 -560 4340 -537
rect 1073 -568 1107 -560
rect 884 -579 912 -568
rect 915 -579 996 -568
rect -17 -589 996 -579
rect 1002 -585 1107 -568
rect -17 -613 983 -589
rect -17 -650 791 -613
rect 854 -648 872 -634
rect 942 -636 947 -613
rect 949 -636 983 -613
rect -17 -675 800 -650
rect -17 -681 837 -675
rect -105 -1135 -71 -685
rect -17 -695 800 -681
rect 832 -695 841 -681
rect 854 -695 905 -648
rect 912 -695 916 -637
rect 949 -641 993 -636
rect 1002 -637 1036 -585
rect 1000 -641 1036 -637
rect 949 -686 1036 -641
rect 949 -695 993 -686
rect -17 -706 852 -695
rect -17 -708 841 -706
rect 854 -708 993 -695
rect -17 -718 993 -708
rect -57 -719 993 -718
rect -17 -720 993 -719
rect 1000 -720 1036 -686
rect -17 -729 1036 -720
rect -17 -748 800 -729
rect 854 -748 859 -729
rect 866 -736 903 -729
rect -17 -781 791 -748
rect 835 -762 869 -758
rect 871 -762 905 -736
rect 825 -767 905 -762
rect 912 -748 916 -729
rect 949 -748 1036 -729
rect 1042 -714 1070 -636
rect 1073 -709 1107 -585
rect 1126 -622 1160 -560
rect 1318 -568 4340 -560
rect 1196 -576 4340 -568
rect 1196 -608 3971 -576
rect 1196 -622 1241 -608
rect 1126 -628 1241 -622
rect 1126 -662 1160 -628
rect 1196 -636 1241 -628
rect 1174 -662 1241 -636
rect 1272 -629 3971 -608
rect 3979 -607 4019 -576
rect 4045 -607 4079 -576
rect 4091 -607 4121 -576
rect 4133 -607 4167 -576
rect 4200 -584 4246 -576
rect 4200 -607 4233 -584
rect 4247 -607 4281 -576
rect 4295 -604 4334 -576
rect 4348 -604 4382 -382
rect 4402 -404 4448 -382
rect 4462 -404 4536 -382
rect 4402 -416 4536 -404
rect 4402 -420 4538 -416
rect 4550 -420 4574 -382
rect 4582 -416 4584 -382
rect 4402 -453 4542 -420
rect 4544 -453 4574 -420
rect 4591 -431 4596 -382
rect 4585 -450 4596 -431
rect 4402 -466 4574 -453
rect 4582 -466 4596 -450
rect 4402 -472 4596 -466
rect 4616 -389 5632 -382
rect 4616 -423 5655 -389
rect 5735 -413 6210 -359
rect 6259 -350 6381 -316
rect 6259 -366 6305 -350
rect 6335 -366 6381 -350
rect 6456 -356 6495 -53
rect 6259 -413 6293 -366
rect 6347 -413 6381 -366
rect 5735 -418 6233 -413
rect 6247 -418 6447 -413
rect 4616 -461 5647 -423
rect 5735 -435 6210 -418
rect 5737 -445 6210 -435
rect 4616 -467 5632 -461
rect 4414 -484 4588 -472
rect 4388 -499 4588 -484
rect 4388 -511 4570 -499
rect 4582 -511 4588 -499
rect 4388 -539 4460 -511
rect 4462 -515 4588 -511
rect 4388 -584 4448 -539
rect 4454 -552 4460 -539
rect 4470 -539 4588 -515
rect 4470 -542 4538 -539
rect 4540 -542 4588 -539
rect 4470 -550 4588 -542
rect 4616 -529 5639 -467
rect 5723 -475 6210 -445
rect 6236 -447 6447 -418
rect 6236 -452 6399 -447
rect 6241 -475 6399 -452
rect 5689 -529 5691 -495
rect 4414 -604 4448 -584
rect 4490 -592 4587 -550
rect 4616 -563 5637 -529
rect 5657 -563 5695 -529
rect 5698 -563 5703 -499
rect 5723 -563 6227 -475
rect 4616 -569 5703 -563
rect 5737 -569 6227 -563
rect 4490 -600 4556 -592
rect 4616 -597 6227 -569
rect 6247 -505 6281 -475
rect 6317 -496 6347 -481
rect 6385 -484 6393 -475
rect 6378 -496 6393 -484
rect 6247 -527 6293 -505
rect 6317 -515 6393 -496
rect 6247 -543 6305 -527
rect 6335 -543 6415 -515
rect 6247 -549 6415 -543
rect 6247 -580 6393 -549
rect 6247 -583 6387 -580
rect 6247 -593 6305 -583
rect 6319 -592 6387 -583
rect 6307 -593 6387 -592
rect 6247 -596 6299 -593
rect 6307 -596 6341 -593
rect 6347 -596 6387 -593
rect 6395 -596 6415 -592
rect 4616 -600 5660 -597
rect 4466 -604 4580 -600
rect 4616 -604 5632 -600
rect 4295 -607 5632 -604
rect 1272 -638 3596 -629
rect 3608 -638 3636 -629
rect 3664 -638 3670 -629
rect 3676 -638 3798 -629
rect 3878 -638 3928 -629
rect 1272 -648 3608 -638
rect 1284 -658 3608 -648
rect 3625 -649 3928 -638
rect 1126 -668 1210 -662
rect 1126 -670 1160 -668
rect 1124 -684 1160 -670
rect 1196 -670 1210 -668
rect 1124 -686 1162 -684
rect 1112 -709 1162 -686
rect 1196 -685 1242 -670
rect 1196 -686 1244 -685
rect 1262 -686 1274 -685
rect 1196 -693 1274 -686
rect 1196 -709 1207 -693
rect 1073 -714 1162 -709
rect 1042 -724 1162 -714
rect 1208 -720 1274 -693
rect 1042 -736 1107 -724
rect 1108 -734 1162 -724
rect 1073 -748 1107 -736
rect 1116 -748 1160 -734
rect 1204 -748 1238 -721
rect 1240 -748 1274 -720
rect 1286 -714 1316 -658
rect 1318 -671 3608 -658
rect 3636 -661 3928 -649
rect 3625 -671 3928 -661
rect 1318 -672 3928 -671
rect 1318 -675 3596 -672
rect 3664 -675 3670 -672
rect 3676 -675 3801 -672
rect 1318 -714 3608 -675
rect 1286 -736 3608 -714
rect 3664 -694 3801 -675
rect 3664 -706 3722 -694
rect 3664 -722 3740 -706
rect 1286 -748 1316 -736
rect 1318 -748 3608 -736
rect 912 -767 917 -748
rect 949 -762 3608 -748
rect 3636 -726 3740 -722
rect 3764 -722 3798 -694
rect 3764 -726 3828 -722
rect 3878 -726 3928 -672
rect 3636 -762 3928 -726
rect 949 -765 3928 -762
rect 949 -767 3608 -765
rect 825 -781 917 -767
rect -17 -797 793 -781
rect 823 -787 917 -781
rect 819 -797 917 -787
rect -17 -816 917 -797
rect 947 -778 3608 -767
rect 3636 -778 3928 -765
rect 947 -782 3928 -778
rect 947 -806 1107 -782
rect 947 -816 1036 -806
rect -17 -820 905 -816
rect 949 -820 993 -816
rect -17 -821 872 -820
rect 949 -821 988 -820
rect 1002 -821 1036 -816
rect -17 -838 1036 -821
rect 1073 -838 1107 -806
rect 1116 -796 3928 -782
rect 3931 -723 3965 -629
rect 3979 -638 4179 -607
rect 4200 -618 5632 -607
rect 4200 -638 4334 -618
rect 4348 -638 4382 -618
rect 4414 -638 4448 -618
rect 4466 -626 4536 -618
rect 4542 -626 4580 -618
rect 4616 -623 5632 -618
rect 5651 -623 5660 -600
rect 5670 -623 5697 -600
rect 5698 -623 5725 -600
rect 5740 -623 6227 -597
rect 6259 -600 6293 -596
rect 6301 -600 6381 -596
rect 6301 -609 6354 -600
rect 6389 -608 6415 -596
rect 6301 -619 6371 -609
rect 6389 -619 6419 -608
rect 6427 -619 6429 -592
rect 4490 -638 4536 -626
rect 4616 -631 6227 -623
rect 6259 -624 6293 -619
rect 6301 -624 6381 -619
rect 4616 -638 5725 -631
rect 3979 -641 5725 -638
rect 4000 -652 4019 -641
rect 4020 -669 4179 -641
rect 4200 -652 5725 -641
rect 4247 -661 4288 -652
rect 4300 -660 4334 -652
rect 4346 -660 4382 -652
rect 4402 -660 4548 -652
rect 4600 -657 5725 -652
rect 5737 -653 6227 -631
rect 6247 -627 6299 -624
rect 6301 -627 6387 -624
rect 6247 -653 6387 -627
rect 6389 -653 6433 -619
rect 6436 -653 6441 -596
rect 5737 -657 6213 -653
rect 4549 -660 5632 -657
rect 4296 -661 5632 -660
rect 4020 -671 4228 -669
rect 4247 -670 5632 -661
rect 4246 -671 5632 -670
rect 4020 -672 5632 -671
rect 4042 -704 4170 -672
rect 4213 -704 4246 -672
rect 4247 -704 4288 -672
rect 4296 -679 5632 -672
rect 5651 -679 5660 -657
rect 5670 -679 5697 -657
rect 5698 -679 6213 -657
rect 4296 -688 5019 -679
rect 4296 -694 4734 -688
rect 4296 -704 4448 -694
rect 4042 -706 4212 -704
rect 4246 -706 4448 -704
rect 4042 -713 4170 -706
rect 4051 -723 4170 -713
rect 4247 -709 4448 -706
rect 4490 -709 4536 -694
rect 4548 -704 4580 -694
rect 4616 -703 4734 -694
rect 4751 -703 5019 -688
rect 4616 -704 4737 -703
rect 4746 -704 4764 -703
rect 4771 -704 4817 -703
rect 4824 -704 4829 -703
rect 4844 -704 4917 -703
rect 4548 -709 4734 -704
rect 4247 -723 4734 -709
rect 4746 -713 4751 -704
rect 4764 -713 4917 -704
rect 4932 -713 4939 -703
rect 4951 -713 4966 -703
rect 4985 -713 5019 -703
rect 5033 -713 5072 -679
rect 3931 -726 3982 -723
rect 3931 -796 3965 -726
rect 4033 -730 4185 -723
rect 4217 -728 4734 -723
rect 4764 -722 4932 -713
rect 4966 -722 5005 -713
rect 4764 -728 5005 -722
rect 4000 -756 4185 -730
rect 4200 -738 4334 -728
rect 4000 -757 4179 -756
rect 4200 -757 4281 -738
rect 4288 -743 4334 -738
rect 4288 -754 4296 -743
rect 4000 -790 4168 -757
rect 1116 -802 3916 -796
rect 1116 -816 1160 -802
rect 1204 -816 1238 -802
rect 1116 -838 1238 -816
rect 1240 -825 1274 -802
rect 1318 -804 3916 -802
rect 1318 -812 3676 -804
rect 3682 -812 3916 -804
rect 1318 -815 3916 -812
rect 3928 -815 3996 -796
rect 1318 -816 3996 -815
rect 4000 -815 4019 -790
rect 4033 -815 4161 -790
rect 4200 -806 4246 -757
rect 4200 -815 4233 -806
rect 4247 -815 4281 -757
rect 1318 -818 3706 -816
rect 1318 -825 3712 -818
rect 1240 -830 3712 -825
rect 1240 -838 3596 -830
rect 3602 -838 3712 -830
rect 3720 -830 3916 -816
rect 3720 -834 3754 -830
rect 3760 -838 3916 -830
rect -17 -846 3793 -838
rect 3838 -846 3916 -838
rect -17 -849 3883 -846
rect -17 -854 3872 -849
rect -17 -872 3870 -854
rect -17 -917 791 -872
rect 835 -876 869 -872
rect -17 -942 815 -917
rect 835 -923 881 -876
rect 899 -889 903 -872
rect 915 -885 928 -872
rect 949 -885 983 -872
rect 915 -889 983 -885
rect 899 -897 983 -889
rect 949 -914 983 -897
rect 915 -923 983 -914
rect 835 -942 869 -923
rect -17 -948 869 -942
rect 899 -931 983 -923
rect 899 -948 903 -931
rect 915 -935 983 -931
rect 915 -948 928 -935
rect 949 -948 983 -935
rect 1002 -948 1036 -872
rect 1073 -877 1107 -872
rect 1116 -873 1272 -872
rect 1116 -877 1241 -873
rect 1073 -889 1250 -877
rect 1268 -882 1272 -873
rect 1284 -878 1297 -872
rect 1318 -874 3596 -872
rect 3636 -873 3816 -872
rect 3840 -873 3870 -872
rect 3897 -872 3916 -846
rect 3931 -849 3966 -816
rect 4000 -820 4281 -815
rect 4033 -840 4281 -820
rect 4033 -844 4191 -840
rect 4200 -844 4281 -840
rect 4300 -776 4334 -743
rect 4402 -740 4548 -728
rect 4565 -737 5005 -728
rect 4565 -738 4703 -737
rect 4565 -740 4600 -738
rect 4402 -754 4600 -740
rect 4402 -760 4588 -754
rect 4338 -776 4346 -760
rect 4376 -772 4588 -760
rect 4376 -776 4548 -772
rect 4554 -776 4570 -772
rect 4582 -776 4588 -772
rect 4616 -776 4703 -738
rect 4717 -747 4978 -737
rect 4730 -776 4737 -747
rect 4749 -776 4764 -747
rect 4783 -776 4798 -747
rect 4810 -776 4817 -747
rect 4824 -754 4829 -747
rect 4832 -754 4905 -747
rect 4833 -756 4905 -754
rect 4844 -769 4905 -756
rect 4844 -776 4878 -769
rect 4898 -776 4905 -769
rect 4932 -776 4939 -747
rect 4300 -781 4737 -776
rect 4764 -781 4783 -776
rect 4817 -781 4878 -776
rect 4905 -781 4932 -776
rect 4300 -810 4703 -781
rect 4730 -790 4737 -781
rect 4832 -785 4899 -781
rect 4300 -844 4334 -810
rect 4338 -826 4346 -810
rect 4376 -816 4460 -810
rect 4490 -814 4530 -810
rect 4542 -814 4548 -810
rect 4376 -826 4448 -816
rect 4402 -844 4448 -826
rect 4490 -844 4548 -814
rect 4616 -844 4703 -810
rect 4720 -830 4758 -808
rect 4777 -810 4911 -785
rect 4832 -813 4899 -810
rect 4951 -811 4978 -747
rect 4815 -819 4899 -813
rect 4033 -846 4703 -844
rect 4718 -846 4758 -830
rect 4033 -849 4758 -846
rect 1318 -878 3579 -874
rect 1284 -880 2495 -878
rect 2569 -880 2615 -878
rect 2657 -880 2691 -878
rect 2771 -880 3579 -878
rect 1284 -882 2714 -880
rect 1073 -948 1107 -889
rect 1116 -893 1162 -889
rect 1126 -900 1162 -893
rect 1192 -893 1238 -889
rect 1192 -900 1210 -893
rect 1126 -909 1160 -900
rect 1268 -904 2714 -882
rect 1318 -906 2714 -904
rect 2748 -906 2771 -880
rect 1126 -914 1184 -909
rect 1318 -914 2495 -906
rect 2569 -914 2615 -906
rect 2657 -914 2691 -906
rect 1116 -931 1194 -914
rect 1204 -929 1238 -914
rect 1284 -916 2714 -914
rect 1268 -929 2714 -916
rect 1204 -931 2714 -929
rect 1116 -940 2714 -931
rect 2748 -940 2771 -914
rect 2788 -940 3579 -880
rect 3625 -880 3816 -873
rect 3829 -874 3878 -873
rect 3625 -882 3797 -880
rect 3829 -882 3881 -874
rect 3596 -884 3881 -882
rect 3752 -918 3796 -884
rect 3686 -936 3796 -918
rect 3878 -936 3881 -884
rect 3897 -936 3912 -872
rect 3931 -936 3965 -849
rect 4051 -858 4758 -849
rect 4811 -820 4899 -819
rect 4920 -820 4978 -811
rect 4985 -747 5005 -737
rect 5038 -726 5053 -713
rect 5038 -747 5072 -726
rect 4985 -820 5019 -747
rect 4811 -853 4877 -820
rect 4051 -859 4776 -858
rect 4815 -859 4873 -853
rect 4051 -880 4091 -859
rect 4112 -880 4113 -859
rect 4121 -865 4776 -859
rect 4890 -865 4919 -820
rect 4951 -865 4966 -820
rect 4985 -865 5000 -820
rect 4121 -867 4931 -865
rect 4045 -896 4091 -880
rect 4121 -896 4985 -867
rect 4045 -902 4088 -896
rect 4058 -918 4088 -902
rect 4132 -899 4985 -896
rect 4132 -908 4776 -899
rect 4132 -912 4703 -908
rect 4133 -914 4196 -912
rect 4045 -924 4088 -918
rect 1116 -942 2615 -940
rect 2657 -942 2691 -940
rect 2771 -942 3579 -940
rect 1116 -948 1308 -942
rect 1318 -946 3579 -942
rect 3596 -946 3996 -936
rect 1318 -948 3996 -946
rect -17 -982 3996 -948
rect 4045 -961 4091 -924
rect 4112 -961 4196 -914
rect 4045 -971 4196 -961
rect 4200 -924 4233 -912
rect 4200 -971 4201 -924
rect 4247 -971 4281 -912
rect -17 -984 1036 -982
rect 1073 -984 1107 -982
rect -17 -999 1107 -984
rect -17 -1000 872 -999
rect 949 -1000 988 -999
rect -17 -1004 905 -1000
rect 949 -1004 993 -1000
rect 1002 -1004 1036 -999
rect -17 -1023 917 -1004
rect -17 -1046 869 -1023
rect -17 -1058 793 -1046
rect 800 -1058 869 -1046
rect -17 -1071 791 -1058
rect 835 -1062 869 -1058
rect 871 -1024 917 -1023
rect 947 -1014 1036 -1004
rect 1073 -1014 1107 -999
rect 947 -1024 1107 -1014
rect -17 -1078 859 -1071
rect 871 -1078 905 -1024
rect -17 -1084 905 -1078
rect 912 -1072 917 -1046
rect -17 -1091 903 -1084
rect 912 -1091 916 -1072
rect 949 -1091 993 -1024
rect 1002 -1038 1107 -1024
rect 1116 -1018 1184 -982
rect 1192 -984 1238 -982
rect 1188 -1018 1238 -984
rect 1240 -1018 1274 -982
rect 1318 -1004 3722 -982
rect 3752 -990 3996 -982
rect 3740 -1004 3996 -990
rect 4027 -1000 4281 -971
rect 1318 -1008 3916 -1004
rect 1318 -1018 3596 -1008
rect 1116 -1024 3596 -1018
rect 3598 -1020 3832 -1008
rect 3856 -1019 3916 -1008
rect 3856 -1020 3872 -1019
rect 3598 -1024 3706 -1020
rect 3722 -1024 3828 -1020
rect 3878 -1024 3916 -1019
rect 3928 -1024 3996 -1004
rect 4000 -1005 4281 -1000
rect 1116 -1038 3928 -1024
rect 1002 -1046 1036 -1038
rect -17 -1125 993 -1091
rect -17 -1139 800 -1125
rect 832 -1139 841 -1125
rect 854 -1139 905 -1125
rect -17 -1145 837 -1139
rect -17 -1170 800 -1145
rect 854 -1170 856 -1139
rect -17 -1207 791 -1170
rect 866 -1172 905 -1139
rect 912 -1172 916 -1125
rect 949 -1184 993 -1125
rect 1000 -1050 1036 -1046
rect 1073 -1042 3928 -1038
rect 1073 -1050 3608 -1042
rect 1000 -1055 3608 -1050
rect 3636 -1055 3928 -1042
rect 1000 -1058 3928 -1055
rect 1000 -1072 3608 -1058
rect 1000 -1172 1036 -1072
rect 1073 -1084 1184 -1072
rect 868 -1207 996 -1184
rect -17 -1241 996 -1207
rect -17 -1267 791 -1241
rect 884 -1252 912 -1241
rect 915 -1252 996 -1241
rect 1002 -1206 1036 -1172
rect 1042 -1099 1184 -1084
rect 1204 -1085 1238 -1072
rect 1240 -1085 1274 -1072
rect 1204 -1099 1274 -1085
rect 1042 -1106 1162 -1099
rect 1042 -1184 1070 -1106
rect 1073 -1111 1162 -1106
rect 1208 -1111 1274 -1099
rect 1073 -1206 1107 -1111
rect 1112 -1134 1162 -1111
rect 1124 -1136 1162 -1134
rect 1196 -1119 1274 -1111
rect 1196 -1134 1242 -1119
rect 1196 -1135 1244 -1134
rect 1262 -1135 1274 -1119
rect 1286 -1084 1316 -1072
rect 1318 -1084 3608 -1072
rect 1286 -1106 3608 -1084
rect 3636 -1094 3928 -1058
rect 3636 -1098 3740 -1094
rect 1286 -1131 1316 -1106
rect 1318 -1115 3608 -1106
rect 1318 -1131 3596 -1115
rect 1124 -1150 1160 -1136
rect 1002 -1237 1107 -1206
rect 1126 -1152 1160 -1150
rect 1196 -1150 1242 -1135
rect 1286 -1148 3596 -1131
rect 3608 -1148 3636 -1122
rect 3664 -1148 3670 -1098
rect 3676 -1110 3740 -1098
rect 3754 -1098 3828 -1094
rect 3676 -1114 3752 -1110
rect 3754 -1114 3801 -1098
rect 3676 -1148 3801 -1114
rect 3878 -1148 3928 -1094
rect 1196 -1152 1241 -1150
rect 1126 -1158 1241 -1152
rect 1126 -1192 1160 -1158
rect 1174 -1184 1241 -1158
rect 1286 -1162 3608 -1148
rect 3625 -1159 3928 -1148
rect 1284 -1172 3608 -1162
rect 3636 -1171 3928 -1159
rect 1196 -1192 1241 -1184
rect 1272 -1173 3608 -1172
rect 3625 -1173 3928 -1171
rect 1272 -1182 3928 -1173
rect 1272 -1191 3596 -1182
rect 3664 -1191 3670 -1182
rect 3676 -1191 3710 -1182
rect 3722 -1191 3752 -1182
rect 3764 -1191 3798 -1182
rect 3878 -1191 3928 -1182
rect 3931 -1094 3965 -1024
rect 4000 -1063 4019 -1005
rect 4033 -1014 4167 -1005
rect 4200 -1014 4233 -1005
rect 4033 -1063 4168 -1014
rect 4200 -1063 4246 -1014
rect 4247 -1063 4281 -1005
rect 4000 -1082 4281 -1063
rect 4300 -918 4334 -912
rect 4406 -918 4502 -912
rect 4542 -918 4543 -912
rect 4616 -918 4758 -912
rect 4300 -921 4758 -918
rect 4951 -921 4966 -899
rect 4985 -921 5000 -899
rect 4300 -933 4932 -921
rect 4966 -933 4985 -921
rect 4300 -952 4776 -933
rect 4300 -1010 4334 -952
rect 4406 -959 4502 -952
rect 4542 -959 4543 -952
rect 4616 -955 4776 -952
rect 4777 -944 4920 -933
rect 4777 -946 4931 -944
rect 5004 -946 5019 -820
rect 4777 -955 5019 -946
rect 4402 -972 4460 -959
rect 4388 -973 4460 -972
rect 4388 -976 4454 -973
rect 4388 -981 4448 -976
rect 4490 -977 4548 -959
rect 4490 -981 4536 -977
rect 4388 -994 4536 -981
rect 4338 -1010 4346 -994
rect 4376 -1010 4536 -994
rect 4542 -1010 4548 -977
rect 4616 -974 4758 -955
rect 4815 -967 4873 -961
rect 4616 -1010 4703 -974
rect 4718 -990 4736 -974
rect 4811 -1000 4877 -967
rect 4890 -1000 4919 -955
rect 4951 -1000 4966 -955
rect 4811 -1001 4899 -1000
rect 4815 -1007 4890 -1001
rect 4832 -1010 4890 -1007
rect 4300 -1039 4703 -1010
rect 4730 -1039 4737 -1030
rect 4300 -1044 4737 -1039
rect 4288 -1077 4296 -1066
rect 4300 -1077 4334 -1044
rect 4338 -1060 4346 -1044
rect 4376 -1048 4548 -1044
rect 4554 -1048 4570 -1044
rect 4582 -1048 4588 -1044
rect 4376 -1054 4588 -1048
rect 4376 -1060 4460 -1054
rect 4388 -1064 4460 -1060
rect 4470 -1064 4588 -1054
rect 4402 -1070 4460 -1064
rect 4402 -1072 4448 -1070
rect 4288 -1082 4334 -1077
rect 4000 -1090 4334 -1082
rect 4027 -1091 4334 -1090
rect 4376 -1091 4448 -1072
rect 4454 -1080 4460 -1070
rect 4027 -1092 4448 -1091
rect 4027 -1094 4201 -1092
rect 4217 -1094 4334 -1092
rect 3931 -1097 4334 -1094
rect 3931 -1191 3965 -1097
rect 4051 -1107 4170 -1097
rect 4051 -1114 4091 -1107
rect 4121 -1114 4161 -1107
rect 4247 -1114 4334 -1097
rect 4045 -1116 4100 -1114
rect 4121 -1116 4212 -1114
rect 4246 -1116 4334 -1114
rect 3994 -1148 4033 -1122
rect 4045 -1123 4091 -1116
rect 4045 -1145 4088 -1123
rect 4100 -1145 4113 -1116
rect 4121 -1123 4167 -1116
rect 4213 -1122 4246 -1116
rect 4247 -1122 4281 -1116
rect 4300 -1122 4334 -1116
rect 4414 -1114 4448 -1092
rect 4490 -1114 4536 -1064
rect 4542 -1066 4588 -1064
rect 4542 -1082 4600 -1066
rect 4616 -1082 4703 -1044
rect 4730 -1073 4737 -1044
rect 4749 -1039 4764 -1030
rect 4777 -1035 4911 -1010
rect 4832 -1039 4905 -1035
rect 4951 -1039 4978 -1000
rect 4749 -1044 4978 -1039
rect 4749 -1063 4764 -1044
rect 4779 -1051 4817 -1044
rect 4749 -1073 4771 -1063
rect 4779 -1073 4798 -1051
rect 4810 -1073 4817 -1051
rect 4844 -1064 4917 -1044
rect 4932 -1063 4978 -1044
rect 4824 -1073 4829 -1066
rect 4844 -1073 4851 -1064
rect 4871 -1066 4917 -1064
rect 4859 -1073 4917 -1066
rect 4920 -1073 4978 -1063
rect 4985 -1073 5019 -955
rect 5038 -812 5073 -747
rect 5086 -766 5120 -679
rect 5150 -688 5154 -679
rect 5206 -681 5230 -679
rect 5244 -681 5268 -679
rect 5201 -688 5294 -681
rect 5308 -688 5336 -679
rect 5150 -689 5336 -688
rect 5180 -695 5294 -689
rect 5308 -695 5336 -689
rect 5180 -698 5337 -695
rect 5180 -705 5294 -698
rect 5308 -705 5336 -698
rect 5180 -706 5336 -705
rect 5201 -714 5336 -706
rect 5201 -722 5246 -714
rect 5262 -722 5327 -714
rect 5150 -726 5184 -722
rect 5201 -723 5228 -722
rect 5259 -723 5327 -722
rect 5150 -738 5196 -726
rect 5243 -732 5327 -723
rect 5240 -738 5327 -732
rect 5354 -726 5388 -679
rect 5354 -738 5396 -726
rect 5150 -740 5327 -738
rect 5150 -744 5196 -740
rect 5240 -744 5327 -740
rect 5150 -766 5186 -744
rect 5228 -759 5327 -744
rect 5240 -766 5327 -759
rect 5350 -766 5396 -738
rect 5402 -759 5441 -679
rect 5455 -726 5489 -679
rect 5508 -691 5538 -679
rect 5623 -683 5632 -679
rect 5689 -683 5691 -679
rect 5563 -691 5632 -683
rect 5508 -698 5632 -691
rect 5508 -709 5538 -698
rect 5563 -704 5584 -698
rect 5563 -709 5618 -704
rect 5698 -707 5725 -679
rect 5549 -711 5618 -709
rect 5549 -725 5659 -711
rect 5723 -717 5725 -707
rect 5737 -687 6213 -679
rect 6225 -687 6227 -653
rect 6241 -687 6441 -653
rect 5737 -719 6227 -687
rect 5549 -726 5663 -725
rect 5450 -759 5495 -726
rect 5538 -741 5663 -726
rect 5549 -751 5663 -741
rect 5723 -745 6227 -719
rect 6247 -693 6387 -687
rect 6247 -721 6299 -693
rect 6301 -721 6341 -693
rect 6247 -732 6341 -721
rect 6347 -732 6387 -693
rect 6247 -745 6387 -732
rect 6389 -711 6419 -687
rect 6427 -711 6429 -687
rect 6389 -745 6433 -711
rect 6436 -745 6441 -687
rect 5549 -759 5618 -751
rect 5402 -765 5709 -759
rect 5723 -765 6213 -745
rect 5402 -766 6213 -765
rect 5086 -772 5396 -766
rect 5407 -772 5441 -766
rect 5450 -772 6213 -766
rect 5086 -779 6213 -772
rect 6225 -779 6227 -745
rect 6241 -776 6441 -745
rect 6241 -779 6393 -776
rect 6399 -779 6415 -776
rect 5086 -793 6227 -779
rect 5086 -800 5441 -793
rect 5150 -808 5222 -800
rect 5150 -809 5226 -808
rect 5138 -812 5226 -809
rect 5240 -812 5296 -800
rect 5354 -806 5396 -800
rect 5407 -806 5441 -800
rect 5450 -797 5596 -793
rect 5609 -797 5643 -793
rect 5450 -804 5584 -797
rect 5450 -806 5561 -804
rect 5354 -812 5561 -806
rect 5567 -809 5584 -804
rect 5575 -810 5584 -809
rect 5038 -819 5561 -812
rect 5572 -819 5589 -810
rect 5597 -818 5655 -797
rect 5609 -819 5643 -818
rect 5723 -819 6227 -793
rect 5038 -827 6227 -819
rect 5038 -834 5441 -827
rect 5038 -846 5396 -834
rect 5038 -860 5073 -846
rect 5138 -859 5218 -846
rect 5138 -860 5196 -859
rect 5038 -872 5196 -860
rect 5250 -860 5268 -846
rect 5354 -860 5396 -846
rect 5038 -876 5226 -872
rect 5038 -880 5230 -876
rect 5250 -880 5396 -860
rect 5038 -894 5396 -880
rect 5038 -906 5246 -894
rect 5250 -906 5396 -894
rect 5038 -914 5072 -906
rect 5262 -914 5280 -906
rect 5038 -974 5073 -914
rect 5165 -926 5246 -914
rect 5250 -926 5280 -914
rect 5165 -929 5280 -926
rect 5180 -940 5280 -929
rect 5354 -914 5388 -906
rect 5180 -944 5230 -940
rect 5180 -945 5226 -944
rect 5138 -948 5226 -945
rect 5228 -948 5230 -944
rect 5250 -948 5268 -940
rect 5138 -961 5196 -948
rect 5138 -974 5198 -961
rect 5250 -974 5261 -948
rect 5354 -974 5396 -914
rect 5038 -975 5396 -974
rect 5038 -985 5239 -975
rect 5038 -986 5228 -985
rect 5250 -986 5396 -975
rect 5407 -986 5441 -834
rect 5455 -853 5655 -827
rect 5461 -856 5643 -853
rect 5487 -857 5584 -856
rect 5597 -857 5643 -856
rect 5487 -872 5643 -857
rect 5509 -875 5643 -872
rect 5723 -861 6227 -827
rect 6247 -789 6393 -779
rect 6395 -780 6415 -779
rect 6427 -780 6429 -779
rect 6247 -805 6305 -789
rect 6311 -795 6393 -789
rect 6247 -861 6293 -805
rect 6317 -823 6393 -795
rect 6335 -857 6415 -823
rect 6335 -861 6393 -857
rect 5723 -871 6233 -861
rect 6247 -871 6435 -861
rect 6461 -871 6495 -356
rect 6509 -413 6548 -34
rect 6847 -53 6918 -19
rect 6994 -53 7122 -19
rect 7218 -43 7233 332
rect 6847 -55 6917 -53
rect 6651 -95 6717 -61
rect 6619 -114 6722 -102
rect 6619 -136 6733 -114
rect 6619 -142 6669 -136
rect 6718 -138 6733 -136
rect 6825 -120 6917 -55
rect 7029 -73 7041 -53
rect 7029 -83 7043 -73
rect 7073 -83 7075 -73
rect 7029 -89 7087 -83
rect 6711 -142 6745 -138
rect 6623 -152 6669 -142
rect 6699 -152 6745 -142
rect 6623 -195 6657 -152
rect 6699 -183 6704 -152
rect 6623 -310 6662 -195
rect 6508 -447 6548 -413
rect 6509 -471 6548 -447
rect 6628 -353 6662 -310
rect 6669 -322 6673 -184
rect 6711 -195 6745 -152
rect 6825 -154 6918 -120
rect 7032 -121 7084 -120
rect 6985 -154 7131 -121
rect 6711 -310 6750 -195
rect 6716 -322 6750 -310
rect 6669 -353 6674 -322
rect 6628 -369 6674 -353
rect 6701 -369 6750 -322
rect 6628 -403 6750 -369
rect 6628 -419 6674 -403
rect 6704 -419 6750 -403
rect 6825 -351 6917 -154
rect 6997 -184 7031 -154
rect 7085 -184 7119 -154
rect 6997 -199 7119 -184
rect 6996 -211 7119 -199
rect 6993 -216 7043 -211
rect 7073 -216 7123 -211
rect 7199 -216 7233 -43
rect 6993 -249 7123 -216
rect 6988 -256 7123 -249
rect 6988 -289 7118 -256
rect 6988 -294 7038 -289
rect 6992 -299 7038 -294
rect 7068 -294 7118 -289
rect 7068 -299 7115 -294
rect 6992 -317 7032 -299
rect 7074 -306 7115 -299
rect 7074 -317 7114 -306
rect 6992 -351 7026 -317
rect 7080 -351 7114 -317
rect 6825 -385 6918 -351
rect 6980 -384 7126 -351
rect 7137 -372 7148 -351
rect 7194 -366 7233 -216
rect 7252 298 7287 332
rect 7252 106 7286 298
rect 7585 236 7655 353
rect 7954 352 8007 388
rect 8359 354 8374 388
rect 8692 335 8762 431
rect 8874 418 8932 424
rect 8874 384 8886 418
rect 8874 378 8932 384
rect 7840 302 7853 319
rect 8692 318 8745 335
rect 7767 285 7825 291
rect 7767 251 7779 285
rect 7813 274 7825 285
rect 7937 262 7971 291
rect 8692 282 8763 318
rect 8824 282 8982 318
rect 7767 245 7825 251
rect 7366 106 7400 162
rect 7420 106 7422 186
rect 7448 106 7450 158
rect 7454 106 7488 162
rect 7568 159 7655 236
rect 7937 226 8007 262
rect 8359 231 8394 265
rect 7735 159 7769 208
rect 7823 159 7857 208
rect 7937 178 8025 226
rect 8086 178 8244 226
rect 7568 125 7656 159
rect 7723 125 7869 159
rect 7252 72 7287 106
rect 7354 72 7500 106
rect 7252 -72 7286 72
rect 7410 -30 7444 30
rect 7332 -72 7522 -46
rect 7252 -106 7287 -72
rect 7332 -80 7500 -72
rect 7348 -106 7500 -80
rect 7506 -106 7522 -72
rect 7252 -298 7286 -106
rect 7420 -186 7422 -106
rect 7448 -158 7450 -106
rect 7568 -125 7655 125
rect 7741 73 7769 95
rect 7813 73 7860 104
rect 7741 57 7781 73
rect 7811 57 7860 73
rect 7741 36 7860 57
rect 7748 30 7860 36
rect 7723 24 7869 30
rect 7763 23 7829 24
rect 7763 7 7781 23
rect 7811 7 7829 23
rect 7812 -23 7825 -17
rect 7763 -24 7829 -23
rect 7840 -24 7853 24
rect 7748 -36 7860 -24
rect 7741 -57 7860 -36
rect 7741 -73 7781 -57
rect 7811 -73 7851 -57
rect 7741 -91 7769 -73
rect 7735 -125 7769 -91
rect 7823 -91 7851 -73
rect 7823 -125 7857 -91
rect 7568 -159 7656 -125
rect 7717 -159 7869 -125
rect 7875 -159 7891 -125
rect 7568 -236 7655 -159
rect 7252 -332 7287 -298
rect 7585 -332 7655 -236
rect 7937 -178 8024 178
rect 8108 144 8164 158
rect 8325 130 8340 226
rect 8136 116 8192 130
rect 8148 90 8182 116
rect 8132 76 8198 90
rect 8136 70 8194 76
rect 8104 52 8138 56
rect 8192 52 8226 56
rect 8104 45 8150 52
rect 8180 45 8226 52
rect 8104 42 8144 45
rect 8186 42 8226 45
rect 8104 -28 8138 40
rect 8192 -28 8226 40
rect 8098 -38 8144 -28
rect 8186 -38 8226 -28
rect 8098 -40 8226 -38
rect 8098 -42 8220 -40
rect 8098 -52 8226 -42
rect 8104 -56 8138 -52
rect 8192 -56 8226 -52
rect 8070 -70 8164 -56
rect 8070 -76 8194 -70
rect 8070 -80 8198 -76
rect 8132 -90 8198 -80
rect 8148 -124 8182 -90
rect 8306 -130 8340 130
rect 7937 -226 8025 -178
rect 8086 -226 8244 -178
rect 8325 -226 8340 -130
rect 8359 173 8393 231
rect 8692 228 8762 282
rect 8852 228 8954 250
rect 8483 173 8585 197
rect 8692 194 8763 228
rect 8848 194 8958 228
rect 9063 222 9078 638
rect 8359 139 8394 173
rect 8470 145 8598 173
rect 8692 169 8762 194
rect 8874 184 8886 194
rect 8407 139 8661 145
rect 8359 -139 8393 139
rect 8505 129 8517 139
rect 8505 123 8563 129
rect 8551 87 8589 91
rect 8501 79 8519 87
rect 8479 71 8519 79
rect 8549 71 8589 87
rect 8479 53 8589 71
rect 8461 1 8607 53
rect 8467 -21 8513 -1
rect 8551 -21 8601 -1
rect 8467 -27 8519 -21
rect 8479 -37 8519 -27
rect 8549 -27 8601 -21
rect 8549 -37 8589 -27
rect 8479 -71 8589 -37
rect 8479 -79 8519 -71
rect 8501 -85 8519 -79
rect 8461 -87 8519 -85
rect 8549 -79 8589 -71
rect 8549 -85 8567 -79
rect 8549 -87 8607 -85
rect 8461 -91 8501 -87
rect 8567 -91 8607 -87
rect 8505 -129 8563 -123
rect 8505 -139 8517 -129
rect 8359 -173 8394 -139
rect 8490 -150 8578 -139
rect 8501 -162 8567 -150
rect 8490 -173 8578 -162
rect 8675 -169 8762 169
rect 8870 182 8888 184
rect 8918 182 8936 184
rect 8870 176 8936 182
rect 8870 166 8888 176
rect 8918 166 8936 176
rect 8855 126 8888 135
rect 8918 126 8967 135
rect 8855 123 8967 126
rect 8842 92 8967 123
rect 8842 76 8888 92
rect 8918 76 8964 92
rect 8842 -76 8876 76
rect 8930 -45 8964 76
rect 8920 -76 8967 -45
rect 8842 -92 8888 -76
rect 8918 -92 8967 -76
rect 8842 -123 8967 -92
rect 8855 -126 8967 -123
rect 8855 -135 8888 -126
rect 8870 -142 8888 -135
rect 8918 -135 8951 -126
rect 8918 -142 8936 -135
rect 8359 -226 8393 -173
rect 8692 -194 8762 -169
rect 8874 -182 8932 -176
rect 8874 -194 8886 -182
rect 7767 -251 7825 -245
rect 7767 -285 7779 -251
rect 7937 -262 8007 -226
rect 8359 -260 8374 -226
rect 8692 -228 8763 -194
rect 8859 -205 8947 -194
rect 8870 -217 8936 -205
rect 8859 -228 8947 -217
rect 9044 -222 9078 222
rect 7813 -285 7825 -270
rect 7767 -291 7825 -285
rect 7937 -291 7971 -262
rect 8692 -265 8762 -228
rect 8692 -282 8745 -265
rect 7840 -319 7853 -298
rect 8692 -318 8763 -282
rect 8824 -318 8982 -282
rect 6989 -385 7117 -384
rect 6825 -409 6912 -385
rect 6628 -466 6662 -419
rect 6716 -466 6750 -419
rect 6830 -430 6912 -409
rect 7024 -422 7082 -416
rect 6562 -471 6602 -466
rect 6616 -471 6816 -466
rect 6509 -528 6549 -471
rect 6605 -500 6816 -471
rect 6605 -505 6768 -500
rect 6610 -528 6768 -505
rect 6509 -600 6548 -528
rect 6509 -634 6549 -600
rect 6562 -623 6596 -528
rect 6616 -543 6662 -528
rect 6674 -543 6762 -528
rect 6628 -547 6662 -543
rect 6716 -547 6750 -543
rect 6708 -568 6766 -562
rect 6704 -580 6770 -568
rect 6690 -581 6770 -580
rect 6830 -573 6948 -430
rect 7024 -456 7036 -422
rect 7024 -462 7082 -456
rect 7194 -462 7228 -366
rect 7585 -368 7638 -332
rect 7937 -352 7971 -334
rect 7937 -353 8007 -352
rect 7936 -387 8007 -353
rect 7954 -388 8007 -387
rect 8359 -369 8394 -335
rect 7954 -422 8025 -388
rect 7621 -458 7656 -441
rect 7198 -494 7228 -462
rect 7585 -475 7656 -458
rect 6974 -547 7132 -524
rect 7218 -547 7228 -494
rect 7252 -528 7287 -494
rect 6974 -558 7137 -547
rect 6979 -573 7137 -558
rect 6830 -581 7199 -573
rect 6690 -584 6708 -581
rect 6672 -600 6706 -590
rect 6720 -600 6744 -581
rect 6830 -600 6948 -581
rect 6610 -623 6948 -600
rect 6562 -627 6948 -623
rect 7218 -627 7233 -547
rect 6562 -634 6971 -627
rect 6509 -692 6548 -634
rect 6509 -726 6549 -692
rect 6509 -863 6548 -726
rect 5509 -879 5637 -875
rect 5509 -887 5655 -879
rect 5521 -891 5546 -887
rect 5549 -890 5611 -887
rect 5549 -891 5599 -890
rect 5604 -891 5611 -890
rect 5549 -895 5615 -891
rect 5549 -901 5611 -895
rect 5549 -919 5580 -901
rect 5549 -925 5611 -919
rect 5632 -925 5639 -887
rect 5723 -895 6509 -871
rect 6514 -895 6548 -863
rect 5723 -925 6227 -895
rect 6247 -925 6293 -895
rect 6347 -925 6381 -895
rect 6385 -925 6393 -916
rect 6461 -925 6495 -895
rect 6509 -925 6548 -895
rect 5549 -929 5643 -925
rect 5723 -929 6509 -925
rect 5521 -933 5546 -929
rect 5549 -930 5599 -929
rect 5604 -930 5611 -929
rect 5549 -933 5611 -930
rect 5632 -933 5639 -929
rect 5509 -948 5643 -933
rect 5487 -959 5643 -948
rect 5487 -964 5567 -959
rect 5575 -964 5584 -959
rect 5597 -964 5643 -959
rect 5461 -967 5567 -964
rect 5584 -965 5643 -964
rect 5572 -967 5643 -965
rect 5723 -959 6233 -929
rect 6247 -959 6435 -929
rect 5038 -993 5441 -986
rect 5455 -973 5655 -967
rect 5723 -973 6227 -959
rect 5455 -993 6227 -973
rect 5038 -1001 6227 -993
rect 5038 -1008 5561 -1001
rect 5572 -1005 5589 -1001
rect 5038 -1073 5073 -1008
rect 5138 -1011 5198 -1008
rect 5150 -1020 5186 -1011
rect 5240 -1020 5296 -1008
rect 5350 -1014 5561 -1008
rect 5350 -1020 5396 -1014
rect 5407 -1020 5441 -1014
rect 5086 -1027 5441 -1020
rect 5450 -1027 5496 -1014
rect 5509 -1023 5561 -1014
rect 5567 -1010 5589 -1005
rect 5567 -1023 5584 -1010
rect 5597 -1023 5655 -1001
rect 5521 -1027 5546 -1023
rect 5567 -1027 5596 -1023
rect 5609 -1027 5618 -1023
rect 5723 -1027 6227 -1001
rect 5086 -1035 6227 -1027
rect 5086 -1048 5697 -1035
rect 5086 -1054 5396 -1048
rect 5407 -1054 5441 -1048
rect 5450 -1054 5697 -1048
rect 4542 -1083 4703 -1082
rect 4717 -1083 5005 -1073
rect 4542 -1092 5005 -1083
rect 4550 -1114 4734 -1092
rect 4751 -1107 5005 -1092
rect 5038 -1107 5072 -1073
rect 4414 -1116 4734 -1114
rect 4746 -1116 4751 -1107
rect 4764 -1110 4805 -1107
rect 4817 -1110 4917 -1107
rect 4764 -1116 4917 -1110
rect 4133 -1145 4167 -1123
rect 4179 -1145 4281 -1122
rect 4045 -1148 4281 -1145
rect 4288 -1148 4346 -1122
rect 4414 -1126 4602 -1116
rect 4616 -1117 4737 -1116
rect 4746 -1117 4764 -1116
rect 4771 -1117 4817 -1116
rect 4824 -1117 4829 -1116
rect 4844 -1117 4851 -1116
rect 4859 -1117 4917 -1116
rect 4932 -1117 4939 -1107
rect 4951 -1117 4966 -1107
rect 4985 -1117 5019 -1107
rect 4616 -1126 4734 -1117
rect 4348 -1148 4388 -1126
rect 4402 -1132 4734 -1126
rect 4764 -1132 4932 -1117
rect 4960 -1132 5019 -1117
rect 4402 -1141 5019 -1132
rect 5033 -1141 5072 -1107
rect 5086 -1141 5120 -1054
rect 5150 -1064 5186 -1054
rect 5221 -1064 5308 -1054
rect 5150 -1076 5184 -1064
rect 5228 -1076 5336 -1064
rect 5150 -1080 5196 -1076
rect 5243 -1080 5336 -1076
rect 5150 -1082 5336 -1080
rect 5150 -1094 5196 -1082
rect 5150 -1098 5184 -1094
rect 5243 -1097 5336 -1082
rect 5262 -1098 5296 -1097
rect 5180 -1116 5278 -1114
rect 5180 -1122 5290 -1116
rect 5308 -1122 5336 -1097
rect 5354 -1094 5396 -1054
rect 5402 -1061 5697 -1054
rect 5723 -1041 6227 -1035
rect 6247 -1015 6293 -959
rect 6317 -963 6393 -959
rect 6317 -972 6415 -963
rect 6335 -997 6415 -972
rect 6335 -1007 6393 -997
rect 6303 -1015 6393 -1007
rect 6247 -1028 6393 -1015
rect 6247 -1041 6387 -1028
rect 6395 -1041 6415 -1040
rect 6427 -1041 6429 -1040
rect 5180 -1125 5337 -1122
rect 5180 -1131 5294 -1125
rect 5308 -1131 5336 -1125
rect 5150 -1132 5336 -1131
rect 5150 -1141 5154 -1132
rect 5206 -1141 5230 -1132
rect 5244 -1141 5268 -1132
rect 5308 -1141 5336 -1132
rect 5354 -1141 5388 -1094
rect 5402 -1141 5441 -1061
rect 5450 -1094 5495 -1061
rect 5549 -1079 5599 -1061
rect 5615 -1069 5631 -1061
rect 5538 -1087 5599 -1079
rect 5508 -1094 5599 -1087
rect 5613 -1094 5663 -1069
rect 5455 -1141 5489 -1094
rect 5549 -1095 5663 -1094
rect 5723 -1075 6213 -1041
rect 6241 -1044 6393 -1041
rect 6241 -1075 6441 -1044
rect 5549 -1101 5659 -1095
rect 5549 -1111 5584 -1101
rect 5597 -1103 5659 -1101
rect 5601 -1109 5659 -1103
rect 5563 -1122 5584 -1111
rect 5723 -1113 6227 -1075
rect 5525 -1129 5632 -1122
rect 5563 -1137 5632 -1129
rect 5698 -1133 6227 -1113
rect 6247 -1081 6387 -1075
rect 6247 -1127 6299 -1081
rect 6301 -1127 6341 -1081
rect 6347 -1127 6387 -1081
rect 6247 -1133 6387 -1127
rect 6389 -1133 6419 -1075
rect 6427 -1133 6429 -1075
rect 6436 -1133 6441 -1075
rect 5623 -1141 5632 -1137
rect 5689 -1141 5691 -1137
rect 4402 -1148 5632 -1141
rect 4020 -1150 4334 -1148
rect 4020 -1159 4299 -1150
rect 4020 -1168 4288 -1159
rect 4300 -1168 4334 -1150
rect 4335 -1159 5632 -1148
rect 4346 -1160 5632 -1159
rect 4346 -1168 4382 -1160
rect 4402 -1168 4548 -1160
rect 4600 -1163 5632 -1160
rect 5651 -1163 5660 -1141
rect 5670 -1163 5697 -1141
rect 5698 -1163 6213 -1133
rect 4600 -1168 5725 -1163
rect 4000 -1179 4019 -1168
rect 4020 -1169 5725 -1168
rect 5737 -1167 6213 -1163
rect 6241 -1167 6441 -1133
rect 5737 -1169 6227 -1167
rect 4020 -1179 6227 -1169
rect 3979 -1182 6227 -1179
rect 1126 -1198 1210 -1192
rect 1126 -1237 1160 -1198
rect 1002 -1252 1160 -1237
rect 1196 -1206 1210 -1198
rect 1196 -1252 1254 -1206
rect 1272 -1218 3971 -1191
rect 1284 -1244 3971 -1218
rect 3979 -1213 4179 -1182
rect 4200 -1202 4334 -1182
rect 4348 -1202 4382 -1182
rect 4414 -1202 4448 -1182
rect 4489 -1194 4587 -1182
rect 4466 -1202 4587 -1194
rect 4616 -1197 6227 -1182
rect 6247 -1177 6387 -1167
rect 6247 -1183 6305 -1177
rect 6307 -1183 6387 -1177
rect 6247 -1193 6387 -1183
rect 6247 -1196 6299 -1193
rect 6301 -1196 6341 -1193
rect 6347 -1196 6387 -1193
rect 4616 -1200 5660 -1197
rect 5670 -1200 5697 -1197
rect 5698 -1200 5725 -1197
rect 4616 -1202 5632 -1200
rect 4200 -1213 5632 -1202
rect 3979 -1244 4019 -1213
rect 4045 -1244 4079 -1213
rect 4091 -1244 4121 -1213
rect 4133 -1244 4167 -1213
rect 4200 -1236 4233 -1213
rect 4200 -1244 4246 -1236
rect 4247 -1244 4281 -1213
rect 4295 -1216 5632 -1213
rect 4295 -1244 4334 -1216
rect 1284 -1252 4340 -1244
rect 0 -1271 791 -1267
rect 0 -1279 774 -1271
rect 121 -1281 139 -1279
rect 119 -1303 124 -1281
rect 187 -1285 209 -1281
rect 136 -1289 261 -1285
rect 187 -1303 209 -1289
rect 161 -1319 166 -1303
rect 187 -1319 227 -1303
rect 161 -1323 227 -1319
rect 161 -1367 166 -1323
rect 195 -1353 227 -1323
rect 161 -1369 227 -1367
rect 229 -1369 269 -1323
rect 229 -1387 261 -1369
rect 229 -1389 295 -1387
rect 106 -1421 208 -1391
rect 354 -1406 370 -1279
rect 388 -1368 422 -1279
rect 530 -1316 566 -1279
rect 618 -1288 774 -1279
rect 899 -1281 912 -1252
rect 942 -1281 965 -1252
rect 1000 -1279 1030 -1252
rect 1073 -1260 1160 -1252
rect 1036 -1271 1318 -1260
rect 1036 -1277 1073 -1271
rect 1098 -1276 1318 -1271
rect 1000 -1281 1073 -1279
rect 670 -1304 700 -1288
rect 704 -1304 774 -1288
rect 1002 -1294 1073 -1281
rect 1098 -1280 1322 -1276
rect 1335 -1280 4340 -1252
rect 1098 -1294 4340 -1280
rect 700 -1338 704 -1334
rect 712 -1338 774 -1304
rect 932 -1333 936 -1304
rect 670 -1368 700 -1338
rect 704 -1368 774 -1338
rect 871 -1342 961 -1333
rect 989 -1338 1041 -1333
rect 972 -1342 1080 -1338
rect 1092 -1342 1107 -1294
rect 1126 -1303 1161 -1294
rect 1212 -1297 4340 -1294
rect 1126 -1314 1169 -1303
rect 1212 -1304 1512 -1297
rect 1212 -1314 1322 -1304
rect 1331 -1313 1514 -1304
rect 1331 -1314 1585 -1313
rect 871 -1344 1107 -1342
rect 882 -1354 950 -1344
rect 912 -1356 942 -1354
rect 901 -1367 953 -1356
rect 958 -1367 1107 -1344
rect 1335 -1324 1585 -1314
rect 1335 -1336 1574 -1324
rect 1335 -1342 1585 -1336
rect 1335 -1347 1586 -1342
rect 1335 -1350 1512 -1347
rect 388 -1372 423 -1368
rect 483 -1372 535 -1368
rect 700 -1372 704 -1368
rect 388 -1379 535 -1372
rect 388 -1391 532 -1379
rect 388 -1402 535 -1391
rect 570 -1402 638 -1388
rect 712 -1391 774 -1368
rect 701 -1402 774 -1391
rect 992 -1401 1141 -1376
rect 1337 -1381 1586 -1376
rect 1668 -1383 4340 -1297
rect 721 -1403 774 -1402
rect 83 -1423 335 -1421
rect 83 -1432 221 -1423
rect 283 -1432 335 -1423
rect 93 -1444 221 -1432
rect 294 -1444 324 -1432
rect 354 -1436 498 -1406
rect 1042 -1410 1044 -1401
rect 570 -1436 604 -1422
rect 1681 -1438 4340 -1383
rect 4348 -1438 4382 -1216
rect 4414 -1236 4448 -1216
rect 4466 -1220 4587 -1216
rect 4489 -1228 4587 -1220
rect 4388 -1239 4448 -1236
rect 4490 -1239 4587 -1228
rect 4388 -1262 4587 -1239
rect 4616 -1220 5632 -1216
rect 4616 -1223 5637 -1220
rect 5740 -1223 6227 -1197
rect 6259 -1200 6293 -1196
rect 4616 -1231 6227 -1223
rect 6259 -1224 6293 -1220
rect 6301 -1224 6383 -1196
rect 6389 -1212 6419 -1167
rect 6389 -1224 6415 -1212
rect 4616 -1257 5703 -1231
rect 5737 -1257 6227 -1231
rect 4388 -1270 4556 -1262
rect 4388 -1278 4588 -1270
rect 4388 -1281 4538 -1278
rect 4388 -1286 4542 -1281
rect 4388 -1309 4460 -1286
rect 4470 -1305 4542 -1286
rect 4554 -1305 4588 -1278
rect 4462 -1307 4542 -1305
rect 4462 -1309 4549 -1307
rect 4550 -1309 4588 -1305
rect 4388 -1320 4588 -1309
rect 4388 -1334 4542 -1320
rect 4388 -1336 4454 -1334
rect 4414 -1348 4454 -1336
rect 4402 -1350 4454 -1348
rect 4456 -1350 4542 -1334
rect 4402 -1360 4542 -1350
rect 4402 -1366 4460 -1360
rect 4462 -1366 4542 -1360
rect 4402 -1400 4542 -1366
rect 4544 -1321 4570 -1320
rect 4544 -1400 4574 -1321
rect 4582 -1348 4588 -1320
rect 4616 -1291 5637 -1257
rect 4582 -1370 4596 -1348
rect 4585 -1389 4596 -1370
rect 4402 -1416 4460 -1400
rect 4462 -1404 4538 -1400
rect 4550 -1404 4574 -1400
rect 4462 -1416 4536 -1404
rect 4402 -1438 4448 -1416
rect 4462 -1438 4496 -1416
rect 4502 -1438 4536 -1416
rect 4550 -1438 4584 -1404
rect 4591 -1438 4596 -1389
rect 4616 -1353 5639 -1291
rect 5689 -1325 5691 -1257
rect 5698 -1321 5703 -1257
rect 5723 -1321 6227 -1257
rect 4616 -1359 5632 -1353
rect 5723 -1359 5725 -1321
rect 5737 -1345 6227 -1321
rect 6247 -1227 6299 -1224
rect 6247 -1237 6305 -1227
rect 6307 -1228 6393 -1224
rect 6395 -1228 6415 -1224
rect 6427 -1228 6429 -1167
rect 6436 -1224 6441 -1167
rect 6335 -1237 6393 -1228
rect 6247 -1271 6393 -1237
rect 6247 -1277 6415 -1271
rect 6247 -1293 6305 -1277
rect 6247 -1345 6293 -1293
rect 6335 -1305 6415 -1277
rect 6335 -1321 6393 -1305
rect 6347 -1336 6393 -1321
rect 6347 -1345 6381 -1336
rect 4616 -1397 5647 -1359
rect 5737 -1385 6210 -1345
rect 6241 -1368 6415 -1345
rect 4616 -1424 5655 -1397
rect 5735 -1402 6210 -1385
rect 6236 -1373 6415 -1368
rect 6236 -1402 6447 -1373
rect 5735 -1407 6233 -1402
rect 6247 -1407 6447 -1402
rect 4616 -1438 5643 -1424
rect 5735 -1427 6210 -1407
rect 83 -1455 221 -1444
rect 283 -1455 335 -1444
rect 816 -1480 820 -1446
rect 1374 -1474 1376 -1446
rect 1342 -1480 1376 -1474
rect 1681 -1461 5643 -1438
rect 1681 -1472 5709 -1461
rect 1640 -1585 1650 -1478
rect 1086 -1628 1088 -1590
rect 1668 -1613 1678 -1478
rect 1681 -1489 4340 -1472
rect 1681 -1506 2200 -1489
rect 2234 -1506 2296 -1489
rect 2322 -1506 4340 -1489
rect 1681 -1510 2120 -1506
rect 1846 -1516 1865 -1510
rect 1850 -1528 1865 -1516
rect 1907 -1538 1918 -1510
rect 1919 -1516 1953 -1510
rect 1919 -1528 1952 -1516
rect 1907 -1550 1933 -1538
rect 2033 -1550 2043 -1510
rect 2050 -1550 2120 -1510
rect 2138 -1514 2158 -1506
rect 2188 -1514 2195 -1506
rect 2276 -1536 2296 -1506
rect 2402 -1536 2436 -1506
rect 2442 -1536 4340 -1506
rect 1124 -1664 1126 -1628
rect 1717 -1693 1751 -1550
rect 1819 -1553 1877 -1550
rect 1907 -1553 1965 -1550
rect 1825 -1659 1838 -1616
rect 1844 -1656 1850 -1604
rect 1859 -1625 1872 -1591
rect 1875 -1598 1888 -1591
rect 1906 -1598 1909 -1591
rect 1875 -1625 1909 -1598
rect 2033 -1604 2120 -1550
rect 2140 -1550 2246 -1536
rect 2266 -1542 4340 -1536
rect 2266 -1546 2615 -1542
rect 2628 -1546 4340 -1542
rect 2266 -1550 2613 -1546
rect 2628 -1548 2657 -1546
rect 2140 -1559 2613 -1550
rect 2663 -1551 4340 -1546
rect 2140 -1582 2628 -1559
rect 2140 -1587 2613 -1582
rect 2140 -1593 2659 -1587
rect 2663 -1593 3212 -1551
rect 2140 -1595 3212 -1593
rect 2140 -1599 2841 -1595
rect 2140 -1604 2246 -1599
rect 2266 -1604 2841 -1599
rect 1884 -1646 1894 -1632
rect 1908 -1641 1918 -1632
rect 1908 -1646 1928 -1641
rect 1804 -1666 1838 -1659
rect 1884 -1659 1928 -1646
rect 1944 -1659 1956 -1604
rect 1884 -1682 1990 -1659
rect 2033 -1666 2112 -1604
rect 2114 -1656 2120 -1604
rect 2208 -1616 2209 -1604
rect 2231 -1616 2266 -1604
rect 2138 -1656 2158 -1632
rect 2166 -1637 2266 -1616
rect 2114 -1666 2158 -1656
rect 2033 -1693 2103 -1666
rect 2132 -1676 2158 -1666
rect 2132 -1682 2148 -1676
rect 1717 -1694 2103 -1693
rect 2208 -1693 2209 -1637
rect 2228 -1640 2266 -1637
rect 2278 -1616 2316 -1608
rect 2342 -1616 2436 -1604
rect 2278 -1632 2436 -1616
rect 2278 -1637 2342 -1632
rect 2278 -1640 2328 -1637
rect 2228 -1679 2328 -1640
rect 2213 -1680 2328 -1679
rect 2213 -1686 2290 -1680
rect 2308 -1682 2328 -1680
rect 2354 -1666 2436 -1632
rect 2440 -1641 2490 -1604
rect 2563 -1641 2574 -1616
rect 2597 -1627 2742 -1604
rect 2601 -1633 2663 -1627
rect 2616 -1641 2663 -1633
rect 2674 -1641 2742 -1627
rect 2771 -1641 2805 -1604
rect 2354 -1682 2422 -1666
rect 2213 -1693 2266 -1686
rect 2354 -1693 2436 -1682
rect 2208 -1694 2436 -1693
rect 2440 -1693 2498 -1641
rect 2528 -1693 2586 -1641
rect 2616 -1693 2805 -1641
rect 2832 -1682 2839 -1616
rect 2841 -1693 2878 -1604
rect 3132 -1632 3144 -1604
rect 3180 -1616 3212 -1595
rect 3216 -1582 3231 -1551
rect 3241 -1582 3275 -1551
rect 3355 -1578 3389 -1551
rect 3400 -1578 3401 -1551
rect 3431 -1578 3434 -1551
rect 3532 -1578 4340 -1551
rect 3277 -1582 3329 -1578
rect 3343 -1582 3489 -1578
rect 3509 -1582 4340 -1578
rect 3216 -1612 4340 -1582
rect 4348 -1610 4382 -1472
rect 4396 -1489 4596 -1472
rect 4396 -1491 4542 -1489
rect 4396 -1498 4549 -1491
rect 4616 -1495 5709 -1472
rect 5723 -1478 6210 -1427
rect 6259 -1454 6293 -1407
rect 6347 -1423 6381 -1407
rect 6259 -1470 6305 -1454
rect 6332 -1470 6381 -1423
rect 6461 -1464 6495 -929
rect 6514 -957 6548 -925
rect 6509 -1094 6548 -957
rect 6562 -808 6596 -634
rect 6660 -636 6718 -634
rect 6676 -649 6710 -645
rect 6722 -649 6746 -646
rect 6764 -649 6798 -645
rect 6664 -658 6722 -649
rect 6628 -668 6662 -658
rect 6664 -664 6750 -658
rect 6752 -659 6810 -649
rect 6670 -668 6710 -664
rect 6628 -677 6710 -668
rect 6616 -686 6710 -677
rect 6716 -677 6750 -664
rect 6716 -686 6756 -677
rect 6616 -692 6756 -686
rect 6758 -692 6802 -659
rect 6805 -692 6810 -659
rect 6610 -726 6810 -692
rect 6616 -752 6756 -726
rect 6616 -808 6668 -752
rect 6670 -808 6710 -752
rect 6716 -808 6756 -752
rect 6758 -774 6788 -726
rect 6796 -774 6798 -726
rect 6758 -808 6798 -774
rect 6805 -808 6810 -726
rect 6830 -661 6971 -634
rect 7025 -650 7091 -633
rect 7165 -643 7185 -627
rect 7252 -643 7286 -528
rect 7014 -661 7102 -650
rect 7199 -661 7219 -643
rect 7246 -661 7286 -643
rect 6830 -755 6965 -661
rect 7029 -683 7041 -661
rect 7073 -683 7091 -671
rect 7029 -689 7091 -683
rect 7073 -699 7091 -689
rect 6997 -721 6999 -717
rect 7089 -721 7153 -699
rect 7213 -721 7233 -661
rect 6985 -733 7031 -721
rect 6985 -755 7019 -733
rect 7051 -755 7153 -721
rect 7199 -755 7233 -721
rect 6830 -781 6971 -755
rect 6985 -781 7233 -755
rect 6830 -789 7233 -781
rect 6830 -808 6965 -789
rect 6562 -842 6602 -808
rect 6616 -829 6810 -808
rect 6816 -817 6965 -808
rect 6985 -811 7037 -789
rect 7057 -797 7079 -789
rect 7045 -801 7079 -797
rect 6997 -815 7031 -811
rect 6616 -838 6762 -829
rect 6830 -835 6965 -817
rect 7039 -818 7079 -801
rect 7085 -811 7125 -789
rect 7133 -801 7167 -797
rect 7085 -815 7119 -811
rect 7127 -814 7179 -801
rect 7033 -833 7079 -818
rect 7127 -823 7167 -814
rect 7033 -835 7091 -833
rect 7127 -835 7161 -823
rect 7165 -835 7167 -823
rect 7174 -835 7179 -814
rect 6616 -842 6792 -838
rect 6562 -978 6596 -842
rect 6616 -857 6668 -842
rect 6616 -963 6662 -857
rect 6716 -860 6762 -842
rect 6704 -876 6762 -860
rect 6830 -849 7179 -835
rect 6704 -944 6784 -876
rect 6704 -960 6762 -944
rect 6616 -978 6668 -963
rect 6716 -975 6762 -960
rect 6830 -955 6965 -849
rect 6979 -869 6999 -849
rect 7025 -858 7179 -849
rect 7014 -869 7179 -858
rect 7033 -875 7161 -869
rect 7165 -875 7167 -869
rect 7174 -875 7179 -869
rect 7033 -879 7179 -875
rect 7025 -891 7179 -879
rect 7199 -835 7233 -789
rect 7199 -869 7201 -835
rect 7213 -869 7233 -835
rect 7025 -895 7091 -891
rect 7121 -895 7167 -891
rect 7025 -897 7139 -895
rect 7025 -899 7091 -897
rect 7073 -907 7091 -899
rect 7121 -907 7139 -897
rect 7011 -925 7075 -907
rect 7089 -923 7123 -917
rect 7077 -925 7135 -923
rect 7011 -929 7079 -925
rect 7089 -929 7123 -925
rect 7133 -929 7167 -925
rect 7011 -941 7161 -929
rect 7033 -951 7161 -941
rect 7165 -951 7167 -929
rect 7174 -951 7179 -929
rect 6979 -955 6999 -951
rect 7014 -955 7179 -951
rect 6716 -978 6756 -975
rect 6830 -977 7179 -955
rect 7199 -951 7233 -869
rect 7199 -977 7201 -951
rect 6562 -1012 6602 -978
rect 6616 -991 6762 -978
rect 6830 -985 7201 -977
rect 7213 -985 7233 -951
rect 6616 -1012 6810 -991
rect 6509 -1128 6549 -1094
rect 6509 -1186 6548 -1128
rect 6509 -1220 6549 -1186
rect 6509 -1292 6548 -1220
rect 6562 -1292 6596 -1012
rect 6616 -1068 6668 -1012
rect 6670 -1037 6710 -1012
rect 6716 -1037 6756 -1012
rect 6670 -1068 6756 -1037
rect 6616 -1094 6756 -1068
rect 6758 -1094 6788 -1012
rect 6796 -1094 6798 -1012
rect 6805 -1094 6810 -1012
rect 6610 -1128 6810 -1094
rect 6616 -1132 6756 -1128
rect 6758 -1132 6788 -1128
rect 6796 -1132 6798 -1128
rect 6805 -1132 6810 -1128
rect 6616 -1134 6810 -1132
rect 6616 -1143 6668 -1134
rect 6628 -1147 6662 -1143
rect 6670 -1156 6710 -1134
rect 6716 -1143 6810 -1134
rect 6716 -1147 6750 -1143
rect 6664 -1159 6719 -1156
rect 6664 -1171 6722 -1159
rect 6752 -1171 6810 -1143
rect 6830 -1031 6965 -985
rect 7033 -987 7091 -985
rect 6993 -1009 7031 -997
rect 7033 -1002 7079 -987
rect 6985 -1031 7037 -1009
rect 7039 -1019 7079 -1002
rect 7045 -1023 7079 -1019
rect 7085 -997 7107 -991
rect 7085 -1009 7119 -997
rect 7085 -1031 7125 -1009
rect 7127 -1019 7179 -985
rect 7133 -1023 7167 -1019
rect 7199 -1031 7233 -985
rect 7247 -888 7286 -661
rect 7420 -680 7422 -640
rect 7585 -644 7655 -475
rect 7767 -543 7825 -537
rect 7767 -577 7779 -543
rect 7767 -583 7825 -577
rect 7585 -646 7686 -644
rect 7448 -680 7450 -668
rect 7454 -680 7488 -664
rect 7300 -736 7340 -680
rect 7354 -736 7554 -680
rect 7568 -736 7686 -646
rect 7247 -932 7287 -888
rect 6830 -1065 6971 -1031
rect 6985 -1057 7219 -1031
rect 6985 -1065 7150 -1057
rect 7199 -1065 7219 -1057
rect 6830 -1159 6965 -1065
rect 6985 -1099 7019 -1065
rect 7051 -1087 7153 -1065
rect 7073 -1099 7131 -1087
rect 6997 -1103 6999 -1099
rect 7073 -1107 7133 -1099
rect 7213 -1125 7233 -1065
rect 7041 -1131 7075 -1125
rect 7029 -1137 7087 -1131
rect 7029 -1159 7041 -1137
rect 7199 -1159 7233 -1125
rect 7247 -1159 7286 -932
rect 7300 -1084 7334 -736
rect 7354 -758 7388 -736
rect 7420 -758 7500 -744
rect 7366 -762 7368 -758
rect 7454 -762 7488 -758
rect 7446 -782 7504 -776
rect 7442 -796 7508 -782
rect 7420 -816 7444 -796
rect 7458 -816 7492 -796
rect 7582 -800 7686 -736
rect 7394 -830 7508 -816
rect 7398 -836 7508 -830
rect 7442 -838 7508 -836
rect 7446 -844 7504 -838
rect 7414 -854 7448 -850
rect 7502 -854 7536 -850
rect 7402 -861 7460 -854
rect 7408 -864 7460 -861
rect 7414 -869 7460 -864
rect 7490 -869 7536 -854
rect 7414 -872 7454 -869
rect 7496 -872 7536 -869
rect 7414 -888 7448 -872
rect 7502 -888 7536 -872
rect 7543 -888 7548 -854
rect 7568 -888 7686 -800
rect 7723 -804 7781 -779
rect 7811 -804 7869 -779
rect 7954 -792 8024 -422
rect 8158 -656 8164 -534
rect 8186 -652 8192 -562
rect 8136 -690 8194 -684
rect 8136 -724 8148 -690
rect 8136 -730 8194 -724
rect 7735 -808 7769 -804
rect 7823 -808 7857 -804
rect 7840 -833 7853 -817
rect 7954 -826 8025 -792
rect 8325 -807 8340 -388
rect 8359 -739 8393 -369
rect 8505 -437 8563 -431
rect 8505 -471 8517 -437
rect 8505 -477 8563 -471
rect 8505 -637 8563 -631
rect 8505 -671 8517 -637
rect 8505 -677 8563 -671
rect 8692 -702 8762 -318
rect 8874 -384 8932 -378
rect 8874 -418 8886 -384
rect 8874 -424 8932 -418
rect 8874 -692 8932 -686
rect 8874 -702 8886 -692
rect 9063 -702 9078 -222
rect 9097 371 9131 638
rect 9177 600 9367 620
rect 9413 614 9483 638
rect 9430 604 9562 614
rect 9642 604 9816 614
rect 10512 604 10794 634
rect 9205 572 9251 592
rect 9293 572 9339 592
rect 9430 580 9501 604
rect 10811 600 10881 638
rect 9199 412 9239 425
rect 9305 412 9345 425
rect 9430 424 9500 580
rect 10811 564 10864 600
rect 11182 547 11197 638
rect 11216 547 11250 638
rect 11358 604 11424 630
rect 11374 600 11408 604
rect 11532 590 11619 638
rect 11787 636 11806 638
rect 11703 600 11817 611
rect 11906 604 11988 638
rect 9580 424 9614 444
rect 9668 424 9702 444
rect 9430 390 9501 424
rect 9568 390 9714 424
rect 9097 337 9132 371
rect 9228 360 9316 371
rect 9239 348 9305 360
rect 9228 337 9316 348
rect 9097 263 9131 337
rect 9243 331 9255 337
rect 9243 327 9301 331
rect 9239 315 9305 327
rect 9255 275 9289 297
rect 9430 275 9500 390
rect 9580 360 9614 390
rect 9668 360 9702 390
rect 9580 350 9702 360
rect 9580 346 9614 350
rect 9668 346 9702 350
rect 9608 312 9674 322
rect 9624 288 9658 312
rect 9608 278 9674 288
rect 9243 269 9301 275
rect 9243 263 9255 269
rect 9097 229 9132 263
rect 9228 252 9316 263
rect 9239 242 9305 252
rect 9145 229 9399 242
rect 9097 175 9131 229
rect 9413 210 9500 275
rect 9580 250 9614 254
rect 9668 250 9702 254
rect 9580 247 9626 250
rect 9656 247 9702 250
rect 9580 238 9614 247
rect 9668 238 9702 247
rect 9211 175 9245 209
rect 9299 175 9333 209
rect 9413 176 9501 210
rect 9568 176 9714 210
rect 9097 141 9132 175
rect 9193 141 9345 175
rect 9351 141 9367 175
rect 9097 -141 9131 141
rect 9217 89 9245 111
rect 9289 89 9336 120
rect 9217 73 9257 89
rect 9287 73 9336 89
rect 9217 46 9336 73
rect 9199 8 9345 46
rect 9413 20 9500 176
rect 9782 82 9816 518
rect 11216 513 11231 547
rect 11549 494 11619 590
rect 11731 572 11789 583
rect 11731 543 11743 572
rect 11731 537 11789 543
rect 11549 458 11602 494
rect 11918 441 11988 604
rect 12122 558 12128 600
rect 12150 562 12156 600
rect 12072 544 12128 558
rect 12100 524 12158 530
rect 12100 516 12156 524
rect 12100 490 12112 516
rect 12100 484 12158 490
rect 12270 484 12304 638
rect 11918 405 11971 441
rect 12289 388 12304 484
rect 12323 388 12357 638
rect 12465 637 12495 638
rect 12524 637 12531 671
rect 12558 638 12565 672
rect 12590 653 12726 672
rect 12800 671 12934 672
rect 12566 639 12726 653
rect 12768 639 12966 671
rect 12974 639 13095 672
rect 13192 661 13280 672
rect 13343 668 13411 672
rect 13447 668 13473 672
rect 13668 670 13701 672
rect 13203 649 13269 661
rect 13192 646 13280 649
rect 13343 646 13506 668
rect 13109 639 13506 646
rect 12566 638 13506 639
rect 13640 653 13834 668
rect 14073 653 15583 672
rect 13640 639 15583 653
rect 15629 639 15780 672
rect 15810 666 15952 702
rect 16064 690 16076 702
rect 16064 684 16122 690
rect 13640 638 15780 639
rect 12403 600 12593 627
rect 12431 572 12477 599
rect 12519 572 12565 599
rect 12469 471 12527 477
rect 12469 437 12481 471
rect 12469 431 12527 437
rect 12639 431 12726 638
rect 12806 600 12840 633
rect 12894 600 12928 633
rect 12323 354 12338 388
rect 12656 335 12726 431
rect 12838 418 12896 424
rect 12838 384 12850 418
rect 12838 378 12896 384
rect 12656 299 12709 335
rect 13027 282 13042 638
rect 13061 282 13095 638
rect 13141 600 13331 620
rect 13377 614 13447 638
rect 13394 604 13526 614
rect 13606 604 13780 614
rect 14476 604 14758 634
rect 13169 572 13215 592
rect 13257 572 13303 592
rect 13394 580 13465 604
rect 14775 600 14845 638
rect 13207 365 13265 371
rect 13207 331 13219 365
rect 13207 325 13265 331
rect 13061 248 13076 282
rect 13394 229 13464 580
rect 14775 564 14828 600
rect 15146 547 15161 638
rect 15180 547 15214 638
rect 15322 604 15388 630
rect 15338 600 15372 604
rect 15496 590 15583 638
rect 15751 636 15770 638
rect 15667 600 15781 611
rect 15180 513 15195 547
rect 15513 494 15583 590
rect 15695 572 15753 583
rect 15695 543 15707 572
rect 15695 537 15753 543
rect 15513 458 15566 494
rect 15882 441 15952 666
rect 16064 524 16122 530
rect 16064 490 16076 524
rect 16064 484 16122 490
rect 15882 405 15935 441
rect 16253 388 16268 773
rect 16287 739 16322 773
rect 16287 388 16321 739
rect 16433 671 16491 677
rect 16433 637 16445 671
rect 16433 631 16491 637
rect 16433 471 16491 477
rect 16433 437 16445 471
rect 16433 431 16491 437
rect 16287 354 16302 388
rect 16620 335 16690 794
rect 16894 793 17411 827
rect 17632 810 17780 844
rect 17490 793 17780 810
rect 17814 842 17872 848
rect 17814 808 17826 842
rect 17814 802 17872 808
rect 16894 776 17780 793
rect 16972 775 17006 776
rect 16802 726 16860 732
rect 16802 692 16814 726
rect 16802 686 16860 692
rect 16802 418 16860 424
rect 16802 384 16814 418
rect 16802 378 16860 384
rect 16620 299 16673 335
rect 16991 282 17006 775
rect 17025 741 17060 775
rect 17263 759 17553 776
rect 17025 282 17059 741
rect 17263 723 17411 759
rect 17632 740 17780 776
rect 17632 723 17685 740
rect 17171 673 17229 679
rect 17171 639 17183 673
rect 17632 670 17665 723
rect 18003 706 18018 1252
rect 18037 706 18071 1253
rect 18183 1243 18195 1253
rect 18183 1237 18241 1243
rect 18183 789 18241 795
rect 18183 755 18195 789
rect 18183 749 18241 755
rect 18037 672 18052 706
rect 17341 650 17375 668
rect 18372 653 18387 1461
rect 18406 1326 18440 1495
rect 18454 1442 18488 1892
rect 18580 1840 18596 1852
rect 18580 1830 18600 1840
rect 18580 1824 18596 1830
rect 18564 1809 18566 1818
rect 18574 1809 18598 1824
rect 18612 1818 18636 1852
rect 18734 1826 18840 1990
rect 18916 1964 18928 1998
rect 18916 1958 18974 1964
rect 18736 1825 18756 1826
rect 18548 1790 18614 1809
rect 18552 1784 18610 1790
rect 18568 1771 18602 1775
rect 18614 1771 18638 1774
rect 18656 1771 18676 1775
rect 18556 1759 18614 1771
rect 18650 1759 18676 1771
rect 18556 1756 18611 1759
rect 18520 1743 18522 1747
rect 18534 1743 18554 1747
rect 18508 1563 18560 1743
rect 18562 1591 18602 1756
rect 18568 1587 18602 1591
rect 18608 1743 18642 1747
rect 18608 1591 18648 1743
rect 18650 1603 18680 1759
rect 18650 1591 18676 1603
rect 18608 1578 18654 1591
rect 18656 1587 18676 1591
rect 18688 1587 18690 1775
rect 18697 1591 18702 1771
rect 18722 1621 18756 1825
rect 18770 1793 18840 1826
rect 18770 1759 18858 1793
rect 18770 1621 18857 1759
rect 18969 1691 19027 1697
rect 18969 1657 18981 1691
rect 18969 1651 19027 1657
rect 18722 1591 18857 1621
rect 18508 1553 18554 1563
rect 18508 1442 18542 1553
rect 18578 1544 18654 1578
rect 18722 1553 18724 1591
rect 18736 1585 18857 1591
rect 18937 1585 18971 1623
rect 18736 1551 18840 1585
rect 18871 1551 18891 1585
rect 18925 1551 19071 1585
rect 18596 1510 18676 1544
rect 18596 1494 18654 1510
rect 18639 1479 18654 1494
rect 18736 1476 18857 1551
rect 18937 1525 18971 1551
rect 19294 1498 19440 1532
rect 18949 1483 18965 1491
rect 18608 1442 18642 1476
rect 18454 1408 18494 1442
rect 18508 1408 18654 1442
rect 18722 1408 18857 1476
rect 18943 1449 18967 1483
rect 18981 1457 19005 1491
rect 18885 1411 18923 1423
rect 18739 1389 18857 1408
rect 18877 1399 18923 1411
rect 18877 1389 18911 1399
rect 18977 1389 19011 1423
rect 18739 1372 18863 1389
rect 18564 1342 18598 1360
rect 18552 1336 18610 1342
rect 18552 1326 18564 1336
rect 18406 1292 18441 1326
rect 18537 1315 18625 1326
rect 18548 1303 18614 1315
rect 18537 1292 18625 1303
rect 18406 1234 18440 1292
rect 18406 1200 18441 1234
rect 18537 1223 18625 1234
rect 18548 1211 18614 1223
rect 18537 1200 18625 1211
rect 18406 653 18440 1200
rect 18552 1190 18564 1200
rect 18552 1184 18610 1190
rect 18739 1181 18809 1372
rect 18823 1355 18863 1372
rect 18877 1355 19023 1389
rect 19246 1302 19392 1336
rect 18921 1283 18979 1289
rect 18921 1249 18933 1283
rect 19477 1266 19578 1623
rect 18921 1243 18979 1249
rect 18739 1147 18810 1181
rect 18739 1111 18792 1147
rect 19477 1058 19530 1266
rect 18722 1021 18756 1039
rect 18722 985 18792 1021
rect 18739 951 18810 985
rect 18552 736 18610 742
rect 18552 702 18564 736
rect 18552 696 18610 702
rect 17171 633 17229 639
rect 17341 614 17411 650
rect 18406 619 18421 653
rect 17358 580 17429 614
rect 18739 600 18809 951
rect 18921 883 18979 889
rect 18921 849 18933 883
rect 18921 843 18979 849
rect 18921 683 18979 689
rect 18921 649 18933 683
rect 18921 643 18979 649
rect 17171 365 17229 371
rect 17171 331 17183 365
rect 17171 325 17229 331
rect 17025 248 17040 282
rect 17358 229 17428 580
rect 18739 564 18792 600
rect 17540 512 17598 518
rect 17540 478 17552 512
rect 17540 472 17598 478
rect 19477 458 19530 968
rect 19846 952 19899 1462
rect 19846 405 19899 862
rect 17540 312 17598 318
rect 17540 278 17552 312
rect 17540 272 17598 278
rect 13394 193 13447 229
rect 17358 193 17411 229
rect 9211 4 9245 8
rect 9299 4 9333 8
rect 9211 -8 9245 -4
rect 9299 -8 9333 -4
rect 9211 -20 9251 -8
rect 9289 -20 9339 -8
rect 9413 -20 9501 20
rect 9562 -20 9720 20
rect 9211 -23 9245 -20
rect 9289 -23 9336 -20
rect 9211 -30 9257 -23
rect 9217 -39 9257 -30
rect 9287 -39 9336 -23
rect 9217 -73 9336 -39
rect 9217 -89 9257 -73
rect 9287 -89 9327 -73
rect 9217 -111 9245 -89
rect 9299 -111 9327 -89
rect 9097 -175 9132 -141
rect 9199 -175 9345 -141
rect 9097 -229 9131 -175
rect 9199 -188 9245 -175
rect 9211 -192 9245 -188
rect 9299 -188 9345 -175
rect 9413 -176 9500 -20
rect 9580 -176 9614 -156
rect 9668 -176 9702 -156
rect 9299 -192 9333 -188
rect 9413 -210 9501 -176
rect 9568 -210 9714 -176
rect 9097 -263 9132 -229
rect 9228 -240 9316 -229
rect 9239 -252 9305 -240
rect 9228 -263 9316 -252
rect 9097 -337 9131 -263
rect 9243 -269 9255 -263
rect 9243 -273 9301 -269
rect 9239 -285 9305 -273
rect 9413 -275 9500 -210
rect 9580 -240 9614 -210
rect 9668 -240 9702 -210
rect 9580 -250 9702 -240
rect 9580 -254 9614 -250
rect 9668 -254 9702 -250
rect 9255 -325 9289 -303
rect 9243 -331 9301 -325
rect 9243 -337 9255 -331
rect 9097 -371 9132 -337
rect 9228 -348 9316 -337
rect 9239 -358 9305 -348
rect 9145 -371 9399 -358
rect 9097 -702 9131 -371
rect 9430 -390 9500 -275
rect 9612 -278 9648 -272
rect 9608 -288 9674 -278
rect 9624 -312 9658 -288
rect 9608 -322 9674 -312
rect 9612 -328 9648 -322
rect 9580 -350 9614 -346
rect 9668 -350 9702 -346
rect 9580 -353 9626 -350
rect 9656 -353 9702 -350
rect 9580 -356 9620 -353
rect 9580 -390 9614 -356
rect 9668 -390 9702 -353
rect 9430 -424 9501 -390
rect 9562 -424 9714 -390
rect 9720 -424 9736 -390
rect 9430 -580 9500 -424
rect 9782 -518 9816 -82
rect 9430 -614 9501 -580
rect 9243 -639 9301 -633
rect 9243 -673 9255 -639
rect 9430 -650 9483 -614
rect 9243 -679 9301 -673
rect 8359 -773 8394 -739
rect 8692 -755 9368 -702
rect 8692 -811 9483 -755
rect 7701 -842 7891 -833
rect 7763 -856 7829 -842
rect 7840 -856 7853 -842
rect 7752 -867 7853 -856
rect 7954 -862 8007 -826
rect 8692 -864 9114 -811
rect 7767 -877 7779 -867
rect 7812 -877 7825 -867
rect 7348 -932 7548 -888
rect 7582 -932 7686 -888
rect 7763 -901 7829 -877
rect 7840 -898 7853 -867
rect 7779 -929 7813 -919
rect 7414 -944 7448 -932
rect 7502 -944 7536 -932
rect 7414 -952 7536 -944
rect 7402 -966 7536 -952
rect 7543 -966 7548 -932
rect 7568 -962 7686 -932
rect 7767 -935 7825 -929
rect 7767 -953 7779 -935
rect 7937 -953 7971 -940
rect 7752 -962 7840 -953
rect 7936 -958 7971 -953
rect 7568 -966 7923 -962
rect 7414 -970 7448 -966
rect 7502 -970 7536 -966
rect 7418 -984 7422 -970
rect 7446 -982 7504 -976
rect 7442 -984 7508 -982
rect 7568 -984 7570 -966
rect 7422 -990 7508 -984
rect 7394 -1004 7508 -990
rect 7582 -987 7923 -966
rect 7936 -987 8007 -958
rect 7420 -1024 7444 -1004
rect 7458 -1024 7492 -1004
rect 7362 -1062 7400 -1050
rect 7354 -1074 7400 -1062
rect 7418 -1072 7422 -1030
rect 7442 -1038 7508 -1024
rect 7446 -1044 7504 -1038
rect 7582 -1050 7686 -987
rect 7937 -994 8007 -987
rect 7735 -1021 7769 -1012
rect 7823 -1021 7857 -1012
rect 7454 -1062 7488 -1050
rect 7442 -1069 7500 -1062
rect 7354 -1084 7388 -1074
rect 7420 -1084 7422 -1072
rect 7448 -1072 7494 -1069
rect 7448 -1084 7450 -1072
rect 7454 -1084 7488 -1072
rect 7300 -1140 7340 -1084
rect 7354 -1140 7554 -1084
rect 7568 -1140 7686 -1050
rect 6676 -1175 6710 -1171
rect 6722 -1174 6746 -1171
rect 6764 -1175 6798 -1171
rect 6660 -1186 6718 -1184
rect 6830 -1185 6971 -1159
rect 7014 -1170 7102 -1159
rect 7025 -1185 7091 -1170
rect 7199 -1177 7219 -1159
rect 6830 -1186 7199 -1185
rect 6610 -1220 6630 -1186
rect 6642 -1193 7199 -1186
rect 6642 -1209 6948 -1193
rect 6645 -1220 6781 -1209
rect 6672 -1230 6706 -1220
rect 6720 -1230 6744 -1220
rect 6720 -1239 6754 -1230
rect 6704 -1252 6770 -1239
rect 6708 -1258 6766 -1252
rect 6628 -1277 6662 -1258
rect 6716 -1277 6750 -1258
rect 6616 -1292 6662 -1277
rect 6704 -1283 6762 -1277
rect 6710 -1286 6756 -1283
rect 6716 -1292 6750 -1286
rect 6509 -1349 6549 -1292
rect 6610 -1315 6784 -1292
rect 6605 -1320 6784 -1315
rect 6605 -1349 6816 -1320
rect 6509 -1373 6548 -1349
rect 6562 -1354 6602 -1349
rect 6616 -1354 6816 -1349
rect 6514 -1407 6548 -1373
rect 5723 -1495 5841 -1478
rect 4396 -1502 4578 -1498
rect 4504 -1508 4580 -1502
rect 4442 -1510 4580 -1508
rect 4616 -1508 5656 -1495
rect 4616 -1510 5632 -1508
rect 4442 -1530 4524 -1510
rect 4616 -1521 4751 -1510
rect 4999 -1513 5019 -1510
rect 4985 -1521 5019 -1513
rect 4442 -1536 4552 -1530
rect 4468 -1542 4492 -1536
rect 4504 -1538 4552 -1536
rect 4506 -1570 4530 -1538
rect 4616 -1548 4734 -1521
rect 4630 -1555 4734 -1548
rect 4751 -1555 5019 -1521
rect 5033 -1527 5072 -1510
rect 5086 -1514 5120 -1510
rect 5354 -1512 5388 -1510
rect 5368 -1514 5388 -1512
rect 5402 -1514 5441 -1510
rect 5086 -1520 5126 -1514
rect 5146 -1520 5340 -1514
rect 5086 -1527 5349 -1520
rect 5553 -1525 5611 -1519
rect 5033 -1555 5349 -1527
rect 5407 -1548 5441 -1536
rect 4630 -1567 4751 -1555
rect 5033 -1567 5053 -1555
rect 5072 -1561 5349 -1555
rect 4630 -1589 5053 -1567
rect 4630 -1591 4752 -1589
rect 3230 -1616 3275 -1612
rect 3343 -1616 3489 -1612
rect 3180 -1632 3276 -1616
rect 2904 -1656 2916 -1632
rect 2928 -1656 2948 -1632
rect 2904 -1666 2948 -1656
rect 3170 -1646 3276 -1632
rect 3330 -1636 3508 -1616
rect 3330 -1646 3376 -1636
rect 3389 -1646 3508 -1636
rect 3170 -1648 3214 -1646
rect 3170 -1656 3182 -1648
rect 3194 -1656 3214 -1648
rect 3170 -1666 3214 -1656
rect 2922 -1676 2948 -1666
rect 3188 -1676 3214 -1666
rect 3230 -1666 3275 -1646
rect 3343 -1648 3376 -1646
rect 3400 -1648 3489 -1646
rect 3376 -1657 3444 -1648
rect 3364 -1661 3444 -1657
rect 3462 -1661 3472 -1648
rect 3364 -1666 3474 -1661
rect 2922 -1682 2938 -1676
rect 3188 -1682 3204 -1676
rect 2440 -1694 2878 -1693
rect 3205 -1694 3212 -1676
rect 3230 -1693 3231 -1666
rect 3241 -1682 3275 -1666
rect 3349 -1682 3483 -1666
rect 3241 -1693 3444 -1682
rect 3230 -1694 3444 -1693
rect 1717 -1727 2120 -1694
rect 2204 -1714 2318 -1710
rect 2421 -1722 2436 -1694
rect 2455 -1695 2489 -1694
rect 2771 -1695 2805 -1694
rect 2455 -1722 2805 -1695
rect 3241 -1695 3387 -1694
rect 3445 -1695 3458 -1682
rect 3462 -1693 3471 -1682
rect 3549 -1693 4340 -1612
rect 4396 -1638 4554 -1610
rect 4630 -1638 4650 -1591
rect 4664 -1601 4752 -1591
rect 5072 -1595 5349 -1574
rect 4664 -1637 4734 -1601
rect 5141 -1608 5275 -1595
rect 5368 -1608 5388 -1548
rect 5402 -1608 5441 -1548
rect 5549 -1559 5615 -1525
rect 5735 -1531 5841 -1495
rect 5891 -1501 5924 -1485
rect 5963 -1501 6010 -1478
rect 5891 -1519 6010 -1501
rect 6092 -1517 6126 -1478
rect 5898 -1531 6010 -1519
rect 5735 -1536 5810 -1531
rect 5553 -1565 5611 -1559
rect 5723 -1565 5810 -1536
rect 5886 -1544 5963 -1531
rect 5966 -1544 6016 -1531
rect 5886 -1557 6016 -1544
rect 5548 -1576 5606 -1570
rect 4664 -1638 4698 -1637
rect 4396 -1644 4602 -1638
rect 5175 -1642 5241 -1629
rect 4348 -1672 4383 -1644
rect 4444 -1672 4602 -1644
rect 3462 -1694 4340 -1693
rect 3241 -1698 3458 -1695
rect 3241 -1710 3275 -1698
rect 3383 -1710 3449 -1698
rect 3549 -1701 4340 -1694
rect 3230 -1722 3486 -1710
rect 3557 -1722 3596 -1701
rect 3610 -1722 3644 -1701
rect 3918 -1710 4340 -1701
rect 3848 -1714 4340 -1710
rect 2050 -1748 2103 -1727
rect 2421 -1748 2841 -1722
rect 3205 -1744 3644 -1722
rect 3706 -1726 4340 -1714
rect 3205 -1748 3645 -1744
rect 3706 -1748 3874 -1726
rect 1748 -1761 1804 -1748
rect 1838 -1761 2540 -1748
rect 2050 -1763 2540 -1761
rect 2574 -1763 2744 -1748
rect 2778 -1763 2839 -1748
rect 2086 -1781 2436 -1763
rect 2841 -1765 2867 -1748
rect 2472 -1781 2498 -1765
rect 2050 -1782 2498 -1781
rect 3205 -1781 3591 -1748
rect 3610 -1778 3888 -1748
rect 3918 -1754 4340 -1726
rect 3945 -1759 3960 -1754
rect 3888 -1781 3914 -1778
rect 3205 -1782 3914 -1781
rect 3205 -1797 3549 -1782
rect 3205 -1804 3557 -1797
rect 3205 -1831 3591 -1804
rect 3205 -1832 3549 -1831
rect 3205 -1858 3627 -1832
rect 5050 -1856 5141 -1848
rect 5187 -1856 5229 -1848
rect 3205 -1865 3625 -1858
rect 3205 -1867 3549 -1865
rect 3627 -1867 3653 -1858
rect 5222 -1876 5229 -1856
rect 5050 -1884 5141 -1876
rect 5187 -1884 5229 -1876
rect 1086 -1976 1088 -1948
rect 1846 -1974 1850 -1946
rect 1902 -1964 1918 -1958
rect 1874 -1974 1928 -1964
rect 1124 -2012 1126 -1976
rect 1868 -1984 1934 -1974
rect 1868 -1990 1894 -1984
rect 1884 -2008 1894 -1990
rect 1908 -1990 1934 -1984
rect 1908 -2008 1928 -1990
rect 1944 -2008 1956 -1946
rect 2076 -1974 2090 -1946
rect 2132 -1964 2148 -1958
rect 2104 -1974 2158 -1964
rect 2342 -1974 2354 -1946
rect 2398 -1964 2414 -1958
rect 2370 -1974 2424 -1964
rect 2098 -1984 2164 -1974
rect 2098 -1990 2128 -1984
rect 2114 -2008 2128 -1990
rect 2138 -1990 2164 -1984
rect 2364 -1984 2430 -1974
rect 2364 -1990 2392 -1984
rect 2138 -2008 2158 -1990
rect 2380 -2008 2392 -1990
rect 2404 -1990 2430 -1984
rect 2404 -2008 2424 -1990
rect 2440 -2008 2452 -1946
rect 2866 -1974 2878 -1946
rect 2922 -1964 2938 -1958
rect 2894 -1974 2948 -1964
rect 2744 -2008 2878 -1977
rect 2888 -1984 2954 -1974
rect 3112 -1977 3144 -1946
rect 3188 -1964 3204 -1958
rect 3160 -1974 3214 -1964
rect 2888 -1990 2916 -1984
rect 2904 -2008 2916 -1990
rect 2928 -1990 2954 -1984
rect 2928 -2008 2948 -1990
rect 2743 -2020 2878 -2008
rect 112 -2056 236 -2048
rect 112 -2084 236 -2076
rect 1304 -2128 1412 -2122
rect 816 -2194 820 -2160
rect 1374 -2194 1376 -2160
rect 1640 -2162 1650 -2055
rect 1668 -2162 1678 -2027
rect 2732 -2036 2878 -2020
rect 2998 -2036 3144 -1977
rect 3154 -1984 3220 -1974
rect 3154 -1990 3182 -1984
rect 3194 -1990 3220 -1984
rect 3170 -1994 3214 -1990
rect 3230 -1992 3376 -1946
rect 3418 -1964 3434 -1958
rect 3390 -1974 3444 -1964
rect 3384 -1984 3450 -1974
rect 3384 -1990 3414 -1984
rect 3400 -1992 3414 -1990
rect 3424 -1990 3450 -1984
rect 3424 -1992 3444 -1990
rect 3230 -1994 3242 -1992
rect 3376 -1994 3444 -1992
rect 3462 -1992 3549 -1946
rect 3598 -1974 3608 -1946
rect 3654 -1964 3670 -1958
rect 3626 -1974 3680 -1964
rect 3620 -1975 3686 -1974
rect 3694 -1975 3708 -1946
rect 3954 -1956 3989 -1922
rect 3585 -1992 3608 -1975
rect 3620 -1990 3935 -1975
rect 3462 -1994 3472 -1992
rect 3170 -2008 3276 -1994
rect 3180 -2024 3276 -2008
rect 3330 -2024 3508 -1994
rect 3549 -2009 3608 -1992
rect 3636 -1998 3935 -1990
rect 3625 -2008 3935 -1998
rect 3625 -2009 3681 -2008
rect 3694 -2009 3935 -2008
rect 3180 -2036 3212 -2024
rect 3230 -2028 3231 -2024
rect 3376 -2028 3444 -2024
rect 3462 -2028 3463 -2024
rect 3549 -2028 3619 -2009
rect 3636 -2024 3653 -2009
rect 2732 -2048 2748 -2042
rect 2714 -2058 2758 -2048
rect 3216 -2058 3619 -2028
rect 3901 -2036 3935 -2009
rect 2714 -2068 2764 -2058
rect 2738 -2074 2764 -2068
rect 2738 -2082 2758 -2074
rect 2904 -2081 2914 -2058
rect 2928 -2081 2948 -2058
rect 2714 -2092 2758 -2082
rect 2732 -2102 2758 -2092
rect 2847 -2098 2882 -2081
rect 2732 -2108 2748 -2102
rect 2811 -2115 2882 -2098
rect 2904 -2092 2976 -2081
rect 3045 -2092 3097 -2081
rect 3159 -2088 3197 -2081
rect 3132 -2092 3197 -2088
rect 2904 -2104 2938 -2092
rect 3056 -2104 3086 -2092
rect 2893 -2115 2949 -2104
rect 3045 -2115 3097 -2104
rect 3120 -2115 3197 -2092
rect 2778 -2126 2790 -2116
rect 2811 -2126 2881 -2115
rect 2114 -2153 2124 -2126
rect 2138 -2153 2158 -2126
rect 2772 -2134 2800 -2126
rect 2810 -2134 2881 -2126
rect 2478 -2145 2539 -2134
rect 2575 -2145 2627 -2134
rect 2772 -2142 2881 -2134
rect 2478 -2147 2528 -2145
rect 2478 -2153 2574 -2147
rect 2098 -2160 2574 -2153
rect 2586 -2157 2616 -2145
rect 2788 -2157 2881 -2142
rect 2575 -2160 2627 -2157
rect 2779 -2160 2881 -2157
rect 1884 -2196 1894 -2162
rect 1908 -2196 1928 -2162
rect 2478 -2168 2881 -2160
rect 2109 -2194 2459 -2187
rect 2109 -2198 2159 -2194
rect 2255 -2198 2307 -2194
rect 2369 -2198 2425 -2194
rect 2109 -2206 2148 -2198
rect 2266 -2206 2296 -2198
rect 2380 -2206 2414 -2198
rect 2444 -2206 2459 -2194
rect 2478 -2194 2512 -2168
rect 2528 -2184 2530 -2178
rect 2528 -2194 2540 -2184
rect 2586 -2194 2616 -2178
rect 2794 -2194 2881 -2168
rect 2478 -2202 2881 -2194
rect 2478 -2206 2546 -2202
rect 2586 -2206 2720 -2202
rect 2794 -2206 2881 -2202
rect 1042 -2264 1044 -2230
rect 1704 -2257 2881 -2206
rect 2993 -2183 3051 -2177
rect 2993 -2217 3005 -2183
rect 3056 -2206 3086 -2125
rect 3163 -2126 3197 -2115
rect 3216 -2088 3231 -2058
rect 3277 -2062 3329 -2058
rect 3389 -2062 3445 -2058
rect 3509 -2062 3619 -2058
rect 3154 -2149 3163 -2126
rect 3170 -2160 3214 -2126
rect 3216 -2160 3242 -2088
rect 3316 -2090 3318 -2072
rect 3258 -2098 3458 -2090
rect 3316 -2114 3318 -2098
rect 3358 -2118 3360 -2114
rect 3258 -2126 3458 -2118
rect 3358 -2160 3360 -2126
rect 2993 -2223 3051 -2217
rect 2927 -2228 3117 -2226
rect 1337 -2264 1586 -2259
rect -88 -2298 0 -2290
rect 1371 -2298 1586 -2293
rect -88 -2326 0 -2318
rect 932 -2336 936 -2302
rect 1371 -2304 1383 -2298
rect 1467 -2304 1585 -2298
rect 1371 -2310 1372 -2304
rect 1335 -2312 1388 -2310
rect 1234 -2336 1388 -2312
rect 1478 -2316 1574 -2304
rect 1668 -2314 2881 -2257
rect 2961 -2262 2995 -2260
rect 3049 -2262 3083 -2260
rect 3170 -2261 3197 -2160
rect 3216 -2261 3231 -2160
rect 3358 -2164 3424 -2160
rect 3358 -2180 3360 -2164
rect 3324 -2198 3458 -2194
rect 3532 -2206 3619 -2062
rect 3727 -2111 3793 -2092
rect 3665 -2125 3855 -2121
rect 3665 -2206 3670 -2125
rect 3693 -2145 3821 -2126
rect 3752 -2149 3755 -2145
rect 3776 -2149 3796 -2145
rect 3693 -2153 3739 -2149
rect 3752 -2153 3833 -2149
rect 3693 -2190 3698 -2153
rect 3752 -2156 3824 -2153
rect 3825 -2156 3833 -2153
rect 3901 -2155 3919 -2147
rect 3920 -2155 3935 -2036
rect 3954 -2155 3988 -1956
rect 4072 -2070 4076 -1990
rect 4100 -2024 4158 -2018
rect 4100 -2058 4112 -2024
rect 5033 -2055 5073 -2031
rect 5129 -2032 5287 -2021
rect 5368 -2032 5383 -1608
rect 5402 -1661 5437 -1608
rect 5544 -1610 5610 -1576
rect 5548 -1616 5606 -1610
rect 5632 -1627 5634 -1600
rect 5510 -1644 5644 -1627
rect 5562 -1648 5592 -1644
rect 5504 -1661 5650 -1648
rect 5735 -1661 5810 -1565
rect 5889 -1578 5898 -1557
rect 5917 -1563 5975 -1557
rect 5922 -1578 5980 -1572
rect 5881 -1591 6011 -1578
rect 5881 -1604 5931 -1591
rect 5903 -1616 5931 -1604
rect 5934 -1604 6011 -1591
rect 5934 -1612 6015 -1604
rect 5896 -1628 5931 -1616
rect 5961 -1616 5999 -1612
rect 5961 -1628 6006 -1616
rect 5896 -1650 5919 -1628
rect 5973 -1650 6006 -1628
rect 5402 -1968 5436 -1661
rect 5735 -1714 5806 -1661
rect 5873 -1714 6019 -1680
rect 6087 -1714 6126 -1517
rect 6140 -1714 6179 -1478
rect 6259 -1504 6381 -1470
rect 6259 -1520 6305 -1504
rect 6335 -1520 6381 -1504
rect 6259 -1547 6293 -1520
rect 6254 -1572 6293 -1547
rect 6300 -1551 6305 -1520
rect 6347 -1547 6381 -1520
rect 6300 -1572 6304 -1551
rect 6331 -1563 6335 -1552
rect 6342 -1572 6381 -1547
rect 6254 -1615 6288 -1572
rect 6342 -1584 6376 -1572
rect 6330 -1615 6335 -1584
rect 6337 -1615 6384 -1584
rect 6254 -1679 6300 -1615
rect 6330 -1631 6384 -1615
rect 6303 -1665 6384 -1631
rect 5548 -1866 5606 -1860
rect 5548 -1900 5560 -1866
rect 5548 -1906 5606 -1900
rect 5735 -1926 5805 -1714
rect 5889 -1899 5898 -1800
rect 5917 -1831 5975 -1825
rect 5917 -1865 5929 -1831
rect 5917 -1871 5975 -1865
rect 6087 -1871 6121 -1714
rect 6106 -1926 6121 -1871
rect 6140 -1767 6175 -1714
rect 6242 -1731 6300 -1679
rect 6330 -1679 6376 -1665
rect 6330 -1731 6388 -1679
rect 6242 -1756 6388 -1733
rect 6248 -1767 6382 -1756
rect 6456 -1767 6495 -1464
rect 6509 -1767 6548 -1407
rect 6628 -1401 6662 -1354
rect 6716 -1370 6750 -1354
rect 6628 -1417 6674 -1401
rect 6701 -1417 6750 -1370
rect 6830 -1390 6948 -1209
rect 6979 -1262 7137 -1239
rect 6974 -1273 7137 -1262
rect 7218 -1273 7233 -1193
rect 7252 -1273 7286 -1159
rect 7585 -1176 7686 -1140
rect 7954 -1028 8025 -994
rect 8305 -1028 8340 -994
rect 8728 -1011 8763 -993
rect 7398 -1190 7456 -1184
rect 7398 -1224 7410 -1190
rect 7398 -1230 7456 -1224
rect 6974 -1296 7132 -1273
rect 7218 -1358 7228 -1273
rect 7252 -1326 7282 -1273
rect 7585 -1326 7655 -1176
rect 7767 -1243 7825 -1237
rect 7767 -1277 7779 -1243
rect 7812 -1277 7825 -1243
rect 7767 -1283 7825 -1277
rect 7840 -1298 7853 -1209
rect 7024 -1364 7082 -1358
rect 7024 -1388 7036 -1364
rect 6830 -1411 6912 -1390
rect 7024 -1398 7038 -1388
rect 7068 -1398 7070 -1388
rect 7024 -1404 7082 -1398
rect 6628 -1451 6750 -1417
rect 6628 -1467 6674 -1451
rect 6704 -1467 6750 -1451
rect 6628 -1510 6662 -1467
rect 6623 -1625 6662 -1510
rect 6669 -1498 6674 -1467
rect 6669 -1625 6673 -1498
rect 6700 -1510 6704 -1499
rect 6716 -1510 6750 -1467
rect 6711 -1625 6750 -1510
rect 6825 -1435 6912 -1411
rect 7194 -1435 7228 -1358
rect 7585 -1362 7638 -1326
rect 7954 -1398 8024 -1028
rect 8306 -1047 8340 -1028
rect 8692 -1026 8763 -1011
rect 9043 -1026 9078 -992
rect 8136 -1096 8194 -1090
rect 8136 -1130 8148 -1096
rect 8136 -1136 8194 -1130
rect 8158 -1286 8164 -1256
rect 8186 -1258 8192 -1228
rect 7954 -1432 8025 -1398
rect 8325 -1432 8340 -1047
rect 8359 -1081 8394 -1047
rect 8359 -1432 8393 -1081
rect 8505 -1149 8563 -1143
rect 8505 -1183 8517 -1149
rect 8505 -1189 8563 -1183
rect 8505 -1349 8563 -1343
rect 8505 -1383 8517 -1349
rect 8505 -1389 8563 -1383
rect 6825 -1469 6918 -1435
rect 7027 -1436 7079 -1435
rect 6980 -1469 7126 -1436
rect 6623 -1637 6657 -1625
rect 6711 -1637 6745 -1625
rect 6623 -1678 6753 -1637
rect 6825 -1666 6917 -1469
rect 6992 -1499 7026 -1469
rect 7080 -1499 7114 -1469
rect 6992 -1514 7114 -1499
rect 6992 -1526 7115 -1514
rect 6988 -1531 7038 -1526
rect 7068 -1531 7118 -1526
rect 6988 -1564 7118 -1531
rect 6988 -1571 7123 -1564
rect 6993 -1604 7123 -1571
rect 7194 -1604 7233 -1435
rect 7621 -1452 7656 -1434
rect 7585 -1467 7656 -1452
rect 6993 -1609 7043 -1604
rect 6996 -1614 7043 -1609
rect 7073 -1609 7123 -1604
rect 7073 -1614 7119 -1609
rect 6996 -1621 7037 -1614
rect 6997 -1632 7037 -1621
rect 7079 -1632 7119 -1614
rect 6997 -1666 7031 -1632
rect 7085 -1666 7119 -1632
rect 6619 -1684 6669 -1678
rect 6711 -1682 6745 -1678
rect 6619 -1718 6722 -1684
rect 6825 -1700 6918 -1666
rect 6985 -1699 7131 -1666
rect 7132 -1687 7153 -1666
rect 6994 -1700 7122 -1699
rect 6651 -1759 6717 -1725
rect 6825 -1765 6917 -1700
rect 6847 -1767 6917 -1765
rect 7029 -1737 7087 -1731
rect 7029 -1767 7041 -1737
rect 6140 -1873 6174 -1767
rect 6286 -1778 6344 -1772
rect 6282 -1801 6348 -1778
rect 6286 -1812 6298 -1801
rect 6286 -1818 6344 -1812
rect 6456 -1818 6490 -1767
rect 6475 -1873 6490 -1818
rect 6509 -1819 6544 -1767
rect 6847 -1785 6918 -1767
rect 7014 -1778 7102 -1767
rect 7199 -1777 7233 -1604
rect 7025 -1785 7091 -1778
rect 6509 -1861 6549 -1819
rect 6610 -1827 6768 -1786
rect 6605 -1854 6768 -1827
rect 6847 -1801 7199 -1785
rect 6847 -1839 6917 -1801
rect 7007 -1839 7109 -1835
rect 6605 -1861 6763 -1854
rect 6140 -1914 6180 -1873
rect 6241 -1880 6399 -1873
rect 6236 -1907 6399 -1880
rect 6475 -1895 6495 -1873
rect 6236 -1914 6394 -1907
rect 5735 -1967 5811 -1926
rect 5872 -1933 6030 -1926
rect 5867 -1960 6030 -1933
rect 6106 -1948 6126 -1926
rect 5867 -1967 6025 -1960
rect 5402 -1978 5437 -1968
rect 5402 -2002 5442 -1978
rect 5498 -1979 5656 -1968
rect 5498 -2002 5661 -1979
rect 5407 -2013 5442 -2002
rect 5503 -2013 5661 -2002
rect 5735 -2003 5810 -1967
rect 5129 -2055 5292 -2032
rect 5368 -2036 5388 -2032
rect 4100 -2064 4158 -2058
rect 5038 -2066 5073 -2055
rect 5134 -2066 5292 -2055
rect 4072 -2080 4090 -2070
rect 4076 -2096 4090 -2080
rect 4669 -2102 4704 -2085
rect 4999 -2089 5019 -2085
rect 4056 -2155 4114 -2137
rect 4144 -2155 4202 -2137
rect 4264 -2155 4340 -2102
rect 3752 -2160 3833 -2156
rect 3752 -2165 3768 -2160
rect 3770 -2164 3833 -2160
rect 3770 -2165 3786 -2164
rect 3687 -2206 3698 -2190
rect 3775 -2206 3782 -2165
rect 3800 -2184 3833 -2164
rect 3870 -2184 3872 -2178
rect 3800 -2192 3840 -2184
rect 3870 -2192 3882 -2184
rect 3800 -2194 3882 -2192
rect 3822 -2206 3888 -2194
rect 3895 -2206 4340 -2155
rect 3318 -2239 3333 -2211
rect 3406 -2226 3449 -2211
rect 3248 -2261 3250 -2248
rect 3318 -2261 3367 -2239
rect 3406 -2261 3434 -2226
rect 3532 -2261 4340 -2206
rect 4633 -2119 4704 -2102
rect 2949 -2314 2953 -2264
rect 2965 -2279 3007 -2264
rect 2980 -2314 3007 -2279
rect 3088 -2286 3095 -2264
rect 3056 -2314 3095 -2286
rect 3157 -2314 4340 -2261
rect 4446 -2240 4504 -2234
rect 4446 -2274 4458 -2240
rect 4446 -2280 4504 -2274
rect 1467 -2327 1585 -2316
rect 1335 -2346 1388 -2336
rect 1002 -2352 1388 -2346
rect 1478 -2352 1544 -2337
rect 1668 -2352 4340 -2314
rect 1002 -2357 4340 -2352
rect 1002 -2388 1030 -2357
rect 1036 -2380 4340 -2357
rect 1318 -2388 4340 -2380
rect 214 -2448 236 -2395
rect 112 -2456 130 -2448
rect 176 -2456 236 -2448
rect 242 -2452 264 -2423
rect 448 -2452 482 -2419
rect 633 -2433 800 -2399
rect 854 -2433 983 -2399
rect 536 -2452 552 -2435
rect 102 -2476 112 -2456
rect 130 -2476 140 -2456
rect 112 -2484 130 -2476
rect 176 -2484 236 -2476
rect 214 -2505 236 -2484
rect 242 -2486 382 -2452
rect 436 -2486 582 -2452
rect 599 -2486 614 -2452
rect 242 -2505 298 -2486
rect 36 -2539 182 -2505
rect 214 -2539 298 -2505
rect 36 -2603 134 -2560
rect 44 -2624 94 -2603
rect 136 -2607 137 -2591
rect 211 -2603 298 -2539
rect 375 -2554 382 -2507
rect 448 -2523 495 -2507
rect 312 -2603 382 -2581
rect 422 -2588 429 -2554
rect 436 -2581 495 -2523
rect 546 -2581 570 -2486
rect 436 -2603 570 -2581
rect 102 -2624 103 -2607
rect 44 -2641 103 -2624
rect 48 -2658 77 -2650
rect 211 -2658 245 -2603
rect 248 -2658 298 -2603
rect 344 -2607 370 -2603
rect 494 -2604 514 -2603
rect 494 -2624 496 -2604
rect 546 -2607 570 -2603
rect 378 -2658 412 -2624
rect 466 -2635 500 -2624
rect 466 -2644 512 -2635
rect 466 -2658 500 -2644
rect 580 -2658 614 -2486
rect 633 -2568 668 -2433
rect 854 -2467 872 -2454
rect 785 -2485 800 -2470
rect 775 -2495 800 -2485
rect 775 -2501 837 -2495
rect 775 -2528 800 -2501
rect 742 -2535 800 -2528
rect 832 -2535 841 -2501
rect 854 -2528 875 -2467
rect 949 -2490 983 -2433
rect 1002 -2405 1088 -2388
rect 1196 -2405 1254 -2388
rect 1284 -2396 4340 -2388
rect 1284 -2405 3971 -2396
rect 742 -2541 837 -2535
rect 742 -2568 800 -2541
rect 854 -2568 935 -2528
rect 633 -2658 667 -2568
rect 735 -2597 757 -2582
rect 835 -2590 869 -2578
rect 735 -2609 750 -2597
rect 819 -2624 835 -2607
rect 747 -2641 781 -2624
rect 819 -2641 869 -2624
rect 949 -2641 988 -2490
rect 1002 -2641 1036 -2405
rect 1196 -2442 1241 -2405
rect 1148 -2448 1241 -2442
rect 1148 -2456 1160 -2448
rect 1196 -2456 1241 -2448
rect 1042 -2475 1070 -2456
rect 1077 -2475 1088 -2459
rect 1042 -2529 1088 -2475
rect 1144 -2482 1241 -2456
rect 1318 -2449 3971 -2405
rect 1318 -2458 3596 -2449
rect 3608 -2458 3636 -2449
rect 3664 -2458 3670 -2449
rect 3676 -2458 3710 -2449
rect 3764 -2458 3798 -2449
rect 3878 -2458 3928 -2449
rect 1148 -2488 1210 -2482
rect 1196 -2490 1210 -2488
rect 1124 -2504 1158 -2490
rect 1112 -2529 1162 -2504
rect 1196 -2513 1242 -2490
rect 1196 -2529 1207 -2513
rect 1042 -2556 1070 -2529
rect 1104 -2554 1162 -2529
rect 1208 -2540 1242 -2513
rect 1318 -2491 3608 -2458
rect 3625 -2469 3928 -2458
rect 3636 -2481 3928 -2469
rect 3625 -2491 3928 -2481
rect 1318 -2492 3928 -2491
rect 1318 -2495 3596 -2492
rect 3664 -2495 3670 -2492
rect 3676 -2495 3710 -2492
rect 1318 -2534 3608 -2495
rect 1104 -2568 1142 -2554
rect 1188 -2588 1238 -2554
rect 1250 -2568 1254 -2534
rect 1284 -2542 3608 -2534
rect 3664 -2542 3717 -2495
rect 3730 -2531 3740 -2526
rect 3722 -2542 3740 -2531
rect 1284 -2546 3596 -2542
rect 3636 -2546 3740 -2542
rect 3764 -2542 3798 -2492
rect 3764 -2546 3828 -2542
rect 3878 -2546 3928 -2492
rect 1284 -2568 3608 -2546
rect 1239 -2588 1250 -2568
rect 1318 -2588 3608 -2568
rect 1126 -2604 3608 -2588
rect 3636 -2604 3928 -2546
rect 3931 -2482 3965 -2449
rect 3994 -2458 4033 -2432
rect 4045 -2458 4079 -2424
rect 4133 -2458 4167 -2424
rect 4266 -2432 4281 -2396
rect 4300 -2432 4334 -2396
rect 4179 -2458 4247 -2432
rect 4266 -2458 4402 -2432
rect 4414 -2458 4448 -2424
rect 4502 -2458 4536 -2424
rect 4548 -2458 4616 -2432
rect 4633 -2458 4703 -2119
rect 4815 -2187 4873 -2181
rect 4815 -2221 4827 -2187
rect 4815 -2227 4873 -2221
rect 5004 -2404 5019 -2089
rect 4827 -2421 4861 -2411
rect 4020 -2480 4179 -2458
rect 4247 -2480 4281 -2458
rect 4300 -2480 4334 -2458
rect 4380 -2480 4548 -2458
rect 4616 -2480 4936 -2458
rect 4020 -2482 4936 -2480
rect 3931 -2492 4936 -2482
rect 4951 -2489 4952 -2458
rect 4985 -2489 5019 -2404
rect 5038 -2436 5072 -2066
rect 5222 -2276 5234 -2268
rect 5038 -2470 5073 -2436
rect 5134 -2458 5292 -2436
rect 5373 -2451 5388 -2036
rect 5407 -2383 5441 -2013
rect 5553 -2081 5611 -2075
rect 5553 -2115 5565 -2081
rect 5604 -2115 5611 -2081
rect 5553 -2121 5611 -2115
rect 5632 -2149 5639 -2047
rect 5553 -2281 5611 -2275
rect 5553 -2315 5565 -2281
rect 5553 -2321 5611 -2315
rect 5407 -2404 5442 -2383
rect 5407 -2417 5645 -2404
rect 5740 -2417 5810 -2003
rect 5894 -2096 5898 -2000
rect 5922 -2028 5980 -2022
rect 5922 -2062 5934 -2028
rect 5922 -2068 5980 -2062
rect 5894 -2400 5898 -2302
rect 5922 -2336 5980 -2330
rect 5922 -2370 5934 -2336
rect 5922 -2376 5980 -2370
rect 5740 -2453 5793 -2417
rect 5004 -2492 5019 -2489
rect 5107 -2492 5567 -2458
rect 6111 -2472 6126 -1948
rect 3931 -2550 4033 -2492
rect 4066 -2524 4079 -2492
rect 4058 -2542 4088 -2524
rect 4045 -2550 4088 -2542
rect 4100 -2550 4113 -2492
rect 4132 -2494 4402 -2492
rect 4548 -2494 4704 -2492
rect 4765 -2494 4923 -2492
rect 4132 -2529 4430 -2494
rect 4546 -2496 4923 -2494
rect 4996 -2496 5019 -2492
rect 4546 -2522 5019 -2496
rect 4546 -2529 4630 -2522
rect 4132 -2548 4630 -2529
rect 4633 -2523 5019 -2522
rect 6145 -2503 6179 -1914
rect 6291 -1975 6349 -1969
rect 6291 -2009 6303 -1975
rect 6291 -2015 6349 -2009
rect 6291 -2463 6349 -2457
rect 6291 -2473 6303 -2463
rect 6276 -2484 6364 -2473
rect 6287 -2496 6353 -2484
rect 6145 -2507 6180 -2503
rect 6276 -2507 6364 -2496
rect 4633 -2548 4686 -2523
rect 5373 -2546 5384 -2545
rect 4133 -2550 4168 -2548
rect 3931 -2574 3950 -2550
rect 4000 -2576 4019 -2550
rect 4033 -2576 4168 -2550
rect 3931 -2604 3950 -2576
rect 1126 -2607 3840 -2604
rect 1116 -2608 3680 -2607
rect 3694 -2608 3708 -2607
rect 1116 -2620 3676 -2608
rect 3694 -2616 3704 -2608
rect 3722 -2616 3752 -2607
rect 3764 -2611 3774 -2607
rect 3782 -2616 3840 -2607
rect 3694 -2620 3840 -2616
rect 1116 -2622 3840 -2620
rect 747 -2658 1036 -2641
rect 1082 -2658 1107 -2641
rect 1116 -2658 1160 -2622
rect 1318 -2624 3840 -2622
rect 1204 -2658 1238 -2624
rect 1318 -2636 3676 -2624
rect 3682 -2635 3840 -2624
rect 3870 -2635 3916 -2604
rect 3928 -2635 3996 -2604
rect 3694 -2636 3996 -2635
rect 4000 -2610 4168 -2576
rect 1318 -2656 3596 -2636
rect 3662 -2638 3670 -2636
rect 1250 -2658 3596 -2656
rect 3704 -2658 3712 -2638
rect 3720 -2654 3754 -2636
rect 3878 -2658 3881 -2636
rect 41 -2669 3793 -2658
rect 3829 -2669 3881 -2658
rect 41 -2675 3782 -2669
rect 41 -2684 85 -2675
rect 14 -2688 85 -2684
rect 93 -2681 3782 -2675
rect 3840 -2681 3870 -2669
rect 93 -2688 3793 -2681
rect 3829 -2688 3881 -2681
rect -88 -2698 0 -2690
rect 14 -2692 3881 -2688
rect 14 -2711 43 -2692
rect 97 -2711 131 -2700
rect 211 -2711 245 -2692
rect 264 -2711 298 -2692
rect 352 -2711 791 -2692
rect 868 -2709 881 -2696
rect 949 -2709 983 -2692
rect -17 -2718 791 -2711
rect -88 -2726 791 -2718
rect -17 -2737 791 -2726
rect 865 -2730 989 -2709
rect -17 -2750 815 -2737
rect 865 -2743 881 -2730
rect 949 -2737 983 -2730
rect 903 -2743 983 -2737
rect -17 -2803 791 -2750
rect 865 -2766 869 -2743
rect 899 -2758 983 -2743
rect 899 -2762 928 -2758
rect 899 -2777 915 -2762
rect 949 -2777 983 -2758
rect 903 -2783 983 -2777
rect -17 -2809 837 -2803
rect -17 -2843 791 -2809
rect 812 -2824 825 -2809
rect 837 -2843 841 -2809
rect 949 -2820 983 -2783
rect 871 -2824 875 -2820
rect 859 -2843 875 -2824
rect -17 -2849 837 -2843
rect -17 -2911 791 -2849
rect 871 -2877 875 -2843
rect 949 -2911 993 -2820
rect 1002 -2824 1036 -2692
rect 1002 -2892 1027 -2824
rect 1073 -2858 1107 -2692
rect 1116 -2697 1184 -2692
rect 1116 -2713 1160 -2697
rect 1234 -2713 1238 -2692
rect 1126 -2722 1160 -2713
rect 1120 -2730 1234 -2722
rect 1268 -2724 1272 -2692
rect 1284 -2709 1297 -2692
rect 1318 -2694 3596 -2692
rect 1318 -2698 3579 -2694
rect 1318 -2730 2495 -2698
rect 1126 -2750 1160 -2730
rect 1318 -2734 1959 -2730
rect 1966 -2734 2024 -2730
rect 2033 -2734 2495 -2730
rect 1126 -2756 1206 -2750
rect 1126 -2758 1210 -2756
rect 1126 -2790 1160 -2758
rect 1181 -2771 1194 -2758
rect 1206 -2790 1210 -2758
rect 1318 -2761 1965 -2734
rect 1966 -2746 2495 -2734
rect 1975 -2750 2495 -2746
rect 1972 -2751 2495 -2750
rect 2586 -2751 2615 -2698
rect 2771 -2726 3579 -2698
rect 3704 -2704 3712 -2692
rect 3782 -2716 3786 -2710
rect 3782 -2726 3796 -2716
rect 1972 -2761 2250 -2751
rect 1318 -2762 2250 -2761
rect 1240 -2771 1244 -2767
rect 1228 -2790 1244 -2771
rect 1126 -2796 1206 -2790
rect 1126 -2858 1160 -2796
rect 1240 -2824 1244 -2790
rect 1318 -2768 1965 -2762
rect 1972 -2768 2250 -2762
rect 1318 -2773 1959 -2768
rect 1318 -2777 1952 -2773
rect 1318 -2796 1932 -2777
rect 2033 -2778 2250 -2768
rect 2010 -2784 2250 -2778
rect 1318 -2806 1918 -2796
rect 2006 -2802 2250 -2784
rect 2006 -2806 2022 -2802
rect 2033 -2806 2250 -2802
rect 1318 -2838 2250 -2806
rect 2276 -2804 2296 -2751
rect 2276 -2819 2311 -2804
rect 2276 -2838 2296 -2819
rect 1318 -2857 2263 -2838
rect 1318 -2858 1352 -2857
rect 1073 -2892 1352 -2858
rect -17 -2926 993 -2911
rect -17 -2945 983 -2926
rect -17 -2981 791 -2945
rect -17 -3034 650 -2981
rect -17 -3087 281 -3034
rect 187 -3129 200 -3087
rect 215 -3101 228 -3087
rect 354 -3256 369 -3034
rect 388 -3188 422 -3034
rect 534 -3086 592 -3080
rect 534 -3120 546 -3086
rect 534 -3126 592 -3120
rect 721 -3153 791 -2981
rect 903 -3051 961 -3045
rect 903 -3085 915 -3051
rect 903 -3091 961 -3085
rect 1073 -3091 1107 -2892
rect 721 -3187 792 -3153
rect 1092 -3168 1107 -3091
rect 1126 -3100 1160 -2892
rect 1272 -2998 1330 -2992
rect 1272 -3032 1284 -2998
rect 1272 -3038 1330 -3032
rect 1126 -3134 1161 -3100
rect 1461 -3115 1476 -2857
rect 1495 -3047 1529 -2857
rect 1640 -2898 1649 -2857
rect 1668 -2920 1677 -2857
rect 1681 -2860 2263 -2857
rect 1681 -2866 2290 -2860
rect 1681 -2876 2298 -2866
rect 1681 -2886 2308 -2876
rect 1681 -2902 2314 -2886
rect 1681 -2906 2308 -2902
rect 1681 -2916 2263 -2906
rect 1681 -2956 2250 -2916
rect 2264 -2920 2308 -2906
rect 2296 -2930 2308 -2920
rect 2402 -2906 2436 -2751
rect 2455 -2784 2489 -2751
rect 2571 -2754 2615 -2751
rect 2557 -2766 2615 -2754
rect 2788 -2730 3579 -2726
rect 2788 -2754 2858 -2730
rect 2788 -2760 2869 -2754
rect 2893 -2760 2949 -2754
rect 3045 -2760 3097 -2754
rect 3170 -2760 3174 -2730
rect 3193 -2735 3251 -2730
rect 3277 -2735 3329 -2730
rect 3389 -2735 3445 -2730
rect 3509 -2735 3579 -2730
rect 3194 -2760 3214 -2735
rect 3526 -2760 3579 -2735
rect 3752 -2756 3762 -2726
rect 3772 -2736 3802 -2726
rect 3776 -2742 3802 -2736
rect 3776 -2756 3796 -2742
rect 3878 -2756 3881 -2692
rect 3897 -2692 3916 -2636
rect 3897 -2756 3912 -2692
rect 3625 -2760 3681 -2756
rect 3752 -2760 3797 -2756
rect 3816 -2760 3912 -2756
rect 2569 -2770 2603 -2766
rect 2657 -2770 2691 -2760
rect 2528 -2784 2530 -2778
rect 2535 -2784 2542 -2782
rect 2455 -2794 2498 -2784
rect 2528 -2794 2542 -2784
rect 2788 -2788 3174 -2760
rect 3526 -2771 3912 -2760
rect 2788 -2794 2841 -2788
rect 3562 -2790 3912 -2771
rect 3828 -2792 3840 -2790
rect 3870 -2792 3882 -2790
rect 3828 -2794 3882 -2792
rect 3931 -2791 3965 -2636
rect 4000 -2639 4019 -2610
rect 4033 -2639 4146 -2610
rect 4000 -2640 4146 -2639
rect 4200 -2626 4246 -2548
rect 4058 -2719 4088 -2640
rect 4091 -2719 4179 -2713
rect 4045 -2722 4179 -2719
rect 4043 -2734 4179 -2722
rect 4200 -2727 4233 -2626
rect 4247 -2727 4281 -2548
rect 4300 -2684 4334 -2548
rect 4402 -2576 4548 -2548
rect 4616 -2559 4686 -2548
rect 4388 -2610 4460 -2576
rect 4402 -2650 4448 -2610
rect 4454 -2626 4460 -2610
rect 4470 -2612 4548 -2576
rect 4554 -2610 4570 -2576
rect 4490 -2626 4520 -2612
rect 4402 -2681 4434 -2650
rect 4490 -2666 4504 -2626
rect 4490 -2681 4519 -2666
rect 4542 -2681 4548 -2612
rect 4582 -2626 4588 -2560
rect 4616 -2649 4650 -2559
rect 4686 -2649 4754 -2559
rect 5353 -2579 5396 -2546
rect 5550 -2579 5584 -2542
rect 5776 -2543 5811 -2526
rect 5740 -2560 5811 -2543
rect 4832 -2640 4890 -2631
rect 4920 -2640 4978 -2631
rect 5373 -2632 5396 -2579
rect 4434 -2684 4502 -2681
rect 4300 -2727 4346 -2684
rect 4376 -2722 4502 -2684
rect 4542 -2684 4543 -2681
rect 4376 -2727 4504 -2722
rect 4200 -2728 4504 -2727
rect 4542 -2727 4600 -2684
rect 4616 -2685 4686 -2649
rect 5038 -2666 5196 -2632
rect 5250 -2666 5396 -2632
rect 4616 -2719 4776 -2685
rect 4879 -2696 4931 -2685
rect 4890 -2708 4920 -2696
rect 4879 -2719 4931 -2708
rect 4616 -2722 4703 -2719
rect 4616 -2727 4758 -2722
rect 4542 -2728 4758 -2727
rect 4091 -2744 4121 -2734
rect 4133 -2738 4167 -2734
rect 4039 -2791 4046 -2747
rect 4112 -2772 4201 -2760
rect 4132 -2775 4157 -2772
rect 4077 -2781 4157 -2775
rect 4073 -2791 4089 -2781
rect 4132 -2791 4157 -2781
rect 4162 -2791 4166 -2772
rect 2455 -2804 2725 -2794
rect 2455 -2810 2546 -2804
rect 2788 -2806 3208 -2794
rect 2455 -2844 2489 -2810
rect 2496 -2828 2540 -2810
rect 2528 -2838 2540 -2828
rect 2601 -2813 2659 -2807
rect 2528 -2844 2530 -2838
rect 2601 -2844 2613 -2813
rect 2616 -2844 2663 -2813
rect 2788 -2824 3210 -2806
rect 2296 -2936 2298 -2930
rect 1681 -2968 2120 -2956
rect 2180 -2964 2191 -2956
rect 2221 -2964 2232 -2956
rect 2174 -2968 2201 -2964
rect 2211 -2968 2238 -2964
rect 2402 -2968 2414 -2906
rect 1681 -2970 2159 -2968
rect 2174 -2970 2238 -2968
rect 2255 -2970 2307 -2968
rect 2369 -2970 2414 -2968
rect 1681 -2979 2414 -2970
rect 1681 -2983 2148 -2979
rect 1716 -3013 1737 -2983
rect 1811 -3047 1845 -2983
rect 2000 -2998 2044 -2983
rect 2032 -3008 2044 -2998
rect 2086 -2991 2148 -2983
rect 2154 -2991 2414 -2979
rect 2415 -2964 2436 -2906
rect 2440 -2915 2490 -2844
rect 2601 -2853 2674 -2844
rect 2616 -2859 2674 -2853
rect 2616 -2863 2663 -2859
rect 2790 -2896 2805 -2824
rect 3528 -2828 3888 -2794
rect 3931 -2825 3982 -2791
rect 4047 -2802 4191 -2791
rect 4058 -2810 4180 -2802
rect 4058 -2814 4139 -2810
rect 4047 -2825 4150 -2814
rect 3870 -2836 3882 -2828
rect 3870 -2842 3872 -2836
rect 3562 -2861 3928 -2844
rect 3157 -2862 3928 -2861
rect 3157 -2867 3670 -2862
rect 3072 -2876 3088 -2870
rect 3046 -2886 3098 -2876
rect 3157 -2878 3681 -2867
rect 3694 -2878 3928 -2862
rect 2771 -2914 2805 -2896
rect 3040 -2896 3104 -2886
rect 3040 -2902 3066 -2896
rect 3056 -2914 3066 -2902
rect 3078 -2902 3104 -2896
rect 3078 -2910 3098 -2902
rect 3076 -2914 3098 -2910
rect 3157 -2914 3596 -2878
rect 2771 -2915 3596 -2914
rect 2440 -2930 2674 -2915
rect 2770 -2920 3596 -2915
rect 2770 -2930 3579 -2920
rect 2440 -2949 3579 -2930
rect 3585 -2931 3596 -2920
rect 2440 -2964 2490 -2949
rect 2788 -2964 3579 -2949
rect 2415 -2970 3579 -2964
rect 3704 -2940 3752 -2930
rect 3754 -2940 3801 -2899
rect 2415 -2991 3596 -2970
rect 2086 -2998 3596 -2991
rect 3704 -2980 3801 -2940
rect 3704 -2986 3766 -2980
rect 3704 -2996 3752 -2986
rect 2086 -3002 2436 -2998
rect 2440 -3003 2490 -2998
rect 2788 -3003 3596 -2998
rect 2032 -3014 2034 -3008
rect 2440 -3024 3596 -3003
rect 2086 -3027 2090 -3024
rect 2208 -3027 2266 -3024
rect 2296 -3027 2354 -3024
rect 1495 -3081 1530 -3047
rect 1704 -3073 1845 -3047
rect 2440 -3032 3608 -3024
rect 3672 -3027 3710 -3018
rect 3722 -3027 3752 -2996
rect 2440 -3037 2674 -3032
rect 2732 -3037 3608 -3032
rect 2086 -3073 2090 -3056
rect 2103 -3067 2159 -3056
rect 1681 -3104 2103 -3073
rect 2114 -3079 2148 -3067
rect 2114 -3090 2159 -3079
rect 2208 -3090 2354 -3056
rect 2369 -3067 2436 -3056
rect 2380 -3079 2414 -3067
rect 2369 -3090 2414 -3079
rect 2114 -3104 2120 -3090
rect 1681 -3117 2120 -3104
rect 1668 -3142 2120 -3117
rect 2210 -3129 2254 -3124
rect 2208 -3142 2254 -3129
rect 2278 -3126 2325 -3111
rect 1668 -3152 2103 -3142
rect 1668 -3170 2112 -3152
rect 1681 -3176 2112 -3170
rect 2114 -3166 2120 -3142
rect 2138 -3166 2158 -3142
rect 2114 -3176 2158 -3166
rect 2208 -3152 2266 -3142
rect 2278 -3152 2328 -3126
rect 2333 -3142 2354 -3095
rect 2402 -3104 2414 -3090
rect 2415 -3104 2436 -3067
rect 2208 -3176 2328 -3152
rect 2380 -3166 2401 -3142
rect 2402 -3152 2436 -3104
rect 2402 -3166 2414 -3152
rect 2380 -3176 2414 -3166
rect 2415 -3176 2436 -3152
rect 388 -3222 423 -3188
rect 721 -3223 774 -3187
rect 1681 -3192 2120 -3176
rect 2132 -3186 2158 -3176
rect 2228 -3185 2328 -3176
rect 2132 -3192 2148 -3186
rect 1668 -3200 2120 -3192
rect 1681 -3220 2120 -3200
rect 2208 -3204 2354 -3185
rect 1668 -3228 2120 -3220
rect 2204 -3224 2318 -3220
rect 1681 -3258 2120 -3228
rect 2200 -3226 2322 -3224
rect 2200 -3258 2234 -3226
rect 2288 -3239 2322 -3226
rect 2276 -3245 2322 -3239
rect 2288 -3258 2322 -3245
rect 2402 -3258 2436 -3176
rect 2440 -3204 2490 -3037
rect 2647 -3089 2674 -3058
rect 2616 -3099 2674 -3089
rect 2601 -3105 2674 -3099
rect 2563 -3158 2574 -3126
rect 2597 -3139 2674 -3105
rect 2601 -3145 2663 -3139
rect 2616 -3155 2663 -3145
rect 2563 -3164 2603 -3158
rect 2540 -3176 2603 -3164
rect 2574 -3182 2603 -3176
rect 2594 -3187 2603 -3182
rect 2616 -3164 2645 -3155
rect 2616 -3176 2662 -3164
rect 2616 -3186 2645 -3176
rect 2586 -3204 2603 -3187
rect 2455 -3258 2489 -3204
rect 2586 -3224 2615 -3204
rect 2569 -3230 2615 -3224
rect 2569 -3258 2603 -3230
rect 2628 -3258 2637 -3186
rect 2732 -3204 2757 -3132
rect 2771 -3204 3608 -3037
rect 3664 -3039 3710 -3027
rect 3764 -3028 3798 -3018
rect 3753 -3039 3798 -3028
rect 3664 -3042 3685 -3039
rect 3664 -3052 3670 -3042
rect 3672 -3052 3676 -3042
rect 3764 -3052 3798 -3039
rect 3878 -3052 3928 -2878
rect 3610 -3086 3928 -3052
rect 3931 -2883 3965 -2825
rect 4055 -2883 4157 -2859
rect 3931 -2917 3982 -2883
rect 4047 -2894 4161 -2883
rect 4258 -2886 4281 -2728
rect 4300 -2768 4315 -2728
rect 4446 -2738 4458 -2728
rect 4616 -2738 4630 -2728
rect 4335 -2749 4387 -2738
rect 4431 -2749 4519 -2738
rect 4589 -2749 4630 -2738
rect 4346 -2761 4376 -2749
rect 4442 -2761 4508 -2749
rect 4600 -2761 4630 -2749
rect 4335 -2772 4387 -2761
rect 4431 -2772 4519 -2761
rect 4589 -2772 4630 -2761
rect 4051 -2906 4161 -2894
rect 4228 -2902 4281 -2886
rect 4300 -2834 4315 -2794
rect 4327 -2830 4334 -2803
rect 4400 -2824 4404 -2814
rect 4424 -2830 4526 -2806
rect 4616 -2830 4630 -2772
rect 4327 -2834 4530 -2830
rect 4300 -2841 4530 -2834
rect 4589 -2841 4630 -2830
rect 4300 -2853 4334 -2841
rect 4338 -2853 4530 -2841
rect 4600 -2853 4630 -2841
rect 4300 -2864 4530 -2853
rect 4589 -2864 4630 -2853
rect 4228 -2906 4298 -2902
rect 4047 -2917 4161 -2906
rect 4217 -2917 4298 -2906
rect 3931 -3086 3965 -2917
rect 4077 -2927 4089 -2917
rect 4077 -2933 4135 -2927
rect 4247 -2936 4298 -2917
rect 4046 -2970 4079 -2965
rect 4041 -2974 4079 -2970
rect 4091 -2974 4121 -2943
rect 4133 -2974 4167 -2965
rect 4041 -2988 4091 -2974
rect 4133 -2988 4179 -2974
rect 4000 -2999 4019 -2988
rect 4041 -2989 4079 -2988
rect 4088 -2989 4121 -2988
rect 4041 -2999 4045 -2989
rect 4058 -2999 4079 -2989
rect 4091 -2999 4121 -2989
rect 4133 -2999 4167 -2988
rect 4200 -2999 4233 -2988
rect 4247 -2999 4281 -2936
rect 4300 -2999 4334 -2864
rect 4442 -2874 4458 -2864
rect 4442 -2880 4504 -2874
rect 4616 -2886 4630 -2864
rect 4633 -2859 4703 -2728
rect 4720 -2781 4722 -2760
rect 4815 -2787 4873 -2781
rect 4815 -2796 4827 -2787
rect 4811 -2821 4877 -2796
rect 4815 -2827 4873 -2821
rect 4890 -2830 4919 -2729
rect 4777 -2837 4919 -2830
rect 4777 -2855 4911 -2837
rect 4890 -2859 4901 -2855
rect 4633 -2864 4932 -2859
rect 4633 -2886 4703 -2864
rect 4580 -2912 4596 -2902
rect 4616 -2910 4703 -2886
rect 4779 -2871 4817 -2864
rect 4779 -2893 4783 -2871
rect 4871 -2886 4917 -2864
rect 4824 -2893 4829 -2886
rect 4859 -2893 4917 -2886
rect 4932 -2893 4939 -2864
rect 4951 -2893 4966 -2719
rect 4985 -2859 5000 -2719
rect 5004 -2859 5019 -2685
rect 4985 -2893 5019 -2859
rect 5038 -2694 5073 -2666
rect 5354 -2694 5396 -2666
rect 5038 -2714 5096 -2694
rect 5158 -2700 5196 -2696
rect 5250 -2700 5268 -2696
rect 5150 -2714 5280 -2700
rect 5350 -2714 5396 -2694
rect 5038 -2716 5073 -2714
rect 5038 -2726 5084 -2716
rect 5150 -2726 5196 -2714
rect 5250 -2726 5280 -2714
rect 5354 -2716 5396 -2714
rect 5342 -2726 5396 -2716
rect 5407 -2613 5596 -2579
rect 4717 -2898 4932 -2893
rect 4717 -2902 4737 -2898
rect 4717 -2904 4729 -2902
rect 4771 -2904 4931 -2898
rect 4717 -2910 4718 -2904
rect 4616 -2912 4734 -2910
rect 4410 -2933 4448 -2912
rect 4502 -2921 4536 -2912
rect 4410 -2946 4414 -2933
rect 4490 -2946 4536 -2921
rect 4580 -2936 4734 -2912
rect 4771 -2916 4920 -2904
rect 4771 -2927 4931 -2916
rect 4985 -2927 5005 -2893
rect 5038 -2927 5072 -2726
rect 5150 -2730 5184 -2726
rect 5262 -2730 5280 -2726
rect 5170 -2748 5246 -2734
rect 5170 -2764 5226 -2748
rect 5228 -2764 5246 -2748
rect 5170 -2765 5180 -2764
rect 5196 -2768 5226 -2764
rect 5373 -2768 5388 -2726
rect 5154 -2806 5198 -2781
rect 5407 -2806 5441 -2613
rect 5450 -2636 5495 -2613
rect 5462 -2640 5475 -2636
rect 5508 -2665 5538 -2623
rect 5549 -2675 5580 -2665
rect 5549 -2681 5611 -2675
rect 5549 -2715 5580 -2681
rect 5740 -2698 5810 -2560
rect 5922 -2628 5980 -2622
rect 5922 -2662 5934 -2628
rect 5922 -2668 5980 -2662
rect 6111 -2698 6126 -2526
rect 6145 -2565 6179 -2507
rect 6269 -2565 6371 -2541
rect 6145 -2599 6180 -2565
rect 6265 -2599 6375 -2565
rect 6145 -2698 6179 -2599
rect 6291 -2609 6303 -2599
rect 6291 -2615 6349 -2609
rect 6480 -2647 6495 -1895
rect 6255 -2668 6293 -2647
rect 6255 -2681 6259 -2668
rect 6347 -2681 6381 -2647
rect 6461 -2681 6495 -2647
rect 6514 -2420 6548 -1861
rect 6847 -1873 6918 -1839
rect 6994 -1873 7122 -1839
rect 6660 -1922 6718 -1916
rect 6660 -1956 6672 -1922
rect 6660 -1962 6718 -1956
rect 6847 -2171 6917 -1873
rect 7029 -1903 7041 -1873
rect 7029 -1909 7087 -1903
rect 7029 -2069 7087 -2063
rect 7029 -2103 7041 -2069
rect 7029 -2109 7087 -2103
rect 6847 -2205 6918 -2171
rect 7218 -2186 7233 -1777
rect 7252 -1522 7287 -1488
rect 7252 -1714 7286 -1522
rect 7585 -1584 7655 -1467
rect 7954 -1468 8007 -1432
rect 8359 -1466 8374 -1432
rect 8692 -1485 8762 -1026
rect 9044 -1045 9078 -1026
rect 8874 -1094 8932 -1088
rect 8874 -1128 8886 -1094
rect 8874 -1134 8932 -1128
rect 8874 -1402 8932 -1396
rect 8874 -1436 8886 -1402
rect 8874 -1442 8932 -1436
rect 7767 -1535 7825 -1529
rect 7767 -1569 7779 -1535
rect 7812 -1569 7825 -1535
rect 7767 -1575 7825 -1569
rect 7398 -1590 7456 -1584
rect 7398 -1624 7410 -1590
rect 7398 -1630 7456 -1624
rect 7366 -1714 7400 -1658
rect 7454 -1714 7488 -1658
rect 7568 -1661 7655 -1584
rect 7840 -1603 7853 -1501
rect 8692 -1502 8745 -1485
rect 7937 -1558 7971 -1529
rect 8692 -1538 8763 -1502
rect 8824 -1538 8982 -1502
rect 7937 -1594 8007 -1558
rect 8359 -1589 8394 -1555
rect 7735 -1661 7769 -1612
rect 7823 -1661 7857 -1612
rect 7937 -1642 8025 -1594
rect 8086 -1642 8244 -1594
rect 7568 -1695 7656 -1661
rect 7723 -1695 7869 -1661
rect 7252 -1748 7287 -1714
rect 7354 -1748 7500 -1714
rect 7252 -1892 7286 -1748
rect 7410 -1850 7444 -1790
rect 7332 -1892 7522 -1866
rect 7252 -1926 7287 -1892
rect 7332 -1900 7500 -1892
rect 7348 -1926 7500 -1900
rect 7506 -1926 7522 -1892
rect 7252 -2118 7286 -1926
rect 7568 -1945 7655 -1695
rect 7741 -1747 7769 -1725
rect 7813 -1747 7860 -1716
rect 7741 -1763 7781 -1747
rect 7811 -1763 7860 -1747
rect 7741 -1784 7860 -1763
rect 7748 -1790 7860 -1784
rect 7723 -1796 7869 -1790
rect 7763 -1797 7829 -1796
rect 7763 -1813 7781 -1797
rect 7811 -1813 7829 -1797
rect 7763 -1844 7829 -1843
rect 7748 -1856 7860 -1844
rect 7741 -1877 7860 -1856
rect 7741 -1893 7781 -1877
rect 7811 -1893 7851 -1877
rect 7741 -1911 7769 -1893
rect 7735 -1945 7769 -1911
rect 7823 -1911 7851 -1893
rect 7823 -1945 7857 -1911
rect 7568 -1979 7656 -1945
rect 7717 -1979 7869 -1945
rect 7875 -1979 7891 -1945
rect 7398 -2016 7456 -2010
rect 7398 -2050 7410 -2016
rect 7398 -2056 7456 -2050
rect 7568 -2056 7655 -1979
rect 7937 -1998 8024 -1642
rect 8325 -1690 8340 -1594
rect 8148 -1730 8182 -1696
rect 8132 -1744 8198 -1730
rect 8158 -1750 8194 -1744
rect 8104 -1768 8138 -1764
rect 8104 -1775 8150 -1768
rect 8104 -1778 8138 -1775
rect 8104 -1858 8138 -1780
rect 8158 -1856 8164 -1750
rect 8192 -1768 8226 -1764
rect 8180 -1775 8226 -1768
rect 8186 -1778 8226 -1775
rect 8186 -1780 8192 -1778
rect 8186 -1858 8226 -1780
rect 8104 -1860 8226 -1858
rect 8110 -1862 8220 -1860
rect 8104 -1872 8226 -1862
rect 8104 -1876 8138 -1872
rect 8192 -1876 8226 -1872
rect 8136 -1896 8194 -1890
rect 8132 -1910 8198 -1896
rect 8148 -1944 8182 -1910
rect 8306 -1950 8340 -1690
rect 7252 -2152 7287 -2118
rect 7585 -2152 7655 -2056
rect 7767 -2071 7825 -2065
rect 7767 -2105 7779 -2071
rect 7812 -2105 7825 -2071
rect 7840 -2098 7853 -2037
rect 7937 -2046 8025 -1998
rect 8086 -2046 8244 -1998
rect 8325 -2046 8340 -1950
rect 8359 -1647 8393 -1589
rect 8692 -1592 8762 -1538
rect 8852 -1592 8954 -1570
rect 8483 -1647 8585 -1623
rect 8692 -1626 8763 -1592
rect 8848 -1626 8958 -1592
rect 9063 -1598 9078 -1045
rect 8359 -1681 8394 -1647
rect 8470 -1675 8598 -1647
rect 8692 -1651 8762 -1626
rect 8874 -1636 8886 -1626
rect 8407 -1681 8661 -1675
rect 8359 -1959 8393 -1681
rect 8505 -1691 8517 -1681
rect 8505 -1697 8563 -1691
rect 8551 -1733 8589 -1729
rect 8501 -1741 8519 -1733
rect 8479 -1749 8519 -1741
rect 8549 -1749 8589 -1733
rect 8479 -1767 8589 -1749
rect 8461 -1819 8607 -1767
rect 8467 -1841 8513 -1821
rect 8551 -1841 8601 -1821
rect 8467 -1847 8519 -1841
rect 8479 -1857 8519 -1847
rect 8549 -1847 8601 -1841
rect 8549 -1857 8589 -1847
rect 8479 -1891 8589 -1857
rect 8479 -1899 8519 -1891
rect 8501 -1905 8519 -1899
rect 8461 -1907 8519 -1905
rect 8549 -1899 8589 -1891
rect 8549 -1905 8567 -1899
rect 8549 -1907 8607 -1905
rect 8461 -1911 8501 -1907
rect 8567 -1911 8607 -1907
rect 8505 -1949 8563 -1943
rect 8505 -1959 8517 -1949
rect 8359 -1993 8394 -1959
rect 8490 -1970 8578 -1959
rect 8501 -1982 8567 -1970
rect 8490 -1993 8578 -1982
rect 8675 -1989 8762 -1651
rect 8870 -1638 8888 -1636
rect 8918 -1638 8936 -1636
rect 8870 -1644 8936 -1638
rect 8870 -1654 8888 -1644
rect 8918 -1654 8936 -1644
rect 8855 -1694 8888 -1685
rect 8918 -1694 8967 -1685
rect 8855 -1697 8967 -1694
rect 8842 -1728 8967 -1697
rect 8842 -1744 8888 -1728
rect 8918 -1744 8964 -1728
rect 8842 -1896 8876 -1744
rect 8930 -1865 8964 -1744
rect 8920 -1896 8967 -1865
rect 8842 -1912 8888 -1896
rect 8918 -1912 8967 -1896
rect 8842 -1943 8967 -1912
rect 8855 -1946 8967 -1943
rect 8855 -1955 8888 -1946
rect 8870 -1962 8888 -1955
rect 8918 -1955 8951 -1946
rect 8918 -1962 8936 -1955
rect 8359 -2046 8393 -1993
rect 8692 -2014 8762 -1989
rect 8874 -2002 8932 -1996
rect 8874 -2014 8886 -2002
rect 7937 -2082 8007 -2046
rect 8359 -2080 8374 -2046
rect 8692 -2048 8763 -2014
rect 8859 -2025 8947 -2014
rect 8870 -2037 8936 -2025
rect 8859 -2048 8947 -2037
rect 9044 -2042 9078 -1598
rect 7767 -2111 7825 -2105
rect 7937 -2111 7971 -2082
rect 8692 -2085 8762 -2048
rect 8692 -2102 8745 -2085
rect 8692 -2138 8763 -2102
rect 8824 -2138 8982 -2102
rect 7585 -2188 7638 -2152
rect 7937 -2172 7971 -2154
rect 7937 -2173 8007 -2172
rect 6847 -2241 6900 -2205
rect 7936 -2207 8007 -2173
rect 7954 -2208 8007 -2207
rect 8359 -2189 8394 -2155
rect 7954 -2242 8025 -2208
rect 7621 -2278 7656 -2261
rect 7585 -2295 7656 -2278
rect 6830 -2331 6864 -2313
rect 6830 -2367 6900 -2331
rect 7252 -2348 7287 -2314
rect 6847 -2401 6918 -2367
rect 6660 -2410 6718 -2404
rect 6660 -2420 6672 -2410
rect 6514 -2454 6549 -2420
rect 6645 -2431 6733 -2420
rect 6656 -2443 6722 -2431
rect 6645 -2454 6733 -2443
rect 6514 -2512 6548 -2454
rect 6638 -2512 6740 -2488
rect 6514 -2546 6549 -2512
rect 6634 -2546 6744 -2512
rect 6193 -2698 6233 -2681
rect 5740 -2715 6233 -2698
rect 6247 -2715 6393 -2681
rect 6461 -2715 6481 -2681
rect 6514 -2715 6548 -2546
rect 6660 -2556 6672 -2546
rect 6660 -2562 6718 -2556
rect 6847 -2592 6917 -2401
rect 7029 -2469 7087 -2463
rect 7029 -2503 7041 -2469
rect 7029 -2509 7087 -2503
rect 7218 -2541 7233 -2367
rect 6993 -2553 7031 -2541
rect 6993 -2575 6997 -2553
rect 7085 -2575 7119 -2541
rect 7199 -2575 7233 -2541
rect 6931 -2592 6971 -2575
rect 6847 -2594 6971 -2592
rect 6624 -2615 6662 -2594
rect 6624 -2628 6628 -2615
rect 6716 -2628 6750 -2594
rect 6830 -2609 6971 -2594
rect 6985 -2609 7131 -2575
rect 7199 -2609 7219 -2575
rect 7252 -2609 7286 -2348
rect 7398 -2416 7456 -2410
rect 7398 -2450 7410 -2416
rect 7398 -2456 7456 -2450
rect 7585 -2486 7655 -2295
rect 7767 -2363 7825 -2357
rect 7767 -2397 7779 -2363
rect 7767 -2403 7825 -2397
rect 7585 -2488 7686 -2486
rect 7362 -2500 7400 -2488
rect 7362 -2522 7366 -2500
rect 7454 -2522 7488 -2488
rect 5549 -2721 5611 -2715
rect 5549 -2731 5584 -2721
rect 5521 -2753 5546 -2749
rect 5567 -2753 5584 -2731
rect 5509 -2768 5561 -2753
rect 5487 -2784 5561 -2768
rect 5575 -2772 5584 -2753
rect 5609 -2753 5618 -2749
rect 5740 -2753 6227 -2715
rect 5461 -2787 5561 -2784
rect 5572 -2784 5589 -2772
rect 5609 -2784 5643 -2753
rect 5572 -2787 5643 -2784
rect 5138 -2815 5226 -2806
rect 5138 -2831 5204 -2815
rect 5140 -2840 5186 -2831
rect 5240 -2840 5274 -2806
rect 5354 -2834 5374 -2806
rect 5388 -2834 5441 -2806
rect 5354 -2840 5388 -2834
rect 5407 -2840 5441 -2834
rect 4616 -2946 4737 -2936
rect 3610 -3142 3644 -3086
rect 3664 -3095 3670 -3086
rect 3676 -3095 3710 -3086
rect 3664 -3142 3717 -3095
rect 3764 -3120 3798 -3086
rect 3734 -3126 3798 -3120
rect 3718 -3138 3798 -3126
rect 3878 -3126 3912 -3086
rect 3718 -3142 3818 -3138
rect 3610 -3166 3655 -3142
rect 3664 -3154 3828 -3142
rect 3664 -3166 3740 -3154
rect 3610 -3176 3740 -3166
rect 2657 -3258 2691 -3224
rect 2771 -3258 3596 -3204
rect 3610 -3220 3644 -3176
rect 3664 -3181 3710 -3176
rect 3718 -3181 3740 -3176
rect 3664 -3192 3740 -3181
rect 3752 -3176 3828 -3154
rect 3752 -3181 3849 -3176
rect 3878 -3181 3916 -3126
rect 3664 -3207 3722 -3192
rect 3752 -3204 3916 -3181
rect 3752 -3207 3810 -3204
rect 3676 -3211 3678 -3207
rect 3690 -3211 3710 -3207
rect 3764 -3211 3798 -3207
rect 3840 -3220 3842 -3207
rect 3610 -3222 3842 -3220
rect 3610 -3224 3832 -3222
rect 3840 -3224 3842 -3222
rect 3610 -3235 3874 -3224
rect 3610 -3258 3644 -3235
rect 3712 -3247 3800 -3235
rect 3712 -3258 3801 -3247
rect 3812 -3258 3874 -3235
rect 1681 -3292 3874 -3258
rect 3878 -3258 3916 -3204
rect 3878 -3292 3880 -3258
rect 3892 -3292 3916 -3258
rect 1681 -3330 2120 -3292
rect 2050 -3547 2120 -3330
rect 2232 -3466 2290 -3460
rect 2232 -3500 2244 -3466
rect 2232 -3506 2290 -3500
rect 2402 -3506 2436 -3292
rect 2050 -3583 2103 -3547
rect 2421 -3583 2436 -3506
rect 2455 -3515 2489 -3292
rect 2771 -3330 3596 -3292
rect 2771 -3354 2858 -3330
rect 2771 -3388 2859 -3354
rect 3159 -3369 3174 -3330
rect 3193 -3335 3596 -3330
rect 3205 -3356 3596 -3335
rect 3205 -3371 3591 -3356
rect 2601 -3413 2659 -3407
rect 2601 -3447 2613 -3413
rect 2771 -3424 2841 -3388
rect 3205 -3424 3210 -3371
rect 2601 -3453 2659 -3447
rect 2771 -3453 2805 -3424
rect 2455 -3549 2490 -3515
rect 3241 -3555 3275 -3371
rect 3557 -3555 3591 -3371
rect 1668 -3600 1734 -3592
rect 1668 -3628 1734 -3620
rect 3576 -3632 3591 -3555
rect 3610 -3564 3644 -3292
rect 3712 -3304 3770 -3292
rect 3712 -3319 3727 -3304
rect 3844 -3356 3846 -3292
rect 3853 -3356 3858 -3292
rect 3878 -3356 3912 -3292
rect 3658 -3390 3678 -3356
rect 3712 -3390 3858 -3356
rect 3892 -3390 3912 -3356
rect 3724 -3419 3758 -3390
rect 3756 -3462 3814 -3456
rect 3756 -3496 3768 -3462
rect 3926 -3483 3965 -3086
rect 3979 -3033 4179 -2999
rect 4200 -3033 4334 -2999
rect 3979 -3106 4019 -3033
rect 4045 -3106 4079 -3033
rect 3979 -3140 4079 -3106
rect 3979 -3168 4019 -3140
rect 4045 -3154 4079 -3140
rect 4091 -3067 4121 -3033
rect 4091 -3085 4133 -3067
rect 4171 -3070 4179 -3054
rect 4164 -3085 4179 -3070
rect 4091 -3101 4179 -3085
rect 4200 -3056 4233 -3033
rect 4200 -3101 4246 -3056
rect 4091 -3128 4246 -3101
rect 4247 -3128 4281 -3033
rect 4091 -3135 4281 -3128
rect 4091 -3151 4179 -3135
rect 4045 -3168 4085 -3154
rect 4091 -3168 4121 -3151
rect 4133 -3166 4179 -3151
rect 3979 -3483 4013 -3168
rect 4033 -3182 4088 -3168
rect 4100 -3178 4113 -3168
rect 4093 -3182 4113 -3178
rect 4033 -3183 4113 -3182
rect 4033 -3194 4121 -3183
rect 4033 -3220 4085 -3194
rect 4087 -3220 4127 -3194
rect 4033 -3258 4079 -3220
rect 4093 -3258 4127 -3220
rect 4133 -3220 4173 -3166
rect 4200 -3168 4281 -3135
rect 4181 -3182 4215 -3178
rect 4175 -3190 4215 -3182
rect 4175 -3194 4201 -3190
rect 4175 -3220 4205 -3194
rect 4133 -3258 4167 -3220
rect 4181 -3224 4205 -3220
rect 4213 -3224 4215 -3190
rect 4181 -3258 4215 -3224
rect 4222 -3258 4227 -3182
rect 4247 -3258 4281 -3168
rect 4295 -3258 4334 -3033
rect 4348 -2952 4737 -2946
rect 4746 -2949 4751 -2927
rect 4771 -2934 4805 -2927
rect 4824 -2934 4829 -2927
rect 4771 -2949 4829 -2934
rect 4840 -2936 4917 -2927
rect 4749 -2952 4751 -2949
rect 4783 -2952 4785 -2949
rect 4824 -2952 4829 -2949
rect 4859 -2949 4917 -2936
rect 4859 -2952 4919 -2949
rect 4932 -2952 4939 -2927
rect 4951 -2952 4966 -2927
rect 4985 -2952 5019 -2927
rect 4348 -2961 5019 -2952
rect 5033 -2961 5072 -2927
rect 5086 -2851 5286 -2840
rect 5297 -2851 5349 -2840
rect 5086 -2863 5338 -2851
rect 5086 -2874 5349 -2863
rect 5354 -2874 5374 -2840
rect 5388 -2868 5441 -2840
rect 5407 -2874 5441 -2868
rect 5086 -2961 5120 -2874
rect 5140 -2896 5154 -2874
rect 5221 -2884 5286 -2874
rect 5293 -2884 5308 -2874
rect 5228 -2896 5336 -2884
rect 5152 -2900 5154 -2896
rect 5243 -2917 5336 -2896
rect 5206 -2942 5246 -2934
rect 5250 -2942 5290 -2936
rect 5206 -2951 5294 -2942
rect 5150 -2961 5154 -2951
rect 5206 -2961 5230 -2951
rect 5244 -2961 5268 -2951
rect 5308 -2961 5336 -2917
rect 5368 -2961 5388 -2874
rect 5402 -2961 5441 -2874
rect 5455 -2821 5655 -2787
rect 5723 -2821 6227 -2753
rect 5455 -2834 5561 -2821
rect 5572 -2830 5589 -2821
rect 5455 -2961 5489 -2834
rect 5509 -2843 5561 -2834
rect 5575 -2843 5584 -2830
rect 5508 -2847 5546 -2843
rect 5508 -2865 5538 -2847
rect 5567 -2865 5584 -2843
rect 5609 -2831 5643 -2821
rect 5609 -2847 5618 -2831
rect 5549 -2881 5584 -2865
rect 5549 -2915 5599 -2881
rect 5604 -2883 5611 -2875
rect 5615 -2889 5631 -2881
rect 5632 -2883 5639 -2847
rect 5613 -2915 5637 -2889
rect 5737 -2907 6227 -2821
rect 5549 -2931 5584 -2915
rect 5597 -2923 5637 -2915
rect 5563 -2957 5584 -2931
rect 5632 -2961 5637 -2933
rect 4348 -2980 5637 -2961
rect 4348 -2988 4382 -2980
rect 4402 -2988 4448 -2980
rect 4348 -3005 4402 -2988
rect 4348 -3258 4382 -3005
rect 4414 -3056 4448 -2988
rect 4490 -3001 4504 -2980
rect 4616 -2983 5637 -2980
rect 5689 -2983 5691 -2957
rect 5698 -2983 5703 -2961
rect 5723 -2983 6227 -2907
rect 4548 -3001 4600 -2988
rect 4489 -3005 4600 -3001
rect 4489 -3014 4587 -3005
rect 4472 -3048 4587 -3014
rect 4388 -3059 4448 -3056
rect 4490 -3059 4587 -3048
rect 4388 -3082 4587 -3059
rect 4616 -3017 5703 -2983
rect 5737 -3017 6227 -2983
rect 6247 -2826 6281 -2715
rect 6317 -2767 6347 -2749
rect 6385 -2752 6393 -2736
rect 6378 -2767 6393 -2752
rect 6317 -2783 6393 -2767
rect 6335 -2817 6415 -2783
rect 6475 -2810 6495 -2715
rect 6247 -2836 6293 -2826
rect 6335 -2833 6393 -2817
rect 6247 -3016 6299 -2836
rect 6347 -2848 6393 -2833
rect 6307 -2864 6341 -2860
rect 6301 -3016 6341 -2864
rect 6347 -3016 6387 -2848
rect 6395 -2864 6415 -2860
rect 6389 -2876 6415 -2864
rect 4388 -3090 4556 -3082
rect 4388 -3098 4588 -3090
rect 4388 -3106 4549 -3098
rect 4388 -3129 4460 -3106
rect 4470 -3125 4549 -3106
rect 4554 -3125 4588 -3098
rect 4462 -3129 4549 -3125
rect 4550 -3129 4588 -3125
rect 4388 -3140 4588 -3129
rect 4388 -3154 4542 -3140
rect 4388 -3156 4454 -3154
rect 4414 -3168 4454 -3156
rect 4402 -3220 4454 -3168
rect 4456 -3220 4496 -3154
rect 4402 -3258 4448 -3220
rect 4462 -3258 4496 -3220
rect 4502 -3220 4542 -3154
rect 4544 -3141 4570 -3140
rect 4544 -3220 4574 -3141
rect 4582 -3168 4588 -3140
rect 4616 -3159 5632 -3017
rect 5740 -3108 6227 -3017
rect 6259 -3020 6261 -3016
rect 6273 -3020 6293 -3016
rect 6295 -3044 6383 -3016
rect 6389 -3032 6419 -2876
rect 6389 -3044 6415 -3032
rect 6307 -3048 6341 -3044
rect 6353 -3047 6377 -3044
rect 6395 -3048 6415 -3044
rect 6427 -3048 6429 -2860
rect 6436 -3044 6441 -2864
rect 6461 -3044 6495 -2810
rect 6291 -3063 6349 -3057
rect 6287 -3082 6369 -3063
rect 6461 -3082 6463 -3044
rect 6313 -3097 6337 -3082
rect 6349 -3085 6369 -3082
rect 6353 -3091 6369 -3085
rect 4582 -3190 4596 -3168
rect 4585 -3209 4596 -3190
rect 4502 -3224 4538 -3220
rect 4550 -3224 4574 -3220
rect 4502 -3258 4536 -3224
rect 4550 -3258 4584 -3224
rect 4591 -3258 4596 -3209
rect 4616 -3258 4650 -3159
rect 4664 -3173 5632 -3159
rect 4664 -3179 5659 -3173
rect 4664 -3203 5643 -3179
rect 4664 -3219 5659 -3203
rect 5790 -3205 5805 -3108
rect 5824 -3205 5858 -3108
rect 5970 -3126 6028 -3120
rect 5970 -3160 5982 -3126
rect 6109 -3152 6227 -3108
rect 6351 -3125 6375 -3091
rect 5970 -3166 6028 -3160
rect 6104 -3165 6227 -3152
rect 6104 -3205 6210 -3165
rect 6241 -3188 6399 -3165
rect 4664 -3258 5632 -3219
rect 4020 -3281 5632 -3258
rect 4020 -3292 5709 -3281
rect 4033 -3330 4079 -3292
rect 4093 -3330 4127 -3292
rect 4033 -3334 4085 -3330
rect 4087 -3334 4127 -3330
rect 4133 -3330 4167 -3292
rect 4181 -3330 4205 -3292
rect 4133 -3334 4173 -3330
rect 4045 -3338 4047 -3334
rect 4059 -3338 4079 -3334
rect 4081 -3362 4169 -3334
rect 4175 -3350 4205 -3330
rect 4175 -3362 4201 -3350
rect 4093 -3366 4127 -3362
rect 4139 -3365 4163 -3362
rect 4181 -3366 4201 -3362
rect 4213 -3366 4215 -3292
rect 4222 -3362 4227 -3292
rect 4077 -3381 4135 -3375
rect 4073 -3400 4155 -3381
rect 4099 -3415 4123 -3400
rect 4135 -3403 4155 -3400
rect 4139 -3409 4155 -3403
rect 4137 -3443 4161 -3409
rect 4247 -3421 4281 -3292
rect 3756 -3502 3814 -3496
rect 3926 -3502 3960 -3483
rect 4027 -3511 4185 -3483
rect 4261 -3511 4281 -3421
rect 4295 -3430 4334 -3292
rect 4348 -3430 4382 -3292
rect 4450 -3309 4538 -3292
rect 4462 -3313 4496 -3309
rect 4508 -3312 4532 -3309
rect 4582 -3313 4584 -3292
rect 4591 -3309 4596 -3292
rect 4504 -3328 4580 -3322
rect 4442 -3330 4580 -3328
rect 4442 -3347 4524 -3330
rect 4468 -3362 4492 -3347
rect 4504 -3350 4524 -3347
rect 4504 -3358 4552 -3350
rect 4506 -3390 4530 -3358
rect 4616 -3368 4650 -3292
rect 4295 -3464 4335 -3430
rect 4396 -3458 4554 -3430
rect 4630 -3458 4650 -3368
rect 4664 -3315 5709 -3292
rect 5735 -3298 6210 -3205
rect 6236 -3193 6399 -3188
rect 6475 -3193 6495 -3044
rect 6509 -3112 6548 -2715
rect 6562 -2662 6602 -2628
rect 6616 -2662 6762 -2628
rect 6830 -2662 6965 -2609
rect 6985 -2631 7019 -2609
rect 6997 -2635 6999 -2631
rect 6562 -3112 6596 -2662
rect 6616 -2773 6650 -2662
rect 6686 -2714 6716 -2696
rect 6754 -2699 6762 -2683
rect 6747 -2714 6762 -2699
rect 6686 -2730 6762 -2714
rect 6704 -2764 6784 -2730
rect 6844 -2757 6965 -2662
rect 7051 -2703 7075 -2669
rect 7091 -2677 7107 -2669
rect 7089 -2711 7113 -2677
rect 7213 -2695 7233 -2609
rect 6616 -2783 6662 -2773
rect 6704 -2780 6762 -2764
rect 6616 -2963 6668 -2783
rect 6716 -2795 6762 -2780
rect 6830 -2771 6965 -2757
rect 7045 -2771 7079 -2745
rect 7165 -2771 7167 -2745
rect 7174 -2771 7179 -2749
rect 7199 -2771 7233 -2695
rect 6676 -2811 6710 -2807
rect 6670 -2963 6710 -2811
rect 6716 -2963 6756 -2795
rect 6830 -2805 6948 -2771
rect 6979 -2805 6999 -2771
rect 7033 -2805 7179 -2771
rect 7213 -2805 7233 -2771
rect 7247 -2718 7286 -2609
rect 7300 -2556 7340 -2522
rect 7354 -2556 7500 -2522
rect 7568 -2556 7686 -2488
rect 7300 -2718 7334 -2556
rect 7354 -2578 7388 -2556
rect 7366 -2582 7368 -2578
rect 7420 -2650 7444 -2616
rect 7460 -2624 7476 -2616
rect 7458 -2658 7482 -2624
rect 7582 -2642 7686 -2556
rect 7414 -2718 7448 -2692
rect 7534 -2718 7536 -2692
rect 7543 -2718 7548 -2696
rect 7568 -2718 7686 -2642
rect 7954 -2612 8024 -2242
rect 8136 -2310 8194 -2304
rect 8136 -2344 8148 -2310
rect 8136 -2350 8194 -2344
rect 8136 -2510 8194 -2504
rect 8136 -2544 8148 -2510
rect 8136 -2550 8194 -2544
rect 7954 -2646 8025 -2612
rect 8325 -2627 8340 -2208
rect 8359 -2559 8393 -2189
rect 8505 -2257 8563 -2251
rect 8505 -2291 8517 -2257
rect 8505 -2297 8563 -2291
rect 8505 -2457 8563 -2451
rect 8505 -2491 8517 -2457
rect 8505 -2497 8563 -2491
rect 8359 -2593 8394 -2559
rect 8692 -2593 8762 -2138
rect 8874 -2204 8932 -2198
rect 8874 -2238 8886 -2204
rect 8874 -2244 8932 -2238
rect 8874 -2512 8932 -2506
rect 8874 -2546 8886 -2512
rect 8874 -2552 8932 -2546
rect 8692 -2629 8745 -2593
rect 9063 -2629 9078 -2042
rect 9097 -1079 9132 -1045
rect 9097 -1449 9131 -1079
rect 9243 -1147 9301 -1141
rect 9243 -1181 9255 -1147
rect 9413 -1170 9447 -1152
rect 9243 -1187 9301 -1181
rect 9413 -1206 9483 -1170
rect 9430 -1240 9501 -1206
rect 9199 -1408 9239 -1395
rect 9305 -1408 9345 -1395
rect 9430 -1396 9500 -1240
rect 9580 -1396 9614 -1376
rect 9668 -1396 9702 -1376
rect 9430 -1430 9501 -1396
rect 9568 -1430 9714 -1396
rect 9097 -1483 9132 -1449
rect 9228 -1460 9316 -1449
rect 9239 -1472 9305 -1460
rect 9228 -1483 9316 -1472
rect 9097 -1557 9131 -1483
rect 9243 -1489 9255 -1483
rect 9243 -1493 9301 -1489
rect 9239 -1505 9305 -1493
rect 9255 -1545 9289 -1523
rect 9430 -1545 9500 -1430
rect 9580 -1460 9614 -1430
rect 9668 -1460 9702 -1430
rect 9580 -1470 9702 -1460
rect 9580 -1474 9614 -1470
rect 9668 -1474 9702 -1470
rect 9612 -1498 9648 -1492
rect 9608 -1508 9674 -1498
rect 9624 -1532 9658 -1508
rect 9608 -1542 9674 -1532
rect 9243 -1551 9301 -1545
rect 9243 -1557 9255 -1551
rect 9097 -1591 9132 -1557
rect 9228 -1568 9316 -1557
rect 9239 -1578 9305 -1568
rect 9145 -1591 9399 -1578
rect 9097 -1645 9131 -1591
rect 9413 -1610 9500 -1545
rect 9612 -1548 9648 -1542
rect 9580 -1570 9614 -1566
rect 9668 -1570 9702 -1566
rect 9580 -1573 9626 -1570
rect 9656 -1573 9702 -1570
rect 9580 -1576 9620 -1573
rect 9580 -1610 9614 -1576
rect 9668 -1610 9702 -1573
rect 9211 -1645 9245 -1611
rect 9299 -1645 9333 -1611
rect 9413 -1644 9501 -1610
rect 9562 -1644 9714 -1610
rect 9720 -1644 9736 -1610
rect 9097 -1679 9132 -1645
rect 9193 -1679 9345 -1645
rect 9351 -1679 9367 -1645
rect 9097 -1961 9131 -1679
rect 9217 -1731 9245 -1709
rect 9289 -1731 9336 -1700
rect 9217 -1747 9257 -1731
rect 9287 -1747 9336 -1731
rect 9217 -1774 9336 -1747
rect 9199 -1812 9345 -1774
rect 9413 -1800 9500 -1644
rect 9782 -1738 9816 -1302
rect 9211 -1816 9245 -1812
rect 9299 -1816 9333 -1812
rect 9211 -1828 9245 -1824
rect 9299 -1828 9333 -1824
rect 9205 -1840 9251 -1828
rect 9289 -1840 9339 -1828
rect 9413 -1840 9501 -1800
rect 9562 -1840 9720 -1800
rect 9211 -1843 9245 -1840
rect 9289 -1843 9336 -1840
rect 9211 -1850 9257 -1843
rect 9217 -1859 9257 -1850
rect 9287 -1859 9336 -1843
rect 9217 -1893 9336 -1859
rect 9217 -1909 9257 -1893
rect 9287 -1909 9327 -1893
rect 9217 -1931 9245 -1909
rect 9299 -1931 9327 -1909
rect 9097 -1995 9132 -1961
rect 9199 -1995 9345 -1961
rect 9097 -2049 9131 -1995
rect 9199 -2008 9245 -1995
rect 9211 -2012 9245 -2008
rect 9299 -2008 9345 -1995
rect 9413 -1996 9500 -1840
rect 9580 -1996 9614 -1976
rect 9668 -1996 9702 -1976
rect 9299 -2012 9333 -2008
rect 9413 -2030 9501 -1996
rect 9568 -2030 9714 -1996
rect 9097 -2083 9132 -2049
rect 9228 -2060 9316 -2049
rect 9239 -2072 9305 -2060
rect 9228 -2083 9316 -2072
rect 9097 -2157 9131 -2083
rect 9243 -2089 9255 -2083
rect 9243 -2093 9301 -2089
rect 9239 -2105 9305 -2093
rect 9413 -2095 9500 -2030
rect 9580 -2060 9614 -2030
rect 9668 -2060 9702 -2030
rect 9580 -2070 9702 -2060
rect 9580 -2074 9614 -2070
rect 9668 -2074 9702 -2070
rect 9255 -2145 9289 -2123
rect 9243 -2151 9301 -2145
rect 9243 -2157 9255 -2151
rect 9097 -2191 9132 -2157
rect 9228 -2168 9316 -2157
rect 9239 -2178 9305 -2168
rect 9145 -2191 9399 -2178
rect 9097 -2561 9131 -2191
rect 9430 -2210 9500 -2095
rect 9608 -2108 9674 -2098
rect 9624 -2132 9658 -2108
rect 9608 -2142 9674 -2132
rect 9580 -2170 9614 -2166
rect 9668 -2170 9702 -2166
rect 9580 -2173 9626 -2170
rect 9656 -2173 9702 -2170
rect 9580 -2210 9614 -2173
rect 9668 -2210 9702 -2173
rect 9430 -2244 9501 -2210
rect 9562 -2244 9714 -2210
rect 9720 -2244 9736 -2210
rect 9430 -2400 9500 -2244
rect 9782 -2338 9816 -1902
rect 9430 -2434 9501 -2400
rect 9243 -2459 9301 -2453
rect 9243 -2493 9255 -2459
rect 9430 -2470 9483 -2434
rect 9243 -2499 9301 -2493
rect 9097 -2595 9132 -2561
rect 7767 -2671 7825 -2665
rect 7767 -2705 7779 -2671
rect 7954 -2682 8007 -2646
rect 7767 -2711 7825 -2705
rect 7247 -2752 7287 -2718
rect 7300 -2752 7315 -2718
rect 7348 -2752 7368 -2718
rect 7402 -2752 7548 -2718
rect 7582 -2752 7686 -2718
rect 6764 -2811 6784 -2807
rect 6758 -2823 6784 -2811
rect 6628 -2967 6630 -2963
rect 6642 -2967 6662 -2963
rect 6664 -2991 6752 -2963
rect 6758 -2979 6788 -2823
rect 6758 -2991 6784 -2979
rect 6676 -2995 6710 -2991
rect 6722 -2994 6746 -2991
rect 6764 -2995 6784 -2991
rect 6796 -2995 6798 -2807
rect 6805 -2991 6810 -2811
rect 6830 -2841 6965 -2805
rect 6830 -2991 6864 -2841
rect 6660 -3010 6718 -3004
rect 6656 -3029 6738 -3010
rect 6830 -3029 6832 -2991
rect 6682 -3044 6706 -3029
rect 6718 -3032 6738 -3029
rect 6722 -3038 6738 -3032
rect 6720 -3072 6744 -3038
rect 6844 -3046 6864 -2991
rect 6878 -2979 6965 -2841
rect 7045 -2843 7079 -2805
rect 7247 -2839 7281 -2752
rect 7077 -2877 7135 -2871
rect 7077 -2911 7089 -2877
rect 7077 -2917 7135 -2911
rect 6878 -3013 6966 -2979
rect 7266 -2994 7281 -2839
rect 7300 -2926 7334 -2752
rect 7414 -2790 7448 -2752
rect 7446 -2824 7504 -2818
rect 7446 -2858 7458 -2824
rect 7585 -2843 7686 -2752
rect 7446 -2864 7504 -2858
rect 7300 -2960 7335 -2926
rect 6878 -3046 6948 -3013
rect 6509 -3169 6549 -3112
rect 6610 -3135 6768 -3112
rect 6605 -3140 6768 -3135
rect 6605 -3169 6816 -3140
rect 6509 -3193 6543 -3169
rect 6562 -3174 6597 -3169
rect 6658 -3174 6816 -3169
rect 6236 -3222 6447 -3193
rect 6528 -3208 6543 -3193
rect 6289 -3227 6447 -3222
rect 6842 -3210 6948 -3046
rect 7024 -3184 7082 -3178
rect 6286 -3290 6344 -3284
rect 4664 -3328 5656 -3315
rect 4664 -3330 5632 -3328
rect 4664 -3387 4751 -3330
rect 5052 -3347 5067 -3330
rect 5086 -3334 5120 -3330
rect 5086 -3347 5121 -3334
rect 5182 -3347 5340 -3334
rect 5129 -3368 5340 -3347
rect 5735 -3351 5841 -3298
rect 5917 -3343 5975 -3337
rect 5129 -3381 5287 -3368
rect 4664 -3421 4752 -3387
rect 4664 -3457 4734 -3421
rect 4664 -3458 4698 -3457
rect 4396 -3464 4602 -3458
rect 4295 -3511 4329 -3464
rect 4348 -3492 4383 -3464
rect 4444 -3492 4602 -3464
rect 4027 -3517 4233 -3511
rect 3610 -3598 3645 -3564
rect 3945 -3579 3960 -3517
rect 3979 -3545 4014 -3517
rect 4075 -3545 4233 -3517
rect 4314 -3526 4329 -3511
rect 5179 -3739 5237 -3733
rect 5179 -3773 5191 -3739
rect 5179 -3779 5237 -3773
rect 5368 -3856 5383 -3368
rect 5402 -3788 5436 -3368
rect 5548 -3396 5606 -3390
rect 5548 -3430 5560 -3396
rect 5548 -3436 5606 -3430
rect 5548 -3686 5606 -3680
rect 5548 -3720 5560 -3686
rect 5548 -3726 5606 -3720
rect 5735 -3753 5805 -3351
rect 5917 -3377 5929 -3343
rect 5917 -3383 5975 -3377
rect 5917 -3651 5975 -3645
rect 5917 -3685 5929 -3651
rect 5917 -3691 5975 -3685
rect 5735 -3787 5806 -3753
rect 6106 -3768 6121 -3298
rect 6140 -3700 6174 -3298
rect 6286 -3324 6298 -3290
rect 6286 -3330 6344 -3324
rect 6286 -3598 6344 -3592
rect 6286 -3632 6298 -3598
rect 6286 -3638 6344 -3632
rect 6140 -3734 6175 -3700
rect 6475 -3715 6490 -3227
rect 6509 -3647 6543 -3227
rect 6655 -3237 6713 -3231
rect 6655 -3271 6667 -3237
rect 6655 -3277 6713 -3271
rect 6842 -3486 6912 -3210
rect 7024 -3218 7036 -3184
rect 7024 -3224 7082 -3218
rect 7024 -3384 7082 -3378
rect 7024 -3418 7036 -3384
rect 7024 -3424 7082 -3418
rect 6842 -3520 6913 -3486
rect 6655 -3545 6713 -3539
rect 6655 -3579 6667 -3545
rect 6842 -3556 6895 -3520
rect 6655 -3585 6713 -3579
rect 6509 -3681 6544 -3647
rect 5402 -3822 5437 -3788
rect 5735 -3823 5788 -3787
<< metal1 >>
rect 0 872 3964 910
rect 0 20 200 200
rect 0 -18 3964 20
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -929 3964 -891
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -1801 200 -1800
rect 0 -1839 3964 -1801
rect 0 -2000 200 -1839
rect 0 -2400 200 -2200
rect 0 -2692 200 -2600
rect 0 -2730 3964 -2692
rect 0 -2800 200 -2730
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
<< metal2 >>
rect 386 429 456 499
rect 1788 448 1858 518
rect 552 -206 622 383
rect 2478 303 2548 373
rect 3894 254 3964 324
rect 386 -276 622 -206
rect 386 -466 456 -276
rect 3894 -324 3964 -254
rect 552 -1251 622 -383
rect 386 -1321 622 -1251
rect 386 -1364 456 -1321
rect 552 -2018 622 -1458
rect 3894 -1566 3964 -1496
rect 386 -2088 622 -2018
rect 386 -2251 456 -2088
rect 3894 -2144 3964 -2074
use counter1b  counter1b_0
timestamp 1624053917
transform 1 0 1668 0 1 0
box -1809 -3600 8184 2091
use counter1b  counter1b_1
timestamp 1624053917
transform 1 0 1668 0 -1 0
box -1809 -3600 8184 2091
use counter1b  counter1b_2
timestamp 1624053917
transform 1 0 1668 0 1 -1820
box -1809 -3600 8184 2091
use counter1b  counter1b_3
timestamp 1624053917
transform 1 0 1668 0 -1 -1820
box -1809 -3600 8184 2091
use counter1b  xCOUNTER1B
timestamp 1624053917
transform 1 0 1668 0 1 600
box -1809 -3600 8184 2091
use counter1b  xCOUNTER1
timestamp 1624053917
transform 1 0 5632 0 1 600
box -1809 -3600 8184 2091
use counter1b  xCOUNTER2
timestamp 1624053917
transform 1 0 9596 0 1 600
box -1809 -3600 8184 2091
use counter1b  xCOUNTER3
timestamp 1624053917
transform 1 0 13560 0 1 600
box -1809 -3600 8184 2091
<< labels >>
rlabel metal2 420 429 420 429 5 CE
rlabel metal1 0 -2710 0 -2710 7 VDD
rlabel metal1 0 -1819 0 -1819 7 VSS
rlabel metal1 0 -907 0 -907 7 VDD
rlabel metal1 0 0 0 0 7 VSS
rlabel metal1 0 891 0 891 7 VDD
rlabel metal2 1823 448 1823 448 5 CLK
rlabel metal2 2513 303 2513 303 5 CLR
rlabel metal2 3929 254 3929 254 5 Q0
rlabel metal2 3930 -1566 3930 -1566 5 Q2
rlabel metal2 3929 -324 3929 -324 5 Q1
rlabel metal2 3929 -2144 3929 -2144 5 Q3
rlabel metal1 0 -2730 0 -2730 7 VDD
rlabel metal1 0 -929 0 -929 7 VDD
rlabel metal1 0 872 0 872 7 VDD
rlabel metal1 0 -18 0 -18 7 VSS
rlabel metal1 0 -1839 0 -1839 7 VSS
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 CE
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Q0
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLR
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLK
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Q1
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 Q2
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Q3
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 VSS
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 {}
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 VDD
port 11 nsew
<< end >>
