magic
tech sky130A
magscale 1 2
timestamp 1624331961
<< poly >>
rect -78 86 -6 102
rect -78 46 -62 86
rect -22 46 -6 86
rect -78 28 -6 46
rect -56 -99 -26 28
rect 88 -3100 118 -3084
rect 88 -3118 190 -3100
rect 88 -3152 122 -3118
rect 156 -3152 190 -3118
rect 88 -3168 190 -3152
rect 160 -3184 190 -3168
rect 88 -3882 190 -3866
rect 88 -3916 122 -3882
rect 156 -3916 190 -3882
rect 88 -3934 190 -3916
rect -56 -5074 -26 -4681
rect -74 -5090 -8 -5074
rect -74 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -74 -5140 -8 -5124
<< polycont >>
rect -62 46 -22 86
rect 122 -3152 156 -3118
rect 122 -3916 156 -3882
rect -58 -5124 -24 -5090
<< locali >>
rect -78 86 -6 102
rect -78 46 -62 86
rect -22 46 -6 86
rect -78 28 -6 46
rect 108 -3118 176 -3100
rect 108 -3152 122 -3118
rect 156 -3152 176 -3118
rect 108 -3168 176 -3152
rect 108 -3882 176 -3866
rect 108 -3916 122 -3882
rect 156 -3916 176 -3882
rect 108 -3934 176 -3916
rect -74 -5090 -8 -5074
rect -74 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -74 -5140 -8 -5124
<< viali >>
rect -62 46 -22 86
rect 122 -3152 156 -3118
rect 122 -3916 156 -3882
rect -58 -5124 -24 -5090
<< metal1 >>
rect -536 98 -10 99
rect -546 30 -536 98
rect -336 86 -10 98
rect -336 46 -62 86
rect -22 46 -10 86
rect -336 30 -10 46
rect 52 -1138 118 -1040
rect 52 -1190 62 -1138
rect 114 -1190 124 -1138
rect 52 -1286 118 -1190
rect -2698 -1764 -2688 -1526
rect -2428 -1531 -2418 -1526
rect -1846 -1531 -1836 -1526
rect -2428 -1760 -1836 -1531
rect -2428 -1764 -2418 -1760
rect -1846 -1764 -1836 -1760
rect -1576 -1764 -1566 -1526
rect -2288 -2134 -2278 -1896
rect -2018 -1901 -2008 -1896
rect -1836 -1901 -1826 -1894
rect -2018 -2130 -1826 -1901
rect -2018 -2134 -2008 -2130
rect -1836 -2132 -1826 -2130
rect -1566 -2132 -1556 -1894
rect -1842 -2496 -1832 -2258
rect -1572 -2262 -1562 -2258
rect -1572 -2263 -1132 -2262
rect -1572 -2491 -1348 -2263
rect -1572 -2496 -1562 -2491
rect -1358 -2492 -1348 -2491
rect -1119 -2492 -1109 -2263
rect -1842 -2888 -1832 -2650
rect -1572 -2659 -1562 -2650
rect -958 -2659 -948 -2657
rect -1572 -2886 -948 -2659
rect -719 -2886 -709 -2657
rect -1572 -2888 -736 -2886
rect -1842 -3314 -1832 -3076
rect -1572 -3081 -1562 -3076
rect -1572 -3310 -550 -3081
rect -321 -3310 -311 -3081
rect 108 -3104 176 -3102
rect 98 -3164 108 -3104
rect 168 -3164 178 -3104
rect 108 -3168 176 -3164
rect -1572 -3314 -1562 -3310
rect 52 -3484 118 -3386
rect 52 -3536 64 -3484
rect 116 -3536 126 -3484
rect 52 -3632 118 -3536
rect 108 -3870 176 -3866
rect 98 -3930 108 -3870
rect 168 -3930 178 -3870
rect 108 -3932 176 -3930
rect -546 -5140 -536 -5074
rect -336 -5090 -8 -5074
rect -336 -5124 -58 -5090
rect -24 -5124 -8 -5090
rect -336 -5140 -8 -5124
rect -2260 -5328 -2250 -5264
rect -2050 -5284 -2040 -5264
rect -2050 -5317 518 -5284
rect -2050 -5328 -2040 -5317
rect 346 -5368 518 -5317
rect 90 -5510 164 -5508
rect -1344 -5562 -1334 -5510
rect -1134 -5562 164 -5510
rect 90 -5564 164 -5562
rect 228 -5564 238 -5508
rect -2664 -6178 -2654 -6118
rect -2454 -6124 -2444 -6118
rect -2454 -6170 -104 -6124
rect -2454 -6178 -2444 -6170
rect -942 -6656 -932 -6596
rect -732 -6656 -182 -6596
rect -122 -6656 -112 -6596
rect -2258 -6974 -2248 -6916
rect -2050 -6919 -2040 -6916
rect -2050 -6922 -198 -6919
rect -2050 -6968 -66 -6922
rect -2050 -6970 -198 -6968
rect -2050 -6974 -2040 -6970
<< via1 >>
rect -536 30 -336 98
rect 62 -1190 114 -1138
rect -2688 -1764 -2428 -1526
rect -1836 -1764 -1576 -1526
rect -2278 -2134 -2018 -1896
rect -1826 -2132 -1566 -1894
rect -1832 -2496 -1572 -2258
rect -1348 -2492 -1119 -2263
rect -1832 -2888 -1572 -2650
rect -948 -2886 -719 -2657
rect -1832 -3314 -1572 -3076
rect -550 -3310 -321 -3081
rect 108 -3118 168 -3104
rect 108 -3152 122 -3118
rect 122 -3152 156 -3118
rect 156 -3152 168 -3118
rect 108 -3164 168 -3152
rect 64 -3536 116 -3484
rect 108 -3882 168 -3870
rect 108 -3916 122 -3882
rect 122 -3916 156 -3882
rect 156 -3916 168 -3882
rect 108 -3930 168 -3916
rect -536 -5140 -336 -5074
rect -2250 -5328 -2050 -5264
rect -1334 -5562 -1134 -5510
rect 164 -5564 228 -5508
rect -2654 -6178 -2454 -6118
rect -932 -6656 -732 -6596
rect -182 -6656 -122 -6596
rect -2248 -6974 -2050 -6916
<< metal2 >>
rect -2652 -1516 -2452 6040
rect -2688 -1526 -2428 -1516
rect -2688 -1774 -2428 -1764
rect -2652 -6108 -2452 -1774
rect -2250 -1886 -2050 6040
rect -1334 -1134 -1134 6084
rect -1836 -1526 -1576 -1516
rect -1836 -1774 -1576 -1764
rect -2278 -1896 -2018 -1886
rect -2278 -2144 -2018 -2134
rect -1826 -1894 -1566 -1884
rect -1826 -2142 -1566 -2132
rect -2654 -6118 -2452 -6108
rect -2454 -6178 -2452 -6118
rect -2654 -6188 -2452 -6178
rect -2652 -6960 -2452 -6188
rect -2250 -5264 -2050 -2144
rect -1832 -2258 -1572 -2248
rect -1334 -2253 -1134 -1194
rect -1832 -2506 -1572 -2496
rect -1348 -2263 -1119 -2253
rect -1348 -2502 -1119 -2492
rect -1832 -2650 -1572 -2640
rect -1832 -2898 -1572 -2888
rect -1832 -3076 -1572 -3066
rect -1832 -3324 -1572 -3314
rect -2250 -6916 -2050 -5328
rect -1334 -3480 -1134 -2502
rect -932 -2647 -732 6084
rect -536 98 -336 6056
rect 8550 5836 8808 5846
rect 8808 5600 8812 5836
rect 8550 5598 8812 5600
rect 9138 5834 9398 5844
rect 8550 5590 8808 5598
rect 9138 5592 9398 5602
rect 9670 5832 9928 5842
rect 9928 5596 9930 5832
rect 9670 5594 9930 5596
rect 9670 5586 9928 5594
rect 17278 3224 17770 3294
rect 17510 3056 17770 3224
rect 6825 2558 6890 2560
rect 7717 2558 7777 2568
rect 12192 2558 12252 2568
rect 6824 2498 7717 2558
rect 7777 2498 12192 2558
rect -948 -2657 -719 -2647
rect -948 -2896 -719 -2886
rect -1334 -5510 -1134 -3540
rect -1334 -6916 -1134 -5562
rect -932 -2948 -732 -2896
rect -932 -3870 -732 -3006
rect -536 -3071 -336 30
rect 58 -1134 118 -1124
rect 58 -1204 118 -1194
rect 6825 -1604 6890 2498
rect 7717 2488 7777 2498
rect 12192 2488 12252 2498
rect 8244 2432 8304 2440
rect 12717 2432 12777 2442
rect 8244 2430 12717 2432
rect 8304 2372 12717 2430
rect 8244 2360 8304 2370
rect 12717 2362 12777 2372
rect 9220 2316 9280 2326
rect 13654 2316 13714 2326
rect 9280 2256 13654 2316
rect 9220 2246 9280 2256
rect 13654 2246 13714 2256
rect 9754 2198 9814 2208
rect 14170 2198 14230 2208
rect 9814 2138 14170 2198
rect 9754 2128 9814 2138
rect 14170 2128 14230 2138
rect 17256 936 17748 1006
rect 17488 768 17748 936
rect 7694 276 7754 286
rect 12170 276 12230 286
rect 6658 -1669 6890 -1604
rect 6968 216 7694 276
rect 7754 216 12170 276
rect -550 -3081 -321 -3071
rect 108 -3104 168 -3094
rect 108 -3174 168 -3164
rect -550 -3320 -321 -3310
rect -932 -6596 -732 -3930
rect -932 -6916 -732 -6656
rect -536 -5074 -336 -3320
rect 60 -3480 120 -3470
rect 60 -3550 120 -3540
rect 108 -3870 168 -3860
rect 108 -3940 168 -3930
rect 2768 -5009 2828 -5002
rect 6658 -5009 6723 -1669
rect 6968 -1792 7028 216
rect 7694 206 7754 216
rect 12170 206 12230 216
rect 8222 144 8282 152
rect 12695 144 12755 154
rect 8222 142 12695 144
rect 8282 84 12695 142
rect 8222 72 8282 82
rect 12695 74 12755 84
rect 9198 28 9258 38
rect 13632 28 13692 38
rect 9258 -32 13632 28
rect 9198 -42 9258 -32
rect 13632 -42 13692 -32
rect 9732 -90 9792 -80
rect 14148 -90 14208 -80
rect 9792 -150 14148 -90
rect 9732 -160 9792 -150
rect 14148 -160 14208 -150
rect 17240 -1428 17732 -1358
rect 17472 -1596 17732 -1428
rect 2766 -5012 6723 -5009
rect 2766 -5072 2768 -5012
rect 2828 -5072 6723 -5012
rect 6802 -1852 7028 -1792
rect 6802 -4998 6870 -1852
rect 7679 -1982 7739 -1972
rect 6802 -5058 6806 -4998
rect 6866 -5058 6870 -4998
rect 6802 -5060 6870 -5058
rect 6960 -2042 7679 -1984
rect 12154 -1984 12214 -1974
rect 7739 -2042 12154 -1984
rect 6960 -2044 12154 -2042
rect 6806 -5068 6866 -5060
rect 2766 -5074 6723 -5072
rect 2768 -5082 2828 -5074
rect -536 -5369 -336 -5140
rect 4502 -5134 4562 -5124
rect 6960 -5134 7020 -2044
rect 7679 -2052 7739 -2044
rect 12154 -2054 12214 -2044
rect 8206 -2118 8266 -2110
rect 12679 -2118 12739 -2108
rect 8206 -2120 12679 -2118
rect 8266 -2178 12679 -2120
rect 8206 -2190 8266 -2180
rect 12679 -2188 12739 -2178
rect 9182 -2234 9242 -2224
rect 13616 -2234 13676 -2224
rect 9242 -2294 13616 -2234
rect 9182 -2304 9242 -2294
rect 13616 -2304 13676 -2294
rect 9716 -2352 9776 -2342
rect 14132 -2352 14192 -2342
rect 9776 -2412 14132 -2352
rect 9716 -2422 9776 -2412
rect 14132 -2422 14192 -2412
rect 8568 -2850 8790 -2840
rect 8568 -2928 8790 -2918
rect 16024 -2992 16104 -2982
rect 16024 -3082 16104 -3072
rect 17250 -3616 17740 -3546
rect 17480 -3784 17740 -3616
rect 7687 -4290 7747 -4280
rect 12162 -4290 12222 -4280
rect 7396 -4350 7687 -4290
rect 7747 -4350 12162 -4290
rect 4562 -5194 7020 -5134
rect 7397 -4360 7460 -4350
rect 7687 -4360 7747 -4350
rect 12162 -4360 12222 -4350
rect 4502 -5204 4562 -5194
rect 738 -5256 798 -5246
rect 7397 -5254 7457 -4360
rect 8214 -4408 8274 -4400
rect 12687 -4408 12747 -4398
rect 8214 -4410 12687 -4408
rect 8274 -4468 12687 -4410
rect 8214 -4480 8274 -4470
rect 12687 -4478 12747 -4468
rect 9190 -4524 9250 -4514
rect 13624 -4524 13684 -4514
rect 9250 -4584 13624 -4524
rect 9190 -4594 9250 -4584
rect 13624 -4594 13684 -4584
rect 9724 -4642 9784 -4632
rect 14140 -4642 14200 -4632
rect 9784 -4702 14140 -4642
rect 9724 -4712 9784 -4702
rect 14140 -4712 14200 -4702
rect 7396 -5256 7458 -5254
rect 798 -5316 7458 -5256
rect 738 -5326 798 -5316
rect -536 -5397 204 -5369
rect -2250 -6960 -2248 -6916
rect -536 -6944 -336 -5397
rect 164 -5508 228 -5498
rect 164 -5574 228 -5564
rect 738 -5720 798 -5710
rect 738 -5790 798 -5780
rect 4500 -5718 4560 -5708
rect 4500 -5788 4560 -5778
rect 2768 -6512 2828 -6502
rect 2768 -6582 2828 -6572
rect 6534 -6514 6594 -6504
rect 6534 -6584 6594 -6574
rect -182 -6596 -122 -6586
rect -122 -6640 -30 -6612
rect -182 -6666 -122 -6656
rect -2248 -6984 -2050 -6974
<< via2 >>
rect -1334 -1194 -1134 -1134
rect 8550 5600 8808 5836
rect 9138 5602 9398 5834
rect 9670 5596 9928 5832
rect 7717 2498 7777 2558
rect 12192 2498 12252 2558
rect -1334 -3540 -1134 -3480
rect -932 -3006 -732 -2948
rect 58 -1138 118 -1134
rect 58 -1190 62 -1138
rect 62 -1190 114 -1138
rect 114 -1190 118 -1138
rect 58 -1194 118 -1190
rect 8244 2370 8304 2430
rect 12717 2372 12777 2432
rect 9220 2256 9280 2316
rect 13654 2256 13714 2316
rect 9754 2138 9814 2198
rect 14170 2138 14230 2198
rect 7694 216 7754 276
rect 12170 216 12230 276
rect 108 -3164 168 -3104
rect -932 -3930 -732 -3870
rect 60 -3484 120 -3480
rect 60 -3536 64 -3484
rect 64 -3536 116 -3484
rect 116 -3536 120 -3484
rect 60 -3540 120 -3536
rect 108 -3930 168 -3870
rect 8222 82 8282 142
rect 12695 84 12755 144
rect 9198 -32 9258 28
rect 13632 -32 13692 28
rect 9732 -150 9792 -90
rect 14148 -150 14208 -90
rect 2768 -5072 2828 -5012
rect 6806 -5058 6866 -4998
rect 7679 -2042 7739 -1982
rect 12154 -2044 12214 -1984
rect 8206 -2180 8266 -2120
rect 12679 -2178 12739 -2118
rect 9182 -2294 9242 -2234
rect 13616 -2294 13676 -2234
rect 9716 -2412 9776 -2352
rect 14132 -2412 14192 -2352
rect 8568 -2918 8790 -2850
rect 16024 -3072 16104 -2992
rect 7687 -4350 7747 -4290
rect 12162 -4350 12222 -4290
rect 4502 -5194 4562 -5134
rect 8214 -4470 8274 -4410
rect 12687 -4468 12747 -4408
rect 9190 -4584 9250 -4524
rect 13624 -4584 13684 -4524
rect 9724 -4702 9784 -4642
rect 14140 -4702 14200 -4642
rect 738 -5316 798 -5256
rect 738 -5780 798 -5720
rect 4500 -5778 4560 -5718
rect 2768 -6572 2828 -6512
rect 6534 -6574 6594 -6514
<< metal3 >>
rect 8540 5836 8818 5841
rect 8540 5600 8550 5836
rect 8808 5600 8818 5836
rect 8540 5595 8818 5600
rect 9128 5834 9408 5839
rect 9128 5602 9138 5834
rect 9398 5602 9408 5834
rect 9128 5597 9408 5602
rect 9660 5832 9938 5837
rect 9660 5596 9670 5832
rect 9928 5596 9938 5832
rect 9660 5591 9938 5596
rect 7717 2563 7777 2671
rect 7707 2558 7787 2563
rect 7707 2498 7717 2558
rect 7777 2498 7787 2558
rect 7707 2493 7787 2498
rect 8246 2435 8306 2722
rect 8234 2430 8314 2435
rect 8234 2370 8244 2430
rect 8304 2370 8314 2430
rect 8234 2365 8314 2370
rect 9223 2321 9283 2602
rect 9210 2316 9290 2321
rect 9210 2256 9220 2316
rect 9280 2256 9290 2316
rect 9210 2251 9290 2256
rect 9756 2203 9816 2608
rect 12182 2558 12262 2563
rect 12182 2498 12192 2558
rect 12252 2498 12262 2558
rect 12182 2493 12262 2498
rect 12717 2437 12777 2580
rect 12707 2432 12787 2437
rect 12707 2372 12717 2432
rect 12777 2372 12787 2432
rect 12707 2367 12787 2372
rect 13657 2321 13717 2638
rect 13644 2316 13724 2321
rect 13644 2256 13654 2316
rect 13714 2256 13724 2316
rect 13644 2251 13724 2256
rect 14172 2203 14232 2802
rect 9744 2198 9824 2203
rect 9744 2138 9754 2198
rect 9814 2138 9824 2198
rect 9744 2133 9824 2138
rect 14160 2198 14240 2203
rect 14160 2138 14170 2198
rect 14230 2138 14240 2198
rect 14160 2133 14240 2138
rect 7695 281 7755 428
rect 7684 276 7764 281
rect 7684 216 7694 276
rect 7754 216 7764 276
rect 7684 211 7764 216
rect 8224 147 8284 424
rect 8212 142 8292 147
rect 8212 82 8222 142
rect 8282 82 8292 142
rect 8212 77 8292 82
rect 9201 33 9261 298
rect 9188 28 9268 33
rect 9188 -32 9198 28
rect 9258 -32 9268 28
rect 9188 -37 9268 -32
rect 9734 -85 9794 296
rect 12160 276 12240 281
rect 12160 216 12170 276
rect 12230 216 12240 276
rect 12160 211 12240 216
rect 12695 149 12755 294
rect 12685 144 12765 149
rect 12685 84 12695 144
rect 12755 84 12765 144
rect 12685 79 12765 84
rect 13635 33 13695 366
rect 13622 28 13702 33
rect 13622 -32 13632 28
rect 13692 -32 13702 28
rect 13622 -37 13702 -32
rect 14150 -85 14210 510
rect 9722 -90 9802 -85
rect 9722 -150 9732 -90
rect 9792 -150 9802 -90
rect 9722 -155 9802 -150
rect 14138 -90 14218 -85
rect 14138 -150 14148 -90
rect 14208 -150 14218 -90
rect 14138 -155 14218 -150
rect -1344 -1134 -1124 -1129
rect 48 -1134 128 -1129
rect -1344 -1194 -1334 -1134
rect -1134 -1194 58 -1134
rect 118 -1194 128 -1134
rect -1344 -1199 -1124 -1194
rect 48 -1199 128 -1194
rect 7679 -1977 7739 -1842
rect 7669 -1982 7749 -1977
rect 7669 -2042 7679 -1982
rect 7739 -2042 7749 -1982
rect 7669 -2047 7749 -2042
rect 8208 -2115 8268 -1836
rect 8196 -2120 8276 -2115
rect 8196 -2180 8206 -2120
rect 8266 -2180 8276 -2120
rect 8196 -2185 8276 -2180
rect 9185 -2229 9245 -1956
rect 12144 -1984 12224 -1979
rect 9172 -2234 9252 -2229
rect 9172 -2294 9182 -2234
rect 9242 -2294 9252 -2234
rect 9172 -2299 9252 -2294
rect 9718 -2347 9778 -1994
rect 12144 -2044 12154 -1984
rect 12214 -2044 12224 -1984
rect 12144 -2049 12224 -2044
rect 12679 -2113 12739 -1982
rect 12669 -2118 12749 -2113
rect 12669 -2178 12679 -2118
rect 12739 -2178 12749 -2118
rect 12669 -2183 12749 -2178
rect 13619 -2229 13679 -1906
rect 13606 -2234 13686 -2229
rect 13606 -2294 13616 -2234
rect 13676 -2294 13686 -2234
rect 13606 -2299 13686 -2294
rect 14134 -2347 14194 -1722
rect 9706 -2352 9786 -2347
rect 9706 -2412 9716 -2352
rect 9776 -2412 9786 -2352
rect 9706 -2417 9786 -2412
rect 14122 -2352 14202 -2347
rect 14122 -2412 14132 -2352
rect 14192 -2412 14202 -2352
rect 14122 -2417 14202 -2412
rect 9682 -2782 9692 -2702
rect 9926 -2782 16104 -2702
rect 8558 -2850 8800 -2845
rect 8558 -2918 8568 -2850
rect 8790 -2918 8800 -2850
rect 8558 -2923 8800 -2918
rect 9136 -2920 9146 -2850
rect 9382 -2851 9392 -2850
rect 10129 -2851 10215 -2848
rect 9382 -2911 10260 -2851
rect 9382 -2920 9392 -2911
rect -942 -2946 -722 -2943
rect -942 -2948 160 -2946
rect -942 -3006 -932 -2948
rect -732 -3006 160 -2948
rect -942 -3011 -722 -3006
rect 88 -3099 160 -3006
rect 88 -3104 178 -3099
rect 88 -3164 108 -3104
rect 168 -3164 178 -3104
rect 10129 -3149 10215 -2911
rect 16024 -2987 16104 -2782
rect 16014 -2992 16114 -2987
rect 16014 -3072 16024 -2992
rect 16104 -3072 16114 -2992
rect 16014 -3077 16114 -3072
rect 88 -3168 178 -3164
rect 98 -3169 178 -3168
rect -1344 -3480 -1124 -3475
rect 50 -3480 130 -3475
rect -1344 -3540 -1334 -3480
rect -1134 -3540 60 -3480
rect 120 -3540 130 -3480
rect -1344 -3545 -1124 -3540
rect 50 -3545 130 -3540
rect -937 -3870 -727 -3865
rect 98 -3870 178 -3865
rect -937 -3930 -932 -3870
rect -732 -3930 108 -3870
rect 168 -3930 178 -3870
rect -937 -3935 -727 -3930
rect 98 -3935 178 -3930
rect 7687 -4285 7747 -4161
rect 7677 -4290 7757 -4285
rect 7677 -4350 7687 -4290
rect 7747 -4350 7757 -4290
rect 7677 -4355 7757 -4350
rect 8216 -4405 8276 -4171
rect 8204 -4410 8284 -4405
rect 8204 -4470 8214 -4410
rect 8274 -4470 8284 -4410
rect 8204 -4475 8284 -4470
rect 9193 -4519 9253 -4254
rect 9180 -4524 9260 -4519
rect 9180 -4584 9190 -4524
rect 9250 -4584 9260 -4524
rect 9180 -4589 9260 -4584
rect 9726 -4637 9786 -4254
rect 12152 -4290 12232 -4285
rect 12152 -4350 12162 -4290
rect 12222 -4350 12232 -4290
rect 12152 -4355 12232 -4350
rect 12687 -4403 12747 -4272
rect 12677 -4408 12757 -4403
rect 12677 -4468 12687 -4408
rect 12747 -4468 12757 -4408
rect 12677 -4473 12757 -4468
rect 13627 -4519 13687 -4132
rect 13614 -4524 13694 -4519
rect 13614 -4584 13624 -4524
rect 13684 -4584 13694 -4524
rect 13614 -4589 13694 -4584
rect 14142 -4637 14202 -4009
rect 9714 -4642 9794 -4637
rect 9714 -4702 9724 -4642
rect 9784 -4702 9794 -4642
rect 9714 -4707 9794 -4702
rect 14130 -4642 14210 -4637
rect 14130 -4702 14140 -4642
rect 14200 -4702 14210 -4642
rect 14130 -4707 14210 -4702
rect 6796 -4998 6876 -4993
rect 2758 -5012 2838 -5007
rect 2758 -5072 2768 -5012
rect 2828 -5072 2838 -5012
rect 6796 -5058 6806 -4998
rect 6866 -5058 6876 -4998
rect 6796 -5063 6876 -5058
rect 2758 -5077 2838 -5072
rect 728 -5256 808 -5251
rect 728 -5316 738 -5256
rect 798 -5316 808 -5256
rect 728 -5321 808 -5316
rect 738 -5715 798 -5321
rect 728 -5720 808 -5715
rect 728 -5780 738 -5720
rect 798 -5780 808 -5720
rect 728 -5785 808 -5780
rect 2766 -6507 2831 -5077
rect 4502 -5129 4562 -5118
rect 4492 -5134 4572 -5129
rect 4492 -5194 4502 -5134
rect 4562 -5194 4572 -5134
rect 4492 -5199 4572 -5194
rect 4502 -5713 4562 -5199
rect 4490 -5718 4570 -5713
rect 4490 -5778 4500 -5718
rect 4560 -5778 4570 -5718
rect 4490 -5783 4570 -5778
rect 2758 -6512 2838 -6507
rect 2758 -6572 2768 -6512
rect 2828 -6572 2838 -6512
rect 2758 -6577 2838 -6572
rect 6524 -6510 6604 -6509
rect 6802 -6510 6870 -5063
rect 6524 -6514 6870 -6510
rect 6524 -6574 6534 -6514
rect 6594 -6574 6870 -6514
rect 2766 -6578 2831 -6577
rect 6524 -6578 6870 -6574
rect 6524 -6579 6604 -6578
<< via3 >>
rect 8550 5600 8808 5836
rect 9138 5602 9398 5834
rect 9670 5596 9928 5832
rect 9692 -2782 9926 -2702
rect 8568 -2918 8790 -2850
rect 9146 -2920 9382 -2850
<< metal4 >>
rect 8549 5836 8809 5837
rect 8549 5600 8550 5836
rect 8808 5600 8809 5836
rect 9137 5834 9399 5835
rect 9137 5606 9138 5834
rect 8549 5599 8809 5600
rect 9136 5602 9138 5606
rect 9398 5602 9399 5834
rect 9136 5601 9399 5602
rect 9669 5832 9929 5833
rect 8552 5378 8808 5599
rect 8571 -2849 8790 5378
rect 9136 5366 9396 5601
rect 9669 5596 9670 5832
rect 9928 5596 9929 5832
rect 9669 5595 9940 5596
rect 9146 -2849 9382 5366
rect 9670 5362 9940 5595
rect 9691 -2701 9925 5362
rect 9691 -2702 9927 -2701
rect 9691 -2782 9692 -2702
rect 9926 -2782 9927 -2702
rect 9691 -2783 9927 -2782
rect 8567 -2850 8791 -2849
rect 8567 -2918 8568 -2850
rect 8790 -2918 8791 -2850
rect 8567 -2919 8791 -2918
rect 9145 -2850 9383 -2849
rect 8571 -2943 8790 -2919
rect 9145 -2920 9146 -2850
rect 9382 -2920 9383 -2850
rect 9145 -2921 9383 -2920
rect 9146 -2936 9382 -2921
rect 9691 -2941 9925 -2783
use contador  contador_0
timestamp 1624067212
transform 1 0 -206 0 1 -6968
box 0 0 7741 1645
use mux_8to1  mux_8to1_2
timestamp 1624074478
transform 1 0 7154 0 1 -3114
box -54 1072 10324 2553
use c4b  c4b_0
timestamp 1624067212
transform 1 0 -56 0 1 -2384
box -120 -2346 3972 2370
use mux_8to1  mux_8to1_0
timestamp 1624074478
transform 1 0 7192 0 1 1436
box -54 1072 10324 2553
use mux_8to1  mux_8to1_1
timestamp 1624074478
transform 1 0 7170 0 1 -852
box -54 1072 10324 2553
use mux_8to1  mux_8to1_3
timestamp 1624074478
transform 1 0 7162 0 1 -5404
box -54 1072 10324 2553
use contador4bits  contador4bits_0
timestamp 1624067212
transform 1 0 -64 0 1 4130
box -56 0 6948 1980
use 4bitc  4bitc_0
timestamp 1624067212
transform 1 0 -63 0 1 1939
box -107 -1605 5377 1735
<< labels >>
rlabel metal2 8552 5598 8812 5836 1 reg2
rlabel metal2 9138 5598 9398 5836 1 reg1
rlabel metal2 9670 5594 9930 5832 1 reg0
rlabel metal2 -1826 -2132 -1566 -1894 1 VSS
rlabel metal2 -1832 -2890 -1572 -2652 1 CE
rlabel metal2 -1832 -2496 -1572 -2258 1 CLK
rlabel metal2 -1836 -1764 -1576 -1526 1 VDD
rlabel metal2 -1832 -3314 -1572 -3076 1 CLR
rlabel poly 132 -3154 190 -3118 1 ce
rlabel metal2 17488 768 17748 1006 1 Q1
rlabel metal2 17472 -1596 17732 -1358 1 Q2
rlabel metal2 17480 -3784 17740 -3546 1 Q3
rlabel metal2 17510 3056 17770 3294 1 Q0
<< end >>
